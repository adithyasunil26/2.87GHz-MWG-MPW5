magic
tech sky130A
timestamp 1640957100
<< nwell >>
rect 965 1061 1081 1192
rect 965 1036 1082 1061
rect 997 760 1073 1036
rect 995 743 1073 760
rect 201 527 277 721
rect 195 459 277 527
rect 195 271 271 459
rect 195 265 353 271
rect 208 260 353 265
rect 995 260 1035 743
<< locali >>
rect 225 1285 245 1310
rect 990 1090 1010 1380
rect 1350 1135 1430 1155
rect 990 1065 1025 1090
rect 1410 1015 1430 1135
rect -155 185 -135 330
rect -155 165 -80 185
rect 225 160 245 255
rect 1015 210 1055 235
rect 1795 210 1825 235
rect 225 140 255 160
rect 1035 140 1055 210
rect 1805 80 1825 210
<< viali >>
rect 200 1285 225 1310
rect 1410 995 1430 1015
rect -155 330 -135 350
rect 1060 140 1080 160
rect 1805 60 1825 80
<< metal1 >>
rect 190 1310 235 1320
rect -155 1295 200 1310
rect -155 360 -140 1295
rect 190 1285 200 1295
rect 225 1285 235 1310
rect 190 1275 235 1285
rect 1350 1095 1795 1110
rect 1400 1015 1440 1025
rect 1400 995 1410 1015
rect 1430 995 1440 1015
rect 1400 985 1440 995
rect 140 770 160 775
rect 130 765 170 770
rect 130 735 135 765
rect 165 755 170 765
rect 1415 755 1430 985
rect 165 740 1430 755
rect 165 735 170 740
rect 130 730 170 735
rect -165 350 -125 360
rect -165 330 -155 350
rect -135 330 -125 350
rect -165 325 -125 330
rect -155 210 -80 225
rect -155 160 -135 210
rect 1050 165 1090 170
rect -165 155 -125 160
rect -165 125 -160 155
rect -130 125 -125 155
rect 1050 135 1055 165
rect 1085 135 1090 165
rect 1780 140 1795 1095
rect 1050 130 1090 135
rect -165 120 -125 125
rect 1795 85 1835 90
rect 1795 55 1800 85
rect 1830 55 1835 85
rect 1795 50 1835 55
<< via1 >>
rect 135 735 165 765
rect -160 125 -130 155
rect 1055 160 1085 165
rect 1055 140 1060 160
rect 1060 140 1080 160
rect 1080 140 1085 160
rect 1055 135 1085 140
rect 1800 80 1830 85
rect 1800 60 1805 80
rect 1805 60 1825 80
rect 1825 60 1830 80
rect 1800 55 1830 60
<< metal2 >>
rect 125 765 175 775
rect 125 755 135 765
rect -210 740 135 755
rect 125 735 135 740
rect 165 735 175 765
rect 125 725 175 735
rect 995 250 1010 1290
rect -210 230 255 250
rect 485 230 1035 250
rect 1045 165 1095 175
rect -170 155 -120 165
rect -170 125 -160 155
rect -130 125 -120 155
rect 1045 135 1055 165
rect 1085 155 1095 165
rect 1085 140 1930 155
rect 1085 135 1095 140
rect 1045 125 1095 135
rect -170 115 -120 125
rect -155 80 -135 115
rect 1790 85 1840 95
rect 1790 80 1800 85
rect -155 60 1800 80
rect 1790 55 1800 60
rect 1830 55 1840 85
rect 1790 45 1840 55
<< metal4 >>
rect 965 1675 1085 1705
rect 1050 1330 1085 1675
rect 1300 1330 1890 1360
rect 175 730 285 790
rect 990 730 1075 790
rect 1365 760 1775 790
rect 175 530 220 730
rect 195 -155 225 -10
rect 1860 -155 1890 1330
rect 195 -160 265 -155
rect 195 -185 270 -160
rect 985 -185 1055 -155
rect 1750 -185 1890 -155
use nand  nand_1
timestamp 1640957032
transform -1 0 1325 0 -1 1050
box -40 -310 300 315
use nand  nand_0
timestamp 1640957032
transform 1 0 -55 0 1 270
box -40 -310 300 315
use tspc  tspc_0
timestamp 1640956963
transform 1 0 325 0 1 295
box -70 -490 690 465
use tspc  tspc_1
timestamp 1640956963
transform 1 0 1105 0 1 295
box -70 -490 690 465
use tspc  tspc_2
timestamp 1640956963
transform -1 0 935 0 -1 1225
box -70 -490 690 465
<< labels >>
rlabel metal2 -210 740 170 755 1 mc1
rlabel metal1 170 740 1430 755 1 mc1
rlabel metal1 1415 740 1430 1015 1 mc1
rlabel metal2 -210 230 255 250 1 clk
rlabel space 255 230 1035 250 1 clk
rlabel metal2 1055 140 1930 155 1 Out
rlabel metal4 1050 1360 1085 1705 1 GND
rlabel metal4 1345 1330 1890 1360 1 GND
rlabel metal4 1860 -185 1890 1330 1 GND
rlabel metal4 1750 -185 1860 -155 1 GND
rlabel space 985 -185 1060 -155 1 GND
rlabel metal4 195 -185 225 -40 1 GND
rlabel space 195 -185 270 -155 1 GND
rlabel metal4 220 -40 225 -10 1 GND
rlabel space 175 560 225 795 1 VDD
rlabel space 175 730 295 790 1 VDD
rlabel metal4 990 730 1070 790 1 VDD
<< end >>
