magic
tech sky130A
magscale 1 2
timestamp 1647888148
<< nwell >>
rect 560 910 7640 2090
rect 1790 -2020 7640 -810
<< nmos >>
rect 90 160 120 660
rect 320 160 350 660
rect 550 160 580 660
rect 780 160 810 660
rect 1010 160 1040 660
rect 1240 160 1270 660
rect 1470 160 1500 660
rect 1700 160 1730 660
rect 1930 160 1960 660
rect 2160 160 2190 660
rect 2390 160 2420 660
rect 2620 160 2650 660
rect 2850 160 2880 660
rect 3080 160 3110 660
rect 3310 160 3340 660
rect 3540 160 3570 660
rect 3770 160 3800 660
rect 4000 160 4030 660
rect 4230 160 4260 660
rect 4460 160 4490 660
rect 4690 160 4720 660
rect 4920 160 4950 660
rect 5150 160 5180 660
rect 5380 160 5410 660
rect 5610 160 5640 660
rect 5840 160 5870 660
rect 6070 160 6100 660
rect 6300 160 6330 660
rect 6530 160 6560 660
rect 6760 160 6790 660
rect 90 -550 120 -50
rect 320 -550 350 -50
rect 550 -550 580 -50
rect 780 -550 810 -50
rect 1010 -550 1040 -50
rect 1240 -550 1270 -50
rect 1470 -550 1500 -50
rect 1700 -550 1730 -50
rect 1930 -550 1960 -50
rect 2160 -550 2190 -50
rect 2390 -550 2420 -50
rect 2620 -550 2650 -50
rect 2850 -550 2880 -50
rect 3080 -550 3110 -50
rect 3310 -550 3340 -50
rect 3540 -550 3570 -50
rect 3770 -550 3800 -50
rect 4000 -550 4030 -50
rect 4230 -550 4260 -50
rect 4460 -550 4490 -50
rect 4690 -550 4720 -50
rect 4920 -550 4950 -50
rect 5150 -550 5180 -50
rect 5380 -550 5410 -50
rect 5610 -550 5640 -50
rect 5840 -550 5870 -50
rect 6070 -550 6100 -50
rect 6300 -550 6330 -50
rect 6530 -550 6560 -50
rect 6760 -550 6790 -50
<< pmos >>
rect 1550 1220 1610 1760
rect 1810 1220 1870 1760
rect 2340 1160 2400 1760
rect 2600 1160 2660 1760
rect 2860 1160 2920 1760
rect 3120 1160 3180 1760
rect 3380 1160 3440 1760
rect 3640 1160 3700 1760
rect 3900 1160 3960 1760
rect 4160 1160 4220 1760
rect 4420 1160 4480 1760
rect 4680 1160 4740 1760
rect 4940 1160 5000 1760
rect 5200 1160 5260 1760
rect 5460 1160 5520 1760
rect 5720 1160 5780 1760
rect 5980 1160 6040 1760
rect 6240 1160 6300 1760
rect 6500 1160 6560 1760
rect 6760 1160 6820 1760
rect 2290 -1650 2350 -1050
rect 2550 -1650 2610 -1050
rect 2810 -1650 2870 -1050
rect 3070 -1650 3130 -1050
rect 3330 -1650 3390 -1050
rect 3590 -1650 3650 -1050
rect 3850 -1650 3910 -1050
rect 4110 -1650 4170 -1050
rect 4370 -1650 4430 -1050
rect 4630 -1650 4690 -1050
rect 4890 -1650 4950 -1050
rect 5150 -1650 5210 -1050
rect 5410 -1650 5470 -1050
rect 5670 -1650 5730 -1050
rect 5930 -1650 5990 -1050
rect 6190 -1650 6250 -1050
rect 6450 -1650 6510 -1050
rect 6710 -1650 6770 -1050
<< ndiff >>
rect -110 610 90 660
rect -110 510 -60 610
rect 40 510 90 610
rect -110 310 90 510
rect -110 210 -60 310
rect 40 210 90 310
rect -110 160 90 210
rect 120 610 320 660
rect 120 510 170 610
rect 270 510 320 610
rect 120 310 320 510
rect 120 210 170 310
rect 270 210 320 310
rect 120 160 320 210
rect 350 610 550 660
rect 350 510 400 610
rect 500 510 550 610
rect 350 310 550 510
rect 350 210 400 310
rect 500 210 550 310
rect 350 160 550 210
rect 580 610 780 660
rect 580 510 630 610
rect 730 510 780 610
rect 580 310 780 510
rect 580 210 630 310
rect 730 210 780 310
rect 580 160 780 210
rect 810 610 1010 660
rect 810 510 860 610
rect 960 510 1010 610
rect 810 310 1010 510
rect 810 210 860 310
rect 960 210 1010 310
rect 810 160 1010 210
rect 1040 610 1240 660
rect 1040 510 1090 610
rect 1190 510 1240 610
rect 1040 310 1240 510
rect 1040 210 1090 310
rect 1190 210 1240 310
rect 1040 160 1240 210
rect 1270 610 1470 660
rect 1270 510 1320 610
rect 1420 510 1470 610
rect 1270 310 1470 510
rect 1270 210 1320 310
rect 1420 210 1470 310
rect 1270 160 1470 210
rect 1500 610 1700 660
rect 1500 510 1550 610
rect 1650 510 1700 610
rect 1500 310 1700 510
rect 1500 210 1550 310
rect 1650 210 1700 310
rect 1500 160 1700 210
rect 1730 610 1930 660
rect 1730 510 1780 610
rect 1880 510 1930 610
rect 1730 310 1930 510
rect 1730 210 1780 310
rect 1880 210 1930 310
rect 1730 160 1930 210
rect 1960 610 2160 660
rect 1960 510 2010 610
rect 2110 510 2160 610
rect 1960 310 2160 510
rect 1960 210 2010 310
rect 2110 210 2160 310
rect 1960 160 2160 210
rect 2190 610 2390 660
rect 2190 510 2240 610
rect 2340 510 2390 610
rect 2190 310 2390 510
rect 2190 210 2240 310
rect 2340 210 2390 310
rect 2190 160 2390 210
rect 2420 610 2620 660
rect 2420 510 2470 610
rect 2570 510 2620 610
rect 2420 310 2620 510
rect 2420 210 2470 310
rect 2570 210 2620 310
rect 2420 160 2620 210
rect 2650 610 2850 660
rect 2650 510 2700 610
rect 2800 510 2850 610
rect 2650 310 2850 510
rect 2650 210 2700 310
rect 2800 210 2850 310
rect 2650 160 2850 210
rect 2880 610 3080 660
rect 2880 510 2930 610
rect 3030 510 3080 610
rect 2880 310 3080 510
rect 2880 210 2930 310
rect 3030 210 3080 310
rect 2880 160 3080 210
rect 3110 610 3310 660
rect 3110 510 3160 610
rect 3260 510 3310 610
rect 3110 310 3310 510
rect 3110 210 3160 310
rect 3260 210 3310 310
rect 3110 160 3310 210
rect 3340 610 3540 660
rect 3340 510 3390 610
rect 3490 510 3540 610
rect 3340 310 3540 510
rect 3340 210 3390 310
rect 3490 210 3540 310
rect 3340 160 3540 210
rect 3570 610 3770 660
rect 3570 510 3620 610
rect 3720 510 3770 610
rect 3570 310 3770 510
rect 3570 210 3620 310
rect 3720 210 3770 310
rect 3570 160 3770 210
rect 3800 610 4000 660
rect 3800 510 3850 610
rect 3950 510 4000 610
rect 3800 310 4000 510
rect 3800 210 3850 310
rect 3950 210 4000 310
rect 3800 160 4000 210
rect 4030 610 4230 660
rect 4030 510 4080 610
rect 4180 510 4230 610
rect 4030 310 4230 510
rect 4030 210 4080 310
rect 4180 210 4230 310
rect 4030 160 4230 210
rect 4260 610 4460 660
rect 4260 510 4310 610
rect 4410 510 4460 610
rect 4260 310 4460 510
rect 4260 210 4310 310
rect 4410 210 4460 310
rect 4260 160 4460 210
rect 4490 610 4690 660
rect 4490 510 4540 610
rect 4640 510 4690 610
rect 4490 310 4690 510
rect 4490 210 4540 310
rect 4640 210 4690 310
rect 4490 160 4690 210
rect 4720 610 4920 660
rect 4720 510 4770 610
rect 4870 510 4920 610
rect 4720 310 4920 510
rect 4720 210 4770 310
rect 4870 210 4920 310
rect 4720 160 4920 210
rect 4950 610 5150 660
rect 4950 510 5000 610
rect 5100 510 5150 610
rect 4950 310 5150 510
rect 4950 210 5000 310
rect 5100 210 5150 310
rect 4950 160 5150 210
rect 5180 610 5380 660
rect 5180 510 5230 610
rect 5330 510 5380 610
rect 5180 310 5380 510
rect 5180 210 5230 310
rect 5330 210 5380 310
rect 5180 160 5380 210
rect 5410 610 5610 660
rect 5410 510 5460 610
rect 5560 510 5610 610
rect 5410 310 5610 510
rect 5410 210 5460 310
rect 5560 210 5610 310
rect 5410 160 5610 210
rect 5640 610 5840 660
rect 5640 510 5690 610
rect 5790 510 5840 610
rect 5640 310 5840 510
rect 5640 210 5690 310
rect 5790 210 5840 310
rect 5640 160 5840 210
rect 5870 610 6070 660
rect 5870 510 5920 610
rect 6020 510 6070 610
rect 5870 310 6070 510
rect 5870 210 5920 310
rect 6020 210 6070 310
rect 5870 160 6070 210
rect 6100 610 6300 660
rect 6100 510 6150 610
rect 6250 510 6300 610
rect 6100 310 6300 510
rect 6100 210 6150 310
rect 6250 210 6300 310
rect 6100 160 6300 210
rect 6330 610 6530 660
rect 6330 510 6380 610
rect 6480 510 6530 610
rect 6330 310 6530 510
rect 6330 210 6380 310
rect 6480 210 6530 310
rect 6330 160 6530 210
rect 6560 610 6760 660
rect 6560 510 6610 610
rect 6710 510 6760 610
rect 6560 310 6760 510
rect 6560 210 6610 310
rect 6710 210 6760 310
rect 6560 160 6760 210
rect 6790 610 6990 660
rect 6790 510 6840 610
rect 6940 510 6990 610
rect 6790 310 6990 510
rect 6790 210 6840 310
rect 6940 210 6990 310
rect 6790 160 6990 210
rect -110 -100 90 -50
rect -110 -200 -60 -100
rect 40 -200 90 -100
rect -110 -400 90 -200
rect -110 -500 -60 -400
rect 40 -500 90 -400
rect -110 -550 90 -500
rect 120 -100 320 -50
rect 120 -200 170 -100
rect 270 -200 320 -100
rect 120 -400 320 -200
rect 120 -500 170 -400
rect 270 -500 320 -400
rect 120 -550 320 -500
rect 350 -100 550 -50
rect 350 -200 400 -100
rect 500 -200 550 -100
rect 350 -400 550 -200
rect 350 -500 400 -400
rect 500 -500 550 -400
rect 350 -550 550 -500
rect 580 -100 780 -50
rect 580 -200 630 -100
rect 730 -200 780 -100
rect 580 -400 780 -200
rect 580 -500 630 -400
rect 730 -500 780 -400
rect 580 -550 780 -500
rect 810 -100 1010 -50
rect 810 -200 860 -100
rect 960 -200 1010 -100
rect 810 -400 1010 -200
rect 810 -500 860 -400
rect 960 -500 1010 -400
rect 810 -550 1010 -500
rect 1040 -100 1240 -50
rect 1040 -200 1090 -100
rect 1190 -200 1240 -100
rect 1040 -400 1240 -200
rect 1040 -500 1090 -400
rect 1190 -500 1240 -400
rect 1040 -550 1240 -500
rect 1270 -100 1470 -50
rect 1270 -200 1320 -100
rect 1420 -200 1470 -100
rect 1270 -400 1470 -200
rect 1270 -500 1320 -400
rect 1420 -500 1470 -400
rect 1270 -550 1470 -500
rect 1500 -100 1700 -50
rect 1500 -200 1550 -100
rect 1650 -200 1700 -100
rect 1500 -400 1700 -200
rect 1500 -500 1550 -400
rect 1650 -500 1700 -400
rect 1500 -550 1700 -500
rect 1730 -100 1930 -50
rect 1730 -200 1780 -100
rect 1880 -200 1930 -100
rect 1730 -400 1930 -200
rect 1730 -500 1780 -400
rect 1880 -500 1930 -400
rect 1730 -550 1930 -500
rect 1960 -100 2160 -50
rect 1960 -200 2010 -100
rect 2110 -200 2160 -100
rect 1960 -400 2160 -200
rect 1960 -500 2010 -400
rect 2110 -500 2160 -400
rect 1960 -550 2160 -500
rect 2190 -100 2390 -50
rect 2190 -200 2240 -100
rect 2340 -200 2390 -100
rect 2190 -400 2390 -200
rect 2190 -500 2240 -400
rect 2340 -500 2390 -400
rect 2190 -550 2390 -500
rect 2420 -100 2620 -50
rect 2420 -200 2470 -100
rect 2570 -200 2620 -100
rect 2420 -400 2620 -200
rect 2420 -500 2470 -400
rect 2570 -500 2620 -400
rect 2420 -550 2620 -500
rect 2650 -100 2850 -50
rect 2650 -200 2700 -100
rect 2800 -200 2850 -100
rect 2650 -400 2850 -200
rect 2650 -500 2700 -400
rect 2800 -500 2850 -400
rect 2650 -550 2850 -500
rect 2880 -100 3080 -50
rect 2880 -200 2930 -100
rect 3030 -200 3080 -100
rect 2880 -400 3080 -200
rect 2880 -500 2930 -400
rect 3030 -500 3080 -400
rect 2880 -550 3080 -500
rect 3110 -100 3310 -50
rect 3110 -200 3160 -100
rect 3260 -200 3310 -100
rect 3110 -400 3310 -200
rect 3110 -500 3160 -400
rect 3260 -500 3310 -400
rect 3110 -550 3310 -500
rect 3340 -100 3540 -50
rect 3340 -200 3390 -100
rect 3490 -200 3540 -100
rect 3340 -400 3540 -200
rect 3340 -500 3390 -400
rect 3490 -500 3540 -400
rect 3340 -550 3540 -500
rect 3570 -100 3770 -50
rect 3570 -200 3620 -100
rect 3720 -200 3770 -100
rect 3570 -400 3770 -200
rect 3570 -500 3620 -400
rect 3720 -500 3770 -400
rect 3570 -550 3770 -500
rect 3800 -100 4000 -50
rect 3800 -200 3850 -100
rect 3950 -200 4000 -100
rect 3800 -400 4000 -200
rect 3800 -500 3850 -400
rect 3950 -500 4000 -400
rect 3800 -550 4000 -500
rect 4030 -100 4230 -50
rect 4030 -200 4080 -100
rect 4180 -200 4230 -100
rect 4030 -400 4230 -200
rect 4030 -500 4080 -400
rect 4180 -500 4230 -400
rect 4030 -550 4230 -500
rect 4260 -100 4460 -50
rect 4260 -200 4310 -100
rect 4410 -200 4460 -100
rect 4260 -400 4460 -200
rect 4260 -500 4310 -400
rect 4410 -500 4460 -400
rect 4260 -550 4460 -500
rect 4490 -100 4690 -50
rect 4490 -200 4540 -100
rect 4640 -200 4690 -100
rect 4490 -400 4690 -200
rect 4490 -500 4540 -400
rect 4640 -500 4690 -400
rect 4490 -550 4690 -500
rect 4720 -100 4920 -50
rect 4720 -200 4770 -100
rect 4870 -200 4920 -100
rect 4720 -400 4920 -200
rect 4720 -500 4770 -400
rect 4870 -500 4920 -400
rect 4720 -550 4920 -500
rect 4950 -100 5150 -50
rect 4950 -200 5000 -100
rect 5100 -200 5150 -100
rect 4950 -400 5150 -200
rect 4950 -500 5000 -400
rect 5100 -500 5150 -400
rect 4950 -550 5150 -500
rect 5180 -100 5380 -50
rect 5180 -200 5230 -100
rect 5330 -200 5380 -100
rect 5180 -400 5380 -200
rect 5180 -500 5230 -400
rect 5330 -500 5380 -400
rect 5180 -550 5380 -500
rect 5410 -100 5610 -50
rect 5410 -200 5460 -100
rect 5560 -200 5610 -100
rect 5410 -400 5610 -200
rect 5410 -500 5460 -400
rect 5560 -500 5610 -400
rect 5410 -550 5610 -500
rect 5640 -100 5840 -50
rect 5640 -200 5690 -100
rect 5790 -200 5840 -100
rect 5640 -400 5840 -200
rect 5640 -500 5690 -400
rect 5790 -500 5840 -400
rect 5640 -550 5840 -500
rect 5870 -100 6070 -50
rect 5870 -200 5920 -100
rect 6020 -200 6070 -100
rect 5870 -400 6070 -200
rect 5870 -500 5920 -400
rect 6020 -500 6070 -400
rect 5870 -550 6070 -500
rect 6100 -100 6300 -50
rect 6100 -200 6150 -100
rect 6250 -200 6300 -100
rect 6100 -400 6300 -200
rect 6100 -500 6150 -400
rect 6250 -500 6300 -400
rect 6100 -550 6300 -500
rect 6330 -100 6530 -50
rect 6330 -200 6380 -100
rect 6480 -200 6530 -100
rect 6330 -400 6530 -200
rect 6330 -500 6380 -400
rect 6480 -500 6530 -400
rect 6330 -550 6530 -500
rect 6560 -100 6760 -50
rect 6560 -200 6610 -100
rect 6710 -200 6760 -100
rect 6560 -400 6760 -200
rect 6560 -500 6610 -400
rect 6710 -500 6760 -400
rect 6560 -550 6760 -500
rect 6790 -100 6990 -50
rect 6790 -200 6840 -100
rect 6940 -200 6990 -100
rect 6790 -400 6990 -200
rect 6790 -500 6840 -400
rect 6940 -500 6990 -400
rect 6790 -550 6990 -500
<< pdiff >>
rect 1350 1680 1550 1760
rect 1350 1580 1400 1680
rect 1500 1580 1550 1680
rect 1350 1400 1550 1580
rect 1350 1300 1400 1400
rect 1500 1300 1550 1400
rect 1350 1220 1550 1300
rect 1610 1680 1810 1760
rect 1610 1580 1660 1680
rect 1760 1580 1810 1680
rect 1610 1400 1810 1580
rect 1610 1300 1660 1400
rect 1760 1300 1810 1400
rect 1610 1220 1810 1300
rect 1870 1680 2070 1760
rect 1870 1580 1920 1680
rect 2020 1580 2070 1680
rect 1870 1400 2070 1580
rect 1870 1300 1920 1400
rect 2020 1300 2070 1400
rect 1870 1220 2070 1300
rect 2140 1680 2340 1760
rect 2140 1580 2190 1680
rect 2290 1580 2340 1680
rect 2140 1340 2340 1580
rect 2140 1240 2190 1340
rect 2290 1240 2340 1340
rect 2140 1160 2340 1240
rect 2400 1680 2600 1760
rect 2400 1580 2450 1680
rect 2550 1580 2600 1680
rect 2400 1340 2600 1580
rect 2400 1240 2450 1340
rect 2550 1240 2600 1340
rect 2400 1160 2600 1240
rect 2660 1680 2860 1760
rect 2660 1580 2710 1680
rect 2810 1580 2860 1680
rect 2660 1340 2860 1580
rect 2660 1240 2710 1340
rect 2810 1240 2860 1340
rect 2660 1160 2860 1240
rect 2920 1680 3120 1760
rect 2920 1580 2970 1680
rect 3070 1580 3120 1680
rect 2920 1340 3120 1580
rect 2920 1240 2970 1340
rect 3070 1240 3120 1340
rect 2920 1160 3120 1240
rect 3180 1680 3380 1760
rect 3180 1580 3230 1680
rect 3330 1580 3380 1680
rect 3180 1340 3380 1580
rect 3180 1240 3230 1340
rect 3330 1240 3380 1340
rect 3180 1160 3380 1240
rect 3440 1680 3640 1760
rect 3440 1580 3490 1680
rect 3590 1580 3640 1680
rect 3440 1340 3640 1580
rect 3440 1240 3490 1340
rect 3590 1240 3640 1340
rect 3440 1160 3640 1240
rect 3700 1680 3900 1760
rect 3700 1580 3750 1680
rect 3850 1580 3900 1680
rect 3700 1340 3900 1580
rect 3700 1240 3750 1340
rect 3850 1240 3900 1340
rect 3700 1160 3900 1240
rect 3960 1680 4160 1760
rect 3960 1580 4010 1680
rect 4110 1580 4160 1680
rect 3960 1340 4160 1580
rect 3960 1240 4010 1340
rect 4110 1240 4160 1340
rect 3960 1160 4160 1240
rect 4220 1680 4420 1760
rect 4220 1580 4270 1680
rect 4370 1580 4420 1680
rect 4220 1340 4420 1580
rect 4220 1240 4270 1340
rect 4370 1240 4420 1340
rect 4220 1160 4420 1240
rect 4480 1680 4680 1760
rect 4480 1580 4530 1680
rect 4630 1580 4680 1680
rect 4480 1340 4680 1580
rect 4480 1240 4530 1340
rect 4630 1240 4680 1340
rect 4480 1160 4680 1240
rect 4740 1680 4940 1760
rect 4740 1580 4790 1680
rect 4890 1580 4940 1680
rect 4740 1340 4940 1580
rect 4740 1240 4790 1340
rect 4890 1240 4940 1340
rect 4740 1160 4940 1240
rect 5000 1680 5200 1760
rect 5000 1580 5050 1680
rect 5150 1580 5200 1680
rect 5000 1340 5200 1580
rect 5000 1240 5050 1340
rect 5150 1240 5200 1340
rect 5000 1160 5200 1240
rect 5260 1680 5460 1760
rect 5260 1580 5310 1680
rect 5410 1580 5460 1680
rect 5260 1340 5460 1580
rect 5260 1240 5310 1340
rect 5410 1240 5460 1340
rect 5260 1160 5460 1240
rect 5520 1680 5720 1760
rect 5520 1580 5570 1680
rect 5670 1580 5720 1680
rect 5520 1340 5720 1580
rect 5520 1240 5570 1340
rect 5670 1240 5720 1340
rect 5520 1160 5720 1240
rect 5780 1680 5980 1760
rect 5780 1580 5830 1680
rect 5930 1580 5980 1680
rect 5780 1340 5980 1580
rect 5780 1240 5830 1340
rect 5930 1240 5980 1340
rect 5780 1160 5980 1240
rect 6040 1680 6240 1760
rect 6040 1580 6090 1680
rect 6190 1580 6240 1680
rect 6040 1340 6240 1580
rect 6040 1240 6090 1340
rect 6190 1240 6240 1340
rect 6040 1160 6240 1240
rect 6300 1680 6500 1760
rect 6300 1580 6350 1680
rect 6450 1580 6500 1680
rect 6300 1340 6500 1580
rect 6300 1240 6350 1340
rect 6450 1240 6500 1340
rect 6300 1160 6500 1240
rect 6560 1680 6760 1760
rect 6560 1580 6610 1680
rect 6710 1580 6760 1680
rect 6560 1340 6760 1580
rect 6560 1240 6610 1340
rect 6710 1240 6760 1340
rect 6560 1160 6760 1240
rect 6820 1680 7020 1760
rect 6820 1580 6870 1680
rect 6970 1580 7020 1680
rect 6820 1340 7020 1580
rect 6820 1240 6870 1340
rect 6970 1240 7020 1340
rect 6820 1160 7020 1240
rect 2090 -1130 2290 -1050
rect 2090 -1230 2140 -1130
rect 2240 -1230 2290 -1130
rect 2090 -1470 2290 -1230
rect 2090 -1570 2140 -1470
rect 2240 -1570 2290 -1470
rect 2090 -1650 2290 -1570
rect 2350 -1130 2550 -1050
rect 2350 -1230 2400 -1130
rect 2500 -1230 2550 -1130
rect 2350 -1470 2550 -1230
rect 2350 -1570 2400 -1470
rect 2500 -1570 2550 -1470
rect 2350 -1650 2550 -1570
rect 2610 -1130 2810 -1050
rect 2610 -1230 2660 -1130
rect 2760 -1230 2810 -1130
rect 2610 -1470 2810 -1230
rect 2610 -1570 2660 -1470
rect 2760 -1570 2810 -1470
rect 2610 -1650 2810 -1570
rect 2870 -1130 3070 -1050
rect 2870 -1230 2920 -1130
rect 3020 -1230 3070 -1130
rect 2870 -1470 3070 -1230
rect 2870 -1570 2920 -1470
rect 3020 -1570 3070 -1470
rect 2870 -1650 3070 -1570
rect 3130 -1130 3330 -1050
rect 3130 -1230 3180 -1130
rect 3280 -1230 3330 -1130
rect 3130 -1470 3330 -1230
rect 3130 -1570 3180 -1470
rect 3280 -1570 3330 -1470
rect 3130 -1650 3330 -1570
rect 3390 -1130 3590 -1050
rect 3390 -1230 3440 -1130
rect 3540 -1230 3590 -1130
rect 3390 -1470 3590 -1230
rect 3390 -1570 3440 -1470
rect 3540 -1570 3590 -1470
rect 3390 -1650 3590 -1570
rect 3650 -1130 3850 -1050
rect 3650 -1230 3700 -1130
rect 3800 -1230 3850 -1130
rect 3650 -1470 3850 -1230
rect 3650 -1570 3700 -1470
rect 3800 -1570 3850 -1470
rect 3650 -1650 3850 -1570
rect 3910 -1130 4110 -1050
rect 3910 -1230 3960 -1130
rect 4060 -1230 4110 -1130
rect 3910 -1470 4110 -1230
rect 3910 -1570 3960 -1470
rect 4060 -1570 4110 -1470
rect 3910 -1650 4110 -1570
rect 4170 -1130 4370 -1050
rect 4170 -1230 4220 -1130
rect 4320 -1230 4370 -1130
rect 4170 -1470 4370 -1230
rect 4170 -1570 4220 -1470
rect 4320 -1570 4370 -1470
rect 4170 -1650 4370 -1570
rect 4430 -1130 4630 -1050
rect 4430 -1230 4480 -1130
rect 4580 -1230 4630 -1130
rect 4430 -1470 4630 -1230
rect 4430 -1570 4480 -1470
rect 4580 -1570 4630 -1470
rect 4430 -1650 4630 -1570
rect 4690 -1130 4890 -1050
rect 4690 -1230 4740 -1130
rect 4840 -1230 4890 -1130
rect 4690 -1470 4890 -1230
rect 4690 -1570 4740 -1470
rect 4840 -1570 4890 -1470
rect 4690 -1650 4890 -1570
rect 4950 -1130 5150 -1050
rect 4950 -1230 5000 -1130
rect 5100 -1230 5150 -1130
rect 4950 -1470 5150 -1230
rect 4950 -1570 5000 -1470
rect 5100 -1570 5150 -1470
rect 4950 -1650 5150 -1570
rect 5210 -1130 5410 -1050
rect 5210 -1230 5260 -1130
rect 5360 -1230 5410 -1130
rect 5210 -1470 5410 -1230
rect 5210 -1570 5260 -1470
rect 5360 -1570 5410 -1470
rect 5210 -1650 5410 -1570
rect 5470 -1130 5670 -1050
rect 5470 -1230 5520 -1130
rect 5620 -1230 5670 -1130
rect 5470 -1470 5670 -1230
rect 5470 -1570 5520 -1470
rect 5620 -1570 5670 -1470
rect 5470 -1650 5670 -1570
rect 5730 -1130 5930 -1050
rect 5730 -1230 5780 -1130
rect 5880 -1230 5930 -1130
rect 5730 -1470 5930 -1230
rect 5730 -1570 5780 -1470
rect 5880 -1570 5930 -1470
rect 5730 -1650 5930 -1570
rect 5990 -1130 6190 -1050
rect 5990 -1230 6040 -1130
rect 6140 -1230 6190 -1130
rect 5990 -1470 6190 -1230
rect 5990 -1570 6040 -1470
rect 6140 -1570 6190 -1470
rect 5990 -1650 6190 -1570
rect 6250 -1130 6450 -1050
rect 6250 -1230 6300 -1130
rect 6400 -1230 6450 -1130
rect 6250 -1470 6450 -1230
rect 6250 -1570 6300 -1470
rect 6400 -1570 6450 -1470
rect 6250 -1650 6450 -1570
rect 6510 -1130 6710 -1050
rect 6510 -1230 6560 -1130
rect 6660 -1230 6710 -1130
rect 6510 -1470 6710 -1230
rect 6510 -1570 6560 -1470
rect 6660 -1570 6710 -1470
rect 6510 -1650 6710 -1570
rect 6770 -1130 6970 -1050
rect 6770 -1230 6820 -1130
rect 6920 -1230 6970 -1130
rect 6770 -1470 6970 -1230
rect 6770 -1570 6820 -1470
rect 6920 -1570 6970 -1470
rect 6770 -1650 6970 -1570
<< ndiffc >>
rect -60 510 40 610
rect -60 210 40 310
rect 170 510 270 610
rect 170 210 270 310
rect 400 510 500 610
rect 400 210 500 310
rect 630 510 730 610
rect 630 210 730 310
rect 860 510 960 610
rect 860 210 960 310
rect 1090 510 1190 610
rect 1090 210 1190 310
rect 1320 510 1420 610
rect 1320 210 1420 310
rect 1550 510 1650 610
rect 1550 210 1650 310
rect 1780 510 1880 610
rect 1780 210 1880 310
rect 2010 510 2110 610
rect 2010 210 2110 310
rect 2240 510 2340 610
rect 2240 210 2340 310
rect 2470 510 2570 610
rect 2470 210 2570 310
rect 2700 510 2800 610
rect 2700 210 2800 310
rect 2930 510 3030 610
rect 2930 210 3030 310
rect 3160 510 3260 610
rect 3160 210 3260 310
rect 3390 510 3490 610
rect 3390 210 3490 310
rect 3620 510 3720 610
rect 3620 210 3720 310
rect 3850 510 3950 610
rect 3850 210 3950 310
rect 4080 510 4180 610
rect 4080 210 4180 310
rect 4310 510 4410 610
rect 4310 210 4410 310
rect 4540 510 4640 610
rect 4540 210 4640 310
rect 4770 510 4870 610
rect 4770 210 4870 310
rect 5000 510 5100 610
rect 5000 210 5100 310
rect 5230 510 5330 610
rect 5230 210 5330 310
rect 5460 510 5560 610
rect 5460 210 5560 310
rect 5690 510 5790 610
rect 5690 210 5790 310
rect 5920 510 6020 610
rect 5920 210 6020 310
rect 6150 510 6250 610
rect 6150 210 6250 310
rect 6380 510 6480 610
rect 6380 210 6480 310
rect 6610 510 6710 610
rect 6610 210 6710 310
rect 6840 510 6940 610
rect 6840 210 6940 310
rect -60 -200 40 -100
rect -60 -500 40 -400
rect 170 -200 270 -100
rect 170 -500 270 -400
rect 400 -200 500 -100
rect 400 -500 500 -400
rect 630 -200 730 -100
rect 630 -500 730 -400
rect 860 -200 960 -100
rect 860 -500 960 -400
rect 1090 -200 1190 -100
rect 1090 -500 1190 -400
rect 1320 -200 1420 -100
rect 1320 -500 1420 -400
rect 1550 -200 1650 -100
rect 1550 -500 1650 -400
rect 1780 -200 1880 -100
rect 1780 -500 1880 -400
rect 2010 -200 2110 -100
rect 2010 -500 2110 -400
rect 2240 -200 2340 -100
rect 2240 -500 2340 -400
rect 2470 -200 2570 -100
rect 2470 -500 2570 -400
rect 2700 -200 2800 -100
rect 2700 -500 2800 -400
rect 2930 -200 3030 -100
rect 2930 -500 3030 -400
rect 3160 -200 3260 -100
rect 3160 -500 3260 -400
rect 3390 -200 3490 -100
rect 3390 -500 3490 -400
rect 3620 -200 3720 -100
rect 3620 -500 3720 -400
rect 3850 -200 3950 -100
rect 3850 -500 3950 -400
rect 4080 -200 4180 -100
rect 4080 -500 4180 -400
rect 4310 -200 4410 -100
rect 4310 -500 4410 -400
rect 4540 -200 4640 -100
rect 4540 -500 4640 -400
rect 4770 -200 4870 -100
rect 4770 -500 4870 -400
rect 5000 -200 5100 -100
rect 5000 -500 5100 -400
rect 5230 -200 5330 -100
rect 5230 -500 5330 -400
rect 5460 -200 5560 -100
rect 5460 -500 5560 -400
rect 5690 -200 5790 -100
rect 5690 -500 5790 -400
rect 5920 -200 6020 -100
rect 5920 -500 6020 -400
rect 6150 -200 6250 -100
rect 6150 -500 6250 -400
rect 6380 -200 6480 -100
rect 6380 -500 6480 -400
rect 6610 -200 6710 -100
rect 6610 -500 6710 -400
rect 6840 -200 6940 -100
rect 6840 -500 6940 -400
<< pdiffc >>
rect 1400 1580 1500 1680
rect 1400 1300 1500 1400
rect 1660 1580 1760 1680
rect 1660 1300 1760 1400
rect 1920 1580 2020 1680
rect 1920 1300 2020 1400
rect 2190 1580 2290 1680
rect 2190 1240 2290 1340
rect 2450 1580 2550 1680
rect 2450 1240 2550 1340
rect 2710 1580 2810 1680
rect 2710 1240 2810 1340
rect 2970 1580 3070 1680
rect 2970 1240 3070 1340
rect 3230 1580 3330 1680
rect 3230 1240 3330 1340
rect 3490 1580 3590 1680
rect 3490 1240 3590 1340
rect 3750 1580 3850 1680
rect 3750 1240 3850 1340
rect 4010 1580 4110 1680
rect 4010 1240 4110 1340
rect 4270 1580 4370 1680
rect 4270 1240 4370 1340
rect 4530 1580 4630 1680
rect 4530 1240 4630 1340
rect 4790 1580 4890 1680
rect 4790 1240 4890 1340
rect 5050 1580 5150 1680
rect 5050 1240 5150 1340
rect 5310 1580 5410 1680
rect 5310 1240 5410 1340
rect 5570 1580 5670 1680
rect 5570 1240 5670 1340
rect 5830 1580 5930 1680
rect 5830 1240 5930 1340
rect 6090 1580 6190 1680
rect 6090 1240 6190 1340
rect 6350 1580 6450 1680
rect 6350 1240 6450 1340
rect 6610 1580 6710 1680
rect 6610 1240 6710 1340
rect 6870 1580 6970 1680
rect 6870 1240 6970 1340
rect 2140 -1230 2240 -1130
rect 2140 -1570 2240 -1470
rect 2400 -1230 2500 -1130
rect 2400 -1570 2500 -1470
rect 2660 -1230 2760 -1130
rect 2660 -1570 2760 -1470
rect 2920 -1230 3020 -1130
rect 2920 -1570 3020 -1470
rect 3180 -1230 3280 -1130
rect 3180 -1570 3280 -1470
rect 3440 -1230 3540 -1130
rect 3440 -1570 3540 -1470
rect 3700 -1230 3800 -1130
rect 3700 -1570 3800 -1470
rect 3960 -1230 4060 -1130
rect 3960 -1570 4060 -1470
rect 4220 -1230 4320 -1130
rect 4220 -1570 4320 -1470
rect 4480 -1230 4580 -1130
rect 4480 -1570 4580 -1470
rect 4740 -1230 4840 -1130
rect 4740 -1570 4840 -1470
rect 5000 -1230 5100 -1130
rect 5000 -1570 5100 -1470
rect 5260 -1230 5360 -1130
rect 5260 -1570 5360 -1470
rect 5520 -1230 5620 -1130
rect 5520 -1570 5620 -1470
rect 5780 -1230 5880 -1130
rect 5780 -1570 5880 -1470
rect 6040 -1230 6140 -1130
rect 6040 -1570 6140 -1470
rect 6300 -1230 6400 -1130
rect 6300 -1570 6400 -1470
rect 6560 -1230 6660 -1130
rect 6560 -1570 6660 -1470
rect 6820 -1230 6920 -1130
rect 6820 -1570 6920 -1470
<< psubdiff >>
rect -690 2484 -430 2514
rect -1990 2324 -1730 2354
rect -1990 2124 -1960 2324
rect -1760 2124 -1730 2324
rect -690 2284 -660 2484
rect -460 2284 -430 2484
rect -690 2254 -430 2284
rect 310 2484 570 2514
rect 310 2284 340 2484
rect 540 2284 570 2484
rect 310 2254 570 2284
rect 1310 2484 1570 2514
rect 1310 2284 1340 2484
rect 1540 2284 1570 2484
rect 1310 2254 1570 2284
rect 2330 2484 2590 2514
rect 2330 2284 2360 2484
rect 2560 2284 2590 2484
rect 2330 2254 2590 2284
rect 3330 2484 3590 2514
rect 3330 2284 3360 2484
rect 3560 2284 3590 2484
rect 3330 2254 3590 2284
rect 4330 2484 4590 2514
rect 4330 2284 4360 2484
rect 4560 2284 4590 2484
rect 4330 2254 4590 2284
rect 5350 2484 5610 2514
rect 5350 2284 5380 2484
rect 5580 2284 5610 2484
rect 5350 2254 5610 2284
rect 6350 2484 6610 2514
rect 6350 2284 6380 2484
rect 6580 2284 6610 2484
rect 6350 2254 6610 2284
rect 7350 2484 7880 2514
rect 7350 2284 7380 2484
rect 7580 2284 7880 2484
rect 7350 2254 7880 2284
rect 7990 2254 8250 2284
rect -1990 2070 -1730 2124
rect 7990 2030 8020 2254
rect 8220 2030 8250 2254
rect 7990 1940 8250 2030
rect -1990 1280 -1730 1310
rect -1990 1080 -1960 1280
rect -1760 1080 -1730 1280
rect 7990 1520 8250 1550
rect 7990 1320 8020 1520
rect 8220 1320 8250 1520
rect 7990 1290 8250 1320
rect -1990 990 -1730 1080
rect 8010 830 8270 860
rect -1990 570 -1730 600
rect -1990 370 -1960 570
rect -1760 370 -1730 570
rect -1990 340 -1730 370
rect 8010 630 8040 830
rect 8240 630 8270 830
rect 8010 600 8270 630
rect 1320 80 1490 100
rect 1320 30 1370 80
rect 1450 30 1490 80
rect 1320 10 1490 30
rect -1990 -450 -1730 -420
rect -1990 -650 -1960 -450
rect -1760 -650 -1730 -450
rect 8010 -190 8270 -160
rect 8010 -390 8040 -190
rect 8240 -390 8270 -190
rect 8010 -420 8270 -390
rect -1990 -680 -1730 -650
rect -1990 -1450 -1730 -1420
rect -1990 -1650 -1960 -1450
rect -1760 -1650 -1730 -1450
rect -1990 -1680 -1730 -1650
rect 8010 -1920 8270 -1890
rect 8010 -2120 8040 -1920
rect 8240 -2120 8270 -1920
rect 8010 -2150 8270 -2120
rect -1800 -2200 -1540 -2170
rect -1800 -2400 -1770 -2200
rect -1570 -2400 -1540 -2200
rect -1800 -2430 -1540 -2400
rect -580 -2200 -320 -2170
rect -580 -2400 -550 -2200
rect -350 -2400 -320 -2200
rect -580 -2430 -320 -2400
rect 280 -2200 540 -2170
rect 280 -2400 310 -2200
rect 510 -2400 540 -2200
rect 280 -2430 540 -2400
rect 1280 -2200 1540 -2170
rect 1280 -2400 1310 -2200
rect 1510 -2400 1540 -2200
rect 1280 -2430 1540 -2400
rect 2300 -2200 2560 -2170
rect 2300 -2400 2330 -2200
rect 2530 -2400 2560 -2200
rect 2300 -2430 2560 -2400
rect 3300 -2200 3560 -2170
rect 3300 -2400 3330 -2200
rect 3530 -2400 3560 -2200
rect 3300 -2430 3560 -2400
rect 4300 -2200 4560 -2170
rect 4300 -2400 4330 -2200
rect 4530 -2400 4560 -2200
rect 4300 -2430 4560 -2400
rect 5320 -2200 5580 -2170
rect 5320 -2400 5350 -2200
rect 5550 -2400 5580 -2200
rect 5320 -2430 5580 -2400
rect 6320 -2200 6580 -2170
rect 6320 -2400 6350 -2200
rect 6550 -2400 6580 -2200
rect 6320 -2430 6580 -2400
rect 7320 -2200 7580 -2170
rect 7320 -2400 7350 -2200
rect 7550 -2400 7580 -2200
rect 7320 -2430 7580 -2400
<< nsubdiff >>
rect 7090 1720 7320 1760
rect 7090 1540 7130 1720
rect 7290 1540 7320 1720
rect 7090 1510 7320 1540
rect 7050 -1100 7280 -1060
rect 7050 -1280 7090 -1100
rect 7250 -1280 7280 -1100
rect 7050 -1310 7280 -1280
<< psubdiffcont >>
rect -1960 2124 -1760 2324
rect -660 2284 -460 2484
rect 340 2284 540 2484
rect 1340 2284 1540 2484
rect 2360 2284 2560 2484
rect 3360 2284 3560 2484
rect 4360 2284 4560 2484
rect 5380 2284 5580 2484
rect 6380 2284 6580 2484
rect 7380 2284 7580 2484
rect 8020 2030 8220 2254
rect -1960 1080 -1760 1280
rect 8020 1320 8220 1520
rect -1960 370 -1760 570
rect 8040 630 8240 830
rect 1370 30 1450 80
rect -1960 -650 -1760 -450
rect 8040 -390 8240 -190
rect -1960 -1650 -1760 -1450
rect 8040 -2120 8240 -1920
rect -1770 -2400 -1570 -2200
rect -550 -2400 -350 -2200
rect 310 -2400 510 -2200
rect 1310 -2400 1510 -2200
rect 2330 -2400 2530 -2200
rect 3330 -2400 3530 -2200
rect 4330 -2400 4530 -2200
rect 5350 -2400 5550 -2200
rect 6350 -2400 6550 -2200
rect 7350 -2400 7550 -2200
<< nsubdiffcont >>
rect 7130 1540 7290 1720
rect 7090 -1280 7250 -1100
<< poly >>
rect 1520 1880 1640 1900
rect 1520 1810 1540 1880
rect 1620 1810 1640 1880
rect 1520 1790 1640 1810
rect 1780 1880 1900 1900
rect 1780 1810 1800 1880
rect 1880 1810 1900 1880
rect 1780 1790 1900 1810
rect 2310 1880 2430 1900
rect 2310 1810 2330 1880
rect 2410 1810 2430 1880
rect 2310 1790 2430 1810
rect 2570 1880 2690 1900
rect 2570 1810 2590 1880
rect 2670 1810 2690 1880
rect 2570 1790 2690 1810
rect 2830 1880 2950 1900
rect 2830 1810 2850 1880
rect 2930 1810 2950 1880
rect 2830 1790 2950 1810
rect 3090 1880 3210 1900
rect 3090 1810 3110 1880
rect 3190 1810 3210 1880
rect 3090 1790 3210 1810
rect 3350 1880 3470 1900
rect 3350 1810 3370 1880
rect 3450 1810 3470 1880
rect 3350 1790 3470 1810
rect 3610 1880 3730 1900
rect 3610 1810 3630 1880
rect 3710 1810 3730 1880
rect 3610 1790 3730 1810
rect 3870 1880 3990 1900
rect 3870 1810 3890 1880
rect 3970 1810 3990 1880
rect 3870 1790 3990 1810
rect 4130 1880 4250 1900
rect 4130 1810 4150 1880
rect 4230 1810 4250 1880
rect 4130 1790 4250 1810
rect 4390 1880 4510 1900
rect 4390 1810 4410 1880
rect 4490 1810 4510 1880
rect 4390 1790 4510 1810
rect 4650 1880 4770 1900
rect 4650 1810 4670 1880
rect 4750 1810 4770 1880
rect 4650 1790 4770 1810
rect 4910 1880 5030 1900
rect 4910 1810 4930 1880
rect 5010 1810 5030 1880
rect 4910 1790 5030 1810
rect 5170 1880 5290 1900
rect 5170 1810 5190 1880
rect 5270 1810 5290 1880
rect 5170 1790 5290 1810
rect 5430 1880 5550 1900
rect 5430 1810 5450 1880
rect 5530 1810 5550 1880
rect 5430 1790 5550 1810
rect 5690 1880 5810 1900
rect 5690 1810 5710 1880
rect 5790 1810 5810 1880
rect 5690 1790 5810 1810
rect 5950 1880 6070 1900
rect 5950 1810 5970 1880
rect 6050 1810 6070 1880
rect 5950 1790 6070 1810
rect 6210 1880 6330 1900
rect 6210 1810 6230 1880
rect 6310 1810 6330 1880
rect 6210 1790 6330 1810
rect 6470 1880 6590 1900
rect 6470 1810 6490 1880
rect 6570 1810 6590 1880
rect 6470 1790 6590 1810
rect 6730 1880 6850 1900
rect 6730 1810 6750 1880
rect 6830 1810 6850 1880
rect 6730 1790 6850 1810
rect 1550 1760 1610 1790
rect 1810 1760 1870 1790
rect 2340 1760 2400 1790
rect 2600 1760 2660 1790
rect 2860 1760 2920 1790
rect 3120 1760 3180 1790
rect 3380 1760 3440 1790
rect 3640 1760 3700 1790
rect 3900 1760 3960 1790
rect 4160 1760 4220 1790
rect 4420 1760 4480 1790
rect 4680 1760 4740 1790
rect 4940 1760 5000 1790
rect 5200 1760 5260 1790
rect 5460 1760 5520 1790
rect 5720 1760 5780 1790
rect 5980 1760 6040 1790
rect 6240 1760 6300 1790
rect 6500 1760 6560 1790
rect 6760 1760 6820 1790
rect 1550 1190 1610 1220
rect 1810 1190 1870 1220
rect 2340 1130 2400 1160
rect 2600 1130 2660 1160
rect 2860 1130 2920 1160
rect 3120 1130 3180 1160
rect 3380 1130 3440 1160
rect 3640 1130 3700 1160
rect 3900 1130 3960 1160
rect 4160 1130 4220 1160
rect 4420 1130 4480 1160
rect 4680 1130 4740 1160
rect 4940 1130 5000 1160
rect 5200 1130 5260 1160
rect 5460 1130 5520 1160
rect 5720 1130 5780 1160
rect 5980 1130 6040 1160
rect 6240 1130 6300 1160
rect 6500 1130 6560 1160
rect 6760 1130 6820 1160
rect 50 770 160 790
rect 50 700 70 770
rect 140 700 160 770
rect 50 680 160 700
rect 280 770 390 790
rect 280 700 300 770
rect 370 700 390 770
rect 280 680 390 700
rect 510 770 620 790
rect 510 700 530 770
rect 600 700 620 770
rect 510 680 620 700
rect 740 770 850 790
rect 740 700 760 770
rect 830 700 850 770
rect 740 680 850 700
rect 970 770 1080 790
rect 970 700 990 770
rect 1060 700 1080 770
rect 970 680 1080 700
rect 1200 770 1310 790
rect 1200 700 1220 770
rect 1290 700 1310 770
rect 1200 680 1310 700
rect 1430 770 1540 790
rect 1430 700 1450 770
rect 1520 700 1540 770
rect 1430 680 1540 700
rect 1660 770 1770 790
rect 1660 700 1680 770
rect 1750 700 1770 770
rect 1660 680 1770 700
rect 1890 770 2000 790
rect 1890 700 1910 770
rect 1980 700 2000 770
rect 1890 680 2000 700
rect 2120 770 2230 790
rect 2120 700 2140 770
rect 2210 700 2230 770
rect 2120 680 2230 700
rect 2350 770 2460 790
rect 2350 700 2370 770
rect 2440 700 2460 770
rect 2350 680 2460 700
rect 2580 770 2690 790
rect 2580 700 2600 770
rect 2670 700 2690 770
rect 2580 680 2690 700
rect 2810 770 2920 790
rect 2810 700 2830 770
rect 2900 700 2920 770
rect 2810 680 2920 700
rect 3040 770 3150 790
rect 3040 700 3060 770
rect 3130 700 3150 770
rect 3040 680 3150 700
rect 3270 770 3380 790
rect 3270 700 3290 770
rect 3360 700 3380 770
rect 3270 680 3380 700
rect 3500 770 3610 790
rect 3500 700 3520 770
rect 3590 700 3610 770
rect 3500 680 3610 700
rect 3730 770 3840 790
rect 3730 700 3750 770
rect 3820 700 3840 770
rect 3730 680 3840 700
rect 3960 770 4070 790
rect 3960 700 3980 770
rect 4050 700 4070 770
rect 3960 680 4070 700
rect 4190 770 4300 790
rect 4190 700 4210 770
rect 4280 700 4300 770
rect 4190 680 4300 700
rect 4420 770 4530 790
rect 4420 700 4440 770
rect 4510 700 4530 770
rect 4420 680 4530 700
rect 4650 770 4760 790
rect 4650 700 4670 770
rect 4740 700 4760 770
rect 4650 680 4760 700
rect 4880 770 4990 790
rect 4880 700 4900 770
rect 4970 700 4990 770
rect 4880 680 4990 700
rect 5110 770 5220 790
rect 5110 700 5130 770
rect 5200 700 5220 770
rect 5110 680 5220 700
rect 5340 770 5450 790
rect 5340 700 5360 770
rect 5430 700 5450 770
rect 5340 680 5450 700
rect 5570 770 5680 790
rect 5570 700 5590 770
rect 5660 700 5680 770
rect 5570 680 5680 700
rect 5800 770 5910 790
rect 5800 700 5820 770
rect 5890 700 5910 770
rect 5800 680 5910 700
rect 6030 770 6140 790
rect 6030 700 6050 770
rect 6120 700 6140 770
rect 6030 680 6140 700
rect 6260 770 6370 790
rect 6260 700 6280 770
rect 6350 700 6370 770
rect 6260 680 6370 700
rect 6490 770 6600 790
rect 6490 700 6510 770
rect 6580 700 6600 770
rect 6490 680 6600 700
rect 6720 770 6830 790
rect 6720 700 6740 770
rect 6810 700 6830 770
rect 6720 680 6830 700
rect 90 660 120 680
rect 320 660 350 680
rect 550 660 580 680
rect 780 660 810 680
rect 1010 660 1040 680
rect 1240 660 1270 680
rect 1470 660 1500 680
rect 1700 660 1730 680
rect 1930 660 1960 680
rect 2160 660 2190 680
rect 2390 660 2420 680
rect 2620 660 2650 680
rect 2850 660 2880 680
rect 3080 660 3110 680
rect 3310 660 3340 680
rect 3540 660 3570 680
rect 3770 660 3800 680
rect 4000 660 4030 680
rect 4230 660 4260 680
rect 4460 660 4490 680
rect 4690 660 4720 680
rect 4920 660 4950 680
rect 5150 660 5180 680
rect 5380 660 5410 680
rect 5610 660 5640 680
rect 5840 660 5870 680
rect 6070 660 6100 680
rect 6300 660 6330 680
rect 6530 660 6560 680
rect 6760 660 6790 680
rect 90 130 120 160
rect 320 130 350 160
rect 550 130 580 160
rect 780 130 810 160
rect 1010 130 1040 160
rect 1240 130 1270 160
rect 1470 130 1500 160
rect 1700 130 1730 160
rect 1930 130 1960 160
rect 2160 130 2190 160
rect 2390 130 2420 160
rect 2620 130 2650 160
rect 2850 130 2880 160
rect 3080 130 3110 160
rect 3310 130 3340 160
rect 3540 130 3570 160
rect 3770 130 3800 160
rect 4000 130 4030 160
rect 4230 130 4260 160
rect 4460 130 4490 160
rect 4690 130 4720 160
rect 4920 130 4950 160
rect 5150 130 5180 160
rect 5380 130 5410 160
rect 5610 130 5640 160
rect 5840 130 5870 160
rect 6070 130 6100 160
rect 6300 130 6330 160
rect 6530 130 6560 160
rect 6760 130 6790 160
rect 90 -50 120 -20
rect 320 -50 350 -20
rect 550 -50 580 -20
rect 780 -50 810 -20
rect 1010 -50 1040 -20
rect 1240 -50 1270 -20
rect 1470 -50 1500 -20
rect 1700 -50 1730 -20
rect 1930 -50 1960 -20
rect 2160 -50 2190 -20
rect 2390 -50 2420 -20
rect 2620 -50 2650 -20
rect 2850 -50 2880 -20
rect 3080 -50 3110 -20
rect 3310 -50 3340 -20
rect 3540 -50 3570 -20
rect 3770 -50 3800 -20
rect 4000 -50 4030 -20
rect 4230 -50 4260 -20
rect 4460 -50 4490 -20
rect 4690 -50 4720 -20
rect 4920 -50 4950 -20
rect 5150 -50 5180 -20
rect 5380 -50 5410 -20
rect 5610 -50 5640 -20
rect 5840 -50 5870 -20
rect 6070 -50 6100 -20
rect 6300 -50 6330 -20
rect 6530 -50 6560 -20
rect 6760 -50 6790 -20
rect 90 -570 120 -550
rect 320 -570 350 -550
rect 550 -570 580 -550
rect 780 -570 810 -550
rect 1010 -570 1040 -550
rect 1240 -570 1270 -550
rect 1470 -570 1500 -550
rect 1700 -570 1730 -550
rect 1930 -570 1960 -550
rect 2160 -570 2190 -550
rect 2390 -570 2420 -550
rect 2620 -570 2650 -550
rect 2850 -570 2880 -550
rect 3080 -570 3110 -550
rect 3310 -570 3340 -550
rect 3540 -570 3570 -550
rect 3770 -570 3800 -550
rect 4000 -570 4030 -550
rect 4230 -570 4260 -550
rect 4460 -570 4490 -550
rect 4690 -570 4720 -550
rect 4920 -570 4950 -550
rect 5150 -570 5180 -550
rect 5380 -570 5410 -550
rect 5610 -570 5640 -550
rect 5840 -570 5870 -550
rect 6070 -570 6100 -550
rect 6300 -570 6330 -550
rect 6530 -570 6560 -550
rect 6760 -570 6790 -550
rect 50 -590 160 -570
rect 50 -660 70 -590
rect 140 -660 160 -590
rect 50 -680 160 -660
rect 280 -590 390 -570
rect 280 -660 300 -590
rect 370 -660 390 -590
rect 280 -680 390 -660
rect 510 -590 620 -570
rect 510 -660 530 -590
rect 600 -660 620 -590
rect 510 -680 620 -660
rect 740 -590 850 -570
rect 740 -660 760 -590
rect 830 -660 850 -590
rect 740 -680 850 -660
rect 970 -590 1080 -570
rect 970 -660 990 -590
rect 1060 -660 1080 -590
rect 970 -680 1080 -660
rect 1200 -590 1310 -570
rect 1200 -660 1220 -590
rect 1290 -660 1310 -590
rect 1200 -680 1310 -660
rect 1430 -590 1540 -570
rect 1430 -660 1450 -590
rect 1520 -660 1540 -590
rect 1430 -680 1540 -660
rect 1660 -590 1770 -570
rect 1660 -660 1680 -590
rect 1750 -660 1770 -590
rect 1660 -680 1770 -660
rect 1890 -590 2000 -570
rect 1890 -660 1910 -590
rect 1980 -660 2000 -590
rect 1890 -680 2000 -660
rect 2120 -590 2230 -570
rect 2120 -660 2140 -590
rect 2210 -660 2230 -590
rect 2120 -680 2230 -660
rect 2350 -590 2460 -570
rect 2350 -660 2370 -590
rect 2440 -660 2460 -590
rect 2350 -680 2460 -660
rect 2580 -590 2690 -570
rect 2580 -660 2600 -590
rect 2670 -660 2690 -590
rect 2580 -680 2690 -660
rect 2810 -590 2920 -570
rect 2810 -660 2830 -590
rect 2900 -660 2920 -590
rect 2810 -680 2920 -660
rect 3040 -590 3150 -570
rect 3040 -660 3060 -590
rect 3130 -660 3150 -590
rect 3040 -680 3150 -660
rect 3270 -590 3380 -570
rect 3270 -660 3290 -590
rect 3360 -660 3380 -590
rect 3270 -680 3380 -660
rect 3500 -590 3610 -570
rect 3500 -660 3520 -590
rect 3590 -660 3610 -590
rect 3500 -680 3610 -660
rect 3730 -590 3840 -570
rect 3730 -660 3750 -590
rect 3820 -660 3840 -590
rect 3730 -680 3840 -660
rect 3960 -590 4070 -570
rect 3960 -660 3980 -590
rect 4050 -660 4070 -590
rect 3960 -680 4070 -660
rect 4190 -590 4300 -570
rect 4190 -660 4210 -590
rect 4280 -660 4300 -590
rect 4190 -680 4300 -660
rect 4420 -590 4530 -570
rect 4420 -660 4440 -590
rect 4510 -660 4530 -590
rect 4420 -680 4530 -660
rect 4650 -590 4760 -570
rect 4650 -660 4670 -590
rect 4740 -660 4760 -590
rect 4650 -680 4760 -660
rect 4880 -590 4990 -570
rect 4880 -660 4900 -590
rect 4970 -660 4990 -590
rect 4880 -680 4990 -660
rect 5110 -590 5220 -570
rect 5110 -660 5130 -590
rect 5200 -660 5220 -590
rect 5110 -680 5220 -660
rect 5340 -590 5450 -570
rect 5340 -660 5360 -590
rect 5430 -660 5450 -590
rect 5340 -680 5450 -660
rect 5570 -590 5680 -570
rect 5570 -660 5590 -590
rect 5660 -660 5680 -590
rect 5570 -680 5680 -660
rect 5800 -590 5910 -570
rect 5800 -660 5820 -590
rect 5890 -660 5910 -590
rect 5800 -680 5910 -660
rect 6030 -590 6140 -570
rect 6030 -660 6050 -590
rect 6120 -660 6140 -590
rect 6030 -680 6140 -660
rect 6260 -590 6370 -570
rect 6260 -660 6280 -590
rect 6350 -660 6370 -590
rect 6260 -680 6370 -660
rect 6490 -590 6600 -570
rect 6490 -660 6510 -590
rect 6580 -660 6600 -590
rect 6490 -680 6600 -660
rect 6720 -590 6830 -570
rect 6720 -660 6740 -590
rect 6810 -660 6830 -590
rect 6720 -680 6830 -660
rect 2290 -1050 2350 -1020
rect 2550 -1050 2610 -1020
rect 2810 -1050 2870 -1020
rect 3070 -1050 3130 -1020
rect 3330 -1050 3390 -1020
rect 3590 -1050 3650 -1020
rect 3850 -1050 3910 -1020
rect 4110 -1050 4170 -1020
rect 4370 -1050 4430 -1020
rect 4630 -1050 4690 -1020
rect 4890 -1050 4950 -1020
rect 5150 -1050 5210 -1020
rect 5410 -1050 5470 -1020
rect 5670 -1050 5730 -1020
rect 5930 -1050 5990 -1020
rect 6190 -1050 6250 -1020
rect 6450 -1050 6510 -1020
rect 6710 -1050 6770 -1020
rect 2290 -1680 2350 -1650
rect 2550 -1680 2610 -1650
rect 2810 -1680 2870 -1650
rect 3070 -1680 3130 -1650
rect 3330 -1680 3390 -1650
rect 3590 -1680 3650 -1650
rect 3850 -1680 3910 -1650
rect 4110 -1680 4170 -1650
rect 4370 -1680 4430 -1650
rect 4630 -1680 4690 -1650
rect 4890 -1680 4950 -1650
rect 5150 -1680 5210 -1650
rect 5410 -1680 5470 -1650
rect 5670 -1680 5730 -1650
rect 5930 -1680 5990 -1650
rect 6190 -1680 6250 -1650
rect 6450 -1680 6510 -1650
rect 6710 -1680 6770 -1650
rect 2260 -1700 2380 -1680
rect 2260 -1770 2280 -1700
rect 2360 -1770 2380 -1700
rect 2260 -1790 2380 -1770
rect 2520 -1700 2640 -1680
rect 2520 -1770 2540 -1700
rect 2620 -1770 2640 -1700
rect 2520 -1790 2640 -1770
rect 2780 -1700 2900 -1680
rect 2780 -1770 2800 -1700
rect 2880 -1770 2900 -1700
rect 2780 -1790 2900 -1770
rect 3040 -1700 3160 -1680
rect 3040 -1770 3060 -1700
rect 3140 -1770 3160 -1700
rect 3040 -1790 3160 -1770
rect 3300 -1700 3420 -1680
rect 3300 -1770 3320 -1700
rect 3400 -1770 3420 -1700
rect 3300 -1790 3420 -1770
rect 3560 -1700 3680 -1680
rect 3560 -1770 3580 -1700
rect 3660 -1770 3680 -1700
rect 3560 -1790 3680 -1770
rect 3820 -1700 3940 -1680
rect 3820 -1770 3840 -1700
rect 3920 -1770 3940 -1700
rect 3820 -1790 3940 -1770
rect 4080 -1700 4200 -1680
rect 4080 -1770 4100 -1700
rect 4180 -1770 4200 -1700
rect 4080 -1790 4200 -1770
rect 4340 -1700 4460 -1680
rect 4340 -1770 4360 -1700
rect 4440 -1770 4460 -1700
rect 4340 -1790 4460 -1770
rect 4600 -1700 4720 -1680
rect 4600 -1770 4620 -1700
rect 4700 -1770 4720 -1700
rect 4600 -1790 4720 -1770
rect 4860 -1700 4980 -1680
rect 4860 -1770 4880 -1700
rect 4960 -1770 4980 -1700
rect 4860 -1790 4980 -1770
rect 5120 -1700 5240 -1680
rect 5120 -1770 5140 -1700
rect 5220 -1770 5240 -1700
rect 5120 -1790 5240 -1770
rect 5380 -1700 5500 -1680
rect 5380 -1770 5400 -1700
rect 5480 -1770 5500 -1700
rect 5380 -1790 5500 -1770
rect 5640 -1700 5760 -1680
rect 5640 -1770 5660 -1700
rect 5740 -1770 5760 -1700
rect 5640 -1790 5760 -1770
rect 5900 -1700 6020 -1680
rect 5900 -1770 5920 -1700
rect 6000 -1770 6020 -1700
rect 5900 -1790 6020 -1770
rect 6160 -1700 6280 -1680
rect 6160 -1770 6180 -1700
rect 6260 -1770 6280 -1700
rect 6160 -1790 6280 -1770
rect 6420 -1700 6540 -1680
rect 6420 -1770 6440 -1700
rect 6520 -1770 6540 -1700
rect 6420 -1790 6540 -1770
rect 6680 -1700 6800 -1680
rect 6680 -1770 6700 -1700
rect 6780 -1770 6800 -1700
rect 6680 -1790 6800 -1770
<< polycont >>
rect 1540 1810 1620 1880
rect 1800 1810 1880 1880
rect 2330 1810 2410 1880
rect 2590 1810 2670 1880
rect 2850 1810 2930 1880
rect 3110 1810 3190 1880
rect 3370 1810 3450 1880
rect 3630 1810 3710 1880
rect 3890 1810 3970 1880
rect 4150 1810 4230 1880
rect 4410 1810 4490 1880
rect 4670 1810 4750 1880
rect 4930 1810 5010 1880
rect 5190 1810 5270 1880
rect 5450 1810 5530 1880
rect 5710 1810 5790 1880
rect 5970 1810 6050 1880
rect 6230 1810 6310 1880
rect 6490 1810 6570 1880
rect 6750 1810 6830 1880
rect 70 700 140 770
rect 300 700 370 770
rect 530 700 600 770
rect 760 700 830 770
rect 990 700 1060 770
rect 1220 700 1290 770
rect 1450 700 1520 770
rect 1680 700 1750 770
rect 1910 700 1980 770
rect 2140 700 2210 770
rect 2370 700 2440 770
rect 2600 700 2670 770
rect 2830 700 2900 770
rect 3060 700 3130 770
rect 3290 700 3360 770
rect 3520 700 3590 770
rect 3750 700 3820 770
rect 3980 700 4050 770
rect 4210 700 4280 770
rect 4440 700 4510 770
rect 4670 700 4740 770
rect 4900 700 4970 770
rect 5130 700 5200 770
rect 5360 700 5430 770
rect 5590 700 5660 770
rect 5820 700 5890 770
rect 6050 700 6120 770
rect 6280 700 6350 770
rect 6510 700 6580 770
rect 6740 700 6810 770
rect 70 -660 140 -590
rect 300 -660 370 -590
rect 530 -660 600 -590
rect 760 -660 830 -590
rect 990 -660 1060 -590
rect 1220 -660 1290 -590
rect 1450 -660 1520 -590
rect 1680 -660 1750 -590
rect 1910 -660 1980 -590
rect 2140 -660 2210 -590
rect 2370 -660 2440 -590
rect 2600 -660 2670 -590
rect 2830 -660 2900 -590
rect 3060 -660 3130 -590
rect 3290 -660 3360 -590
rect 3520 -660 3590 -590
rect 3750 -660 3820 -590
rect 3980 -660 4050 -590
rect 4210 -660 4280 -590
rect 4440 -660 4510 -590
rect 4670 -660 4740 -590
rect 4900 -660 4970 -590
rect 5130 -660 5200 -590
rect 5360 -660 5430 -590
rect 5590 -660 5660 -590
rect 5820 -660 5890 -590
rect 6050 -660 6120 -590
rect 6280 -660 6350 -590
rect 6510 -660 6580 -590
rect 6740 -660 6810 -590
rect 2280 -1770 2360 -1700
rect 2540 -1770 2620 -1700
rect 2800 -1770 2880 -1700
rect 3060 -1770 3140 -1700
rect 3320 -1770 3400 -1700
rect 3580 -1770 3660 -1700
rect 3840 -1770 3920 -1700
rect 4100 -1770 4180 -1700
rect 4360 -1770 4440 -1700
rect 4620 -1770 4700 -1700
rect 4880 -1770 4960 -1700
rect 5140 -1770 5220 -1700
rect 5400 -1770 5480 -1700
rect 5660 -1770 5740 -1700
rect 5920 -1770 6000 -1700
rect 6180 -1770 6260 -1700
rect 6440 -1770 6520 -1700
rect 6700 -1770 6780 -1700
<< locali >>
rect -2100 2484 8350 2594
rect -2100 2324 -660 2484
rect -2100 2124 -1960 2324
rect -1760 2284 -660 2324
rect -460 2284 340 2484
rect 540 2284 1340 2484
rect 1540 2284 2360 2484
rect 2560 2284 3360 2484
rect 3560 2284 4360 2484
rect 4560 2284 5380 2484
rect 5580 2284 6380 2484
rect 6580 2284 7380 2484
rect 7580 2284 8350 2484
rect -1760 2254 8350 2284
rect -1760 2144 8020 2254
rect -1760 2124 -1650 2144
rect -2100 1280 -1650 2124
rect 7900 2030 8020 2144
rect 8220 2030 8350 2254
rect 1520 1880 1640 1900
rect 1520 1810 1540 1880
rect 1620 1810 1640 1880
rect 1520 1790 1640 1810
rect 1780 1880 1900 1900
rect 1780 1810 1800 1880
rect 1880 1810 1900 1880
rect 1780 1790 1900 1810
rect 2310 1880 2430 1900
rect 2310 1810 2330 1880
rect 2410 1810 2430 1880
rect 2310 1790 2430 1810
rect 2570 1880 2690 1900
rect 2570 1810 2590 1880
rect 2670 1810 2690 1880
rect 2570 1790 2690 1810
rect 2830 1880 2950 1900
rect 2830 1810 2850 1880
rect 2930 1810 2950 1880
rect 2830 1790 2950 1810
rect 3090 1880 3210 1900
rect 3090 1810 3110 1880
rect 3190 1810 3210 1880
rect 3090 1790 3210 1810
rect 3350 1880 3470 1900
rect 3350 1810 3370 1880
rect 3450 1810 3470 1880
rect 3350 1790 3470 1810
rect 3610 1880 3730 1900
rect 3610 1810 3630 1880
rect 3710 1810 3730 1880
rect 3610 1790 3730 1810
rect 3870 1880 3990 1900
rect 3870 1810 3890 1880
rect 3970 1810 3990 1880
rect 3870 1790 3990 1810
rect 4130 1880 4250 1900
rect 4130 1810 4150 1880
rect 4230 1810 4250 1880
rect 4130 1790 4250 1810
rect 4390 1880 4510 1900
rect 4390 1810 4410 1880
rect 4490 1810 4510 1880
rect 4390 1790 4510 1810
rect 4650 1880 4770 1900
rect 4650 1810 4670 1880
rect 4750 1810 4770 1880
rect 4650 1790 4770 1810
rect 4910 1880 5030 1900
rect 4910 1810 4930 1880
rect 5010 1810 5030 1880
rect 4910 1790 5030 1810
rect 5170 1880 5290 1900
rect 5170 1810 5190 1880
rect 5270 1810 5290 1880
rect 5170 1790 5290 1810
rect 5430 1880 5550 1900
rect 5430 1810 5450 1880
rect 5530 1810 5550 1880
rect 5430 1790 5550 1810
rect 5690 1880 5810 1900
rect 5690 1810 5710 1880
rect 5790 1810 5810 1880
rect 5690 1790 5810 1810
rect 5950 1880 6070 1900
rect 5950 1810 5970 1880
rect 6050 1810 6070 1880
rect 5950 1790 6070 1810
rect 6210 1880 6330 1900
rect 6210 1810 6230 1880
rect 6310 1810 6330 1880
rect 6210 1790 6330 1810
rect 6470 1880 6590 1900
rect 6470 1810 6490 1880
rect 6570 1810 6590 1880
rect 6470 1790 6590 1810
rect 6730 1880 6850 1900
rect 6730 1810 6750 1880
rect 6830 1810 6850 1880
rect 6730 1790 6850 1810
rect 7090 1720 7320 1760
rect 1380 1680 1520 1700
rect 1380 1580 1400 1680
rect 1500 1580 1520 1680
rect 1380 1560 1520 1580
rect 1640 1680 1780 1700
rect 1640 1580 1660 1680
rect 1760 1580 1780 1680
rect 1640 1560 1780 1580
rect 1900 1680 2040 1700
rect 1900 1580 1920 1680
rect 2020 1580 2040 1680
rect 1900 1560 2040 1580
rect 2170 1680 2310 1700
rect 2170 1580 2190 1680
rect 2290 1580 2310 1680
rect 2170 1560 2310 1580
rect 2430 1680 2570 1700
rect 2430 1580 2450 1680
rect 2550 1580 2570 1680
rect 2430 1560 2570 1580
rect 2690 1680 2830 1700
rect 2690 1580 2710 1680
rect 2810 1580 2830 1680
rect 2690 1560 2830 1580
rect 2950 1680 3090 1700
rect 2950 1580 2970 1680
rect 3070 1580 3090 1680
rect 2950 1560 3090 1580
rect 3210 1680 3350 1700
rect 3210 1580 3230 1680
rect 3330 1580 3350 1680
rect 3210 1560 3350 1580
rect 3470 1680 3610 1700
rect 3470 1580 3490 1680
rect 3590 1580 3610 1680
rect 3470 1560 3610 1580
rect 3730 1680 3870 1700
rect 3730 1580 3750 1680
rect 3850 1580 3870 1680
rect 3730 1560 3870 1580
rect 3990 1680 4130 1700
rect 3990 1580 4010 1680
rect 4110 1580 4130 1680
rect 3990 1560 4130 1580
rect 4250 1680 4390 1700
rect 4250 1580 4270 1680
rect 4370 1580 4390 1680
rect 4250 1560 4390 1580
rect 4510 1680 4650 1700
rect 4510 1580 4530 1680
rect 4630 1580 4650 1680
rect 4510 1560 4650 1580
rect 4770 1680 4910 1700
rect 4770 1580 4790 1680
rect 4890 1580 4910 1680
rect 4770 1560 4910 1580
rect 5030 1680 5170 1700
rect 5030 1580 5050 1680
rect 5150 1580 5170 1680
rect 5030 1560 5170 1580
rect 5290 1680 5430 1700
rect 5290 1580 5310 1680
rect 5410 1580 5430 1680
rect 5290 1560 5430 1580
rect 5550 1680 5690 1700
rect 5550 1580 5570 1680
rect 5670 1580 5690 1680
rect 5550 1560 5690 1580
rect 5810 1680 5950 1700
rect 5810 1580 5830 1680
rect 5930 1580 5950 1680
rect 5810 1560 5950 1580
rect 6070 1680 6210 1700
rect 6070 1580 6090 1680
rect 6190 1580 6210 1680
rect 6070 1560 6210 1580
rect 6330 1680 6470 1700
rect 6330 1580 6350 1680
rect 6450 1580 6470 1680
rect 6330 1560 6470 1580
rect 6590 1680 6730 1700
rect 6590 1580 6610 1680
rect 6710 1580 6730 1680
rect 6590 1560 6730 1580
rect 6850 1680 6990 1700
rect 6850 1580 6870 1680
rect 6970 1580 6990 1680
rect 6850 1560 6990 1580
rect 7090 1540 7130 1720
rect 7290 1540 7320 1720
rect 7090 1510 7320 1540
rect 7900 1520 8350 2030
rect 1380 1400 1520 1420
rect 1380 1300 1400 1400
rect 1500 1300 1520 1400
rect 1380 1280 1520 1300
rect 1640 1400 1780 1420
rect 1640 1300 1660 1400
rect 1760 1300 1780 1400
rect 1640 1280 1780 1300
rect 1900 1400 2040 1420
rect 1900 1300 1920 1400
rect 2020 1300 2040 1400
rect 1900 1280 2040 1300
rect 2170 1340 2310 1360
rect -2100 1080 -1960 1280
rect -1760 1080 -1650 1280
rect 2170 1240 2190 1340
rect 2290 1240 2310 1340
rect 2170 1220 2310 1240
rect 2430 1340 2570 1360
rect 2430 1240 2450 1340
rect 2550 1240 2570 1340
rect 2430 1220 2570 1240
rect 2690 1340 2830 1360
rect 2690 1240 2710 1340
rect 2810 1240 2830 1340
rect 2690 1220 2830 1240
rect 2950 1340 3090 1360
rect 2950 1240 2970 1340
rect 3070 1240 3090 1340
rect 2950 1220 3090 1240
rect 3210 1340 3350 1360
rect 3210 1240 3230 1340
rect 3330 1240 3350 1340
rect 3210 1220 3350 1240
rect 3470 1340 3610 1360
rect 3470 1240 3490 1340
rect 3590 1240 3610 1340
rect 3470 1220 3610 1240
rect 3730 1340 3870 1360
rect 3730 1240 3750 1340
rect 3850 1240 3870 1340
rect 3730 1220 3870 1240
rect 3990 1340 4130 1360
rect 3990 1240 4010 1340
rect 4110 1240 4130 1340
rect 3990 1220 4130 1240
rect 4250 1340 4390 1360
rect 4250 1240 4270 1340
rect 4370 1240 4390 1340
rect 4250 1220 4390 1240
rect 4510 1340 4650 1360
rect 4510 1240 4530 1340
rect 4630 1240 4650 1340
rect 4510 1220 4650 1240
rect 4770 1340 4910 1360
rect 4770 1240 4790 1340
rect 4890 1240 4910 1340
rect 4770 1220 4910 1240
rect 5030 1340 5170 1360
rect 5030 1240 5050 1340
rect 5150 1240 5170 1340
rect 5030 1220 5170 1240
rect 5290 1340 5430 1360
rect 5290 1240 5310 1340
rect 5410 1240 5430 1340
rect 5290 1220 5430 1240
rect 5550 1340 5690 1360
rect 5550 1240 5570 1340
rect 5670 1240 5690 1340
rect 5550 1220 5690 1240
rect 5810 1340 5950 1360
rect 5810 1240 5830 1340
rect 5930 1240 5950 1340
rect 5810 1220 5950 1240
rect 6070 1340 6210 1360
rect 6070 1240 6090 1340
rect 6190 1240 6210 1340
rect 6070 1220 6210 1240
rect 6330 1340 6470 1360
rect 6330 1240 6350 1340
rect 6450 1240 6470 1340
rect 6330 1220 6470 1240
rect 6590 1340 6730 1360
rect 6590 1240 6610 1340
rect 6710 1240 6730 1340
rect 6590 1220 6730 1240
rect 6850 1340 6990 1360
rect 6850 1240 6870 1340
rect 6970 1240 6990 1340
rect 6850 1220 6990 1240
rect 7900 1320 8020 1520
rect 8220 1320 8350 1520
rect -2100 570 -1650 1080
rect 7900 830 8350 1320
rect 50 770 160 790
rect 50 700 70 770
rect 140 700 160 770
rect 50 680 160 700
rect 280 770 390 790
rect 280 700 300 770
rect 370 700 390 770
rect 280 680 390 700
rect 510 770 620 790
rect 510 700 530 770
rect 600 700 620 770
rect 510 680 620 700
rect 740 770 850 790
rect 740 700 760 770
rect 830 700 850 770
rect 740 680 850 700
rect 970 770 1080 790
rect 970 700 990 770
rect 1060 700 1080 770
rect 970 680 1080 700
rect 1200 770 1310 790
rect 1200 700 1220 770
rect 1290 700 1310 770
rect 1200 680 1310 700
rect 1430 770 1540 790
rect 1430 700 1450 770
rect 1520 700 1540 770
rect 1430 680 1540 700
rect 1660 770 1770 790
rect 1660 700 1680 770
rect 1750 700 1770 770
rect 1660 680 1770 700
rect 1890 770 2000 790
rect 1890 700 1910 770
rect 1980 700 2000 770
rect 1890 680 2000 700
rect 2120 770 2230 790
rect 2120 700 2140 770
rect 2210 700 2230 770
rect 2120 680 2230 700
rect 2350 770 2460 790
rect 2350 700 2370 770
rect 2440 700 2460 770
rect 2350 680 2460 700
rect 2580 770 2690 790
rect 2580 700 2600 770
rect 2670 700 2690 770
rect 2580 680 2690 700
rect 2810 770 2920 790
rect 2810 700 2830 770
rect 2900 700 2920 770
rect 2810 680 2920 700
rect 3040 770 3150 790
rect 3040 700 3060 770
rect 3130 700 3150 770
rect 3040 680 3150 700
rect 3270 770 3380 790
rect 3270 700 3290 770
rect 3360 700 3380 770
rect 3270 680 3380 700
rect 3500 770 3610 790
rect 3500 700 3520 770
rect 3590 700 3610 770
rect 3500 680 3610 700
rect 3730 770 3840 790
rect 3730 700 3750 770
rect 3820 700 3840 770
rect 3730 680 3840 700
rect 3960 770 4070 790
rect 3960 700 3980 770
rect 4050 700 4070 770
rect 3960 680 4070 700
rect 4190 770 4300 790
rect 4190 700 4210 770
rect 4280 700 4300 770
rect 4190 680 4300 700
rect 4420 770 4530 790
rect 4420 700 4440 770
rect 4510 700 4530 770
rect 4420 680 4530 700
rect 4650 770 4760 790
rect 4650 700 4670 770
rect 4740 700 4760 770
rect 4650 680 4760 700
rect 4880 770 4990 790
rect 4880 700 4900 770
rect 4970 700 4990 770
rect 4880 680 4990 700
rect 5110 770 5220 790
rect 5110 700 5130 770
rect 5200 700 5220 770
rect 5110 680 5220 700
rect 5340 770 5450 790
rect 5340 700 5360 770
rect 5430 700 5450 770
rect 5340 680 5450 700
rect 5570 770 5680 790
rect 5570 700 5590 770
rect 5660 700 5680 770
rect 5570 680 5680 700
rect 5800 770 5910 790
rect 5800 700 5820 770
rect 5890 700 5910 770
rect 5800 680 5910 700
rect 6030 770 6140 790
rect 6030 700 6050 770
rect 6120 700 6140 770
rect 6030 680 6140 700
rect 6260 770 6370 790
rect 6260 700 6280 770
rect 6350 700 6370 770
rect 6260 680 6370 700
rect 6490 770 6600 790
rect 6490 700 6510 770
rect 6580 700 6600 770
rect 6490 680 6600 700
rect 6720 770 6830 790
rect 6720 700 6740 770
rect 6810 700 6830 770
rect 6720 680 6830 700
rect 7900 630 8040 830
rect 8240 630 8350 830
rect -2100 370 -1960 570
rect -1760 370 -1650 570
rect -80 610 60 630
rect -80 510 -60 610
rect 40 510 60 610
rect -80 490 60 510
rect 150 610 290 630
rect 150 510 170 610
rect 270 510 290 610
rect 150 490 290 510
rect 380 610 520 630
rect 380 510 400 610
rect 500 510 520 610
rect 380 490 520 510
rect 610 610 750 630
rect 610 510 630 610
rect 730 510 750 610
rect 610 490 750 510
rect 840 610 980 630
rect 840 510 860 610
rect 960 510 980 610
rect 840 490 980 510
rect 1070 610 1210 630
rect 1070 510 1090 610
rect 1190 510 1210 610
rect 1070 490 1210 510
rect 1300 610 1440 630
rect 1300 510 1320 610
rect 1420 510 1440 610
rect 1300 490 1440 510
rect 1530 610 1670 630
rect 1530 510 1550 610
rect 1650 510 1670 610
rect 1530 490 1670 510
rect 1760 610 1900 630
rect 1760 510 1780 610
rect 1880 510 1900 610
rect 1760 490 1900 510
rect 1990 610 2130 630
rect 1990 510 2010 610
rect 2110 510 2130 610
rect 1990 490 2130 510
rect 2220 610 2360 630
rect 2220 510 2240 610
rect 2340 510 2360 610
rect 2220 490 2360 510
rect 2450 610 2590 630
rect 2450 510 2470 610
rect 2570 510 2590 610
rect 2450 490 2590 510
rect 2680 610 2820 630
rect 2680 510 2700 610
rect 2800 510 2820 610
rect 2680 490 2820 510
rect 2910 610 3050 630
rect 2910 510 2930 610
rect 3030 510 3050 610
rect 2910 490 3050 510
rect 3140 610 3280 630
rect 3140 510 3160 610
rect 3260 510 3280 610
rect 3140 490 3280 510
rect 3370 610 3510 630
rect 3370 510 3390 610
rect 3490 510 3510 610
rect 3370 490 3510 510
rect 3600 610 3740 630
rect 3600 510 3620 610
rect 3720 510 3740 610
rect 3600 490 3740 510
rect 3830 610 3970 630
rect 3830 510 3850 610
rect 3950 510 3970 610
rect 3830 490 3970 510
rect 4060 610 4200 630
rect 4060 510 4080 610
rect 4180 510 4200 610
rect 4060 490 4200 510
rect 4290 610 4430 630
rect 4290 510 4310 610
rect 4410 510 4430 610
rect 4290 490 4430 510
rect 4520 610 4660 630
rect 4520 510 4540 610
rect 4640 510 4660 610
rect 4520 490 4660 510
rect 4750 610 4890 630
rect 4750 510 4770 610
rect 4870 510 4890 610
rect 4750 490 4890 510
rect 4980 610 5120 630
rect 4980 510 5000 610
rect 5100 510 5120 610
rect 4980 490 5120 510
rect 5210 610 5350 630
rect 5210 510 5230 610
rect 5330 510 5350 610
rect 5210 490 5350 510
rect 5440 610 5580 630
rect 5440 510 5460 610
rect 5560 510 5580 610
rect 5440 490 5580 510
rect 5670 610 5810 630
rect 5670 510 5690 610
rect 5790 510 5810 610
rect 5670 490 5810 510
rect 5900 610 6040 630
rect 5900 510 5920 610
rect 6020 510 6040 610
rect 5900 490 6040 510
rect 6130 610 6270 630
rect 6130 510 6150 610
rect 6250 510 6270 610
rect 6130 490 6270 510
rect 6360 610 6500 630
rect 6360 510 6380 610
rect 6480 510 6500 610
rect 6360 490 6500 510
rect 6590 610 6730 630
rect 6590 510 6610 610
rect 6710 510 6730 610
rect 6590 490 6730 510
rect 6820 610 6960 630
rect 6820 510 6840 610
rect 6940 510 6960 610
rect 6820 490 6960 510
rect -2100 -450 -1650 370
rect -80 310 60 330
rect -80 210 -60 310
rect 40 210 60 310
rect -80 190 60 210
rect 150 310 290 330
rect 150 210 170 310
rect 270 210 290 310
rect 150 190 290 210
rect 380 310 520 330
rect 380 210 400 310
rect 500 210 520 310
rect 380 190 520 210
rect 610 310 750 330
rect 610 210 630 310
rect 730 210 750 310
rect 610 190 750 210
rect 840 310 980 330
rect 840 210 860 310
rect 960 210 980 310
rect 840 190 980 210
rect 1070 310 1210 330
rect 1070 210 1090 310
rect 1190 210 1210 310
rect 1070 190 1210 210
rect 1300 310 1440 330
rect 1300 210 1320 310
rect 1420 210 1440 310
rect 1300 190 1440 210
rect 1530 310 1670 330
rect 1530 210 1550 310
rect 1650 210 1670 310
rect 1530 190 1670 210
rect 1760 310 1900 330
rect 1760 210 1780 310
rect 1880 210 1900 310
rect 1760 190 1900 210
rect 1990 310 2130 330
rect 1990 210 2010 310
rect 2110 210 2130 310
rect 1990 190 2130 210
rect 2220 310 2360 330
rect 2220 210 2240 310
rect 2340 210 2360 310
rect 2220 190 2360 210
rect 2450 310 2590 330
rect 2450 210 2470 310
rect 2570 210 2590 310
rect 2450 190 2590 210
rect 2680 310 2820 330
rect 2680 210 2700 310
rect 2800 210 2820 310
rect 2680 190 2820 210
rect 2910 310 3050 330
rect 2910 210 2930 310
rect 3030 210 3050 310
rect 2910 190 3050 210
rect 3140 310 3280 330
rect 3140 210 3160 310
rect 3260 210 3280 310
rect 3140 190 3280 210
rect 3370 310 3510 330
rect 3370 210 3390 310
rect 3490 210 3510 310
rect 3370 190 3510 210
rect 3600 310 3740 330
rect 3600 210 3620 310
rect 3720 210 3740 310
rect 3600 190 3740 210
rect 3830 310 3970 330
rect 3830 210 3850 310
rect 3950 210 3970 310
rect 3830 190 3970 210
rect 4060 310 4200 330
rect 4060 210 4080 310
rect 4180 210 4200 310
rect 4060 190 4200 210
rect 4290 310 4430 330
rect 4290 210 4310 310
rect 4410 210 4430 310
rect 4290 190 4430 210
rect 4520 310 4660 330
rect 4520 210 4540 310
rect 4640 210 4660 310
rect 4520 190 4660 210
rect 4750 310 4890 330
rect 4750 210 4770 310
rect 4870 210 4890 310
rect 4750 190 4890 210
rect 4980 310 5120 330
rect 4980 210 5000 310
rect 5100 210 5120 310
rect 4980 190 5120 210
rect 5210 310 5350 330
rect 5210 210 5230 310
rect 5330 210 5350 310
rect 5210 190 5350 210
rect 5440 310 5580 330
rect 5440 210 5460 310
rect 5560 210 5580 310
rect 5440 190 5580 210
rect 5670 310 5810 330
rect 5670 210 5690 310
rect 5790 210 5810 310
rect 5670 190 5810 210
rect 5900 310 6040 330
rect 5900 210 5920 310
rect 6020 210 6040 310
rect 5900 190 6040 210
rect 6130 310 6270 330
rect 6130 210 6150 310
rect 6250 210 6270 310
rect 6130 190 6270 210
rect 6360 310 6500 330
rect 6360 210 6380 310
rect 6480 210 6500 310
rect 6360 190 6500 210
rect 6590 310 6730 330
rect 6590 210 6610 310
rect 6710 210 6730 310
rect 6590 190 6730 210
rect 6820 310 6960 330
rect 6820 210 6840 310
rect 6940 210 6960 310
rect 6820 190 6960 210
rect 1320 90 1490 100
rect 1320 20 1340 90
rect 1470 20 1490 90
rect 1320 10 1490 20
rect -80 -100 60 -80
rect -80 -200 -60 -100
rect 40 -200 60 -100
rect -80 -220 60 -200
rect 150 -100 290 -80
rect 150 -200 170 -100
rect 270 -200 290 -100
rect 150 -220 290 -200
rect 380 -100 520 -80
rect 380 -200 400 -100
rect 500 -200 520 -100
rect 380 -220 520 -200
rect 610 -100 750 -80
rect 610 -200 630 -100
rect 730 -200 750 -100
rect 610 -220 750 -200
rect 840 -100 980 -80
rect 840 -200 860 -100
rect 960 -200 980 -100
rect 840 -220 980 -200
rect 1070 -100 1210 -80
rect 1070 -200 1090 -100
rect 1190 -200 1210 -100
rect 1070 -220 1210 -200
rect 1300 -100 1440 -80
rect 1300 -200 1320 -100
rect 1420 -200 1440 -100
rect 1300 -220 1440 -200
rect 1530 -100 1670 -80
rect 1530 -200 1550 -100
rect 1650 -200 1670 -100
rect 1530 -220 1670 -200
rect 1760 -100 1900 -80
rect 1760 -200 1780 -100
rect 1880 -200 1900 -100
rect 1760 -220 1900 -200
rect 1990 -100 2130 -80
rect 1990 -200 2010 -100
rect 2110 -200 2130 -100
rect 1990 -220 2130 -200
rect 2220 -100 2360 -80
rect 2220 -200 2240 -100
rect 2340 -200 2360 -100
rect 2220 -220 2360 -200
rect 2450 -100 2590 -80
rect 2450 -200 2470 -100
rect 2570 -200 2590 -100
rect 2450 -220 2590 -200
rect 2680 -100 2820 -80
rect 2680 -200 2700 -100
rect 2800 -200 2820 -100
rect 2680 -220 2820 -200
rect 2910 -100 3050 -80
rect 2910 -200 2930 -100
rect 3030 -200 3050 -100
rect 2910 -220 3050 -200
rect 3140 -100 3280 -80
rect 3140 -200 3160 -100
rect 3260 -200 3280 -100
rect 3140 -220 3280 -200
rect 3370 -100 3510 -80
rect 3370 -200 3390 -100
rect 3490 -200 3510 -100
rect 3370 -220 3510 -200
rect 3600 -100 3740 -80
rect 3600 -200 3620 -100
rect 3720 -200 3740 -100
rect 3600 -220 3740 -200
rect 3830 -100 3970 -80
rect 3830 -200 3850 -100
rect 3950 -200 3970 -100
rect 3830 -220 3970 -200
rect 4060 -100 4200 -80
rect 4060 -200 4080 -100
rect 4180 -200 4200 -100
rect 4060 -220 4200 -200
rect 4290 -100 4430 -80
rect 4290 -200 4310 -100
rect 4410 -200 4430 -100
rect 4290 -220 4430 -200
rect 4520 -100 4660 -80
rect 4520 -200 4540 -100
rect 4640 -200 4660 -100
rect 4520 -220 4660 -200
rect 4750 -100 4890 -80
rect 4750 -200 4770 -100
rect 4870 -200 4890 -100
rect 4750 -220 4890 -200
rect 4980 -100 5120 -80
rect 4980 -200 5000 -100
rect 5100 -200 5120 -100
rect 4980 -220 5120 -200
rect 5210 -100 5350 -80
rect 5210 -200 5230 -100
rect 5330 -200 5350 -100
rect 5210 -220 5350 -200
rect 5440 -100 5580 -80
rect 5440 -200 5460 -100
rect 5560 -200 5580 -100
rect 5440 -220 5580 -200
rect 5670 -100 5810 -80
rect 5670 -200 5690 -100
rect 5790 -200 5810 -100
rect 5670 -220 5810 -200
rect 5900 -100 6040 -80
rect 5900 -200 5920 -100
rect 6020 -200 6040 -100
rect 5900 -220 6040 -200
rect 6130 -100 6270 -80
rect 6130 -200 6150 -100
rect 6250 -200 6270 -100
rect 6130 -220 6270 -200
rect 6360 -100 6500 -80
rect 6360 -200 6380 -100
rect 6480 -200 6500 -100
rect 6360 -220 6500 -200
rect 6590 -100 6730 -80
rect 6590 -200 6610 -100
rect 6710 -200 6730 -100
rect 6590 -220 6730 -200
rect 6820 -100 6960 -80
rect 6820 -200 6840 -100
rect 6940 -200 6960 -100
rect 6820 -220 6960 -200
rect 7900 -190 8350 630
rect -2100 -650 -1960 -450
rect -1760 -650 -1650 -450
rect -80 -400 60 -380
rect -80 -500 -60 -400
rect 40 -500 60 -400
rect -80 -520 60 -500
rect 150 -400 290 -380
rect 150 -500 170 -400
rect 270 -500 290 -400
rect 150 -520 290 -500
rect 380 -400 520 -380
rect 380 -500 400 -400
rect 500 -500 520 -400
rect 380 -520 520 -500
rect 610 -400 750 -380
rect 610 -500 630 -400
rect 730 -500 750 -400
rect 610 -520 750 -500
rect 840 -400 980 -380
rect 840 -500 860 -400
rect 960 -500 980 -400
rect 840 -520 980 -500
rect 1070 -400 1210 -380
rect 1070 -500 1090 -400
rect 1190 -500 1210 -400
rect 1070 -520 1210 -500
rect 1300 -400 1440 -380
rect 1300 -500 1320 -400
rect 1420 -500 1440 -400
rect 1300 -520 1440 -500
rect 1530 -400 1670 -380
rect 1530 -500 1550 -400
rect 1650 -500 1670 -400
rect 1530 -520 1670 -500
rect 1760 -400 1900 -380
rect 1760 -500 1780 -400
rect 1880 -500 1900 -400
rect 1760 -520 1900 -500
rect 1990 -400 2130 -380
rect 1990 -500 2010 -400
rect 2110 -500 2130 -400
rect 1990 -520 2130 -500
rect 2220 -400 2360 -380
rect 2220 -500 2240 -400
rect 2340 -500 2360 -400
rect 2220 -520 2360 -500
rect 2450 -400 2590 -380
rect 2450 -500 2470 -400
rect 2570 -500 2590 -400
rect 2450 -520 2590 -500
rect 2680 -400 2820 -380
rect 2680 -500 2700 -400
rect 2800 -500 2820 -400
rect 2680 -520 2820 -500
rect 2910 -400 3050 -380
rect 2910 -500 2930 -400
rect 3030 -500 3050 -400
rect 2910 -520 3050 -500
rect 3140 -400 3280 -380
rect 3140 -500 3160 -400
rect 3260 -500 3280 -400
rect 3140 -520 3280 -500
rect 3370 -400 3510 -380
rect 3370 -500 3390 -400
rect 3490 -500 3510 -400
rect 3370 -520 3510 -500
rect 3600 -400 3740 -380
rect 3600 -500 3620 -400
rect 3720 -500 3740 -400
rect 3600 -520 3740 -500
rect 3830 -400 3970 -380
rect 3830 -500 3850 -400
rect 3950 -500 3970 -400
rect 3830 -520 3970 -500
rect 4060 -400 4200 -380
rect 4060 -500 4080 -400
rect 4180 -500 4200 -400
rect 4060 -520 4200 -500
rect 4290 -400 4430 -380
rect 4290 -500 4310 -400
rect 4410 -500 4430 -400
rect 4290 -520 4430 -500
rect 4520 -400 4660 -380
rect 4520 -500 4540 -400
rect 4640 -500 4660 -400
rect 4520 -520 4660 -500
rect 4750 -400 4890 -380
rect 4750 -500 4770 -400
rect 4870 -500 4890 -400
rect 4750 -520 4890 -500
rect 4980 -400 5120 -380
rect 4980 -500 5000 -400
rect 5100 -500 5120 -400
rect 4980 -520 5120 -500
rect 5210 -400 5350 -380
rect 5210 -500 5230 -400
rect 5330 -500 5350 -400
rect 5210 -520 5350 -500
rect 5440 -400 5580 -380
rect 5440 -500 5460 -400
rect 5560 -500 5580 -400
rect 5440 -520 5580 -500
rect 5670 -400 5810 -380
rect 5670 -500 5690 -400
rect 5790 -500 5810 -400
rect 5670 -520 5810 -500
rect 5900 -400 6040 -380
rect 5900 -500 5920 -400
rect 6020 -500 6040 -400
rect 5900 -520 6040 -500
rect 6130 -400 6270 -380
rect 6130 -500 6150 -400
rect 6250 -500 6270 -400
rect 6130 -520 6270 -500
rect 6360 -400 6500 -380
rect 6360 -500 6380 -400
rect 6480 -500 6500 -400
rect 6360 -520 6500 -500
rect 6590 -400 6730 -380
rect 6590 -500 6610 -400
rect 6710 -500 6730 -400
rect 6590 -520 6730 -500
rect 6820 -400 6960 -380
rect 6820 -500 6840 -400
rect 6940 -500 6960 -400
rect 6820 -520 6960 -500
rect 7900 -390 8040 -190
rect 8240 -390 8350 -190
rect -2100 -1450 -1650 -650
rect 50 -590 160 -570
rect 50 -660 70 -590
rect 140 -660 160 -590
rect 50 -680 160 -660
rect 280 -590 390 -570
rect 280 -660 300 -590
rect 370 -660 390 -590
rect 280 -680 390 -660
rect 510 -590 620 -570
rect 510 -660 530 -590
rect 600 -660 620 -590
rect 510 -680 620 -660
rect 740 -590 850 -570
rect 740 -660 760 -590
rect 830 -660 850 -590
rect 740 -680 850 -660
rect 970 -590 1080 -570
rect 970 -660 990 -590
rect 1060 -660 1080 -590
rect 970 -680 1080 -660
rect 1200 -590 1310 -570
rect 1200 -660 1220 -590
rect 1290 -660 1310 -590
rect 1200 -680 1310 -660
rect 1430 -590 1540 -570
rect 1430 -660 1450 -590
rect 1520 -660 1540 -590
rect 1430 -680 1540 -660
rect 1660 -590 1770 -570
rect 1660 -660 1680 -590
rect 1750 -660 1770 -590
rect 1660 -680 1770 -660
rect 1890 -590 2000 -570
rect 1890 -660 1910 -590
rect 1980 -660 2000 -590
rect 1890 -680 2000 -660
rect 2120 -590 2230 -570
rect 2120 -660 2140 -590
rect 2210 -660 2230 -590
rect 2120 -680 2230 -660
rect 2350 -590 2460 -570
rect 2350 -660 2370 -590
rect 2440 -660 2460 -590
rect 2350 -680 2460 -660
rect 2580 -590 2690 -570
rect 2580 -660 2600 -590
rect 2670 -660 2690 -590
rect 2580 -680 2690 -660
rect 2810 -590 2920 -570
rect 2810 -660 2830 -590
rect 2900 -660 2920 -590
rect 2810 -680 2920 -660
rect 3040 -590 3150 -570
rect 3040 -660 3060 -590
rect 3130 -660 3150 -590
rect 3040 -680 3150 -660
rect 3270 -590 3380 -570
rect 3270 -660 3290 -590
rect 3360 -660 3380 -590
rect 3270 -680 3380 -660
rect 3500 -590 3610 -570
rect 3500 -660 3520 -590
rect 3590 -660 3610 -590
rect 3500 -680 3610 -660
rect 3730 -590 3840 -570
rect 3730 -660 3750 -590
rect 3820 -660 3840 -590
rect 3730 -680 3840 -660
rect 3960 -590 4070 -570
rect 3960 -660 3980 -590
rect 4050 -660 4070 -590
rect 3960 -680 4070 -660
rect 4190 -590 4300 -570
rect 4190 -660 4210 -590
rect 4280 -660 4300 -590
rect 4190 -680 4300 -660
rect 4420 -590 4530 -570
rect 4420 -660 4440 -590
rect 4510 -660 4530 -590
rect 4420 -680 4530 -660
rect 4650 -590 4760 -570
rect 4650 -660 4670 -590
rect 4740 -660 4760 -590
rect 4650 -680 4760 -660
rect 4880 -590 4990 -570
rect 4880 -660 4900 -590
rect 4970 -660 4990 -590
rect 4880 -680 4990 -660
rect 5110 -590 5220 -570
rect 5110 -660 5130 -590
rect 5200 -660 5220 -590
rect 5110 -680 5220 -660
rect 5340 -590 5450 -570
rect 5340 -660 5360 -590
rect 5430 -660 5450 -590
rect 5340 -680 5450 -660
rect 5570 -590 5680 -570
rect 5570 -660 5590 -590
rect 5660 -660 5680 -590
rect 5570 -680 5680 -660
rect 5800 -590 5910 -570
rect 5800 -660 5820 -590
rect 5890 -660 5910 -590
rect 5800 -680 5910 -660
rect 6030 -590 6140 -570
rect 6030 -660 6050 -590
rect 6120 -660 6140 -590
rect 6030 -680 6140 -660
rect 6260 -590 6370 -570
rect 6260 -660 6280 -590
rect 6350 -660 6370 -590
rect 6260 -680 6370 -660
rect 6490 -590 6600 -570
rect 6490 -660 6510 -590
rect 6580 -660 6600 -590
rect 6490 -680 6600 -660
rect 6720 -590 6830 -570
rect 6720 -660 6740 -590
rect 6810 -660 6830 -590
rect 6720 -680 6830 -660
rect 7050 -1100 7280 -1060
rect 2120 -1130 2260 -1110
rect 2120 -1230 2140 -1130
rect 2240 -1230 2260 -1130
rect 2120 -1250 2260 -1230
rect 2380 -1130 2520 -1110
rect 2380 -1230 2400 -1130
rect 2500 -1230 2520 -1130
rect 2380 -1250 2520 -1230
rect 2640 -1130 2780 -1110
rect 2640 -1230 2660 -1130
rect 2760 -1230 2780 -1130
rect 2640 -1250 2780 -1230
rect 2900 -1130 3040 -1110
rect 2900 -1230 2920 -1130
rect 3020 -1230 3040 -1130
rect 2900 -1250 3040 -1230
rect 3160 -1130 3300 -1110
rect 3160 -1230 3180 -1130
rect 3280 -1230 3300 -1130
rect 3160 -1250 3300 -1230
rect 3420 -1130 3560 -1110
rect 3420 -1230 3440 -1130
rect 3540 -1230 3560 -1130
rect 3420 -1250 3560 -1230
rect 3680 -1130 3820 -1110
rect 3680 -1230 3700 -1130
rect 3800 -1230 3820 -1130
rect 3680 -1250 3820 -1230
rect 3940 -1130 4080 -1110
rect 3940 -1230 3960 -1130
rect 4060 -1230 4080 -1130
rect 3940 -1250 4080 -1230
rect 4200 -1130 4340 -1110
rect 4200 -1230 4220 -1130
rect 4320 -1230 4340 -1130
rect 4200 -1250 4340 -1230
rect 4460 -1130 4600 -1110
rect 4460 -1230 4480 -1130
rect 4580 -1230 4600 -1130
rect 4460 -1250 4600 -1230
rect 4720 -1130 4860 -1110
rect 4720 -1230 4740 -1130
rect 4840 -1230 4860 -1130
rect 4720 -1250 4860 -1230
rect 4980 -1130 5120 -1110
rect 4980 -1230 5000 -1130
rect 5100 -1230 5120 -1130
rect 4980 -1250 5120 -1230
rect 5240 -1130 5380 -1110
rect 5240 -1230 5260 -1130
rect 5360 -1230 5380 -1130
rect 5240 -1250 5380 -1230
rect 5500 -1130 5640 -1110
rect 5500 -1230 5520 -1130
rect 5620 -1230 5640 -1130
rect 5500 -1250 5640 -1230
rect 5760 -1130 5900 -1110
rect 5760 -1230 5780 -1130
rect 5880 -1230 5900 -1130
rect 5760 -1250 5900 -1230
rect 6020 -1130 6160 -1110
rect 6020 -1230 6040 -1130
rect 6140 -1230 6160 -1130
rect 6020 -1250 6160 -1230
rect 6280 -1130 6420 -1110
rect 6280 -1230 6300 -1130
rect 6400 -1230 6420 -1130
rect 6280 -1250 6420 -1230
rect 6540 -1130 6680 -1110
rect 6540 -1230 6560 -1130
rect 6660 -1230 6680 -1130
rect 6540 -1250 6680 -1230
rect 6800 -1130 6940 -1110
rect 6800 -1230 6820 -1130
rect 6920 -1230 6940 -1130
rect 6800 -1250 6940 -1230
rect 7050 -1280 7090 -1100
rect 7250 -1280 7280 -1100
rect 7050 -1310 7280 -1280
rect -2100 -1650 -1960 -1450
rect -1760 -1650 -1650 -1450
rect 2120 -1470 2260 -1450
rect 2120 -1570 2140 -1470
rect 2240 -1570 2260 -1470
rect 2120 -1590 2260 -1570
rect 2380 -1470 2520 -1450
rect 2380 -1570 2400 -1470
rect 2500 -1570 2520 -1470
rect 2380 -1590 2520 -1570
rect 2640 -1470 2780 -1450
rect 2640 -1570 2660 -1470
rect 2760 -1570 2780 -1470
rect 2640 -1590 2780 -1570
rect 2900 -1470 3040 -1450
rect 2900 -1570 2920 -1470
rect 3020 -1570 3040 -1470
rect 2900 -1590 3040 -1570
rect 3160 -1470 3300 -1450
rect 3160 -1570 3180 -1470
rect 3280 -1570 3300 -1470
rect 3160 -1590 3300 -1570
rect 3420 -1470 3560 -1450
rect 3420 -1570 3440 -1470
rect 3540 -1570 3560 -1470
rect 3420 -1590 3560 -1570
rect 3680 -1470 3820 -1450
rect 3680 -1570 3700 -1470
rect 3800 -1570 3820 -1470
rect 3680 -1590 3820 -1570
rect 3940 -1470 4080 -1450
rect 3940 -1570 3960 -1470
rect 4060 -1570 4080 -1470
rect 3940 -1590 4080 -1570
rect 4200 -1470 4340 -1450
rect 4200 -1570 4220 -1470
rect 4320 -1570 4340 -1470
rect 4200 -1590 4340 -1570
rect 4460 -1470 4600 -1450
rect 4460 -1570 4480 -1470
rect 4580 -1570 4600 -1470
rect 4460 -1590 4600 -1570
rect 4720 -1470 4860 -1450
rect 4720 -1570 4740 -1470
rect 4840 -1570 4860 -1470
rect 4720 -1590 4860 -1570
rect 4980 -1470 5120 -1450
rect 4980 -1570 5000 -1470
rect 5100 -1570 5120 -1470
rect 4980 -1590 5120 -1570
rect 5240 -1470 5380 -1450
rect 5240 -1570 5260 -1470
rect 5360 -1570 5380 -1470
rect 5240 -1590 5380 -1570
rect 5500 -1470 5640 -1450
rect 5500 -1570 5520 -1470
rect 5620 -1570 5640 -1470
rect 5500 -1590 5640 -1570
rect 5760 -1470 5900 -1450
rect 5760 -1570 5780 -1470
rect 5880 -1570 5900 -1470
rect 5760 -1590 5900 -1570
rect 6020 -1470 6160 -1450
rect 6020 -1570 6040 -1470
rect 6140 -1570 6160 -1470
rect 6020 -1590 6160 -1570
rect 6280 -1470 6420 -1450
rect 6280 -1570 6300 -1470
rect 6400 -1570 6420 -1470
rect 6280 -1590 6420 -1570
rect 6540 -1470 6680 -1450
rect 6540 -1570 6560 -1470
rect 6660 -1570 6680 -1470
rect 6540 -1590 6680 -1570
rect 6800 -1470 6940 -1450
rect 6800 -1570 6820 -1470
rect 6920 -1570 6940 -1470
rect 6800 -1590 6940 -1570
rect -2100 -2090 -1650 -1650
rect 2260 -1700 2380 -1680
rect 2260 -1770 2280 -1700
rect 2360 -1770 2380 -1700
rect 2260 -1790 2380 -1770
rect 2520 -1700 2640 -1680
rect 2520 -1770 2540 -1700
rect 2620 -1770 2640 -1700
rect 2520 -1790 2640 -1770
rect 2780 -1700 2900 -1680
rect 2780 -1770 2800 -1700
rect 2880 -1770 2900 -1700
rect 2780 -1790 2900 -1770
rect 3040 -1700 3160 -1680
rect 3040 -1770 3060 -1700
rect 3140 -1770 3160 -1700
rect 3040 -1790 3160 -1770
rect 3300 -1700 3420 -1680
rect 3300 -1770 3320 -1700
rect 3400 -1770 3420 -1700
rect 3300 -1790 3420 -1770
rect 3560 -1700 3680 -1680
rect 3560 -1770 3580 -1700
rect 3660 -1770 3680 -1700
rect 3560 -1790 3680 -1770
rect 3820 -1700 3940 -1680
rect 3820 -1770 3840 -1700
rect 3920 -1770 3940 -1700
rect 3820 -1790 3940 -1770
rect 4080 -1700 4200 -1680
rect 4080 -1770 4100 -1700
rect 4180 -1770 4200 -1700
rect 4080 -1790 4200 -1770
rect 4340 -1700 4460 -1680
rect 4340 -1770 4360 -1700
rect 4440 -1770 4460 -1700
rect 4340 -1790 4460 -1770
rect 4600 -1700 4720 -1680
rect 4600 -1770 4620 -1700
rect 4700 -1770 4720 -1700
rect 4600 -1790 4720 -1770
rect 4860 -1700 4980 -1680
rect 4860 -1770 4880 -1700
rect 4960 -1770 4980 -1700
rect 4860 -1790 4980 -1770
rect 5120 -1700 5240 -1680
rect 5120 -1770 5140 -1700
rect 5220 -1770 5240 -1700
rect 5120 -1790 5240 -1770
rect 5380 -1700 5500 -1680
rect 5380 -1770 5400 -1700
rect 5480 -1770 5500 -1700
rect 5380 -1790 5500 -1770
rect 5640 -1700 5760 -1680
rect 5640 -1770 5660 -1700
rect 5740 -1770 5760 -1700
rect 5640 -1790 5760 -1770
rect 5900 -1700 6020 -1680
rect 5900 -1770 5920 -1700
rect 6000 -1770 6020 -1700
rect 5900 -1790 6020 -1770
rect 6160 -1700 6280 -1680
rect 6160 -1770 6180 -1700
rect 6260 -1770 6280 -1700
rect 6160 -1790 6280 -1770
rect 6420 -1700 6540 -1680
rect 6420 -1770 6440 -1700
rect 6520 -1770 6540 -1700
rect 6420 -1790 6540 -1770
rect 6680 -1700 6800 -1680
rect 6680 -1770 6700 -1700
rect 6780 -1770 6800 -1700
rect 6680 -1790 6800 -1770
rect 7900 -1920 8350 -390
rect 7900 -2090 8040 -1920
rect -2100 -2120 8040 -2090
rect 8240 -2120 8350 -1920
rect -2100 -2198 8350 -2120
rect -2100 -2200 -554 -2198
rect -352 -2200 8350 -2198
rect -2100 -2400 -1770 -2200
rect -1570 -2400 -554 -2200
rect -350 -2400 310 -2200
rect 510 -2400 1310 -2200
rect 1510 -2400 2330 -2200
rect 2530 -2400 3330 -2200
rect 3530 -2400 4330 -2200
rect 4530 -2400 5350 -2200
rect 5550 -2400 6350 -2200
rect 6550 -2400 7350 -2200
rect 7550 -2400 8350 -2200
rect -2100 -2540 8350 -2400
<< viali >>
rect 1540 1810 1620 1880
rect 1800 1810 1880 1880
rect 2330 1810 2410 1880
rect 2590 1810 2670 1880
rect 2850 1810 2930 1880
rect 3110 1810 3190 1880
rect 3370 1810 3450 1880
rect 3630 1810 3710 1880
rect 3890 1810 3970 1880
rect 4150 1810 4230 1880
rect 4410 1810 4490 1880
rect 4670 1810 4750 1880
rect 4930 1810 5010 1880
rect 5190 1810 5270 1880
rect 5450 1810 5530 1880
rect 5710 1810 5790 1880
rect 5970 1810 6050 1880
rect 6230 1810 6310 1880
rect 6490 1810 6570 1880
rect 6750 1810 6830 1880
rect 1400 1580 1500 1680
rect 1920 1580 2020 1680
rect 2190 1580 2290 1680
rect 2710 1580 2810 1680
rect 3230 1580 3330 1680
rect 3750 1580 3850 1680
rect 4270 1580 4370 1680
rect 4790 1580 4890 1680
rect 5310 1580 5410 1680
rect 5830 1580 5930 1680
rect 6350 1580 6450 1680
rect 6870 1580 6970 1680
rect 7130 1540 7290 1720
rect 1660 1300 1760 1400
rect 2450 1240 2550 1340
rect 2970 1240 3070 1340
rect 3490 1240 3590 1340
rect 4010 1240 4110 1340
rect 4530 1240 4630 1340
rect 5050 1240 5150 1340
rect 5570 1240 5670 1340
rect 6090 1240 6190 1340
rect 6610 1240 6710 1340
rect 70 700 140 770
rect 300 700 370 770
rect 530 700 600 770
rect 760 700 830 770
rect 990 700 1060 770
rect 1220 700 1290 770
rect 1450 700 1520 770
rect 1680 700 1750 770
rect 1910 700 1980 770
rect 2140 700 2210 770
rect 2370 700 2440 770
rect 2600 700 2670 770
rect 2830 700 2900 770
rect 3060 700 3130 770
rect 3290 700 3360 770
rect 3520 700 3590 770
rect 3750 700 3820 770
rect 3980 700 4050 770
rect 4210 700 4280 770
rect 4440 700 4510 770
rect 4670 700 4740 770
rect 4900 700 4970 770
rect 5130 700 5200 770
rect 5360 700 5430 770
rect 5590 700 5660 770
rect 5820 700 5890 770
rect 6050 700 6120 770
rect 6280 700 6350 770
rect 6510 700 6580 770
rect 6740 700 6810 770
rect -60 510 40 610
rect 400 510 500 610
rect 860 510 960 610
rect 1320 510 1420 610
rect 1780 510 1880 610
rect 2240 510 2340 610
rect 2700 510 2800 610
rect 3160 510 3260 610
rect 3620 510 3720 610
rect 4080 510 4180 610
rect 4540 510 4640 610
rect 5000 510 5100 610
rect 5460 510 5560 610
rect 5920 510 6020 610
rect 6380 510 6480 610
rect 6840 510 6940 610
rect 170 210 270 310
rect 630 210 730 310
rect 1090 210 1190 310
rect 1550 210 1650 310
rect 2010 210 2110 310
rect 2470 210 2570 310
rect 2930 210 3030 310
rect 3390 210 3490 310
rect 3850 210 3950 310
rect 4310 210 4410 310
rect 4770 210 4870 310
rect 5230 210 5330 310
rect 5690 210 5790 310
rect 6150 210 6250 310
rect 6610 210 6710 310
rect 1340 80 1470 90
rect 1340 30 1370 80
rect 1370 30 1450 80
rect 1450 30 1470 80
rect 1340 20 1470 30
rect 170 -200 270 -100
rect 630 -200 730 -100
rect 1090 -200 1190 -100
rect 1550 -200 1650 -100
rect 2010 -200 2110 -100
rect 2470 -200 2570 -100
rect 2930 -200 3030 -100
rect 3390 -200 3490 -100
rect 3850 -200 3950 -100
rect 4310 -200 4410 -100
rect 4770 -200 4870 -100
rect 5230 -200 5330 -100
rect 5690 -200 5790 -100
rect 6150 -200 6250 -100
rect 6610 -200 6710 -100
rect -60 -500 40 -400
rect 400 -500 500 -400
rect 860 -500 960 -400
rect 1320 -500 1420 -400
rect 1780 -500 1880 -400
rect 2240 -500 2340 -400
rect 2700 -500 2800 -400
rect 3160 -500 3260 -400
rect 3620 -500 3720 -400
rect 4080 -500 4180 -400
rect 4540 -500 4640 -400
rect 5000 -500 5100 -400
rect 5460 -500 5560 -400
rect 5920 -500 6020 -400
rect 6380 -500 6480 -400
rect 6840 -500 6940 -400
rect 70 -660 140 -590
rect 300 -660 370 -590
rect 530 -660 600 -590
rect 760 -660 830 -590
rect 990 -660 1060 -590
rect 1220 -660 1290 -590
rect 1450 -660 1520 -590
rect 1680 -660 1750 -590
rect 1910 -660 1980 -590
rect 2140 -660 2210 -590
rect 2370 -660 2440 -590
rect 2600 -660 2670 -590
rect 2830 -660 2900 -590
rect 3060 -660 3130 -590
rect 3290 -660 3360 -590
rect 3520 -660 3590 -590
rect 3750 -660 3820 -590
rect 3980 -660 4050 -590
rect 4210 -660 4280 -590
rect 4440 -660 4510 -590
rect 4670 -660 4740 -590
rect 4900 -660 4970 -590
rect 5130 -660 5200 -590
rect 5360 -660 5430 -590
rect 5590 -660 5660 -590
rect 5820 -660 5890 -590
rect 6050 -660 6120 -590
rect 6280 -660 6350 -590
rect 6510 -660 6580 -590
rect 6740 -660 6810 -590
rect 2140 -1230 2240 -1130
rect 2660 -1230 2760 -1130
rect 3180 -1230 3280 -1130
rect 3700 -1230 3800 -1130
rect 4220 -1230 4320 -1130
rect 4740 -1230 4840 -1130
rect 5260 -1230 5360 -1130
rect 5780 -1230 5880 -1130
rect 6300 -1230 6400 -1130
rect 6820 -1230 6920 -1130
rect 7090 -1280 7250 -1100
rect 2400 -1570 2500 -1470
rect 2920 -1570 3020 -1470
rect 3440 -1570 3540 -1470
rect 3960 -1570 4060 -1470
rect 4480 -1570 4580 -1470
rect 5000 -1570 5100 -1470
rect 5520 -1570 5620 -1470
rect 6040 -1570 6140 -1470
rect 6560 -1570 6660 -1470
rect 2280 -1770 2360 -1700
rect 2540 -1770 2620 -1700
rect 2800 -1770 2880 -1700
rect 3060 -1770 3140 -1700
rect 3320 -1770 3400 -1700
rect 3580 -1770 3660 -1700
rect 3840 -1770 3920 -1700
rect 4100 -1770 4180 -1700
rect 4360 -1770 4440 -1700
rect 4620 -1770 4700 -1700
rect 4880 -1770 4960 -1700
rect 5140 -1770 5220 -1700
rect 5400 -1770 5480 -1700
rect 5660 -1770 5740 -1700
rect 5920 -1770 6000 -1700
rect 6180 -1770 6260 -1700
rect 6440 -1770 6520 -1700
rect 6700 -1770 6780 -1700
rect -554 -2200 -352 -2198
rect -554 -2400 -550 -2200
rect -550 -2400 -352 -2200
<< metal1 >>
rect 1520 1880 1640 1900
rect 1520 1810 1540 1880
rect 1620 1810 1640 1880
rect 1520 1790 1640 1810
rect 1780 1880 1900 1900
rect 1780 1810 1800 1880
rect 1880 1810 1900 1880
rect 1780 1790 1900 1810
rect 2310 1880 2430 1900
rect 2310 1810 2330 1880
rect 2410 1810 2430 1880
rect 2310 1790 2430 1810
rect 2570 1880 2690 1900
rect 2570 1810 2590 1880
rect 2670 1810 2690 1880
rect 2570 1790 2690 1810
rect 2830 1880 2950 1900
rect 2830 1810 2850 1880
rect 2930 1810 2950 1880
rect 2830 1790 2950 1810
rect 3090 1880 3210 1900
rect 3090 1810 3110 1880
rect 3190 1810 3210 1880
rect 3090 1790 3210 1810
rect 3350 1880 3470 1900
rect 3350 1810 3370 1880
rect 3450 1810 3470 1880
rect 3350 1790 3470 1810
rect 3610 1880 3730 1900
rect 3610 1810 3630 1880
rect 3710 1810 3730 1880
rect 3610 1790 3730 1810
rect 3870 1880 3990 1900
rect 3870 1810 3890 1880
rect 3970 1810 3990 1880
rect 3870 1790 3990 1810
rect 4130 1880 4250 1900
rect 4130 1810 4150 1880
rect 4230 1810 4250 1880
rect 4130 1790 4250 1810
rect 4390 1880 4510 1900
rect 4390 1810 4410 1880
rect 4490 1810 4510 1880
rect 4390 1790 4510 1810
rect 4650 1880 4770 1900
rect 4650 1810 4670 1880
rect 4750 1810 4770 1880
rect 4650 1790 4770 1810
rect 4910 1880 5030 1900
rect 4910 1810 4930 1880
rect 5010 1810 5030 1880
rect 4910 1790 5030 1810
rect 5170 1880 5290 1900
rect 5170 1810 5190 1880
rect 5270 1810 5290 1880
rect 5170 1790 5290 1810
rect 5430 1880 5550 1900
rect 5430 1810 5450 1880
rect 5530 1810 5550 1880
rect 5430 1790 5550 1810
rect 5690 1880 5810 1900
rect 5690 1810 5710 1880
rect 5790 1810 5810 1880
rect 5690 1790 5810 1810
rect 5950 1880 6070 1900
rect 5950 1810 5970 1880
rect 6050 1810 6070 1880
rect 5950 1790 6070 1810
rect 6210 1880 6330 1900
rect 6210 1810 6230 1880
rect 6310 1810 6330 1880
rect 6210 1790 6330 1810
rect 6470 1880 6590 1900
rect 6470 1810 6490 1880
rect 6570 1810 6590 1880
rect 6470 1790 6590 1810
rect 6730 1880 6850 1900
rect 6730 1810 6750 1880
rect 6830 1810 6850 1880
rect 6730 1790 6850 1810
rect 7090 1720 7320 1760
rect 1380 1680 1520 1700
rect 1380 1580 1400 1680
rect 1500 1580 1520 1680
rect 1380 1560 1520 1580
rect 1900 1680 2040 1700
rect 1900 1580 1920 1680
rect 2020 1580 2040 1680
rect 1900 1560 2040 1580
rect 2170 1680 2310 1700
rect 2170 1580 2190 1680
rect 2290 1580 2310 1680
rect 2170 1560 2310 1580
rect 2690 1680 2830 1700
rect 2690 1580 2710 1680
rect 2810 1580 2830 1680
rect 2690 1560 2830 1580
rect 3210 1680 3350 1700
rect 3210 1580 3230 1680
rect 3330 1580 3350 1680
rect 3210 1560 3350 1580
rect 3730 1680 3870 1700
rect 3730 1580 3750 1680
rect 3850 1580 3870 1680
rect 3730 1560 3870 1580
rect 4250 1680 4390 1700
rect 4250 1580 4270 1680
rect 4370 1580 4390 1680
rect 4250 1560 4390 1580
rect 4770 1680 4910 1700
rect 4770 1580 4790 1680
rect 4890 1580 4910 1680
rect 4770 1560 4910 1580
rect 5290 1680 5430 1700
rect 5290 1580 5310 1680
rect 5410 1580 5430 1680
rect 5290 1560 5430 1580
rect 5810 1680 5950 1700
rect 5810 1580 5830 1680
rect 5930 1580 5950 1680
rect 5810 1560 5950 1580
rect 6330 1680 6470 1700
rect 6330 1580 6350 1680
rect 6450 1580 6470 1680
rect 6330 1560 6470 1580
rect 6850 1680 6990 1700
rect 6850 1580 6870 1680
rect 6970 1580 6990 1680
rect 6850 1560 6990 1580
rect 7090 1540 7130 1720
rect 7290 1540 7320 1720
rect 7090 1510 7320 1540
rect 1640 1400 1780 1420
rect 1640 1300 1660 1400
rect 1760 1300 1780 1400
rect 1640 1280 1780 1300
rect 2430 1340 2570 1360
rect 2430 1240 2450 1340
rect 2550 1240 2570 1340
rect 2430 1220 2570 1240
rect 2950 1340 3090 1360
rect 2950 1240 2970 1340
rect 3070 1240 3090 1340
rect 2950 1220 3090 1240
rect 3470 1340 3610 1360
rect 3470 1240 3490 1340
rect 3590 1240 3610 1340
rect 3470 1220 3610 1240
rect 3990 1340 4130 1360
rect 3990 1240 4010 1340
rect 4110 1240 4130 1340
rect 3990 1220 4130 1240
rect 4510 1340 4650 1360
rect 4510 1240 4530 1340
rect 4630 1240 4650 1340
rect 4510 1220 4650 1240
rect 5030 1340 5170 1360
rect 5030 1240 5050 1340
rect 5150 1240 5170 1340
rect 5030 1220 5170 1240
rect 5550 1340 5690 1360
rect 5550 1240 5570 1340
rect 5670 1240 5690 1340
rect 5550 1220 5690 1240
rect 6070 1340 6210 1360
rect 6070 1240 6090 1340
rect 6190 1240 6210 1340
rect 6070 1220 6210 1240
rect 6590 1340 6730 1360
rect 6590 1240 6610 1340
rect 6710 1240 6730 1340
rect 6590 1220 6730 1240
rect 50 770 160 790
rect 50 700 70 770
rect 140 700 160 770
rect 50 680 160 700
rect 280 770 390 790
rect 280 700 300 770
rect 370 700 390 770
rect 280 680 390 700
rect 510 770 620 790
rect 510 700 530 770
rect 600 700 620 770
rect 510 680 620 700
rect 740 770 850 790
rect 740 700 760 770
rect 830 700 850 770
rect 740 680 850 700
rect 970 770 1080 790
rect 970 700 990 770
rect 1060 700 1080 770
rect 970 680 1080 700
rect 1200 770 1310 790
rect 1200 700 1220 770
rect 1290 700 1310 770
rect 1200 680 1310 700
rect 1430 770 1540 790
rect 1430 700 1450 770
rect 1520 700 1540 770
rect 1430 680 1540 700
rect 1660 770 1770 790
rect 1660 700 1680 770
rect 1750 700 1770 770
rect 1660 680 1770 700
rect 1890 770 2000 790
rect 1890 700 1910 770
rect 1980 700 2000 770
rect 1890 680 2000 700
rect 2120 770 2230 790
rect 2120 700 2140 770
rect 2210 700 2230 770
rect 2120 680 2230 700
rect 2350 770 2460 790
rect 2350 700 2370 770
rect 2440 700 2460 770
rect 2350 680 2460 700
rect 2580 770 2690 790
rect 2580 700 2600 770
rect 2670 700 2690 770
rect 2580 680 2690 700
rect 2810 770 2920 790
rect 2810 700 2830 770
rect 2900 700 2920 770
rect 2810 680 2920 700
rect 3040 770 3150 790
rect 3040 700 3060 770
rect 3130 700 3150 770
rect 3040 680 3150 700
rect 3270 770 3380 790
rect 3270 700 3290 770
rect 3360 700 3380 770
rect 3270 680 3380 700
rect 3500 770 3610 790
rect 3500 700 3520 770
rect 3590 700 3610 770
rect 3500 680 3610 700
rect 3730 770 3840 790
rect 3730 700 3750 770
rect 3820 700 3840 770
rect 3730 680 3840 700
rect 3960 770 4070 790
rect 3960 700 3980 770
rect 4050 700 4070 770
rect 3960 680 4070 700
rect 4190 770 4300 790
rect 4190 700 4210 770
rect 4280 700 4300 770
rect 4190 680 4300 700
rect 4420 770 4530 790
rect 4420 700 4440 770
rect 4510 700 4530 770
rect 4420 680 4530 700
rect 4650 770 4760 790
rect 4650 700 4670 770
rect 4740 700 4760 770
rect 4650 680 4760 700
rect 4880 770 4990 790
rect 4880 700 4900 770
rect 4970 700 4990 770
rect 4880 680 4990 700
rect 5110 770 5220 790
rect 5110 700 5130 770
rect 5200 700 5220 770
rect 5110 680 5220 700
rect 5340 770 5450 790
rect 5340 700 5360 770
rect 5430 700 5450 770
rect 5340 680 5450 700
rect 5570 770 5680 790
rect 5570 700 5590 770
rect 5660 700 5680 770
rect 5570 680 5680 700
rect 5800 770 5910 790
rect 5800 700 5820 770
rect 5890 700 5910 770
rect 5800 680 5910 700
rect 6030 770 6140 790
rect 6030 700 6050 770
rect 6120 700 6140 770
rect 6030 680 6140 700
rect 6260 770 6370 790
rect 6260 700 6280 770
rect 6350 700 6370 770
rect 6260 680 6370 700
rect 6490 770 6600 790
rect 6490 700 6510 770
rect 6580 700 6600 770
rect 6490 680 6600 700
rect 6720 770 6830 790
rect 6720 700 6740 770
rect 6810 700 6830 770
rect 6720 680 6830 700
rect -80 610 60 630
rect -80 510 -60 610
rect 40 510 60 610
rect -80 490 60 510
rect 380 610 520 630
rect 380 510 400 610
rect 500 510 520 610
rect 380 490 520 510
rect 840 610 980 630
rect 840 510 860 610
rect 960 510 980 610
rect 840 490 980 510
rect 1300 610 1440 630
rect 1300 510 1320 610
rect 1420 510 1440 610
rect 1300 490 1440 510
rect 1760 610 1900 630
rect 1760 510 1780 610
rect 1880 510 1900 610
rect 1760 490 1900 510
rect 2220 610 2360 630
rect 2220 510 2240 610
rect 2340 510 2360 610
rect 2220 490 2360 510
rect 2680 610 2820 630
rect 2680 510 2700 610
rect 2800 510 2820 610
rect 2680 490 2820 510
rect 3140 610 3280 630
rect 3140 510 3160 610
rect 3260 510 3280 610
rect 3140 490 3280 510
rect 3600 610 3740 630
rect 3600 510 3620 610
rect 3720 510 3740 610
rect 3600 490 3740 510
rect 4060 610 4200 630
rect 4060 510 4080 610
rect 4180 510 4200 610
rect 4060 490 4200 510
rect 4520 610 4660 630
rect 4520 510 4540 610
rect 4640 510 4660 610
rect 4520 490 4660 510
rect 4980 610 5120 630
rect 4980 510 5000 610
rect 5100 510 5120 610
rect 4980 490 5120 510
rect 5440 610 5580 630
rect 5440 510 5460 610
rect 5560 510 5580 610
rect 5440 490 5580 510
rect 5900 610 6040 630
rect 5900 510 5920 610
rect 6020 510 6040 610
rect 5900 490 6040 510
rect 6360 610 6500 630
rect 6360 510 6380 610
rect 6480 510 6500 610
rect 6360 490 6500 510
rect 6820 610 6960 630
rect 6820 510 6840 610
rect 6940 510 6960 610
rect 6820 490 6960 510
rect 150 310 290 330
rect 150 210 170 310
rect 270 210 290 310
rect 150 190 290 210
rect 610 310 750 330
rect 610 210 630 310
rect 730 210 750 310
rect 610 190 750 210
rect 1070 310 1210 330
rect 1070 210 1090 310
rect 1190 210 1210 310
rect 1070 190 1210 210
rect 1530 310 1670 330
rect 1530 210 1550 310
rect 1650 210 1670 310
rect 1530 190 1670 210
rect 1990 310 2130 330
rect 1990 210 2010 310
rect 2110 210 2130 310
rect 1990 190 2130 210
rect 2450 310 2590 330
rect 2450 210 2470 310
rect 2570 210 2590 310
rect 2450 190 2590 210
rect 2910 310 3050 330
rect 2910 210 2930 310
rect 3030 210 3050 310
rect 2910 190 3050 210
rect 3370 310 3510 330
rect 3370 210 3390 310
rect 3490 210 3510 310
rect 3370 190 3510 210
rect 3830 310 3970 330
rect 3830 210 3850 310
rect 3950 210 3970 310
rect 3830 190 3970 210
rect 4290 310 4430 330
rect 4290 210 4310 310
rect 4410 210 4430 310
rect 4290 190 4430 210
rect 4750 310 4890 330
rect 4750 210 4770 310
rect 4870 210 4890 310
rect 4750 190 4890 210
rect 5210 310 5350 330
rect 5210 210 5230 310
rect 5330 210 5350 310
rect 5210 190 5350 210
rect 5670 310 5810 330
rect 5670 210 5690 310
rect 5790 210 5810 310
rect 5670 190 5810 210
rect 6130 310 6270 330
rect 6130 210 6150 310
rect 6250 210 6270 310
rect 6130 190 6270 210
rect 6590 310 6730 330
rect 6590 210 6610 310
rect 6710 210 6730 310
rect 6590 190 6730 210
rect 1320 90 1490 100
rect 1320 20 1340 90
rect 1470 20 1490 90
rect 1320 10 1490 20
rect 150 -100 290 -80
rect 150 -200 170 -100
rect 270 -200 290 -100
rect 150 -220 290 -200
rect 610 -100 750 -80
rect 610 -200 630 -100
rect 730 -200 750 -100
rect 610 -220 750 -200
rect 1070 -100 1210 -80
rect 1070 -200 1090 -100
rect 1190 -200 1210 -100
rect 1070 -220 1210 -200
rect 1530 -100 1670 -80
rect 1530 -200 1550 -100
rect 1650 -200 1670 -100
rect 1530 -220 1670 -200
rect 1990 -100 2130 -80
rect 1990 -200 2010 -100
rect 2110 -200 2130 -100
rect 1990 -220 2130 -200
rect 2450 -100 2590 -80
rect 2450 -200 2470 -100
rect 2570 -200 2590 -100
rect 2450 -220 2590 -200
rect 2910 -100 3050 -80
rect 2910 -200 2930 -100
rect 3030 -200 3050 -100
rect 2910 -220 3050 -200
rect 3370 -100 3510 -80
rect 3370 -200 3390 -100
rect 3490 -200 3510 -100
rect 3370 -220 3510 -200
rect 3830 -100 3970 -80
rect 3830 -200 3850 -100
rect 3950 -200 3970 -100
rect 3830 -220 3970 -200
rect 4290 -100 4430 -80
rect 4290 -200 4310 -100
rect 4410 -200 4430 -100
rect 4290 -220 4430 -200
rect 4750 -100 4890 -80
rect 4750 -200 4770 -100
rect 4870 -200 4890 -100
rect 4750 -220 4890 -200
rect 5210 -100 5350 -80
rect 5210 -200 5230 -100
rect 5330 -200 5350 -100
rect 5210 -220 5350 -200
rect 5670 -100 5810 -80
rect 5670 -200 5690 -100
rect 5790 -200 5810 -100
rect 5670 -220 5810 -200
rect 6130 -100 6270 -80
rect 6130 -200 6150 -100
rect 6250 -200 6270 -100
rect 6130 -220 6270 -200
rect 6590 -100 6730 -80
rect 6590 -200 6610 -100
rect 6710 -200 6730 -100
rect 6590 -220 6730 -200
rect -80 -400 60 -380
rect -80 -500 -60 -400
rect 40 -500 60 -400
rect -80 -520 60 -500
rect 380 -400 520 -380
rect 380 -500 400 -400
rect 500 -500 520 -400
rect 380 -520 520 -500
rect 840 -400 980 -380
rect 840 -500 860 -400
rect 960 -500 980 -400
rect 840 -520 980 -500
rect 1300 -400 1440 -380
rect 1300 -500 1320 -400
rect 1420 -500 1440 -400
rect 1300 -520 1440 -500
rect 1760 -400 1900 -380
rect 1760 -500 1780 -400
rect 1880 -500 1900 -400
rect 1760 -520 1900 -500
rect 2220 -400 2360 -380
rect 2220 -500 2240 -400
rect 2340 -500 2360 -400
rect 2220 -520 2360 -500
rect 2680 -400 2820 -380
rect 2680 -500 2700 -400
rect 2800 -500 2820 -400
rect 2680 -520 2820 -500
rect 3140 -400 3280 -380
rect 3140 -500 3160 -400
rect 3260 -500 3280 -400
rect 3140 -520 3280 -500
rect 3600 -400 3740 -380
rect 3600 -500 3620 -400
rect 3720 -500 3740 -400
rect 3600 -520 3740 -500
rect 4060 -400 4200 -380
rect 4060 -500 4080 -400
rect 4180 -500 4200 -400
rect 4060 -520 4200 -500
rect 4520 -400 4660 -380
rect 4520 -500 4540 -400
rect 4640 -500 4660 -400
rect 4520 -520 4660 -500
rect 4980 -400 5120 -380
rect 4980 -500 5000 -400
rect 5100 -500 5120 -400
rect 4980 -520 5120 -500
rect 5440 -400 5580 -380
rect 5440 -500 5460 -400
rect 5560 -500 5580 -400
rect 5440 -520 5580 -500
rect 5900 -400 6040 -380
rect 5900 -500 5920 -400
rect 6020 -500 6040 -400
rect 5900 -520 6040 -500
rect 6360 -400 6500 -380
rect 6360 -500 6380 -400
rect 6480 -500 6500 -400
rect 6360 -520 6500 -500
rect 6820 -400 6960 -380
rect 6820 -500 6840 -400
rect 6940 -500 6960 -400
rect 6820 -520 6960 -500
rect 50 -590 160 -570
rect 50 -660 70 -590
rect 140 -660 160 -590
rect 50 -680 160 -660
rect 280 -590 390 -570
rect 280 -660 300 -590
rect 370 -660 390 -590
rect 280 -680 390 -660
rect 510 -590 620 -570
rect 510 -660 530 -590
rect 600 -660 620 -590
rect 510 -680 620 -660
rect 740 -590 850 -570
rect 740 -660 760 -590
rect 830 -660 850 -590
rect 740 -680 850 -660
rect 970 -590 1080 -570
rect 970 -660 990 -590
rect 1060 -660 1080 -590
rect 970 -680 1080 -660
rect 1200 -590 1310 -570
rect 1200 -660 1220 -590
rect 1290 -660 1310 -590
rect 1200 -680 1310 -660
rect 1430 -590 1540 -570
rect 1430 -660 1450 -590
rect 1520 -660 1540 -590
rect 1430 -680 1540 -660
rect 1660 -590 1770 -570
rect 1660 -660 1680 -590
rect 1750 -660 1770 -590
rect 1660 -680 1770 -660
rect 1890 -590 2000 -570
rect 1890 -660 1910 -590
rect 1980 -660 2000 -590
rect 1890 -680 2000 -660
rect 2120 -590 2230 -570
rect 2120 -660 2140 -590
rect 2210 -660 2230 -590
rect 2120 -680 2230 -660
rect 2350 -590 2460 -570
rect 2350 -660 2370 -590
rect 2440 -660 2460 -590
rect 2350 -680 2460 -660
rect 2580 -590 2690 -570
rect 2580 -660 2600 -590
rect 2670 -660 2690 -590
rect 2580 -680 2690 -660
rect 2810 -590 2920 -570
rect 2810 -660 2830 -590
rect 2900 -660 2920 -590
rect 2810 -680 2920 -660
rect 3040 -590 3150 -570
rect 3040 -660 3060 -590
rect 3130 -660 3150 -590
rect 3040 -680 3150 -660
rect 3270 -590 3380 -570
rect 3270 -660 3290 -590
rect 3360 -660 3380 -590
rect 3270 -680 3380 -660
rect 3500 -590 3610 -570
rect 3500 -660 3520 -590
rect 3590 -660 3610 -590
rect 3500 -680 3610 -660
rect 3730 -590 3840 -570
rect 3730 -660 3750 -590
rect 3820 -660 3840 -590
rect 3730 -680 3840 -660
rect 3960 -590 4070 -570
rect 3960 -660 3980 -590
rect 4050 -660 4070 -590
rect 3960 -680 4070 -660
rect 4190 -590 4300 -570
rect 4190 -660 4210 -590
rect 4280 -660 4300 -590
rect 4190 -680 4300 -660
rect 4420 -590 4530 -570
rect 4420 -660 4440 -590
rect 4510 -660 4530 -590
rect 4420 -680 4530 -660
rect 4650 -590 4760 -570
rect 4650 -660 4670 -590
rect 4740 -660 4760 -590
rect 4650 -680 4760 -660
rect 4880 -590 4990 -570
rect 4880 -660 4900 -590
rect 4970 -660 4990 -590
rect 4880 -680 4990 -660
rect 5110 -590 5220 -570
rect 5110 -660 5130 -590
rect 5200 -660 5220 -590
rect 5110 -680 5220 -660
rect 5340 -590 5450 -570
rect 5340 -660 5360 -590
rect 5430 -660 5450 -590
rect 5340 -680 5450 -660
rect 5570 -590 5680 -570
rect 5570 -660 5590 -590
rect 5660 -660 5680 -590
rect 5570 -680 5680 -660
rect 5800 -590 5910 -570
rect 5800 -660 5820 -590
rect 5890 -660 5910 -590
rect 5800 -680 5910 -660
rect 6030 -590 6140 -570
rect 6030 -660 6050 -590
rect 6120 -660 6140 -590
rect 6030 -680 6140 -660
rect 6260 -590 6370 -570
rect 6260 -660 6280 -590
rect 6350 -660 6370 -590
rect 6260 -680 6370 -660
rect 6490 -590 6600 -570
rect 6490 -660 6510 -590
rect 6580 -660 6600 -590
rect 6490 -680 6600 -660
rect 6720 -590 6830 -570
rect 6720 -660 6740 -590
rect 6810 -660 6830 -590
rect 6720 -680 6830 -660
rect 7050 -1100 7280 -1060
rect 2120 -1130 2260 -1110
rect 2120 -1230 2140 -1130
rect 2240 -1230 2260 -1130
rect 2120 -1250 2260 -1230
rect 2640 -1130 2780 -1110
rect 2640 -1230 2660 -1130
rect 2760 -1230 2780 -1130
rect 2640 -1250 2780 -1230
rect 3160 -1130 3300 -1110
rect 3160 -1230 3180 -1130
rect 3280 -1230 3300 -1130
rect 3160 -1250 3300 -1230
rect 3680 -1130 3820 -1110
rect 3680 -1230 3700 -1130
rect 3800 -1230 3820 -1130
rect 3680 -1250 3820 -1230
rect 4200 -1130 4340 -1110
rect 4200 -1230 4220 -1130
rect 4320 -1230 4340 -1130
rect 4200 -1250 4340 -1230
rect 4720 -1130 4860 -1110
rect 4720 -1230 4740 -1130
rect 4840 -1230 4860 -1130
rect 4720 -1250 4860 -1230
rect 5240 -1130 5380 -1110
rect 5240 -1230 5260 -1130
rect 5360 -1230 5380 -1130
rect 5240 -1250 5380 -1230
rect 5760 -1130 5900 -1110
rect 5760 -1230 5780 -1130
rect 5880 -1230 5900 -1130
rect 5760 -1250 5900 -1230
rect 6280 -1130 6420 -1110
rect 6280 -1230 6300 -1130
rect 6400 -1230 6420 -1130
rect 6280 -1250 6420 -1230
rect 6800 -1130 6940 -1110
rect 6800 -1230 6820 -1130
rect 6920 -1230 6940 -1130
rect 6800 -1250 6940 -1230
rect 7050 -1280 7090 -1100
rect 7250 -1280 7280 -1100
rect 7050 -1310 7280 -1280
rect 2380 -1470 2520 -1450
rect 2380 -1570 2400 -1470
rect 2500 -1570 2520 -1470
rect 2380 -1590 2520 -1570
rect 2900 -1470 3040 -1450
rect 2900 -1570 2920 -1470
rect 3020 -1570 3040 -1470
rect 2900 -1590 3040 -1570
rect 3420 -1470 3560 -1450
rect 3420 -1570 3440 -1470
rect 3540 -1570 3560 -1470
rect 3420 -1590 3560 -1570
rect 3940 -1470 4080 -1450
rect 3940 -1570 3960 -1470
rect 4060 -1570 4080 -1470
rect 3940 -1590 4080 -1570
rect 4460 -1470 4600 -1450
rect 4460 -1570 4480 -1470
rect 4580 -1570 4600 -1470
rect 4460 -1590 4600 -1570
rect 4980 -1470 5120 -1450
rect 4980 -1570 5000 -1470
rect 5100 -1570 5120 -1470
rect 4980 -1590 5120 -1570
rect 5500 -1470 5640 -1450
rect 5500 -1570 5520 -1470
rect 5620 -1570 5640 -1470
rect 5500 -1590 5640 -1570
rect 6020 -1470 6160 -1450
rect 6020 -1570 6040 -1470
rect 6140 -1570 6160 -1470
rect 6020 -1590 6160 -1570
rect 6540 -1470 6680 -1450
rect 6540 -1570 6560 -1470
rect 6660 -1570 6680 -1470
rect 6540 -1590 6680 -1570
rect 2260 -1700 2380 -1680
rect 2260 -1770 2280 -1700
rect 2360 -1770 2380 -1700
rect 2260 -1790 2380 -1770
rect 2520 -1700 2640 -1680
rect 2520 -1770 2540 -1700
rect 2620 -1770 2640 -1700
rect 2520 -1790 2640 -1770
rect 2780 -1700 2900 -1680
rect 2780 -1770 2800 -1700
rect 2880 -1770 2900 -1700
rect 2780 -1790 2900 -1770
rect 3040 -1700 3160 -1680
rect 3040 -1770 3060 -1700
rect 3140 -1770 3160 -1700
rect 3040 -1790 3160 -1770
rect 3300 -1700 3420 -1680
rect 3300 -1770 3320 -1700
rect 3400 -1770 3420 -1700
rect 3300 -1790 3420 -1770
rect 3560 -1700 3680 -1680
rect 3560 -1770 3580 -1700
rect 3660 -1770 3680 -1700
rect 3560 -1790 3680 -1770
rect 3820 -1700 3940 -1680
rect 3820 -1770 3840 -1700
rect 3920 -1770 3940 -1700
rect 3820 -1790 3940 -1770
rect 4080 -1700 4200 -1680
rect 4080 -1770 4100 -1700
rect 4180 -1770 4200 -1700
rect 4080 -1790 4200 -1770
rect 4340 -1700 4460 -1680
rect 4340 -1770 4360 -1700
rect 4440 -1770 4460 -1700
rect 4340 -1790 4460 -1770
rect 4600 -1700 4720 -1680
rect 4600 -1770 4620 -1700
rect 4700 -1770 4720 -1700
rect 4600 -1790 4720 -1770
rect 4860 -1700 4980 -1680
rect 4860 -1770 4880 -1700
rect 4960 -1770 4980 -1700
rect 4860 -1790 4980 -1770
rect 5120 -1700 5240 -1680
rect 5120 -1770 5140 -1700
rect 5220 -1770 5240 -1700
rect 5120 -1790 5240 -1770
rect 5380 -1700 5500 -1680
rect 5380 -1770 5400 -1700
rect 5480 -1770 5500 -1700
rect 5380 -1790 5500 -1770
rect 5640 -1700 5760 -1680
rect 5640 -1770 5660 -1700
rect 5740 -1770 5760 -1700
rect 5640 -1790 5760 -1770
rect 5900 -1700 6020 -1680
rect 5900 -1770 5920 -1700
rect 6000 -1770 6020 -1700
rect 5900 -1790 6020 -1770
rect 6160 -1700 6280 -1680
rect 6160 -1770 6180 -1700
rect 6260 -1770 6280 -1700
rect 6160 -1790 6280 -1770
rect 6420 -1700 6540 -1680
rect 6420 -1770 6440 -1700
rect 6520 -1770 6540 -1700
rect 6420 -1790 6540 -1770
rect 6680 -1700 6800 -1680
rect 6680 -1770 6700 -1700
rect 6780 -1770 6800 -1700
rect 6680 -1790 6800 -1770
rect -584 -2198 -312 -2172
rect -584 -2400 -554 -2198
rect -352 -2400 -312 -2198
rect -584 -2430 -312 -2400
<< via1 >>
rect 1540 1810 1620 1880
rect 1800 1810 1880 1880
rect 2330 1810 2410 1880
rect 2590 1810 2670 1880
rect 2850 1810 2930 1880
rect 3110 1810 3190 1880
rect 3370 1810 3450 1880
rect 3630 1810 3710 1880
rect 3890 1810 3970 1880
rect 4150 1810 4230 1880
rect 4410 1810 4490 1880
rect 4670 1810 4750 1880
rect 4930 1810 5010 1880
rect 5190 1810 5270 1880
rect 5450 1810 5530 1880
rect 5710 1810 5790 1880
rect 5970 1810 6050 1880
rect 6230 1810 6310 1880
rect 6490 1810 6570 1880
rect 6750 1810 6830 1880
rect 1400 1580 1500 1680
rect 1920 1580 2020 1680
rect 2190 1580 2290 1680
rect 2710 1580 2810 1680
rect 3230 1580 3330 1680
rect 3750 1580 3850 1680
rect 4270 1580 4370 1680
rect 4790 1580 4890 1680
rect 5310 1580 5410 1680
rect 5830 1580 5930 1680
rect 6350 1580 6450 1680
rect 6870 1580 6970 1680
rect 7130 1540 7290 1720
rect 1660 1300 1760 1400
rect 2450 1240 2550 1340
rect 2970 1240 3070 1340
rect 3490 1240 3590 1340
rect 4010 1240 4110 1340
rect 4530 1240 4630 1340
rect 5050 1240 5150 1340
rect 5570 1240 5670 1340
rect 6090 1240 6190 1340
rect 6610 1240 6710 1340
rect 70 700 140 770
rect 300 700 370 770
rect 530 700 600 770
rect 760 700 830 770
rect 990 700 1060 770
rect 1220 700 1290 770
rect 1450 700 1520 770
rect 1680 700 1750 770
rect 1910 700 1980 770
rect 2140 700 2210 770
rect 2370 700 2440 770
rect 2600 700 2670 770
rect 2830 700 2900 770
rect 3060 700 3130 770
rect 3290 700 3360 770
rect 3520 700 3590 770
rect 3750 700 3820 770
rect 3980 700 4050 770
rect 4210 700 4280 770
rect 4440 700 4510 770
rect 4670 700 4740 770
rect 4900 700 4970 770
rect 5130 700 5200 770
rect 5360 700 5430 770
rect 5590 700 5660 770
rect 5820 700 5890 770
rect 6050 700 6120 770
rect 6280 700 6350 770
rect 6510 700 6580 770
rect 6740 700 6810 770
rect -60 510 40 610
rect 400 510 500 610
rect 860 510 960 610
rect 1320 510 1420 610
rect 1780 510 1880 610
rect 2240 510 2340 610
rect 2700 510 2800 610
rect 3160 510 3260 610
rect 3620 510 3720 610
rect 4080 510 4180 610
rect 4540 510 4640 610
rect 5000 510 5100 610
rect 5460 510 5560 610
rect 5920 510 6020 610
rect 6380 510 6480 610
rect 6840 510 6940 610
rect 170 210 270 310
rect 630 210 730 310
rect 1090 210 1190 310
rect 1550 210 1650 310
rect 2010 210 2110 310
rect 2470 210 2570 310
rect 2930 210 3030 310
rect 3390 210 3490 310
rect 3850 210 3950 310
rect 4310 210 4410 310
rect 4770 210 4870 310
rect 5230 210 5330 310
rect 5690 210 5790 310
rect 6150 210 6250 310
rect 6610 210 6710 310
rect 1340 20 1470 90
rect 170 -200 270 -100
rect 630 -200 730 -100
rect 1090 -200 1190 -100
rect 1550 -200 1650 -100
rect 2010 -200 2110 -100
rect 2470 -200 2570 -100
rect 2930 -200 3030 -100
rect 3390 -200 3490 -100
rect 3850 -200 3950 -100
rect 4310 -200 4410 -100
rect 4770 -200 4870 -100
rect 5230 -200 5330 -100
rect 5690 -200 5790 -100
rect 6150 -200 6250 -100
rect 6610 -200 6710 -100
rect -60 -500 40 -400
rect 400 -500 500 -400
rect 860 -500 960 -400
rect 1320 -500 1420 -400
rect 1780 -500 1880 -400
rect 2240 -500 2340 -400
rect 2700 -500 2800 -400
rect 3160 -500 3260 -400
rect 3620 -500 3720 -400
rect 4080 -500 4180 -400
rect 4540 -500 4640 -400
rect 5000 -500 5100 -400
rect 5460 -500 5560 -400
rect 5920 -500 6020 -400
rect 6380 -500 6480 -400
rect 6840 -500 6940 -400
rect 70 -660 140 -590
rect 300 -660 370 -590
rect 530 -660 600 -590
rect 760 -660 830 -590
rect 990 -660 1060 -590
rect 1220 -660 1290 -590
rect 1450 -660 1520 -590
rect 1680 -660 1750 -590
rect 1910 -660 1980 -590
rect 2140 -660 2210 -590
rect 2370 -660 2440 -590
rect 2600 -660 2670 -590
rect 2830 -660 2900 -590
rect 3060 -660 3130 -590
rect 3290 -660 3360 -590
rect 3520 -660 3590 -590
rect 3750 -660 3820 -590
rect 3980 -660 4050 -590
rect 4210 -660 4280 -590
rect 4440 -660 4510 -590
rect 4670 -660 4740 -590
rect 4900 -660 4970 -590
rect 5130 -660 5200 -590
rect 5360 -660 5430 -590
rect 5590 -660 5660 -590
rect 5820 -660 5890 -590
rect 6050 -660 6120 -590
rect 6280 -660 6350 -590
rect 6510 -660 6580 -590
rect 6740 -660 6810 -590
rect 2140 -1230 2240 -1130
rect 2660 -1230 2760 -1130
rect 3180 -1230 3280 -1130
rect 3700 -1230 3800 -1130
rect 4220 -1230 4320 -1130
rect 4740 -1230 4840 -1130
rect 5260 -1230 5360 -1130
rect 5780 -1230 5880 -1130
rect 6300 -1230 6400 -1130
rect 6820 -1230 6920 -1130
rect 7090 -1280 7250 -1100
rect 2400 -1570 2500 -1470
rect 2920 -1570 3020 -1470
rect 3440 -1570 3540 -1470
rect 3960 -1570 4060 -1470
rect 4480 -1570 4580 -1470
rect 5000 -1570 5100 -1470
rect 5520 -1570 5620 -1470
rect 6040 -1570 6140 -1470
rect 6560 -1570 6660 -1470
rect 2280 -1770 2360 -1700
rect 2540 -1770 2620 -1700
rect 2800 -1770 2880 -1700
rect 3060 -1770 3140 -1700
rect 3320 -1770 3400 -1700
rect 3580 -1770 3660 -1700
rect 3840 -1770 3920 -1700
rect 4100 -1770 4180 -1700
rect 4360 -1770 4440 -1700
rect 4620 -1770 4700 -1700
rect 4880 -1770 4960 -1700
rect 5140 -1770 5220 -1700
rect 5400 -1770 5480 -1700
rect 5660 -1770 5740 -1700
rect 5920 -1770 6000 -1700
rect 6180 -1770 6260 -1700
rect 6440 -1770 6520 -1700
rect 6700 -1770 6780 -1700
rect -554 -2400 -352 -2198
<< metal2 >>
rect 2010 1920 2200 1950
rect 1520 1880 1900 1900
rect 2010 1880 2040 1920
rect 1400 1810 1540 1880
rect 1620 1810 1660 1880
rect 1760 1810 1800 1880
rect 1880 1810 2040 1880
rect 1520 1790 1900 1810
rect 2010 1800 2040 1810
rect 2170 1880 2200 1920
rect 2310 1880 2430 1900
rect 2570 1880 2690 1900
rect 2830 1880 2950 1900
rect 3090 1880 3210 1900
rect 3350 1880 3470 1900
rect 3610 1880 3730 1900
rect 3870 1880 3990 1900
rect 4130 1880 4250 1900
rect 4390 1880 4510 1900
rect 4650 1880 4770 1900
rect 4910 1880 5030 1900
rect 5170 1880 5290 1900
rect 5430 1880 5550 1900
rect 5690 1880 5810 1900
rect 5950 1880 6070 1900
rect 6210 1880 6330 1900
rect 6470 1880 6590 1900
rect 6730 1880 6850 1900
rect 2170 1810 2330 1880
rect 2410 1810 2590 1880
rect 2670 1810 2850 1880
rect 2930 1810 3110 1880
rect 3190 1810 3370 1880
rect 3450 1810 3630 1880
rect 3710 1810 3890 1880
rect 3970 1810 4150 1880
rect 4230 1810 4410 1880
rect 4490 1810 4670 1880
rect 4750 1810 4930 1880
rect 5010 1810 5190 1880
rect 5270 1810 5450 1880
rect 5530 1810 5710 1880
rect 5790 1810 5970 1880
rect 6050 1810 6230 1880
rect 6310 1810 6490 1880
rect 6570 1810 6750 1880
rect 6830 1810 6850 1880
rect 2170 1800 2200 1810
rect 2010 1770 2200 1800
rect 2310 1790 2430 1810
rect 2570 1790 2690 1810
rect 2830 1790 2950 1810
rect 3090 1790 3210 1810
rect 3350 1790 3470 1810
rect 3610 1790 3730 1810
rect 3870 1790 3990 1810
rect 4130 1790 4250 1810
rect 4390 1790 4510 1810
rect 4650 1790 4770 1810
rect 4910 1790 5030 1810
rect 5170 1790 5290 1810
rect 5430 1790 5550 1810
rect 5690 1790 5810 1810
rect 5950 1790 6070 1810
rect 6210 1790 6330 1810
rect 6470 1790 6590 1810
rect 6730 1790 6850 1810
rect 7090 1720 7320 1760
rect 1380 1680 1520 1700
rect 1900 1680 2040 1700
rect 2170 1680 2310 1700
rect 2690 1680 2830 1700
rect 3210 1680 3350 1700
rect 3730 1680 3870 1700
rect 4250 1680 4390 1700
rect 4770 1680 4910 1700
rect 5290 1680 5430 1700
rect 5810 1680 5950 1700
rect 6330 1680 6470 1700
rect 6850 1680 6990 1700
rect 7090 1680 7130 1720
rect 1350 1580 1400 1680
rect 1500 1580 1920 1680
rect 2020 1580 2190 1680
rect 2290 1580 2710 1680
rect 2810 1580 3230 1680
rect 3330 1580 3750 1680
rect 3850 1580 4270 1680
rect 4370 1580 4790 1680
rect 4890 1580 5310 1680
rect 5410 1580 5830 1680
rect 5930 1580 6350 1680
rect 6450 1580 6870 1680
rect 6970 1580 7130 1680
rect 1380 1560 1520 1580
rect 1900 1560 2040 1580
rect 2170 1560 2310 1580
rect 2690 1560 2830 1580
rect 3210 1560 3350 1580
rect 3730 1560 3870 1580
rect 4250 1560 4390 1580
rect 4770 1560 4910 1580
rect 5290 1560 5430 1580
rect 5810 1560 5950 1580
rect 6330 1560 6470 1580
rect 6850 1560 6990 1580
rect 7090 1540 7130 1580
rect 7290 1680 7320 1720
rect 7360 1700 7580 1730
rect 7360 1680 7410 1700
rect 7290 1580 7410 1680
rect 7540 1580 7580 1700
rect 7290 1540 7320 1580
rect 7360 1540 7580 1580
rect 7090 1510 7320 1540
rect 1640 1400 1780 1420
rect 1640 1300 1660 1400
rect 1760 1300 1780 1400
rect 1640 1280 1780 1300
rect 2430 1340 2570 1360
rect 2950 1340 3090 1360
rect 3470 1340 3610 1360
rect 3990 1340 4130 1360
rect 4510 1340 4650 1360
rect 5030 1340 5170 1360
rect 5550 1340 5690 1360
rect 6070 1340 6210 1360
rect 6590 1340 6730 1360
rect 7100 1340 7240 1360
rect 2430 1240 2450 1340
rect 2550 1240 2970 1340
rect 3070 1240 3490 1340
rect 3590 1240 4010 1340
rect 4110 1240 4530 1340
rect 4630 1240 5050 1340
rect 5150 1240 5570 1340
rect 5670 1240 6090 1340
rect 6190 1240 6610 1340
rect 6710 1250 7120 1340
rect 7220 1250 7240 1340
rect 6710 1240 7240 1250
rect 2430 1220 2570 1240
rect 2950 1220 3090 1240
rect 3470 1220 3610 1240
rect 3990 1220 4130 1240
rect 4510 1220 4650 1240
rect 5030 1220 5170 1240
rect 5550 1220 5690 1240
rect 6070 1220 6210 1240
rect 6590 1220 6730 1240
rect 7100 1230 7240 1240
rect 50 770 160 790
rect 280 770 390 790
rect 510 770 620 790
rect 740 770 850 790
rect 970 770 1080 790
rect 1200 770 1310 790
rect 50 700 70 770
rect 140 700 300 770
rect 370 700 530 770
rect 600 700 650 770
rect 710 700 760 770
rect 830 700 990 770
rect 1060 700 1220 770
rect 1290 700 1310 770
rect 50 680 160 700
rect 280 680 390 700
rect 510 680 620 700
rect 740 680 850 700
rect 970 680 1080 700
rect 1200 680 1310 700
rect 1430 770 1540 790
rect 1660 770 1770 790
rect 1890 770 2000 790
rect 2120 770 2230 790
rect 2350 770 2460 790
rect 2580 770 2690 790
rect 2810 780 3150 790
rect 2810 770 2940 780
rect 1430 700 1450 770
rect 1520 700 1680 770
rect 1750 700 1910 770
rect 1980 700 2140 770
rect 2210 700 2370 770
rect 2440 700 2600 770
rect 2670 700 2830 770
rect 2900 700 2940 770
rect 1430 680 1540 700
rect 1660 680 1770 700
rect 1890 680 2000 700
rect 2120 680 2230 700
rect 2350 680 2460 700
rect 2580 680 2690 700
rect 2810 690 2940 700
rect 3020 770 3150 780
rect 3270 770 3380 790
rect 3500 770 3610 790
rect 3730 770 3840 790
rect 3960 770 4070 790
rect 4190 780 4530 790
rect 4190 770 4320 780
rect 3020 700 3060 770
rect 3130 700 3290 770
rect 3360 700 3520 770
rect 3590 700 3750 770
rect 3820 700 3980 770
rect 4050 700 4210 770
rect 4280 700 4320 770
rect 3020 690 3150 700
rect 2810 680 3150 690
rect 3270 680 3380 700
rect 3500 680 3610 700
rect 3730 680 3840 700
rect 3960 680 4070 700
rect 4190 690 4320 700
rect 4400 770 4530 780
rect 4650 770 4760 790
rect 4880 770 4990 790
rect 5110 770 5220 790
rect 5340 770 5450 790
rect 5570 770 5680 790
rect 5800 770 5910 790
rect 6030 770 6140 790
rect 6260 770 6370 790
rect 6490 770 6600 790
rect 6720 770 6830 790
rect 4400 700 4440 770
rect 4510 700 4670 770
rect 4740 700 4900 770
rect 4970 700 5130 770
rect 5200 700 5360 770
rect 5430 700 5590 770
rect 5660 700 5820 770
rect 5890 700 6050 770
rect 6120 700 6280 770
rect 6350 700 6510 770
rect 6580 700 6740 770
rect 6810 700 6830 770
rect 4400 690 4530 700
rect 4190 680 4530 690
rect 4650 680 4760 700
rect 4880 680 4990 700
rect 5110 680 5220 700
rect 5340 680 5450 700
rect 5570 680 5680 700
rect 5800 680 5910 700
rect 6030 680 6140 700
rect 6260 680 6370 700
rect 6490 680 6600 700
rect 6720 680 6830 700
rect -80 610 60 630
rect -80 510 -60 610
rect 40 590 60 610
rect 380 610 520 630
rect 380 590 400 610
rect 40 530 400 590
rect 40 510 60 530
rect -80 490 60 510
rect 380 510 400 530
rect 500 590 520 610
rect 840 610 980 630
rect 840 590 860 610
rect 500 530 860 590
rect 500 510 520 530
rect 380 490 520 510
rect 840 510 860 530
rect 960 590 980 610
rect 1300 610 1440 630
rect 1300 590 1320 610
rect 960 530 1320 590
rect 960 510 980 530
rect 840 490 980 510
rect 1300 510 1320 530
rect 1420 590 1440 610
rect 1760 610 1900 630
rect 1760 590 1780 610
rect 1420 530 1780 590
rect 1420 510 1440 530
rect 1300 490 1440 510
rect 1760 510 1780 530
rect 1880 590 1900 610
rect 2220 610 2360 630
rect 2220 590 2240 610
rect 1880 530 2240 590
rect 1880 510 1900 530
rect 1760 490 1900 510
rect 2220 510 2240 530
rect 2340 590 2360 610
rect 2680 610 2820 630
rect 2680 590 2700 610
rect 2340 530 2700 590
rect 2340 510 2360 530
rect 2220 490 2360 510
rect 2680 510 2700 530
rect 2800 590 2820 610
rect 3140 610 3280 630
rect 3140 590 3160 610
rect 2800 530 3160 590
rect 2800 510 2820 530
rect 2680 490 2820 510
rect 3140 510 3160 530
rect 3260 590 3280 610
rect 3600 610 3740 630
rect 3600 590 3620 610
rect 3260 530 3620 590
rect 3260 510 3280 530
rect 3140 490 3280 510
rect 3600 510 3620 530
rect 3720 590 3740 610
rect 4060 610 4200 630
rect 4060 590 4080 610
rect 3720 530 4080 590
rect 3720 510 3740 530
rect 3600 490 3740 510
rect 4060 510 4080 530
rect 4180 590 4200 610
rect 4520 610 4660 630
rect 4520 590 4540 610
rect 4180 530 4540 590
rect 4180 510 4200 530
rect 4060 490 4200 510
rect 4520 510 4540 530
rect 4640 590 4660 610
rect 4980 610 5120 630
rect 4980 590 5000 610
rect 4640 530 5000 590
rect 4640 510 4660 530
rect 4520 490 4660 510
rect 4980 510 5000 530
rect 5100 590 5120 610
rect 5440 610 5580 630
rect 5440 590 5460 610
rect 5100 530 5460 590
rect 5100 510 5120 530
rect 4980 490 5120 510
rect 5440 510 5460 530
rect 5560 590 5580 610
rect 5900 610 6040 630
rect 5900 590 5920 610
rect 5560 530 5920 590
rect 5560 510 5580 530
rect 5440 490 5580 510
rect 5900 510 5920 530
rect 6020 590 6040 610
rect 6360 610 6500 630
rect 6360 590 6380 610
rect 6020 530 6380 590
rect 6020 510 6040 530
rect 5900 490 6040 510
rect 6360 510 6380 530
rect 6480 590 6500 610
rect 6820 610 6960 630
rect 6820 590 6840 610
rect 6480 530 6840 590
rect 6480 510 6500 530
rect 6360 490 6500 510
rect 6820 510 6840 530
rect 6940 510 6960 610
rect 6820 490 6960 510
rect 150 310 290 330
rect 150 210 170 310
rect 270 290 290 310
rect 610 310 750 330
rect 610 290 630 310
rect 270 230 630 290
rect 270 210 290 230
rect 150 190 290 210
rect 610 210 630 230
rect 730 290 750 310
rect 1070 310 1210 330
rect 1070 290 1090 310
rect 730 230 1090 290
rect 730 210 750 230
rect 610 190 750 210
rect 1070 210 1090 230
rect 1190 210 1210 310
rect 1530 310 1670 330
rect 1530 290 1550 310
rect 1470 230 1550 290
rect 1070 190 1210 210
rect 1530 210 1550 230
rect 1650 290 1670 310
rect 1990 310 2130 330
rect 1990 290 2010 310
rect 1650 230 2010 290
rect 1650 210 1670 230
rect 1530 190 1670 210
rect 1990 210 2010 230
rect 2110 290 2130 310
rect 2450 310 2590 330
rect 2450 290 2470 310
rect 2110 230 2470 290
rect 2110 210 2130 230
rect 1990 190 2130 210
rect 2450 210 2470 230
rect 2570 290 2590 310
rect 2910 310 3050 330
rect 2910 290 2930 310
rect 2570 230 2930 290
rect 2570 210 2590 230
rect 2450 190 2590 210
rect 2910 210 2930 230
rect 3030 290 3050 310
rect 3370 310 3510 330
rect 3370 290 3390 310
rect 3030 230 3390 290
rect 3030 210 3050 230
rect 2910 190 3050 210
rect 3370 210 3390 230
rect 3490 290 3510 310
rect 3830 310 3970 330
rect 3830 290 3850 310
rect 3490 230 3850 290
rect 3490 210 3510 230
rect 3370 190 3510 210
rect 3830 210 3850 230
rect 3950 290 3970 310
rect 4290 310 4430 330
rect 4290 290 4310 310
rect 3950 230 4310 290
rect 3950 210 3970 230
rect 3830 190 3970 210
rect 4290 210 4310 230
rect 4410 290 4430 310
rect 4750 310 4890 330
rect 4750 290 4770 310
rect 4410 230 4770 290
rect 4410 210 4430 230
rect 4290 190 4430 210
rect 4750 210 4770 230
rect 4870 290 4890 310
rect 5210 310 5350 330
rect 5210 290 5230 310
rect 4870 230 5230 290
rect 4870 210 4890 230
rect 4750 190 4890 210
rect 5210 210 5230 230
rect 5330 290 5350 310
rect 5670 310 5810 330
rect 5670 290 5690 310
rect 5330 230 5690 290
rect 5330 210 5350 230
rect 5210 190 5350 210
rect 5670 210 5690 230
rect 5790 290 5810 310
rect 6130 310 6270 330
rect 6130 290 6150 310
rect 5790 230 6150 290
rect 5790 210 5810 230
rect 5670 190 5810 210
rect 6130 210 6150 230
rect 6250 290 6270 310
rect 6590 310 6730 330
rect 6590 290 6610 310
rect 6250 230 6610 290
rect 6250 210 6270 230
rect 6130 190 6270 210
rect 6590 210 6610 230
rect 6710 290 6730 310
rect 6710 230 6790 290
rect 6710 210 6730 230
rect 6590 190 6730 210
rect 1320 90 1490 100
rect 1320 20 1340 90
rect 1470 20 1490 90
rect 1320 10 1490 20
rect 150 -100 290 -80
rect 150 -200 170 -100
rect 270 -120 290 -100
rect 610 -100 750 -80
rect 610 -120 630 -100
rect 270 -180 630 -120
rect 270 -200 290 -180
rect 150 -220 290 -200
rect 610 -200 630 -180
rect 730 -120 750 -100
rect 1070 -100 1210 -80
rect 1070 -120 1090 -100
rect 730 -180 1090 -120
rect 730 -200 750 -180
rect 610 -220 750 -200
rect 1070 -200 1090 -180
rect 1190 -200 1210 -100
rect 1530 -100 1670 -80
rect 1530 -120 1550 -100
rect 1470 -180 1550 -120
rect 1070 -220 1210 -200
rect 1530 -200 1550 -180
rect 1650 -120 1670 -100
rect 1990 -100 2130 -80
rect 1990 -120 2010 -100
rect 1650 -180 2010 -120
rect 1650 -200 1670 -180
rect 1530 -220 1670 -200
rect 1990 -200 2010 -180
rect 2110 -120 2130 -100
rect 2450 -100 2590 -80
rect 2450 -120 2470 -100
rect 2110 -180 2470 -120
rect 2110 -200 2130 -180
rect 1990 -220 2130 -200
rect 2450 -200 2470 -180
rect 2570 -120 2590 -100
rect 2910 -100 3050 -80
rect 2910 -120 2930 -100
rect 2570 -180 2930 -120
rect 2570 -200 2590 -180
rect 2450 -220 2590 -200
rect 2910 -200 2930 -180
rect 3030 -120 3050 -100
rect 3370 -100 3510 -80
rect 3370 -120 3390 -100
rect 3030 -180 3390 -120
rect 3030 -200 3050 -180
rect 2910 -220 3050 -200
rect 3370 -200 3390 -180
rect 3490 -120 3510 -100
rect 3830 -100 3970 -80
rect 3830 -120 3850 -100
rect 3490 -180 3850 -120
rect 3490 -200 3510 -180
rect 3370 -220 3510 -200
rect 3830 -200 3850 -180
rect 3950 -120 3970 -100
rect 4290 -100 4430 -80
rect 4290 -120 4310 -100
rect 3950 -180 4310 -120
rect 3950 -200 3970 -180
rect 3830 -220 3970 -200
rect 4290 -200 4310 -180
rect 4410 -120 4430 -100
rect 4750 -100 4890 -80
rect 4750 -120 4770 -100
rect 4410 -180 4770 -120
rect 4410 -200 4430 -180
rect 4290 -220 4430 -200
rect 4750 -200 4770 -180
rect 4870 -120 4890 -100
rect 5210 -100 5350 -80
rect 5210 -120 5230 -100
rect 4870 -180 5230 -120
rect 4870 -200 4890 -180
rect 4750 -220 4890 -200
rect 5210 -200 5230 -180
rect 5330 -120 5350 -100
rect 5670 -100 5810 -80
rect 5670 -120 5690 -100
rect 5330 -180 5690 -120
rect 5330 -200 5350 -180
rect 5210 -220 5350 -200
rect 5670 -200 5690 -180
rect 5790 -120 5810 -100
rect 6130 -100 6270 -80
rect 6130 -120 6150 -100
rect 5790 -180 6150 -120
rect 5790 -200 5810 -180
rect 5670 -220 5810 -200
rect 6130 -200 6150 -180
rect 6250 -120 6270 -100
rect 6590 -100 6730 -80
rect 6590 -120 6610 -100
rect 6250 -180 6610 -120
rect 6250 -200 6270 -180
rect 6130 -220 6270 -200
rect 6590 -200 6610 -180
rect 6710 -120 6730 -100
rect 6710 -180 6790 -120
rect 6710 -200 6730 -180
rect 6590 -220 6730 -200
rect -80 -400 60 -380
rect -80 -500 -60 -400
rect 40 -420 60 -400
rect 380 -400 520 -380
rect 380 -420 400 -400
rect 40 -480 400 -420
rect 40 -500 60 -480
rect -80 -520 60 -500
rect 380 -500 400 -480
rect 500 -420 520 -400
rect 840 -400 980 -380
rect 840 -420 860 -400
rect 500 -480 860 -420
rect 500 -500 520 -480
rect 380 -520 520 -500
rect 840 -500 860 -480
rect 960 -420 980 -400
rect 1300 -400 1440 -380
rect 1300 -420 1320 -400
rect 960 -480 1320 -420
rect 960 -500 980 -480
rect 840 -520 980 -500
rect 1300 -500 1320 -480
rect 1420 -420 1440 -400
rect 1760 -400 1900 -380
rect 1760 -420 1780 -400
rect 1420 -480 1780 -420
rect 1420 -500 1440 -480
rect 1300 -520 1440 -500
rect 1760 -500 1780 -480
rect 1880 -420 1900 -400
rect 2220 -400 2360 -380
rect 2220 -420 2240 -400
rect 1880 -480 2240 -420
rect 1880 -500 1900 -480
rect 1760 -520 1900 -500
rect 2220 -500 2240 -480
rect 2340 -420 2360 -400
rect 2680 -400 2820 -380
rect 2680 -420 2700 -400
rect 2340 -480 2700 -420
rect 2340 -500 2360 -480
rect 2220 -520 2360 -500
rect 2680 -500 2700 -480
rect 2800 -420 2820 -400
rect 3140 -400 3280 -380
rect 3140 -420 3160 -400
rect 2800 -480 3160 -420
rect 2800 -500 2820 -480
rect 2680 -520 2820 -500
rect 3140 -500 3160 -480
rect 3260 -420 3280 -400
rect 3600 -400 3740 -380
rect 3600 -420 3620 -400
rect 3260 -480 3620 -420
rect 3260 -500 3280 -480
rect 3140 -520 3280 -500
rect 3600 -500 3620 -480
rect 3720 -420 3740 -400
rect 4060 -400 4200 -380
rect 4060 -420 4080 -400
rect 3720 -480 4080 -420
rect 3720 -500 3740 -480
rect 3600 -520 3740 -500
rect 4060 -500 4080 -480
rect 4180 -420 4200 -400
rect 4520 -400 4660 -380
rect 4520 -420 4540 -400
rect 4180 -480 4540 -420
rect 4180 -500 4200 -480
rect 4060 -520 4200 -500
rect 4520 -500 4540 -480
rect 4640 -420 4660 -400
rect 4980 -400 5120 -380
rect 4980 -420 5000 -400
rect 4640 -480 5000 -420
rect 4640 -500 4660 -480
rect 4520 -520 4660 -500
rect 4980 -500 5000 -480
rect 5100 -420 5120 -400
rect 5440 -400 5580 -380
rect 5440 -420 5460 -400
rect 5100 -480 5460 -420
rect 5100 -500 5120 -480
rect 4980 -520 5120 -500
rect 5440 -500 5460 -480
rect 5560 -420 5580 -400
rect 5900 -400 6040 -380
rect 5900 -420 5920 -400
rect 5560 -480 5920 -420
rect 5560 -500 5580 -480
rect 5440 -520 5580 -500
rect 5900 -500 5920 -480
rect 6020 -420 6040 -400
rect 6360 -400 6500 -380
rect 6360 -420 6380 -400
rect 6020 -480 6380 -420
rect 6020 -500 6040 -480
rect 5900 -520 6040 -500
rect 6360 -500 6380 -480
rect 6480 -420 6500 -400
rect 6820 -400 6960 -380
rect 6820 -420 6840 -400
rect 6480 -480 6840 -420
rect 6480 -500 6500 -480
rect 6360 -520 6500 -500
rect 6820 -500 6840 -480
rect 6940 -500 6960 -400
rect 6820 -520 6960 -500
rect 50 -590 160 -570
rect 280 -590 390 -570
rect 510 -590 620 -570
rect 740 -590 850 -570
rect 970 -590 1080 -570
rect 1200 -590 1310 -570
rect 50 -660 70 -590
rect 140 -660 300 -590
rect 370 -660 530 -590
rect 600 -660 650 -590
rect 710 -660 760 -590
rect 830 -660 990 -590
rect 1060 -660 1220 -590
rect 1290 -660 1310 -590
rect 50 -680 160 -660
rect 280 -680 390 -660
rect 510 -680 620 -660
rect 740 -680 850 -660
rect 970 -680 1080 -660
rect 1200 -680 1310 -660
rect 1430 -590 1540 -570
rect 1660 -590 1770 -570
rect 1890 -590 2000 -570
rect 2120 -590 2230 -570
rect 2350 -590 2460 -570
rect 2580 -590 2690 -570
rect 2810 -590 2920 -570
rect 3040 -590 3150 -570
rect 3270 -580 3610 -570
rect 3270 -590 3400 -580
rect 1430 -660 1450 -590
rect 1520 -660 1680 -590
rect 1750 -660 1910 -590
rect 1980 -660 2140 -590
rect 2210 -660 2370 -590
rect 2440 -660 2600 -590
rect 2670 -660 2830 -590
rect 2900 -660 3060 -590
rect 3130 -660 3290 -590
rect 3360 -660 3400 -590
rect 1430 -680 1540 -660
rect 1660 -680 1770 -660
rect 1890 -680 2000 -660
rect 2120 -680 2230 -660
rect 2350 -680 2460 -660
rect 2580 -680 2690 -660
rect 2810 -680 2920 -660
rect 3040 -680 3150 -660
rect 3270 -670 3400 -660
rect 3480 -590 3610 -580
rect 3730 -590 3840 -570
rect 3960 -590 4070 -570
rect 4190 -590 4300 -570
rect 4420 -590 4530 -570
rect 4650 -580 4990 -570
rect 4650 -590 4780 -580
rect 3480 -660 3520 -590
rect 3590 -660 3750 -590
rect 3820 -660 3980 -590
rect 4050 -660 4210 -590
rect 4280 -660 4440 -590
rect 4510 -660 4670 -590
rect 4740 -660 4780 -590
rect 3480 -670 3610 -660
rect 3270 -680 3610 -670
rect 3730 -680 3840 -660
rect 3960 -680 4070 -660
rect 4190 -680 4300 -660
rect 4420 -680 4530 -660
rect 4650 -670 4780 -660
rect 4860 -590 4990 -580
rect 5110 -590 5220 -570
rect 5340 -590 5450 -570
rect 5570 -590 5680 -570
rect 5800 -590 5910 -570
rect 6030 -590 6140 -570
rect 6260 -590 6370 -570
rect 6490 -590 6600 -570
rect 6720 -590 6830 -570
rect 4860 -660 4900 -590
rect 4970 -660 5130 -590
rect 5200 -660 5360 -590
rect 5430 -660 5590 -590
rect 5660 -660 5820 -590
rect 5890 -660 6050 -590
rect 6120 -660 6280 -590
rect 6350 -660 6510 -590
rect 6580 -660 6740 -590
rect 6810 -660 6830 -590
rect 4860 -670 4990 -660
rect 4650 -680 4990 -670
rect 5110 -680 5220 -660
rect 5340 -680 5450 -660
rect 5570 -680 5680 -660
rect 5800 -680 5910 -660
rect 6030 -680 6140 -660
rect 6260 -680 6370 -660
rect 6490 -680 6600 -660
rect 6720 -680 6830 -660
rect 7050 -1100 7280 -1060
rect 2120 -1130 2260 -1110
rect 2640 -1130 2780 -1110
rect 3160 -1130 3300 -1110
rect 3680 -1130 3820 -1110
rect 4200 -1130 4340 -1110
rect 4720 -1130 4860 -1110
rect 5240 -1130 5380 -1110
rect 5760 -1130 5900 -1110
rect 6280 -1130 6420 -1110
rect 6800 -1130 6940 -1110
rect 7050 -1130 7090 -1100
rect 2120 -1230 2140 -1130
rect 2240 -1230 2660 -1130
rect 2760 -1230 3180 -1130
rect 3280 -1230 3700 -1130
rect 3800 -1230 4220 -1130
rect 4320 -1230 4740 -1130
rect 4840 -1230 5260 -1130
rect 5360 -1230 5780 -1130
rect 5880 -1230 6300 -1130
rect 6400 -1230 6820 -1130
rect 6920 -1230 7090 -1130
rect 2120 -1250 2260 -1230
rect 2640 -1250 2780 -1230
rect 3160 -1250 3300 -1230
rect 3680 -1250 3820 -1230
rect 4200 -1250 4340 -1230
rect 4720 -1250 4860 -1230
rect 5240 -1250 5380 -1230
rect 5760 -1250 5900 -1230
rect 6280 -1250 6420 -1230
rect 6800 -1250 6940 -1230
rect 7050 -1280 7090 -1230
rect 7250 -1130 7280 -1100
rect 7370 -1100 7590 -1070
rect 7370 -1130 7420 -1100
rect 7250 -1220 7420 -1130
rect 7550 -1220 7590 -1100
rect 7250 -1230 7590 -1220
rect 7250 -1280 7280 -1230
rect 7370 -1260 7590 -1230
rect 7050 -1310 7280 -1280
rect 2380 -1470 2520 -1450
rect 2900 -1470 3040 -1450
rect 3420 -1470 3560 -1450
rect 3940 -1470 4080 -1450
rect 4460 -1470 4600 -1450
rect 4980 -1470 5120 -1450
rect 5500 -1470 5640 -1450
rect 6020 -1470 6160 -1450
rect 6540 -1470 6680 -1450
rect 7100 -1470 7240 -1450
rect 2380 -1570 2400 -1470
rect 2500 -1570 2920 -1470
rect 3020 -1570 3440 -1470
rect 3540 -1570 3960 -1470
rect 4060 -1570 4480 -1470
rect 4580 -1570 5000 -1470
rect 5100 -1570 5520 -1470
rect 5620 -1570 6040 -1470
rect 6140 -1570 6560 -1470
rect 6660 -1560 7120 -1470
rect 7220 -1560 7240 -1470
rect 6660 -1570 7240 -1560
rect 2380 -1590 2520 -1570
rect 2900 -1590 3040 -1570
rect 3420 -1590 3560 -1570
rect 3940 -1590 4080 -1570
rect 4460 -1590 4600 -1570
rect 4980 -1590 5120 -1570
rect 5500 -1590 5640 -1570
rect 6020 -1590 6160 -1570
rect 6540 -1590 6680 -1570
rect 7100 -1580 7240 -1570
rect 2000 -1680 2210 -1650
rect 2000 -1690 2380 -1680
rect 2000 -1800 2040 -1690
rect 2180 -1700 2380 -1690
rect 2520 -1700 2640 -1680
rect 2780 -1700 2900 -1680
rect 3040 -1700 3160 -1680
rect 3300 -1700 3420 -1680
rect 3560 -1700 3680 -1680
rect 3820 -1700 3940 -1680
rect 4080 -1700 4200 -1680
rect 4340 -1700 4460 -1680
rect 4600 -1700 4720 -1680
rect 4860 -1700 4980 -1680
rect 5120 -1700 5240 -1680
rect 5380 -1700 5500 -1680
rect 5640 -1700 5760 -1680
rect 5900 -1700 6020 -1680
rect 6160 -1700 6280 -1680
rect 6420 -1700 6540 -1680
rect 6680 -1700 6800 -1680
rect 2180 -1770 2280 -1700
rect 2360 -1770 2540 -1700
rect 2620 -1770 2800 -1700
rect 2880 -1770 3060 -1700
rect 3140 -1770 3320 -1700
rect 3400 -1770 3580 -1700
rect 3660 -1770 3840 -1700
rect 3920 -1770 4100 -1700
rect 4180 -1770 4360 -1700
rect 4440 -1770 4620 -1700
rect 4700 -1770 4880 -1700
rect 4960 -1770 5140 -1700
rect 5220 -1770 5400 -1700
rect 5480 -1770 5660 -1700
rect 5740 -1770 5920 -1700
rect 6000 -1770 6180 -1700
rect 6260 -1770 6440 -1700
rect 6520 -1770 6700 -1700
rect 6780 -1770 6800 -1700
rect 2180 -1790 2380 -1770
rect 2520 -1790 2640 -1770
rect 2780 -1790 2900 -1770
rect 3040 -1790 3160 -1770
rect 3300 -1790 3420 -1770
rect 3560 -1790 3680 -1770
rect 3820 -1790 3940 -1770
rect 4080 -1790 4200 -1770
rect 4340 -1790 4460 -1770
rect 4600 -1790 4720 -1770
rect 4860 -1790 4980 -1770
rect 5120 -1790 5240 -1770
rect 5380 -1790 5500 -1770
rect 5640 -1790 5760 -1770
rect 5900 -1790 6020 -1770
rect 6160 -1790 6280 -1770
rect 6420 -1790 6540 -1770
rect 6680 -1790 6800 -1770
rect 2180 -1800 2210 -1790
rect 2000 -1830 2210 -1800
rect -584 -2198 -312 -2172
rect -584 -2400 -554 -2198
rect -352 -2400 -312 -2198
rect -584 -2430 -312 -2400
<< via2 >>
rect 1660 1810 1760 1880
rect 2040 1800 2170 1920
rect 7410 1580 7540 1700
rect 1660 1300 1760 1400
rect 7120 1250 7220 1340
rect 650 700 710 770
rect 2940 690 3020 780
rect 4320 690 4400 780
rect -60 510 40 610
rect 170 210 270 310
rect 630 210 730 310
rect 1090 210 1190 310
rect 1550 210 1650 310
rect 3390 210 3490 310
rect 3850 210 3950 310
rect 4770 210 4870 310
rect 6610 210 6710 310
rect 1340 20 1470 90
rect 170 -200 270 -100
rect 630 -200 730 -100
rect 1090 -200 1190 -100
rect 1550 -200 1650 -100
rect 2930 -200 3030 -100
rect 3850 -200 3950 -100
rect 4310 -200 4410 -100
rect 6610 -200 6710 -100
rect -60 -500 40 -400
rect 650 -660 710 -590
rect 3400 -670 3480 -580
rect 4780 -670 4860 -580
rect 7420 -1220 7550 -1100
rect 7120 -1560 7220 -1470
rect 2040 -1800 2180 -1690
rect -554 -2400 -352 -2198
<< metal3 >>
rect 2000 1920 2210 1960
rect 1640 1880 1780 1900
rect 1640 1810 1660 1880
rect 1760 1810 1780 1880
rect 1640 1400 1780 1810
rect 1640 1300 1660 1400
rect 1760 1300 1780 1400
rect 1640 1220 1780 1300
rect 2000 1800 2040 1920
rect 2170 1800 2210 1920
rect 560 950 800 980
rect 560 870 590 950
rect 670 870 690 950
rect 770 870 800 950
rect 560 840 800 870
rect 1470 960 1710 990
rect 1470 880 1500 960
rect 1580 880 1600 960
rect 1680 880 1710 960
rect 1470 850 1710 880
rect 650 780 710 840
rect -1540 -400 -300 780
rect 640 770 720 780
rect 640 700 650 770
rect 710 700 720 770
rect 640 690 720 700
rect -80 610 60 630
rect -80 510 -60 610
rect 40 510 60 610
rect -80 490 60 510
rect 1560 330 1640 850
rect 150 310 290 330
rect 150 210 170 310
rect 270 210 290 310
rect 150 190 290 210
rect 610 310 750 330
rect 610 210 630 310
rect 730 210 750 310
rect 610 190 750 210
rect 1070 310 1210 330
rect 1070 210 1090 310
rect 1190 210 1210 310
rect 1070 190 1210 210
rect 1530 310 1670 330
rect 1530 210 1550 310
rect 1650 210 1670 310
rect 1530 190 1670 210
rect 190 110 250 190
rect 650 110 710 190
rect 1110 110 1170 190
rect 170 100 270 110
rect 170 10 180 100
rect 260 10 270 100
rect 170 0 270 10
rect 630 100 730 110
rect 630 10 640 100
rect 720 10 730 100
rect 630 0 730 10
rect 1090 100 1190 110
rect 1090 10 1100 100
rect 1180 10 1190 100
rect 1320 90 1490 100
rect 1320 20 1340 90
rect 1470 20 1490 90
rect 1320 10 1490 20
rect 1090 0 1190 10
rect 190 -80 250 0
rect 650 -80 710 0
rect 1110 -80 1170 0
rect 150 -100 290 -80
rect 150 -200 170 -100
rect 270 -200 290 -100
rect 150 -220 290 -200
rect 610 -100 750 -80
rect 610 -200 630 -100
rect 730 -200 750 -100
rect 610 -220 750 -200
rect 1070 -100 1210 -80
rect 1070 -200 1090 -100
rect 1190 -200 1210 -100
rect 1070 -220 1210 -200
rect 1530 -100 1670 -80
rect 1530 -200 1550 -100
rect 1650 -200 1670 -100
rect 1530 -220 1670 -200
rect -80 -400 60 -380
rect -1540 -500 -60 -400
rect 40 -500 60 -400
rect -1540 -1820 -300 -500
rect -80 -520 60 -500
rect 640 -590 720 -580
rect 640 -660 650 -590
rect 710 -660 720 -590
rect 640 -670 720 -660
rect 650 -730 710 -670
rect 560 -760 800 -730
rect 1560 -740 1640 -220
rect 560 -840 590 -760
rect 670 -840 690 -760
rect 770 -840 800 -760
rect 560 -870 800 -840
rect 1480 -770 1720 -740
rect 1480 -850 1510 -770
rect 1590 -850 1610 -770
rect 1690 -850 1720 -770
rect 1480 -880 1720 -850
rect 2000 -1690 2210 1800
rect 7140 1510 7280 1760
rect 7400 1730 7530 1740
rect 7360 1700 7580 1730
rect 7360 1580 7410 1700
rect 7540 1580 7580 1700
rect 7360 1540 7580 1580
rect 7100 1340 7240 1360
rect 7100 1250 7120 1340
rect 7220 1250 7240 1340
rect 3770 960 4010 990
rect 3770 880 3800 960
rect 3880 880 3900 960
rect 3980 880 4010 960
rect 3770 850 4010 880
rect 6530 960 6770 990
rect 6530 880 6560 960
rect 6640 880 6660 960
rect 6740 880 6770 960
rect 6530 850 6770 880
rect 2930 780 3030 790
rect 2930 690 2940 780
rect 3020 690 3030 780
rect 2930 -80 3030 690
rect 3860 330 3940 850
rect 4310 780 4410 790
rect 4310 690 4320 780
rect 4400 690 4410 780
rect 3370 310 3510 330
rect 3370 210 3390 310
rect 3490 210 3510 310
rect 3370 190 3510 210
rect 3830 310 3970 330
rect 3830 210 3850 310
rect 3950 210 3970 310
rect 3830 190 3970 210
rect 2910 -100 3050 -80
rect 2910 -200 2930 -100
rect 3030 -200 3050 -100
rect 2910 -220 3050 -200
rect 3390 -580 3490 190
rect 4310 -80 4410 690
rect 6620 330 6700 850
rect 4750 310 4890 330
rect 4750 210 4770 310
rect 4870 210 4890 310
rect 4750 190 4890 210
rect 6590 310 6730 330
rect 6590 210 6610 310
rect 6710 210 6730 310
rect 7100 320 7240 1250
rect 7100 230 7120 320
rect 7220 230 7240 320
rect 7100 210 7240 230
rect 6590 190 6730 210
rect 3830 -100 3970 -80
rect 3830 -200 3850 -100
rect 3950 -200 3970 -100
rect 3830 -220 3970 -200
rect 4290 -100 4430 -80
rect 4290 -200 4310 -100
rect 4410 -200 4430 -100
rect 4290 -220 4430 -200
rect 3390 -670 3400 -580
rect 3480 -670 3490 -580
rect 3390 -680 3490 -670
rect 3860 -740 3940 -220
rect 4770 -580 4870 190
rect 6590 -100 6730 -80
rect 6590 -200 6610 -100
rect 6710 -200 6730 -100
rect 6590 -220 6730 -200
rect 7100 -120 7240 -100
rect 7100 -210 7120 -120
rect 7220 -210 7240 -120
rect 4770 -670 4780 -580
rect 4860 -670 4870 -580
rect 4770 -680 4870 -670
rect 6620 -740 6700 -220
rect 3780 -770 4020 -740
rect 6540 -770 6780 -740
rect 3780 -850 3810 -770
rect 3890 -850 3910 -770
rect 3990 -840 6570 -770
rect 3990 -850 4020 -840
rect 3780 -880 4020 -850
rect 6540 -850 6570 -840
rect 6650 -850 6670 -770
rect 6750 -850 6780 -770
rect 6540 -880 6780 -850
rect 7100 -1470 7240 -210
rect 7400 -1070 7530 1540
rect 7370 -1100 7590 -1070
rect 7370 -1220 7420 -1100
rect 7550 -1220 7590 -1100
rect 7370 -1260 7590 -1220
rect 7400 -1280 7530 -1260
rect 7100 -1560 7120 -1470
rect 7220 -1560 7240 -1470
rect 7100 -1580 7240 -1560
rect 2000 -1800 2040 -1690
rect 2180 -1800 2210 -1690
rect 2000 -1830 2210 -1800
rect -584 -2198 -312 -2172
rect -584 -2400 -554 -2198
rect -352 -2400 -312 -2198
rect -584 -2430 -312 -2400
<< via3 >>
rect 590 870 670 950
rect 690 870 770 950
rect 1500 880 1580 960
rect 1600 880 1680 960
rect -60 510 40 610
rect 180 10 260 100
rect 640 10 720 100
rect 1100 10 1180 100
rect 1340 20 1470 90
rect 590 -840 670 -760
rect 690 -840 770 -760
rect 1510 -850 1590 -770
rect 1610 -850 1690 -770
rect 3800 880 3880 960
rect 3900 880 3980 960
rect 6560 880 6640 960
rect 6660 880 6740 960
rect 6610 210 6710 310
rect 7120 230 7220 320
rect 6610 -200 6710 -100
rect 7120 -210 7220 -120
rect 3810 -850 3890 -770
rect 3910 -850 3990 -770
rect 6570 -850 6650 -770
rect 6670 -850 6750 -770
rect -554 -2400 -352 -2198
<< mimcap >>
rect -1440 640 -398 680
rect -1440 -1680 -1400 640
rect -438 -1680 -398 640
rect -1440 -1720 -398 -1680
<< mimcapcontact >>
rect -1400 -1680 -438 640
<< metal4 >>
rect 560 950 800 980
rect 1470 960 1710 990
rect 1470 950 1500 960
rect 560 870 590 950
rect 670 870 690 950
rect 770 880 1500 950
rect 1580 880 1600 960
rect 1680 950 1710 960
rect 3770 960 4010 990
rect 3770 950 3800 960
rect 1680 880 3800 950
rect 3880 880 3900 960
rect 3980 950 4010 960
rect 6530 960 6770 990
rect 6530 950 6560 960
rect 3980 880 6560 950
rect 6640 880 6660 960
rect 6740 880 6770 960
rect 770 870 800 880
rect 560 840 800 870
rect 1470 850 1710 880
rect 3770 850 4010 880
rect 6530 850 6770 880
rect -1401 640 -437 641
rect -1401 -1680 -1400 640
rect -438 610 -437 640
rect -80 610 60 630
rect -438 510 -60 610
rect 40 510 60 610
rect -438 -1680 -437 510
rect -80 490 60 510
rect 6590 310 6730 330
rect 6590 210 6610 310
rect 6710 290 6730 310
rect 7100 320 7240 340
rect 7100 290 7120 320
rect 6710 230 7120 290
rect 7220 230 7240 320
rect 6710 210 6730 230
rect 7100 210 7240 230
rect 6590 190 6730 210
rect -1401 -1681 -437 -1680
rect -240 100 -50 102
rect 170 100 270 110
rect 630 100 730 110
rect 1090 100 1190 110
rect 1310 100 1500 120
rect -240 10 180 100
rect 260 10 640 100
rect 720 10 1100 100
rect 1180 90 1500 100
rect 1180 20 1340 90
rect 1470 20 1500 90
rect 1180 10 1500 20
rect -240 -600 -152 10
rect 170 0 270 10
rect 630 0 730 10
rect 1090 0 1190 10
rect 1310 -10 1500 10
rect 6590 -100 6730 -80
rect 6590 -200 6610 -100
rect 6710 -120 6730 -100
rect 7100 -120 7240 -100
rect 6710 -180 7120 -120
rect 6710 -200 6730 -180
rect 6590 -220 6730 -200
rect 7100 -210 7120 -180
rect 7220 -210 7240 -120
rect 7100 -230 7240 -210
rect -240 -2172 -148 -600
rect 560 -760 800 -730
rect 560 -840 590 -760
rect 670 -840 690 -760
rect 770 -770 800 -760
rect 1480 -770 1720 -740
rect 3780 -770 4020 -740
rect 6540 -770 6780 -740
rect 770 -840 1510 -770
rect 560 -870 800 -840
rect 1480 -850 1510 -840
rect 1590 -850 1610 -770
rect 1690 -840 3810 -770
rect 1690 -850 1720 -840
rect 1480 -880 1720 -850
rect 3780 -850 3810 -840
rect 3890 -850 3910 -770
rect 3990 -840 6570 -770
rect 3990 -850 4020 -840
rect 3780 -880 4020 -850
rect 6540 -850 6570 -840
rect 6650 -850 6670 -770
rect 6750 -850 6780 -770
rect 6540 -880 6780 -850
rect -584 -2198 -148 -2172
rect -584 -2400 -554 -2198
rect -352 -2254 -148 -2198
rect -352 -2400 -150 -2254
rect -584 -2430 -150 -2400
<< labels >>
rlabel via3 7170 260 7170 260 1 von
rlabel via3 7170 -160 7170 -160 1 vop
rlabel metal4 -330 560 -330 560 1 a
rlabel metal3 -340 -450 -340 -450 1 b
rlabel metal2 1460 1840 1460 1840 1 cm
rlabel via3 210 50 210 50 1 gnd!
rlabel metal3 7240 1630 7240 1630 1 vdd!
<< end >>
