magic
tech sky130A
timestamp 1647885906
<< locali >>
rect -1357 11918 -1166 11948
rect -1357 11807 -1330 11918
rect -1212 11807 -1166 11918
rect -1357 11681 -1166 11807
rect -1357 11655 1527 11681
rect -1357 11535 1376 11655
rect 1500 11535 1527 11655
rect -1357 11490 1527 11535
rect -1357 11481 -1166 11490
rect -12 3222 513 3263
rect -12 3100 1 3222
rect 118 3100 513 3222
rect -12 3082 513 3100
<< viali >>
rect -1330 11807 -1212 11918
rect 1376 11535 1500 11655
rect 1 3100 118 3222
<< metal1 >>
rect -1346 20113 -13 20126
rect -1346 20035 -109 20113
rect -34 20035 -13 20113
rect -1346 20026 -13 20035
rect -1346 18419 -1225 20026
rect -1346 12029 -1225 18283
rect -359 13707 -100 13710
rect -359 13696 -9 13707
rect -359 13599 -119 13696
rect -15 13599 -9 13696
rect -359 13590 -9 13599
rect -359 13581 -100 13590
rect -1348 11918 -1181 12029
rect -1348 11807 -1330 11918
rect -1212 11807 -1181 11918
rect -1348 11790 -1181 11807
rect -353 5828 -256 13581
rect 8180 11701 11053 11702
rect 8180 11697 13702 11701
rect 8180 11694 13725 11697
rect 2496 11693 13725 11694
rect 1347 11655 13725 11693
rect 1347 11535 1376 11655
rect 1500 11535 13725 11655
rect 1347 11513 13725 11535
rect 1347 11505 8206 11513
rect 10829 11512 13725 11513
rect 1347 11504 4220 11505
rect 13566 9837 13725 11512
rect -353 5808 -255 5828
rect -350 4402 -255 5808
rect -183 4402 829 4414
rect -350 4383 829 4402
rect -350 4303 712 4383
rect 800 4303 829 4383
rect -350 4276 829 4303
rect -350 4273 -88 4276
rect -12 3222 142 3249
rect -12 3100 1 3222
rect 118 3100 142 3222
rect -12 3082 142 3100
<< via1 >>
rect -109 20035 -34 20113
rect -119 13599 -15 13696
rect 712 4303 800 4383
rect 1 3100 118 3222
<< metal2 >>
rect -121 20113 35 20128
rect -121 20035 -109 20113
rect -34 20035 35 20113
rect -121 20026 35 20035
rect -227 18620 58 18641
rect -227 18515 -210 18620
rect -98 18515 58 18620
rect -227 18495 58 18515
rect -203 17142 35 17175
rect -203 17016 -170 17142
rect -32 17016 35 17142
rect -203 16983 35 17016
rect -338 15634 62 15684
rect -338 15525 -312 15634
rect -196 15525 62 15634
rect -338 15506 62 15525
rect -130 13696 -9 13707
rect -130 13599 -119 13696
rect -15 13599 -9 13696
rect -130 13590 -9 13599
rect -233 12250 -112 12265
rect -233 12155 -220 12250
rect -123 12155 -112 12250
rect -233 12144 -112 12155
rect -683 11821 -555 11848
rect -683 11738 -662 11821
rect -581 11738 -555 11821
rect -683 11716 -555 11738
rect -673 2806 -565 11716
rect -211 11497 -134 12144
rect -213 6196 -132 11497
rect -213 6096 740 6196
rect 694 4383 818 4403
rect 694 4303 712 4383
rect 800 4303 818 4383
rect 694 4283 818 4303
rect -12 3222 142 3249
rect -12 3100 1 3222
rect 118 3100 142 3222
rect -12 3082 142 3100
rect -673 2799 143 2806
rect -673 2603 582 2799
rect -512 2596 582 2603
<< via2 >>
rect -210 18515 -98 18620
rect -170 17016 -32 17142
rect -312 15525 -196 15634
rect -119 13599 -15 13696
rect -220 12155 -123 12250
rect -662 11738 -581 11821
rect 4248 5088 4335 5168
rect 1 3100 118 3222
<< metal3 >>
rect -1136 18620 -65 18640
rect -1136 18515 -210 18620
rect -98 18515 -65 18620
rect -1136 18499 -65 18515
rect -1123 18419 -1024 18499
rect -1123 4862 -1024 18283
rect -186 17162 -2 17167
rect -889 17142 -2 17162
rect -889 17016 -170 17142
rect -32 17016 -2 17142
rect -889 17015 -2 17016
rect -890 16999 -2 17015
rect -890 6634 -761 16999
rect -696 15634 -123 15677
rect -696 15525 -312 15634
rect -196 15525 -123 15634
rect -696 15490 -123 15525
rect -693 11821 -537 15490
rect -130 13696 -9 13707
rect -130 13599 -119 13696
rect -15 13599 -9 13696
rect -130 13590 -9 13599
rect -233 12250 -112 12265
rect -233 12155 -220 12250
rect -123 12155 -112 12250
rect -233 12144 -112 12155
rect -693 11738 -662 11821
rect -581 11738 -537 11821
rect -693 11717 -537 11738
rect -683 11716 -555 11717
rect -890 6500 4442 6634
rect 4240 5168 4350 5183
rect 4240 5088 4248 5168
rect 4335 5088 4350 5168
rect 4240 4950 4350 5088
rect -975 4863 924 4865
rect -975 4862 2420 4863
rect -1123 4857 2420 4862
rect 4234 4857 4353 4950
rect -1123 4791 4353 4857
rect -1123 4785 -875 4791
rect 521 4789 4353 4791
rect 4234 4787 4353 4789
rect -12 3222 142 3249
rect -12 3100 1 3222
rect 118 3100 142 3222
rect -12 3082 142 3100
<< via3 >>
rect -119 13599 -15 13696
rect -220 12155 -123 12250
rect 1 3100 118 3222
<< metal4 >>
rect -1620 19958 -1457 19967
rect -1620 19827 377 19958
rect -1620 18419 -1457 19827
rect 2125 19180 2333 19294
rect 2111 19019 2345 19180
rect -1620 18283 351 18419
rect -1620 16932 -1457 18283
rect 2128 17672 2336 17786
rect 2114 17511 2348 17672
rect -1620 16796 337 16932
rect -1620 15935 -1457 16796
rect 2128 16178 2336 16292
rect 2114 16017 2348 16178
rect -1629 15436 -1457 15935
rect -1629 15300 314 15436
rect -1629 14008 -1457 15300
rect 2126 14698 2334 14812
rect 2112 14379 2346 14698
rect -1629 13872 360 14008
rect -1629 12562 -1457 13872
rect -139 13696 32 13710
rect -139 13599 -119 13696
rect -15 13599 32 13696
rect -139 13578 32 13599
rect 2125 12915 2333 13361
rect -1629 12426 382 12562
rect -1629 3241 -1457 12426
rect -246 12250 20 12274
rect -246 12155 -220 12250
rect -123 12155 20 12250
rect -246 12131 20 12155
rect 822 11186 1055 11881
rect -12 3241 142 3249
rect -1629 3222 142 3241
rect -1629 3100 1 3222
rect 118 3100 142 3222
rect -1629 3083 142 3100
rect -12 3082 142 3083
<< metal5 >>
rect 194 19057 428 19203
rect 186 18859 431 19057
rect 197 17570 431 17695
rect 192 17372 437 17570
rect 197 16080 431 16201
rect 186 15882 431 16080
rect 195 14402 429 14721
rect 201 13035 421 13264
use tapered_buf  tapered_buf_5
timestamp 1647818295
transform 1 0 483 0 1 20036
box -470 -910 43675 401
use tapered_buf  tapered_buf_4
timestamp 1647818295
transform 1 0 486 0 1 18528
box -470 -910 43675 401
use tapered_buf  tapered_buf_3
timestamp 1647818295
transform 1 0 486 0 1 17034
box -470 -910 43675 401
use tapered_buf  tapered_buf_2
timestamp 1647818295
transform 1 0 484 0 1 15554
box -470 -910 43675 401
use tapered_buf  tapered_buf_1
timestamp 1647818295
transform 1 0 483 0 1 14103
box -470 -910 43675 401
use tapered_buf  tapered_buf_0
timestamp 1647818295
transform 1 0 482 0 1 12660
box -470 -910 43675 401
use pll_full  pll_full_0
timestamp 1647878380
transform 1 0 5793 0 1 555
box -5794 -555 13278 10840
<< labels >>
rlabel space 29 12701 29 12701 1 ref
rlabel space 51 14137 51 14137 1 mc2
rlabel space 56 15087 56 15087 1 div_out
rlabel space 61 16574 61 16574 1 down
rlabel space 38 18042 38 18042 1 upbar
rlabel space 61 19583 61 19583 1 vcont
rlabel metal4 -1568 12076 -1568 12076 1 gnd!
rlabel metal4 2225 13074 2225 13074 1 vdd!
<< end >>
