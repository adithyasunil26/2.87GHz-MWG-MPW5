magic
tech sky130A
magscale 1 2
timestamp 1647912062
<< psubdiff >>
rect 193788 665794 196518 666014
rect 193788 663430 194026 665794
rect 196274 663430 196518 665794
rect 193788 663224 196518 663430
rect 207718 665796 210448 666016
rect 207718 663432 207956 665796
rect 210204 663432 210448 665796
rect 207718 663226 210448 663432
rect 277154 665808 279884 666028
rect 277154 663444 277392 665808
rect 279640 663444 279884 665808
rect 277154 663238 279884 663444
rect 291084 665810 293814 666030
rect 291084 663446 291322 665810
rect 293570 663446 293814 665810
rect 291084 663240 293814 663446
rect 305000 665812 307730 666032
rect 305000 663448 305238 665812
rect 307486 663448 307730 665812
rect 305000 663242 307730 663448
rect 318834 665808 321564 666028
rect 318834 663444 319072 665808
rect 321320 663444 321564 665808
rect 318834 663238 321564 663444
rect 332764 665810 335494 666030
rect 332764 663446 333002 665810
rect 335250 663446 335494 665810
rect 332764 663240 335494 663446
rect 346680 665812 349410 666032
rect 346680 663448 346918 665812
rect 349166 663448 349410 665812
rect 346680 663242 349410 663448
rect 360290 665798 363020 666018
rect 360290 663434 360528 665798
rect 362776 663434 363020 665798
rect 360290 663228 363020 663434
rect 374220 665800 376950 666020
rect 374220 663436 374458 665800
rect 376706 663436 376950 665800
rect 374220 663230 376950 663436
rect 388136 665802 390866 666022
rect 388136 663438 388374 665802
rect 390622 663438 390866 665802
rect 388136 663232 390866 663438
rect 401976 665800 404706 666020
rect 401976 663436 402214 665800
rect 404462 663436 404706 665800
rect 401976 663230 404706 663436
rect 415906 665802 418636 666022
rect 415906 663438 416144 665802
rect 418392 663438 418636 665802
rect 415906 663232 418636 663438
rect 194336 653138 197066 653358
rect 194336 650774 194574 653138
rect 196822 650774 197066 653138
rect 194336 650568 197066 650774
rect 208266 653140 210996 653360
rect 208266 650776 208504 653140
rect 210752 650776 210996 653140
rect 208266 650570 210996 650776
rect 277702 653152 280432 653372
rect 277702 650788 277940 653152
rect 280188 650788 280432 653152
rect 277702 650582 280432 650788
rect 291632 653154 294362 653374
rect 291632 650790 291870 653154
rect 294118 650790 294362 653154
rect 291632 650584 294362 650790
rect 305548 653156 308278 653376
rect 305548 650792 305786 653156
rect 308034 650792 308278 653156
rect 305548 650586 308278 650792
rect 319382 653152 322112 653372
rect 319382 650788 319620 653152
rect 321868 650788 322112 653152
rect 319382 650582 322112 650788
rect 333312 653154 336042 653374
rect 333312 650790 333550 653154
rect 335798 650790 336042 653154
rect 333312 650584 336042 650790
rect 347228 653156 349958 653376
rect 347228 650792 347466 653156
rect 349714 650792 349958 653156
rect 347228 650586 349958 650792
rect 360838 653142 363568 653362
rect 360838 650778 361076 653142
rect 363324 650778 363568 653142
rect 360838 650572 363568 650778
rect 374768 653144 377498 653364
rect 374768 650780 375006 653144
rect 377254 650780 377498 653144
rect 374768 650574 377498 650780
rect 388684 653146 391414 653366
rect 388684 650782 388922 653146
rect 391170 650782 391414 653146
rect 388684 650576 391414 650782
rect 402524 653144 405254 653364
rect 402524 650780 402762 653144
rect 405010 650780 405254 653144
rect 402524 650574 405254 650780
rect 416454 653146 419184 653366
rect 416454 650782 416692 653146
rect 418940 650782 419184 653146
rect 416454 650576 419184 650782
rect 193788 638878 196518 639098
rect 193788 636514 194026 638878
rect 196274 636514 196518 638878
rect 193788 636308 196518 636514
rect 207718 638880 210448 639100
rect 207718 636516 207956 638880
rect 210204 636516 210448 638880
rect 207718 636310 210448 636516
rect 277154 638892 279884 639112
rect 277154 636528 277392 638892
rect 279640 636528 279884 638892
rect 277154 636322 279884 636528
rect 291084 638894 293814 639114
rect 291084 636530 291322 638894
rect 293570 636530 293814 638894
rect 291084 636324 293814 636530
rect 305000 638896 307730 639116
rect 305000 636532 305238 638896
rect 307486 636532 307730 638896
rect 305000 636326 307730 636532
rect 318834 638892 321564 639112
rect 318834 636528 319072 638892
rect 321320 636528 321564 638892
rect 318834 636322 321564 636528
rect 332764 638894 335494 639114
rect 332764 636530 333002 638894
rect 335250 636530 335494 638894
rect 332764 636324 335494 636530
rect 346680 638896 349410 639116
rect 346680 636532 346918 638896
rect 349166 636532 349410 638896
rect 346680 636326 349410 636532
rect 360290 638882 363020 639102
rect 360290 636518 360528 638882
rect 362776 636518 363020 638882
rect 360290 636312 363020 636518
rect 374220 638884 376950 639104
rect 374220 636520 374458 638884
rect 376706 636520 376950 638884
rect 374220 636314 376950 636520
rect 388136 638886 390866 639106
rect 388136 636522 388374 638886
rect 390622 636522 390866 638886
rect 388136 636316 390866 636522
rect 401976 638884 404706 639104
rect 401976 636520 402214 638884
rect 404462 636520 404706 638884
rect 401976 636314 404706 636520
rect 415906 638886 418636 639106
rect 415906 636522 416144 638886
rect 418392 636522 418636 638886
rect 415906 636316 418636 636522
rect 194348 624616 197078 624836
rect 194348 622252 194586 624616
rect 196834 622252 197078 624616
rect 194348 622046 197078 622252
rect 208278 624618 211008 624838
rect 208278 622254 208516 624618
rect 210764 622254 211008 624618
rect 208278 622048 211008 622254
rect 277714 624630 280444 624850
rect 277714 622266 277952 624630
rect 280200 622266 280444 624630
rect 277714 622060 280444 622266
rect 291644 624632 294374 624852
rect 291644 622268 291882 624632
rect 294130 622268 294374 624632
rect 291644 622062 294374 622268
rect 305560 624634 308290 624854
rect 305560 622270 305798 624634
rect 308046 622270 308290 624634
rect 305560 622064 308290 622270
rect 319394 624630 322124 624850
rect 319394 622266 319632 624630
rect 321880 622266 322124 624630
rect 319394 622060 322124 622266
rect 333324 624632 336054 624852
rect 333324 622268 333562 624632
rect 335810 622268 336054 624632
rect 333324 622062 336054 622268
rect 347240 624634 349970 624854
rect 347240 622270 347478 624634
rect 349726 622270 349970 624634
rect 347240 622064 349970 622270
rect 360850 624620 363580 624840
rect 360850 622256 361088 624620
rect 363336 622256 363580 624620
rect 360850 622050 363580 622256
rect 374780 624622 377510 624842
rect 374780 622258 375018 624622
rect 377266 622258 377510 624622
rect 374780 622052 377510 622258
rect 388696 624624 391426 624844
rect 388696 622260 388934 624624
rect 391182 622260 391426 624624
rect 388696 622054 391426 622260
rect 402536 624622 405266 624842
rect 402536 622258 402774 624622
rect 405022 622258 405266 624622
rect 402536 622052 405266 622258
rect 416466 624624 419196 624844
rect 416466 622260 416704 624624
rect 418952 622260 419196 624624
rect 416466 622054 419196 622260
rect 166248 610396 168978 610616
rect 166248 608032 166486 610396
rect 168734 608032 168978 610396
rect 166248 607826 168978 608032
rect 180164 610398 182894 610618
rect 180164 608034 180402 610398
rect 182650 608034 182894 610398
rect 180164 607828 182894 608034
rect 193800 610356 196530 610576
rect 193800 607992 194038 610356
rect 196286 607992 196530 610356
rect 193800 607786 196530 607992
rect 207730 610358 210460 610578
rect 207730 607994 207968 610358
rect 210216 607994 210460 610358
rect 207730 607788 210460 607994
rect 221646 610360 224376 610580
rect 221646 607996 221884 610360
rect 224132 607996 224376 610360
rect 221646 607790 224376 607996
rect 235486 610358 238216 610578
rect 235486 607994 235724 610358
rect 237972 607994 238216 610358
rect 235486 607788 238216 607994
rect 249416 610360 252146 610580
rect 249416 607996 249654 610360
rect 251902 607996 252146 610360
rect 249416 607790 252146 607996
rect 263332 610362 266062 610582
rect 263332 607998 263570 610362
rect 265818 607998 266062 610362
rect 263332 607792 266062 607998
rect 277166 610370 279896 610590
rect 277166 608006 277404 610370
rect 279652 608006 279896 610370
rect 277166 607800 279896 608006
rect 291096 610372 293826 610592
rect 291096 608008 291334 610372
rect 293582 608008 293826 610372
rect 291096 607802 293826 608008
rect 305012 610374 307742 610594
rect 305012 608010 305250 610374
rect 307498 608010 307742 610374
rect 305012 607804 307742 608010
rect 318846 610370 321576 610590
rect 318846 608006 319084 610370
rect 321332 608006 321576 610370
rect 318846 607800 321576 608006
rect 332776 610372 335506 610592
rect 332776 608008 333014 610372
rect 335262 608008 335506 610372
rect 332776 607802 335506 608008
rect 346692 610374 349422 610594
rect 346692 608010 346930 610374
rect 349178 608010 349422 610374
rect 346692 607804 349422 608010
rect 360302 610360 363032 610580
rect 360302 607996 360540 610360
rect 362788 607996 363032 610360
rect 360302 607790 363032 607996
rect 374232 610362 376962 610582
rect 374232 607998 374470 610362
rect 376718 607998 376962 610362
rect 374232 607792 376962 607998
rect 388148 610364 390878 610584
rect 388148 608000 388386 610364
rect 390634 608000 390878 610364
rect 388148 607794 390878 608000
rect 401988 610362 404718 610582
rect 401988 607998 402226 610362
rect 404474 607998 404718 610362
rect 401988 607792 404718 607998
rect 415918 610364 418648 610584
rect 415918 608000 416156 610364
rect 418404 608000 418648 610364
rect 415918 607794 418648 608000
rect 194526 591898 197256 592118
rect 194526 589534 194764 591898
rect 197012 589534 197256 591898
rect 194526 589328 197256 589534
rect 208456 591900 211186 592120
rect 208456 589536 208694 591900
rect 210942 589536 211186 591900
rect 208456 589330 211186 589536
rect 277892 591912 280622 592132
rect 277892 589548 278130 591912
rect 280378 589548 280622 591912
rect 277892 589342 280622 589548
rect 291822 591914 294552 592134
rect 291822 589550 292060 591914
rect 294308 589550 294552 591914
rect 291822 589344 294552 589550
rect 305738 591916 308468 592136
rect 305738 589552 305976 591916
rect 308224 589552 308468 591916
rect 305738 589346 308468 589552
rect 319572 591912 322302 592132
rect 319572 589548 319810 591912
rect 322058 589548 322302 591912
rect 319572 589342 322302 589548
rect 333502 591914 336232 592134
rect 333502 589550 333740 591914
rect 335988 589550 336232 591914
rect 333502 589344 336232 589550
rect 374958 591904 377688 592124
rect 374958 589540 375196 591904
rect 377444 589540 377688 591904
rect 374958 589334 377688 589540
rect 388874 591906 391604 592126
rect 388874 589542 389112 591906
rect 391360 589542 391604 591906
rect 388874 589336 391604 589542
rect 193978 577638 196708 577858
rect 193978 575274 194216 577638
rect 196464 575274 196708 577638
rect 193978 575068 196708 575274
rect 207908 577640 210638 577860
rect 207908 575276 208146 577640
rect 210394 575276 210638 577640
rect 207908 575070 210638 575276
rect 277344 577652 280074 577872
rect 277344 575288 277582 577652
rect 279830 575288 280074 577652
rect 277344 575082 280074 575288
rect 291274 577654 294004 577874
rect 291274 575290 291512 577654
rect 293760 575290 294004 577654
rect 291274 575084 294004 575290
rect 305190 577656 307920 577876
rect 305190 575292 305428 577656
rect 307676 575292 307920 577656
rect 305190 575086 307920 575292
rect 319024 577652 321754 577872
rect 319024 575288 319262 577652
rect 321510 575288 321754 577652
rect 319024 575082 321754 575288
rect 332954 577654 335684 577874
rect 332954 575290 333192 577654
rect 335440 575290 335684 577654
rect 332954 575084 335684 575290
rect 374410 577644 377140 577864
rect 374410 575280 374648 577644
rect 376896 575280 377140 577644
rect 374410 575074 377140 575280
rect 388326 577646 391056 577866
rect 388326 575282 388564 577646
rect 390812 575282 391056 577646
rect 388326 575076 391056 575282
rect 194194 564812 196924 565032
rect 194194 562448 194432 564812
rect 196680 562448 196924 564812
rect 194194 562242 196924 562448
rect 208124 564814 210854 565034
rect 208124 562450 208362 564814
rect 210610 562450 210854 564814
rect 208124 562244 210854 562450
rect 277560 564826 280290 565046
rect 277560 562462 277798 564826
rect 280046 562462 280290 564826
rect 277560 562256 280290 562462
rect 291490 564828 294220 565048
rect 291490 562464 291728 564828
rect 293976 562464 294220 564828
rect 291490 562258 294220 562464
rect 305406 564830 308136 565050
rect 305406 562466 305644 564830
rect 307892 562466 308136 564830
rect 305406 562260 308136 562466
rect 319240 564826 321970 565046
rect 319240 562462 319478 564826
rect 321726 562462 321970 564826
rect 319240 562256 321970 562462
rect 333170 564828 335900 565048
rect 333170 562464 333408 564828
rect 335656 562464 335900 564828
rect 333170 562258 335900 562464
rect 374626 564818 377356 565038
rect 374626 562454 374864 564818
rect 377112 562454 377356 564818
rect 374626 562248 377356 562454
rect 388542 564820 391272 565040
rect 388542 562456 388780 564820
rect 391028 562456 391272 564820
rect 388542 562250 391272 562456
rect 194628 547082 197358 547302
rect 194628 544718 194866 547082
rect 197114 544718 197358 547082
rect 194628 544512 197358 544718
rect 208558 547084 211288 547304
rect 208558 544720 208796 547084
rect 211044 544720 211288 547084
rect 208558 544514 211288 544720
rect 222474 547086 225204 547306
rect 222474 544722 222712 547086
rect 224960 544722 225204 547086
rect 222474 544516 225204 544722
rect 236314 547084 239044 547304
rect 236314 544720 236552 547084
rect 238800 544720 239044 547084
rect 236314 544514 239044 544720
rect 250244 547086 252974 547306
rect 250244 544722 250482 547086
rect 252730 544722 252974 547086
rect 250244 544516 252974 544722
rect 264160 547088 266890 547308
rect 264160 544724 264398 547088
rect 266646 544724 266890 547088
rect 264160 544518 266890 544724
rect 277994 547096 280724 547316
rect 277994 544732 278232 547096
rect 280480 544732 280724 547096
rect 277994 544526 280724 544732
rect 291924 547098 294654 547318
rect 291924 544734 292162 547098
rect 294410 544734 294654 547098
rect 291924 544528 294654 544734
rect 305840 547100 308570 547320
rect 305840 544736 306078 547100
rect 308326 544736 308570 547100
rect 305840 544530 308570 544736
rect 319674 547096 322404 547316
rect 319674 544732 319912 547096
rect 322160 544732 322404 547096
rect 319674 544526 322404 544732
rect 333604 547098 336334 547318
rect 333604 544734 333842 547098
rect 336090 544734 336334 547098
rect 333604 544528 336334 544734
rect 347520 547100 350250 547320
rect 347520 544736 347758 547100
rect 350006 544736 350250 547100
rect 347520 544530 350250 544736
rect 361130 547086 363860 547306
rect 361130 544722 361368 547086
rect 363616 544722 363860 547086
rect 361130 544516 363860 544722
rect 375060 547088 377790 547308
rect 375060 544724 375298 547088
rect 377546 544724 377790 547088
rect 375060 544518 377790 544724
rect 388976 547090 391706 547310
rect 388976 544726 389214 547090
rect 391462 544726 391706 547090
rect 388976 544520 391706 544726
rect 402816 547088 405546 547308
rect 402816 544724 403054 547088
rect 405302 544724 405546 547088
rect 402816 544518 405546 544724
rect 416746 547090 419476 547310
rect 416746 544726 416984 547090
rect 419232 544726 419476 547090
rect 416746 544520 419476 544726
rect 194080 532822 196810 533042
rect 194080 530458 194318 532822
rect 196566 530458 196810 532822
rect 194080 530252 196810 530458
rect 208010 532824 210740 533044
rect 208010 530460 208248 532824
rect 210496 530460 210740 532824
rect 208010 530254 210740 530460
rect 221926 532826 224656 533046
rect 221926 530462 222164 532826
rect 224412 530462 224656 532826
rect 221926 530256 224656 530462
rect 235766 532824 238496 533044
rect 235766 530460 236004 532824
rect 238252 530460 238496 532824
rect 235766 530254 238496 530460
rect 249696 532826 252426 533046
rect 249696 530462 249934 532826
rect 252182 530462 252426 532826
rect 249696 530256 252426 530462
rect 263612 532828 266342 533048
rect 263612 530464 263850 532828
rect 266098 530464 266342 532828
rect 263612 530258 266342 530464
rect 277446 532836 280176 533056
rect 277446 530472 277684 532836
rect 279932 530472 280176 532836
rect 277446 530266 280176 530472
rect 291376 532838 294106 533058
rect 291376 530474 291614 532838
rect 293862 530474 294106 532838
rect 291376 530268 294106 530474
rect 305292 532840 308022 533060
rect 305292 530476 305530 532840
rect 307778 530476 308022 532840
rect 305292 530270 308022 530476
rect 319126 532836 321856 533056
rect 319126 530472 319364 532836
rect 321612 530472 321856 532836
rect 319126 530266 321856 530472
rect 333056 532838 335786 533058
rect 333056 530474 333294 532838
rect 335542 530474 335786 532838
rect 333056 530268 335786 530474
rect 346972 532840 349702 533060
rect 346972 530476 347210 532840
rect 349458 530476 349702 532840
rect 346972 530270 349702 530476
rect 360582 532826 363312 533046
rect 360582 530462 360820 532826
rect 363068 530462 363312 532826
rect 360582 530256 363312 530462
rect 374512 532828 377242 533048
rect 374512 530464 374750 532828
rect 376998 530464 377242 532828
rect 374512 530258 377242 530464
rect 388428 532830 391158 533050
rect 388428 530466 388666 532830
rect 390914 530466 391158 532830
rect 388428 530260 391158 530466
rect 402268 532828 404998 533048
rect 402268 530464 402506 532828
rect 404754 530464 404998 532828
rect 402268 530258 404998 530464
rect 416198 532830 418928 533050
rect 416198 530466 416436 532830
rect 418684 530466 418928 532830
rect 416198 530260 418928 530466
rect 194296 519996 197026 520216
rect 194296 517632 194534 519996
rect 196782 517632 197026 519996
rect 194296 517426 197026 517632
rect 208226 519998 210956 520218
rect 208226 517634 208464 519998
rect 210712 517634 210956 519998
rect 208226 517428 210956 517634
rect 222142 520000 224872 520220
rect 222142 517636 222380 520000
rect 224628 517636 224872 520000
rect 222142 517430 224872 517636
rect 235982 519998 238712 520218
rect 235982 517634 236220 519998
rect 238468 517634 238712 519998
rect 235982 517428 238712 517634
rect 249912 520000 252642 520220
rect 249912 517636 250150 520000
rect 252398 517636 252642 520000
rect 249912 517430 252642 517636
rect 263828 520002 266558 520222
rect 263828 517638 264066 520002
rect 266314 517638 266558 520002
rect 263828 517432 266558 517638
rect 277662 520010 280392 520230
rect 277662 517646 277900 520010
rect 280148 517646 280392 520010
rect 277662 517440 280392 517646
rect 291592 520012 294322 520232
rect 291592 517648 291830 520012
rect 294078 517648 294322 520012
rect 291592 517442 294322 517648
rect 305508 520014 308238 520234
rect 305508 517650 305746 520014
rect 307994 517650 308238 520014
rect 305508 517444 308238 517650
rect 319342 520010 322072 520230
rect 319342 517646 319580 520010
rect 321828 517646 322072 520010
rect 319342 517440 322072 517646
rect 333272 520012 336002 520232
rect 333272 517648 333510 520012
rect 335758 517648 336002 520012
rect 333272 517442 336002 517648
rect 347188 520014 349918 520234
rect 347188 517650 347426 520014
rect 349674 517650 349918 520014
rect 347188 517444 349918 517650
rect 360798 520000 363528 520220
rect 360798 517636 361036 520000
rect 363284 517636 363528 520000
rect 360798 517430 363528 517636
rect 374728 520002 377458 520222
rect 374728 517638 374966 520002
rect 377214 517638 377458 520002
rect 374728 517432 377458 517638
rect 388644 520004 391374 520224
rect 388644 517640 388882 520004
rect 391130 517640 391374 520004
rect 388644 517434 391374 517640
rect 402484 520002 405214 520222
rect 402484 517638 402722 520002
rect 404970 517638 405214 520002
rect 402484 517432 405214 517638
rect 416414 520004 419144 520224
rect 416414 517640 416652 520004
rect 418900 517640 419144 520004
rect 416414 517434 419144 517640
rect 194690 498574 197420 498794
rect 194690 496210 194928 498574
rect 197176 496210 197420 498574
rect 194690 496004 197420 496210
rect 208620 498576 211350 498796
rect 208620 496212 208858 498576
rect 211106 496212 211350 498576
rect 208620 496006 211350 496212
rect 222536 498578 225266 498798
rect 222536 496214 222774 498578
rect 225022 496214 225266 498578
rect 222536 496008 225266 496214
rect 236376 498576 239106 498796
rect 236376 496212 236614 498576
rect 238862 496212 239106 498576
rect 236376 496006 239106 496212
rect 250306 498578 253036 498798
rect 250306 496214 250544 498578
rect 252792 496214 253036 498578
rect 250306 496008 253036 496214
rect 264222 498580 266952 498800
rect 264222 496216 264460 498580
rect 266708 496216 266952 498580
rect 264222 496010 266952 496216
rect 278056 498588 280786 498808
rect 278056 496224 278294 498588
rect 280542 496224 280786 498588
rect 278056 496018 280786 496224
rect 291986 498590 294716 498810
rect 291986 496226 292224 498590
rect 294472 496226 294716 498590
rect 291986 496020 294716 496226
rect 305902 498592 308632 498812
rect 305902 496228 306140 498592
rect 308388 496228 308632 498592
rect 305902 496022 308632 496228
rect 319736 498588 322466 498808
rect 319736 496224 319974 498588
rect 322222 496224 322466 498588
rect 319736 496018 322466 496224
rect 333666 498590 336396 498810
rect 333666 496226 333904 498590
rect 336152 496226 336396 498590
rect 333666 496020 336396 496226
rect 347582 498592 350312 498812
rect 347582 496228 347820 498592
rect 350068 496228 350312 498592
rect 347582 496022 350312 496228
rect 361192 498578 363922 498798
rect 361192 496214 361430 498578
rect 363678 496214 363922 498578
rect 361192 496008 363922 496214
rect 375122 498580 377852 498800
rect 375122 496216 375360 498580
rect 377608 496216 377852 498580
rect 375122 496010 377852 496216
rect 389038 498582 391768 498802
rect 389038 496218 389276 498582
rect 391524 496218 391768 498582
rect 389038 496012 391768 496218
rect 402878 498580 405608 498800
rect 402878 496216 403116 498580
rect 405364 496216 405608 498580
rect 402878 496010 405608 496216
rect 416808 498582 419538 498802
rect 416808 496218 417046 498582
rect 419294 496218 419538 498582
rect 416808 496012 419538 496218
rect 194142 484314 196872 484534
rect 194142 481950 194380 484314
rect 196628 481950 196872 484314
rect 194142 481744 196872 481950
rect 208072 484316 210802 484536
rect 208072 481952 208310 484316
rect 210558 481952 210802 484316
rect 208072 481746 210802 481952
rect 221988 484318 224718 484538
rect 221988 481954 222226 484318
rect 224474 481954 224718 484318
rect 221988 481748 224718 481954
rect 235828 484316 238558 484536
rect 235828 481952 236066 484316
rect 238314 481952 238558 484316
rect 235828 481746 238558 481952
rect 249758 484318 252488 484538
rect 249758 481954 249996 484318
rect 252244 481954 252488 484318
rect 249758 481748 252488 481954
rect 263674 484320 266404 484540
rect 263674 481956 263912 484320
rect 266160 481956 266404 484320
rect 263674 481750 266404 481956
rect 277508 484328 280238 484548
rect 277508 481964 277746 484328
rect 279994 481964 280238 484328
rect 277508 481758 280238 481964
rect 291438 484330 294168 484550
rect 291438 481966 291676 484330
rect 293924 481966 294168 484330
rect 291438 481760 294168 481966
rect 305354 484332 308084 484552
rect 305354 481968 305592 484332
rect 307840 481968 308084 484332
rect 305354 481762 308084 481968
rect 319188 484328 321918 484548
rect 319188 481964 319426 484328
rect 321674 481964 321918 484328
rect 319188 481758 321918 481964
rect 333118 484330 335848 484550
rect 333118 481966 333356 484330
rect 335604 481966 335848 484330
rect 333118 481760 335848 481966
rect 347034 484332 349764 484552
rect 347034 481968 347272 484332
rect 349520 481968 349764 484332
rect 347034 481762 349764 481968
rect 360644 484318 363374 484538
rect 360644 481954 360882 484318
rect 363130 481954 363374 484318
rect 360644 481748 363374 481954
rect 374574 484320 377304 484540
rect 374574 481956 374812 484320
rect 377060 481956 377304 484320
rect 374574 481750 377304 481956
rect 388490 484322 391220 484542
rect 388490 481958 388728 484322
rect 390976 481958 391220 484322
rect 388490 481752 391220 481958
rect 402330 484320 405060 484540
rect 402330 481956 402568 484320
rect 404816 481956 405060 484320
rect 402330 481750 405060 481956
rect 416260 484322 418990 484542
rect 416260 481958 416498 484322
rect 418746 481958 418990 484322
rect 416260 481752 418990 481958
rect 194358 471488 197088 471708
rect 194358 469124 194596 471488
rect 196844 469124 197088 471488
rect 194358 468918 197088 469124
rect 208288 471490 211018 471710
rect 208288 469126 208526 471490
rect 210774 469126 211018 471490
rect 208288 468920 211018 469126
rect 222204 471492 224934 471712
rect 222204 469128 222442 471492
rect 224690 469128 224934 471492
rect 222204 468922 224934 469128
rect 236044 471490 238774 471710
rect 236044 469126 236282 471490
rect 238530 469126 238774 471490
rect 236044 468920 238774 469126
rect 249974 471492 252704 471712
rect 249974 469128 250212 471492
rect 252460 469128 252704 471492
rect 249974 468922 252704 469128
rect 263890 471494 266620 471714
rect 263890 469130 264128 471494
rect 266376 469130 266620 471494
rect 263890 468924 266620 469130
rect 277724 471502 280454 471722
rect 277724 469138 277962 471502
rect 280210 469138 280454 471502
rect 277724 468932 280454 469138
rect 291654 471504 294384 471724
rect 291654 469140 291892 471504
rect 294140 469140 294384 471504
rect 291654 468934 294384 469140
rect 305570 471506 308300 471726
rect 305570 469142 305808 471506
rect 308056 469142 308300 471506
rect 305570 468936 308300 469142
rect 319404 471502 322134 471722
rect 319404 469138 319642 471502
rect 321890 469138 322134 471502
rect 319404 468932 322134 469138
rect 333334 471504 336064 471724
rect 333334 469140 333572 471504
rect 335820 469140 336064 471504
rect 333334 468934 336064 469140
rect 347250 471506 349980 471726
rect 347250 469142 347488 471506
rect 349736 469142 349980 471506
rect 347250 468936 349980 469142
rect 360860 471492 363590 471712
rect 360860 469128 361098 471492
rect 363346 469128 363590 471492
rect 360860 468922 363590 469128
rect 374790 471494 377520 471714
rect 374790 469130 375028 471494
rect 377276 469130 377520 471494
rect 374790 468924 377520 469130
rect 388706 471496 391436 471716
rect 388706 469132 388944 471496
rect 391192 469132 391436 471496
rect 388706 468926 391436 469132
rect 402546 471494 405276 471714
rect 402546 469130 402784 471494
rect 405032 469130 405276 471494
rect 402546 468924 405276 469130
rect 416476 471496 419206 471716
rect 416476 469132 416714 471496
rect 418962 469132 419206 471496
rect 416476 468926 419206 469132
rect 194938 458042 197668 458262
rect 194938 455678 195176 458042
rect 197424 455678 197668 458042
rect 194938 455472 197668 455678
rect 208868 458044 211598 458264
rect 208868 455680 209106 458044
rect 211354 455680 211598 458044
rect 208868 455474 211598 455680
rect 222784 458046 225514 458266
rect 222784 455682 223022 458046
rect 225270 455682 225514 458046
rect 222784 455476 225514 455682
rect 236624 458044 239354 458264
rect 236624 455680 236862 458044
rect 239110 455680 239354 458044
rect 236624 455474 239354 455680
rect 250554 458046 253284 458266
rect 250554 455682 250792 458046
rect 253040 455682 253284 458046
rect 250554 455476 253284 455682
rect 264470 458048 267200 458268
rect 264470 455684 264708 458048
rect 266956 455684 267200 458048
rect 264470 455478 267200 455684
rect 278304 458056 281034 458276
rect 278304 455692 278542 458056
rect 280790 455692 281034 458056
rect 278304 455486 281034 455692
rect 292234 458058 294964 458278
rect 292234 455694 292472 458058
rect 294720 455694 294964 458058
rect 292234 455488 294964 455694
rect 306150 458060 308880 458280
rect 306150 455696 306388 458060
rect 308636 455696 308880 458060
rect 306150 455490 308880 455696
rect 319984 458056 322714 458276
rect 319984 455692 320222 458056
rect 322470 455692 322714 458056
rect 319984 455486 322714 455692
rect 333914 458058 336644 458278
rect 333914 455694 334152 458058
rect 336400 455694 336644 458058
rect 333914 455488 336644 455694
rect 347830 458060 350560 458280
rect 347830 455696 348068 458060
rect 350316 455696 350560 458060
rect 347830 455490 350560 455696
rect 361440 458046 364170 458266
rect 361440 455682 361678 458046
rect 363926 455682 364170 458046
rect 361440 455476 364170 455682
rect 375370 458048 378100 458268
rect 375370 455684 375608 458048
rect 377856 455684 378100 458048
rect 375370 455478 378100 455684
rect 389286 458050 392016 458270
rect 389286 455686 389524 458050
rect 391772 455686 392016 458050
rect 389286 455480 392016 455686
rect 403126 458048 405856 458268
rect 403126 455684 403364 458048
rect 405612 455684 405856 458048
rect 403126 455478 405856 455684
rect 417056 458050 419786 458270
rect 417056 455686 417294 458050
rect 419542 455686 419786 458050
rect 417056 455480 419786 455686
rect 194898 446318 197628 446538
rect 194898 443954 195136 446318
rect 197384 443954 197628 446318
rect 194898 443748 197628 443954
rect 208828 446320 211558 446540
rect 208828 443956 209066 446320
rect 211314 443956 211558 446320
rect 208828 443750 211558 443956
rect 222744 446322 225474 446542
rect 222744 443958 222982 446322
rect 225230 443958 225474 446322
rect 222744 443752 225474 443958
rect 236584 446320 239314 446540
rect 236584 443956 236822 446320
rect 239070 443956 239314 446320
rect 236584 443750 239314 443956
rect 250514 446322 253244 446542
rect 250514 443958 250752 446322
rect 253000 443958 253244 446322
rect 250514 443752 253244 443958
rect 264430 446324 267160 446544
rect 264430 443960 264668 446324
rect 266916 443960 267160 446324
rect 264430 443754 267160 443960
rect 278264 446332 280994 446552
rect 278264 443968 278502 446332
rect 280750 443968 280994 446332
rect 278264 443762 280994 443968
rect 292194 446334 294924 446554
rect 292194 443970 292432 446334
rect 294680 443970 294924 446334
rect 292194 443764 294924 443970
rect 306110 446336 308840 446556
rect 306110 443972 306348 446336
rect 308596 443972 308840 446336
rect 306110 443766 308840 443972
rect 319944 446332 322674 446552
rect 319944 443968 320182 446332
rect 322430 443968 322674 446332
rect 319944 443762 322674 443968
rect 333874 446334 336604 446554
rect 333874 443970 334112 446334
rect 336360 443970 336604 446334
rect 333874 443764 336604 443970
rect 347790 446336 350520 446556
rect 347790 443972 348028 446336
rect 350276 443972 350520 446336
rect 347790 443766 350520 443972
rect 361400 446322 364130 446542
rect 361400 443958 361638 446322
rect 363886 443958 364130 446322
rect 361400 443752 364130 443958
rect 375330 446324 378060 446544
rect 375330 443960 375568 446324
rect 377816 443960 378060 446324
rect 375330 443754 378060 443960
rect 389246 446326 391976 446546
rect 389246 443962 389484 446326
rect 391732 443962 391976 446326
rect 389246 443756 391976 443962
rect 403086 446324 405816 446544
rect 403086 443960 403324 446324
rect 405572 443960 405816 446324
rect 403086 443754 405816 443960
rect 417016 446326 419746 446546
rect 417016 443962 417254 446326
rect 419502 443962 419746 446326
rect 417016 443756 419746 443962
rect 194978 422192 197708 422412
rect 194978 419828 195216 422192
rect 197464 419828 197708 422192
rect 194978 419622 197708 419828
rect 208908 422194 211638 422414
rect 208908 419830 209146 422194
rect 211394 419830 211638 422194
rect 208908 419624 211638 419830
rect 278344 422206 281074 422426
rect 278344 419842 278582 422206
rect 280830 419842 281074 422206
rect 278344 419636 281074 419842
rect 292274 422208 295004 422428
rect 292274 419844 292512 422208
rect 294760 419844 295004 422208
rect 292274 419638 295004 419844
rect 306190 422210 308920 422430
rect 306190 419846 306428 422210
rect 308676 419846 308920 422210
rect 306190 419640 308920 419846
rect 320024 422206 322754 422426
rect 320024 419842 320262 422206
rect 322510 419842 322754 422206
rect 320024 419636 322754 419842
rect 333954 422208 336684 422428
rect 333954 419844 334192 422208
rect 336440 419844 336684 422208
rect 333954 419638 336684 419844
rect 194430 407932 197160 408152
rect 194430 405568 194668 407932
rect 196916 405568 197160 407932
rect 194430 405362 197160 405568
rect 208360 407934 211090 408154
rect 208360 405570 208598 407934
rect 210846 405570 211090 407934
rect 208360 405364 211090 405570
rect 277796 407946 280526 408166
rect 277796 405582 278034 407946
rect 280282 405582 280526 407946
rect 277796 405376 280526 405582
rect 291726 407948 294456 408168
rect 291726 405584 291964 407948
rect 294212 405584 294456 407948
rect 291726 405378 294456 405584
rect 305642 407950 308372 408170
rect 305642 405586 305880 407950
rect 308128 405586 308372 407950
rect 305642 405380 308372 405586
rect 319476 407946 322206 408166
rect 319476 405582 319714 407946
rect 321962 405582 322206 407946
rect 319476 405376 322206 405582
rect 333406 407948 336136 408168
rect 333406 405584 333644 407948
rect 335892 405584 336136 407948
rect 333406 405378 336136 405584
rect 194646 395106 197376 395326
rect 194646 392742 194884 395106
rect 197132 392742 197376 395106
rect 194646 392536 197376 392742
rect 208576 395108 211306 395328
rect 208576 392744 208814 395108
rect 211062 392744 211306 395108
rect 208576 392538 211306 392744
rect 278012 395120 280742 395340
rect 278012 392756 278250 395120
rect 280498 392756 280742 395120
rect 278012 392550 280742 392756
rect 291942 395122 294672 395342
rect 291942 392758 292180 395122
rect 294428 392758 294672 395122
rect 291942 392552 294672 392758
rect 305858 395124 308588 395344
rect 305858 392760 306096 395124
rect 308344 392760 308588 395124
rect 305858 392554 308588 392760
rect 319692 395120 322422 395340
rect 319692 392756 319930 395120
rect 322178 392756 322422 395120
rect 319692 392550 322422 392756
rect 333622 395122 336352 395342
rect 333622 392758 333860 395122
rect 336108 392758 336352 395122
rect 333622 392552 336352 392758
rect 194952 386406 197682 386626
rect 194952 384042 195190 386406
rect 197438 384042 197682 386406
rect 194952 383836 197682 384042
rect 208882 386408 211612 386628
rect 208882 384044 209120 386408
rect 211368 384044 211612 386408
rect 208882 383838 211612 384044
rect 278318 386420 281048 386640
rect 278318 384056 278556 386420
rect 280804 384056 281048 386420
rect 278318 383850 281048 384056
rect 292248 386422 294978 386642
rect 292248 384058 292486 386422
rect 294734 384058 294978 386422
rect 292248 383852 294978 384058
rect 306164 386424 308894 386644
rect 306164 384060 306402 386424
rect 308650 384060 308894 386424
rect 306164 383854 308894 384060
rect 319998 386420 322728 386640
rect 319998 384056 320236 386420
rect 322484 384056 322728 386420
rect 319998 383850 322728 384056
rect 333928 386422 336658 386642
rect 333928 384058 334166 386422
rect 336414 384058 336658 386422
rect 333928 383852 336658 384058
rect 277770 372160 280500 372380
rect 277770 369796 278008 372160
rect 280256 369796 280500 372160
rect 277770 369590 280500 369796
rect 291700 372162 294430 372382
rect 291700 369798 291938 372162
rect 294186 369798 294430 372162
rect 291700 369592 294430 369798
rect 305616 372164 308346 372384
rect 305616 369800 305854 372164
rect 308102 369800 308346 372164
rect 305616 369594 308346 369800
rect 319450 372160 322180 372380
rect 319450 369796 319688 372160
rect 321936 369796 322180 372160
rect 319450 369590 322180 369796
rect 333380 372162 336110 372382
rect 333380 369798 333618 372162
rect 335866 369798 336110 372162
rect 333380 369592 336110 369798
rect 347296 372164 350026 372384
rect 347296 369800 347534 372164
rect 349782 369800 350026 372164
rect 347296 369594 350026 369800
rect 360906 372150 363636 372370
rect 360906 369786 361144 372150
rect 363392 369786 363636 372150
rect 360906 369580 363636 369786
rect 374836 372152 377566 372372
rect 374836 369788 375074 372152
rect 377322 369788 377566 372152
rect 374836 369582 377566 369788
rect 388752 372154 391482 372374
rect 388752 369790 388990 372154
rect 391238 369790 391482 372154
rect 388752 369584 391482 369790
rect 222466 359324 225196 359544
rect 222466 356960 222704 359324
rect 224952 356960 225196 359324
rect 222466 356754 225196 356960
rect 236306 359322 239036 359542
rect 236306 356958 236544 359322
rect 238792 356958 239036 359322
rect 236306 356752 239036 356958
rect 250236 359324 252966 359544
rect 250236 356960 250474 359324
rect 252722 356960 252966 359324
rect 250236 356754 252966 356960
rect 264152 359326 266882 359546
rect 264152 356962 264390 359326
rect 266638 356962 266882 359326
rect 264152 356756 266882 356962
rect 277986 359334 280716 359554
rect 277986 356970 278224 359334
rect 280472 356970 280716 359334
rect 277986 356764 280716 356970
rect 291916 359336 294646 359556
rect 291916 356972 292154 359336
rect 294402 356972 294646 359336
rect 291916 356766 294646 356972
rect 305832 359338 308562 359558
rect 305832 356974 306070 359338
rect 308318 356974 308562 359338
rect 305832 356768 308562 356974
rect 319666 359334 322396 359554
rect 319666 356970 319904 359334
rect 322152 356970 322396 359334
rect 319666 356764 322396 356970
rect 333596 359336 336326 359556
rect 333596 356972 333834 359336
rect 336082 356972 336326 359336
rect 333596 356766 336326 356972
rect 347512 359338 350242 359558
rect 347512 356974 347750 359338
rect 349998 356974 350242 359338
rect 347512 356768 350242 356974
rect 361122 359324 363852 359544
rect 361122 356960 361360 359324
rect 363608 356960 363852 359324
rect 361122 356754 363852 356960
rect 375052 359326 377782 359546
rect 375052 356962 375290 359326
rect 377538 356962 377782 359326
rect 375052 356756 377782 356962
rect 388968 359328 391698 359548
rect 388968 356964 389206 359328
rect 391454 356964 391698 359328
rect 388968 356758 391698 356964
rect 221896 347496 224626 347716
rect 221896 345132 222134 347496
rect 224382 345132 224626 347496
rect 221896 344926 224626 345132
rect 235736 347494 238466 347714
rect 235736 345130 235974 347494
rect 238222 345130 238466 347494
rect 235736 344924 238466 345130
rect 249666 347496 252396 347716
rect 249666 345132 249904 347496
rect 252152 345132 252396 347496
rect 249666 344926 252396 345132
rect 263582 347498 266312 347718
rect 263582 345134 263820 347498
rect 266068 345134 266312 347498
rect 263582 344928 266312 345134
rect 277416 347506 280146 347726
rect 277416 345142 277654 347506
rect 279902 345142 280146 347506
rect 277416 344936 280146 345142
rect 291346 347508 294076 347728
rect 291346 345144 291584 347508
rect 293832 345144 294076 347508
rect 291346 344938 294076 345144
rect 305262 347510 307992 347730
rect 305262 345146 305500 347510
rect 307748 345146 307992 347510
rect 305262 344940 307992 345146
rect 319096 347506 321826 347726
rect 319096 345142 319334 347506
rect 321582 345142 321826 347506
rect 319096 344936 321826 345142
rect 333026 347508 335756 347728
rect 333026 345144 333264 347508
rect 335512 345144 335756 347508
rect 333026 344938 335756 345144
rect 346942 347510 349672 347730
rect 346942 345146 347180 347510
rect 349428 345146 349672 347510
rect 346942 344940 349672 345146
rect 360552 347496 363282 347716
rect 360552 345132 360790 347496
rect 363038 345132 363282 347496
rect 360552 344926 363282 345132
rect 374482 347498 377212 347718
rect 374482 345134 374720 347498
rect 376968 345134 377212 347498
rect 374482 344928 377212 345134
rect 388398 347500 391128 347720
rect 388398 345136 388636 347500
rect 390884 345136 391128 347500
rect 388398 344930 391128 345136
rect 222112 334670 224842 334890
rect 222112 332306 222350 334670
rect 224598 332306 224842 334670
rect 222112 332100 224842 332306
rect 235952 334668 238682 334888
rect 235952 332304 236190 334668
rect 238438 332304 238682 334668
rect 235952 332098 238682 332304
rect 249882 334670 252612 334890
rect 249882 332306 250120 334670
rect 252368 332306 252612 334670
rect 249882 332100 252612 332306
rect 263798 334672 266528 334892
rect 263798 332308 264036 334672
rect 266284 332308 266528 334672
rect 263798 332102 266528 332308
rect 277632 334680 280362 334900
rect 277632 332316 277870 334680
rect 280118 332316 280362 334680
rect 277632 332110 280362 332316
rect 291562 334682 294292 334902
rect 291562 332318 291800 334682
rect 294048 332318 294292 334682
rect 291562 332112 294292 332318
rect 305478 334684 308208 334904
rect 305478 332320 305716 334684
rect 307964 332320 308208 334684
rect 305478 332114 308208 332320
rect 319312 334680 322042 334900
rect 319312 332316 319550 334680
rect 321798 332316 322042 334680
rect 319312 332110 322042 332316
rect 333242 334682 335972 334902
rect 333242 332318 333480 334682
rect 335728 332318 335972 334682
rect 333242 332112 335972 332318
rect 347158 334684 349888 334904
rect 347158 332320 347396 334684
rect 349644 332320 349888 334684
rect 347158 332114 349888 332320
rect 360768 334670 363498 334890
rect 360768 332306 361006 334670
rect 363254 332306 363498 334670
rect 360768 332100 363498 332306
rect 374698 334672 377428 334892
rect 374698 332308 374936 334672
rect 377184 332308 377428 334672
rect 374698 332102 377428 332308
rect 388614 334674 391344 334894
rect 388614 332310 388852 334674
rect 391100 332310 391344 334674
rect 388614 332104 391344 332310
rect 195800 319988 198530 320208
rect 195800 317624 196038 319988
rect 198286 317624 198530 319988
rect 195800 317418 198530 317624
rect 209730 319990 212460 320210
rect 209730 317626 209968 319990
rect 212216 317626 212460 319990
rect 209730 317420 212460 317626
rect 279166 320002 281896 320222
rect 279166 317638 279404 320002
rect 281652 317638 281896 320002
rect 279166 317432 281896 317638
rect 293096 320004 295826 320224
rect 293096 317640 293334 320004
rect 295582 317640 295826 320004
rect 293096 317434 295826 317640
rect 307012 320006 309742 320226
rect 307012 317642 307250 320006
rect 309498 317642 309742 320006
rect 307012 317436 309742 317642
rect 320846 320002 323576 320222
rect 320846 317638 321084 320002
rect 323332 317638 323576 320002
rect 320846 317432 323576 317638
rect 334776 320004 337506 320224
rect 334776 317640 335014 320004
rect 337262 317640 337506 320004
rect 334776 317434 337506 317640
rect 196370 310322 199100 310542
rect 196370 307958 196608 310322
rect 198856 307958 199100 310322
rect 196370 307752 199100 307958
rect 210300 310324 213030 310544
rect 210300 307960 210538 310324
rect 212786 307960 213030 310324
rect 210300 307754 213030 307960
rect 279736 310336 282466 310556
rect 279736 307972 279974 310336
rect 282222 307972 282466 310336
rect 279736 307766 282466 307972
rect 293666 310338 296396 310558
rect 293666 307974 293904 310338
rect 296152 307974 296396 310338
rect 293666 307768 296396 307974
rect 307582 310340 310312 310560
rect 307582 307976 307820 310340
rect 310068 307976 310312 310340
rect 307582 307770 310312 307976
rect 321416 310336 324146 310556
rect 321416 307972 321654 310336
rect 323902 307972 324146 310336
rect 321416 307766 324146 307972
rect 335346 310338 338076 310558
rect 335346 307974 335584 310338
rect 337832 307974 338076 310338
rect 335346 307768 338076 307974
rect 196512 299802 199242 300022
rect 196512 297438 196750 299802
rect 198998 297438 199242 299802
rect 196512 297232 199242 297438
rect 210442 299804 213172 300024
rect 210442 297440 210680 299804
rect 212928 297440 213172 299804
rect 210442 297234 213172 297440
rect 279878 299816 282608 300036
rect 279878 297452 280116 299816
rect 282364 297452 282608 299816
rect 279878 297246 282608 297452
rect 293808 299818 296538 300038
rect 293808 297454 294046 299818
rect 296294 297454 296538 299818
rect 293808 297248 296538 297454
rect 307724 299820 310454 300040
rect 307724 297456 307962 299820
rect 310210 297456 310454 299820
rect 307724 297250 310454 297456
rect 321558 299816 324288 300036
rect 321558 297452 321796 299816
rect 324044 297452 324288 299816
rect 321558 297246 324288 297452
rect 335488 299818 338218 300038
rect 335488 297454 335726 299818
rect 337974 297454 338218 299818
rect 335488 297248 338218 297454
rect 196370 288854 199100 289074
rect 196370 286490 196608 288854
rect 198856 286490 199100 288854
rect 196370 286284 199100 286490
rect 210300 288856 213030 289076
rect 210300 286492 210538 288856
rect 212786 286492 213030 288856
rect 210300 286286 213030 286492
rect 279736 288868 282466 289088
rect 279736 286504 279974 288868
rect 282222 286504 282466 288868
rect 279736 286298 282466 286504
rect 293666 288870 296396 289090
rect 293666 286506 293904 288870
rect 296152 286506 296396 288870
rect 293666 286300 296396 286506
rect 307582 288872 310312 289092
rect 307582 286508 307820 288872
rect 310068 286508 310312 288872
rect 307582 286302 310312 286508
rect 321416 288868 324146 289088
rect 321416 286504 321654 288868
rect 323902 286504 324146 288868
rect 321416 286298 324146 286504
rect 335346 288870 338076 289090
rect 335346 286506 335584 288870
rect 337832 286506 338076 288870
rect 335346 286300 338076 286506
rect 196654 276630 199384 276850
rect 196654 274266 196892 276630
rect 199140 274266 199384 276630
rect 196654 274060 199384 274266
rect 210584 276632 213314 276852
rect 210584 274268 210822 276632
rect 213070 274268 213314 276632
rect 210584 274062 213314 274268
rect 280020 276644 282750 276864
rect 280020 274280 280258 276644
rect 282506 274280 282750 276644
rect 280020 274074 282750 274280
rect 293950 276646 296680 276866
rect 293950 274282 294188 276646
rect 296436 274282 296680 276646
rect 293950 274076 296680 274282
rect 307866 276648 310596 276868
rect 307866 274284 308104 276648
rect 310352 274284 310596 276648
rect 307866 274078 310596 274284
rect 321700 276644 324430 276864
rect 321700 274280 321938 276644
rect 324186 274280 324430 276644
rect 321700 274074 324430 274280
rect 335630 276646 338360 276866
rect 335630 274282 335868 276646
rect 338116 274282 338360 276646
rect 335630 274076 338360 274282
rect 196234 260882 198964 261102
rect 196234 258518 196472 260882
rect 198720 258518 198964 260882
rect 196234 258312 198964 258518
rect 210164 260884 212894 261104
rect 210164 258520 210402 260884
rect 212650 258520 212894 260884
rect 210164 258314 212894 258520
rect 224080 260886 226810 261106
rect 224080 258522 224318 260886
rect 226566 258522 226810 260886
rect 224080 258316 226810 258522
rect 237920 260884 240650 261104
rect 237920 258520 238158 260884
rect 240406 258520 240650 260884
rect 237920 258314 240650 258520
rect 251850 260886 254580 261106
rect 251850 258522 252088 260886
rect 254336 258522 254580 260886
rect 251850 258316 254580 258522
rect 265766 260888 268496 261108
rect 265766 258524 266004 260888
rect 268252 258524 268496 260888
rect 265766 258318 268496 258524
rect 279600 260896 282330 261116
rect 279600 258532 279838 260896
rect 282086 258532 282330 260896
rect 279600 258326 282330 258532
rect 293530 260898 296260 261118
rect 293530 258534 293768 260898
rect 296016 258534 296260 260898
rect 293530 258328 296260 258534
rect 307446 260900 310176 261120
rect 307446 258536 307684 260900
rect 309932 258536 310176 260900
rect 307446 258330 310176 258536
rect 321280 260896 324010 261116
rect 321280 258532 321518 260896
rect 323766 258532 324010 260896
rect 321280 258326 324010 258532
rect 335210 260898 337940 261118
rect 335210 258534 335448 260898
rect 337696 258534 337940 260898
rect 335210 258328 337940 258534
rect 195268 238250 197998 238470
rect 195268 235886 195506 238250
rect 197754 235886 197998 238250
rect 195268 235680 197998 235886
rect 209198 238252 211928 238472
rect 209198 235888 209436 238252
rect 211684 235888 211928 238252
rect 209198 235682 211928 235888
rect 278634 238264 281364 238484
rect 278634 235900 278872 238264
rect 281120 235900 281364 238264
rect 278634 235694 281364 235900
rect 292564 238266 295294 238486
rect 292564 235902 292802 238266
rect 295050 235902 295294 238266
rect 292564 235696 295294 235902
rect 306480 238268 309210 238488
rect 306480 235904 306718 238268
rect 308966 235904 309210 238268
rect 306480 235698 309210 235904
rect 320314 238264 323044 238484
rect 320314 235900 320552 238264
rect 322800 235900 323044 238264
rect 320314 235694 323044 235900
rect 334244 238266 336974 238486
rect 334244 235902 334482 238266
rect 336730 235902 336974 238266
rect 334244 235696 336974 235902
rect 195678 222346 198408 222566
rect 195678 219982 195916 222346
rect 198164 219982 198408 222346
rect 195678 219776 198408 219982
rect 209608 222348 212338 222568
rect 209608 219984 209846 222348
rect 212094 219984 212338 222348
rect 209608 219778 212338 219984
rect 279044 222360 281774 222580
rect 279044 219996 279282 222360
rect 281530 219996 281774 222360
rect 279044 219790 281774 219996
rect 292974 222362 295704 222582
rect 292974 219998 293212 222362
rect 295460 219998 295704 222362
rect 292974 219792 295704 219998
rect 306890 222364 309620 222584
rect 306890 220000 307128 222364
rect 309376 220000 309620 222364
rect 306890 219794 309620 220000
rect 320724 222360 323454 222580
rect 320724 219996 320962 222360
rect 323210 219996 323454 222360
rect 320724 219790 323454 219996
rect 334654 222362 337384 222582
rect 334654 219998 334892 222362
rect 337140 219998 337384 222362
rect 334654 219792 337384 219998
rect 195678 205894 198408 206114
rect 195678 203530 195916 205894
rect 198164 203530 198408 205894
rect 195678 203324 198408 203530
rect 209608 205896 212338 206116
rect 209608 203532 209846 205896
rect 212094 203532 212338 205896
rect 209608 203326 212338 203532
rect 279044 205908 281774 206128
rect 279044 203544 279282 205908
rect 281530 203544 281774 205908
rect 279044 203338 281774 203544
rect 292974 205910 295704 206130
rect 292974 203546 293212 205910
rect 295460 203546 295704 205910
rect 292974 203340 295704 203546
rect 306890 205912 309620 206132
rect 306890 203548 307128 205912
rect 309376 203548 309620 205912
rect 306890 203342 309620 203548
rect 320724 205908 323454 206128
rect 320724 203544 320962 205908
rect 323210 203544 323454 205908
rect 320724 203338 323454 203544
rect 334654 205910 337384 206130
rect 334654 203546 334892 205910
rect 337140 203546 337384 205910
rect 334654 203340 337384 203546
rect 195268 191086 197998 191306
rect 195268 188722 195506 191086
rect 197754 188722 197998 191086
rect 195268 188516 197998 188722
rect 209198 191088 211928 191308
rect 209198 188724 209436 191088
rect 211684 188724 211928 191088
rect 209198 188518 211928 188724
rect 278634 191100 281364 191320
rect 278634 188736 278872 191100
rect 281120 188736 281364 191100
rect 278634 188530 281364 188736
rect 292564 191102 295294 191322
rect 292564 188738 292802 191102
rect 295050 188738 295294 191102
rect 292564 188532 295294 188738
rect 306480 191104 309210 191324
rect 306480 188740 306718 191104
rect 308966 188740 309210 191104
rect 306480 188534 309210 188740
rect 320314 191100 323044 191320
rect 320314 188736 320552 191100
rect 322800 188736 323044 191100
rect 320314 188530 323044 188736
rect 334244 191102 336974 191322
rect 334244 188738 334482 191102
rect 336730 188738 336974 191102
rect 334244 188532 336974 188738
rect 194720 176826 197450 177046
rect 194720 174462 194958 176826
rect 197206 174462 197450 176826
rect 194720 174256 197450 174462
rect 208650 176828 211380 177048
rect 208650 174464 208888 176828
rect 211136 174464 211380 176828
rect 208650 174258 211380 174464
rect 222566 176830 225296 177050
rect 222566 174466 222804 176830
rect 225052 174466 225296 176830
rect 222566 174260 225296 174466
rect 236406 176828 239136 177048
rect 236406 174464 236644 176828
rect 238892 174464 239136 176828
rect 236406 174258 239136 174464
rect 250336 176830 253066 177050
rect 250336 174466 250574 176830
rect 252822 174466 253066 176830
rect 250336 174260 253066 174466
rect 264252 176832 266982 177052
rect 264252 174468 264490 176832
rect 266738 174468 266982 176832
rect 264252 174262 266982 174468
rect 278086 176840 280816 177060
rect 278086 174476 278324 176840
rect 280572 174476 280816 176840
rect 278086 174270 280816 174476
rect 292016 176842 294746 177062
rect 292016 174478 292254 176842
rect 294502 174478 294746 176842
rect 292016 174272 294746 174478
rect 305932 176844 308662 177064
rect 305932 174480 306170 176844
rect 308418 174480 308662 176844
rect 305932 174274 308662 174480
rect 319766 176840 322496 177060
rect 319766 174476 320004 176840
rect 322252 174476 322496 176840
rect 319766 174270 322496 174476
rect 333696 176842 336426 177062
rect 333696 174478 333934 176842
rect 336182 174478 336426 176842
rect 333696 174272 336426 174478
rect 194936 164000 197666 164220
rect 194936 161636 195174 164000
rect 197422 161636 197666 164000
rect 194936 161430 197666 161636
rect 208866 164002 211596 164222
rect 208866 161638 209104 164002
rect 211352 161638 211596 164002
rect 208866 161432 211596 161638
rect 222782 164004 225512 164224
rect 222782 161640 223020 164004
rect 225268 161640 225512 164004
rect 222782 161434 225512 161640
rect 236622 164002 239352 164222
rect 236622 161638 236860 164002
rect 239108 161638 239352 164002
rect 236622 161432 239352 161638
rect 250552 164004 253282 164224
rect 250552 161640 250790 164004
rect 253038 161640 253282 164004
rect 250552 161434 253282 161640
rect 264468 164006 267198 164226
rect 264468 161642 264706 164006
rect 266954 161642 267198 164006
rect 264468 161436 267198 161642
rect 278302 164014 281032 164234
rect 278302 161650 278540 164014
rect 280788 161650 281032 164014
rect 278302 161444 281032 161650
rect 292232 164016 294962 164236
rect 292232 161652 292470 164016
rect 294718 161652 294962 164016
rect 292232 161446 294962 161652
rect 306148 164018 308878 164238
rect 306148 161654 306386 164018
rect 308634 161654 308878 164018
rect 306148 161448 308878 161654
rect 319982 164014 322712 164234
rect 319982 161650 320220 164014
rect 322468 161650 322712 164014
rect 319982 161444 322712 161650
rect 333912 164016 336642 164236
rect 333912 161652 334150 164016
rect 336398 161652 336642 164016
rect 333912 161446 336642 161652
rect 194668 141640 197398 141860
rect 194668 139276 194906 141640
rect 197154 139276 197398 141640
rect 194668 139070 197398 139276
rect 208598 141642 211328 141862
rect 208598 139278 208836 141642
rect 211084 139278 211328 141642
rect 208598 139072 211328 139278
rect 222514 141644 225244 141864
rect 222514 139280 222752 141644
rect 225000 139280 225244 141644
rect 222514 139074 225244 139280
rect 236354 141642 239084 141862
rect 236354 139278 236592 141642
rect 238840 139278 239084 141642
rect 236354 139072 239084 139278
rect 250284 141644 253014 141864
rect 250284 139280 250522 141644
rect 252770 139280 253014 141644
rect 250284 139074 253014 139280
rect 264200 141646 266930 141866
rect 264200 139282 264438 141646
rect 266686 139282 266930 141646
rect 264200 139076 266930 139282
rect 278034 141654 280764 141874
rect 278034 139290 278272 141654
rect 280520 139290 280764 141654
rect 278034 139084 280764 139290
rect 291964 141656 294694 141876
rect 291964 139292 292202 141656
rect 294450 139292 294694 141656
rect 291964 139086 294694 139292
rect 305880 141658 308610 141878
rect 305880 139294 306118 141658
rect 308366 139294 308610 141658
rect 305880 139088 308610 139294
rect 319714 141654 322444 141874
rect 319714 139290 319952 141654
rect 322200 139290 322444 141654
rect 319714 139084 322444 139290
rect 333644 141656 336374 141876
rect 333644 139292 333882 141656
rect 336130 139292 336374 141656
rect 333644 139086 336374 139292
rect 347560 141658 350290 141878
rect 347560 139294 347798 141658
rect 350046 139294 350290 141658
rect 347560 139088 350290 139294
rect 194598 129160 197328 129380
rect 194598 126796 194836 129160
rect 197084 126796 197328 129160
rect 194598 126590 197328 126796
rect 208528 129162 211258 129382
rect 208528 126798 208766 129162
rect 211014 126798 211258 129162
rect 208528 126592 211258 126798
rect 222444 129164 225174 129384
rect 222444 126800 222682 129164
rect 224930 126800 225174 129164
rect 222444 126594 225174 126800
rect 236284 129162 239014 129382
rect 236284 126798 236522 129162
rect 238770 126798 239014 129162
rect 236284 126592 239014 126798
rect 250214 129164 252944 129384
rect 250214 126800 250452 129164
rect 252700 126800 252944 129164
rect 250214 126594 252944 126800
rect 264130 129166 266860 129386
rect 264130 126802 264368 129166
rect 266616 126802 266860 129166
rect 264130 126596 266860 126802
rect 277964 129174 280694 129394
rect 277964 126810 278202 129174
rect 280450 126810 280694 129174
rect 277964 126604 280694 126810
rect 291894 129176 294624 129396
rect 291894 126812 292132 129176
rect 294380 126812 294624 129176
rect 291894 126606 294624 126812
rect 305810 129178 308540 129398
rect 305810 126814 306048 129178
rect 308296 126814 308540 129178
rect 305810 126608 308540 126814
rect 319644 129174 322374 129394
rect 319644 126810 319882 129174
rect 322130 126810 322374 129174
rect 319644 126604 322374 126810
rect 333574 129176 336304 129396
rect 333574 126812 333812 129176
rect 336060 126812 336304 129176
rect 333574 126606 336304 126812
rect 347490 129178 350220 129398
rect 347490 126814 347728 129178
rect 349976 126814 350220 129178
rect 347490 126608 350220 126814
rect 194528 117726 197258 117946
rect 194528 115362 194766 117726
rect 197014 115362 197258 117726
rect 194528 115156 197258 115362
rect 208458 117728 211188 117948
rect 208458 115364 208696 117728
rect 210944 115364 211188 117728
rect 208458 115158 211188 115364
rect 222374 117730 225104 117950
rect 222374 115366 222612 117730
rect 224860 115366 225104 117730
rect 222374 115160 225104 115366
rect 236214 117728 238944 117948
rect 236214 115364 236452 117728
rect 238700 115364 238944 117728
rect 236214 115158 238944 115364
rect 250144 117730 252874 117950
rect 250144 115366 250382 117730
rect 252630 115366 252874 117730
rect 250144 115160 252874 115366
rect 264060 117732 266790 117952
rect 264060 115368 264298 117732
rect 266546 115368 266790 117732
rect 264060 115162 266790 115368
rect 277894 117740 280624 117960
rect 277894 115376 278132 117740
rect 280380 115376 280624 117740
rect 277894 115170 280624 115376
rect 291824 117742 294554 117962
rect 291824 115378 292062 117742
rect 294310 115378 294554 117742
rect 291824 115172 294554 115378
rect 305740 117744 308470 117964
rect 305740 115380 305978 117744
rect 308226 115380 308470 117744
rect 305740 115174 308470 115380
rect 319574 117740 322304 117960
rect 319574 115376 319812 117740
rect 322060 115376 322304 117740
rect 319574 115170 322304 115376
rect 333504 117742 336234 117962
rect 333504 115378 333742 117742
rect 335990 115378 336234 117742
rect 333504 115172 336234 115378
rect 347420 117744 350150 117964
rect 347420 115380 347658 117744
rect 349906 115380 350150 117744
rect 347420 115174 350150 115380
rect 194390 105316 197120 105536
rect 194390 102952 194628 105316
rect 196876 102952 197120 105316
rect 194390 102746 197120 102952
rect 208320 105318 211050 105538
rect 208320 102954 208558 105318
rect 210806 102954 211050 105318
rect 208320 102748 211050 102954
rect 222236 105320 224966 105540
rect 222236 102956 222474 105320
rect 224722 102956 224966 105320
rect 222236 102750 224966 102956
rect 236076 105318 238806 105538
rect 236076 102954 236314 105318
rect 238562 102954 238806 105318
rect 236076 102748 238806 102954
rect 250006 105320 252736 105540
rect 250006 102956 250244 105320
rect 252492 102956 252736 105320
rect 250006 102750 252736 102956
rect 263922 105322 266652 105542
rect 263922 102958 264160 105322
rect 266408 102958 266652 105322
rect 263922 102752 266652 102958
rect 277756 105330 280486 105550
rect 277756 102966 277994 105330
rect 280242 102966 280486 105330
rect 277756 102760 280486 102966
rect 291686 105332 294416 105552
rect 291686 102968 291924 105332
rect 294172 102968 294416 105332
rect 291686 102762 294416 102968
rect 305602 105334 308332 105554
rect 305602 102970 305840 105334
rect 308088 102970 308332 105334
rect 305602 102764 308332 102970
rect 319436 105330 322166 105550
rect 319436 102966 319674 105330
rect 321922 102966 322166 105330
rect 319436 102760 322166 102966
rect 333366 105332 336096 105552
rect 333366 102968 333604 105332
rect 335852 102968 336096 105332
rect 333366 102762 336096 102968
rect 347282 105334 350012 105554
rect 347282 102970 347520 105334
rect 349768 102970 350012 105334
rect 347282 102764 350012 102970
rect 277180 89614 279910 89834
rect 277180 87250 277418 89614
rect 279666 87250 279910 89614
rect 277180 87044 279910 87250
rect 291110 89616 293840 89836
rect 291110 87252 291348 89616
rect 293596 87252 293840 89616
rect 291110 87046 293840 87252
rect 305026 89618 307756 89838
rect 305026 87254 305264 89618
rect 307512 87254 307756 89618
rect 305026 87048 307756 87254
rect 318860 89614 321590 89834
rect 318860 87250 319098 89614
rect 321346 87250 321590 89614
rect 318860 87044 321590 87250
rect 332790 89616 335520 89836
rect 332790 87252 333028 89616
rect 335276 87252 335520 89616
rect 332790 87046 335520 87252
rect 346706 89618 349436 89838
rect 346706 87254 346944 89618
rect 349192 87254 349436 89618
rect 346706 87048 349436 87254
rect 277180 77026 279910 77246
rect 277180 74662 277418 77026
rect 279666 74662 279910 77026
rect 277180 74456 279910 74662
rect 291110 77028 293840 77248
rect 291110 74664 291348 77028
rect 293596 74664 293840 77028
rect 291110 74458 293840 74664
rect 305026 77030 307756 77250
rect 305026 74666 305264 77030
rect 307512 74666 307756 77030
rect 305026 74460 307756 74666
rect 318860 77026 321590 77246
rect 318860 74662 319098 77026
rect 321346 74662 321590 77026
rect 318860 74456 321590 74662
rect 332790 77028 335520 77248
rect 332790 74664 333028 77028
rect 335276 74664 335520 77028
rect 332790 74458 335520 74664
rect 346706 77030 349436 77250
rect 346706 74666 346944 77030
rect 349192 74666 349436 77030
rect 346706 74460 349436 74666
rect 277180 64438 279910 64658
rect 277180 62074 277418 64438
rect 279666 62074 279910 64438
rect 277180 61868 279910 62074
rect 291110 64440 293840 64660
rect 291110 62076 291348 64440
rect 293596 62076 293840 64440
rect 291110 61870 293840 62076
rect 305026 64442 307756 64662
rect 305026 62078 305264 64442
rect 307512 62078 307756 64442
rect 305026 61872 307756 62078
rect 318860 64438 321590 64658
rect 318860 62074 319098 64438
rect 321346 62074 321590 64438
rect 318860 61868 321590 62074
rect 332790 64440 335520 64660
rect 332790 62076 333028 64440
rect 335276 62076 335520 64440
rect 332790 61870 335520 62076
rect 346706 64442 349436 64662
rect 346706 62078 346944 64442
rect 349192 62078 349436 64442
rect 346706 61872 349436 62078
<< psubdiffcont >>
rect 194026 663430 196274 665794
rect 207956 663432 210204 665796
rect 277392 663444 279640 665808
rect 291322 663446 293570 665810
rect 305238 663448 307486 665812
rect 319072 663444 321320 665808
rect 333002 663446 335250 665810
rect 346918 663448 349166 665812
rect 360528 663434 362776 665798
rect 374458 663436 376706 665800
rect 388374 663438 390622 665802
rect 402214 663436 404462 665800
rect 416144 663438 418392 665802
rect 194574 650774 196822 653138
rect 208504 650776 210752 653140
rect 277940 650788 280188 653152
rect 291870 650790 294118 653154
rect 305786 650792 308034 653156
rect 319620 650788 321868 653152
rect 333550 650790 335798 653154
rect 347466 650792 349714 653156
rect 361076 650778 363324 653142
rect 375006 650780 377254 653144
rect 388922 650782 391170 653146
rect 402762 650780 405010 653144
rect 416692 650782 418940 653146
rect 194026 636514 196274 638878
rect 207956 636516 210204 638880
rect 277392 636528 279640 638892
rect 291322 636530 293570 638894
rect 305238 636532 307486 638896
rect 319072 636528 321320 638892
rect 333002 636530 335250 638894
rect 346918 636532 349166 638896
rect 360528 636518 362776 638882
rect 374458 636520 376706 638884
rect 388374 636522 390622 638886
rect 402214 636520 404462 638884
rect 416144 636522 418392 638886
rect 194586 622252 196834 624616
rect 208516 622254 210764 624618
rect 277952 622266 280200 624630
rect 291882 622268 294130 624632
rect 305798 622270 308046 624634
rect 319632 622266 321880 624630
rect 333562 622268 335810 624632
rect 347478 622270 349726 624634
rect 361088 622256 363336 624620
rect 375018 622258 377266 624622
rect 388934 622260 391182 624624
rect 402774 622258 405022 624622
rect 416704 622260 418952 624624
rect 166486 608032 168734 610396
rect 180402 608034 182650 610398
rect 194038 607992 196286 610356
rect 207968 607994 210216 610358
rect 221884 607996 224132 610360
rect 235724 607994 237972 610358
rect 249654 607996 251902 610360
rect 263570 607998 265818 610362
rect 277404 608006 279652 610370
rect 291334 608008 293582 610372
rect 305250 608010 307498 610374
rect 319084 608006 321332 610370
rect 333014 608008 335262 610372
rect 346930 608010 349178 610374
rect 360540 607996 362788 610360
rect 374470 607998 376718 610362
rect 388386 608000 390634 610364
rect 402226 607998 404474 610362
rect 416156 608000 418404 610364
rect 194764 589534 197012 591898
rect 208694 589536 210942 591900
rect 278130 589548 280378 591912
rect 292060 589550 294308 591914
rect 305976 589552 308224 591916
rect 319810 589548 322058 591912
rect 333740 589550 335988 591914
rect 375196 589540 377444 591904
rect 389112 589542 391360 591906
rect 194216 575274 196464 577638
rect 208146 575276 210394 577640
rect 277582 575288 279830 577652
rect 291512 575290 293760 577654
rect 305428 575292 307676 577656
rect 319262 575288 321510 577652
rect 333192 575290 335440 577654
rect 374648 575280 376896 577644
rect 388564 575282 390812 577646
rect 194432 562448 196680 564812
rect 208362 562450 210610 564814
rect 277798 562462 280046 564826
rect 291728 562464 293976 564828
rect 305644 562466 307892 564830
rect 319478 562462 321726 564826
rect 333408 562464 335656 564828
rect 374864 562454 377112 564818
rect 388780 562456 391028 564820
rect 194866 544718 197114 547082
rect 208796 544720 211044 547084
rect 222712 544722 224960 547086
rect 236552 544720 238800 547084
rect 250482 544722 252730 547086
rect 264398 544724 266646 547088
rect 278232 544732 280480 547096
rect 292162 544734 294410 547098
rect 306078 544736 308326 547100
rect 319912 544732 322160 547096
rect 333842 544734 336090 547098
rect 347758 544736 350006 547100
rect 361368 544722 363616 547086
rect 375298 544724 377546 547088
rect 389214 544726 391462 547090
rect 403054 544724 405302 547088
rect 416984 544726 419232 547090
rect 194318 530458 196566 532822
rect 208248 530460 210496 532824
rect 222164 530462 224412 532826
rect 236004 530460 238252 532824
rect 249934 530462 252182 532826
rect 263850 530464 266098 532828
rect 277684 530472 279932 532836
rect 291614 530474 293862 532838
rect 305530 530476 307778 532840
rect 319364 530472 321612 532836
rect 333294 530474 335542 532838
rect 347210 530476 349458 532840
rect 360820 530462 363068 532826
rect 374750 530464 376998 532828
rect 388666 530466 390914 532830
rect 402506 530464 404754 532828
rect 416436 530466 418684 532830
rect 194534 517632 196782 519996
rect 208464 517634 210712 519998
rect 222380 517636 224628 520000
rect 236220 517634 238468 519998
rect 250150 517636 252398 520000
rect 264066 517638 266314 520002
rect 277900 517646 280148 520010
rect 291830 517648 294078 520012
rect 305746 517650 307994 520014
rect 319580 517646 321828 520010
rect 333510 517648 335758 520012
rect 347426 517650 349674 520014
rect 361036 517636 363284 520000
rect 374966 517638 377214 520002
rect 388882 517640 391130 520004
rect 402722 517638 404970 520002
rect 416652 517640 418900 520004
rect 194928 496210 197176 498574
rect 208858 496212 211106 498576
rect 222774 496214 225022 498578
rect 236614 496212 238862 498576
rect 250544 496214 252792 498578
rect 264460 496216 266708 498580
rect 278294 496224 280542 498588
rect 292224 496226 294472 498590
rect 306140 496228 308388 498592
rect 319974 496224 322222 498588
rect 333904 496226 336152 498590
rect 347820 496228 350068 498592
rect 361430 496214 363678 498578
rect 375360 496216 377608 498580
rect 389276 496218 391524 498582
rect 403116 496216 405364 498580
rect 417046 496218 419294 498582
rect 194380 481950 196628 484314
rect 208310 481952 210558 484316
rect 222226 481954 224474 484318
rect 236066 481952 238314 484316
rect 249996 481954 252244 484318
rect 263912 481956 266160 484320
rect 277746 481964 279994 484328
rect 291676 481966 293924 484330
rect 305592 481968 307840 484332
rect 319426 481964 321674 484328
rect 333356 481966 335604 484330
rect 347272 481968 349520 484332
rect 360882 481954 363130 484318
rect 374812 481956 377060 484320
rect 388728 481958 390976 484322
rect 402568 481956 404816 484320
rect 416498 481958 418746 484322
rect 194596 469124 196844 471488
rect 208526 469126 210774 471490
rect 222442 469128 224690 471492
rect 236282 469126 238530 471490
rect 250212 469128 252460 471492
rect 264128 469130 266376 471494
rect 277962 469138 280210 471502
rect 291892 469140 294140 471504
rect 305808 469142 308056 471506
rect 319642 469138 321890 471502
rect 333572 469140 335820 471504
rect 347488 469142 349736 471506
rect 361098 469128 363346 471492
rect 375028 469130 377276 471494
rect 388944 469132 391192 471496
rect 402784 469130 405032 471494
rect 416714 469132 418962 471496
rect 195176 455678 197424 458042
rect 209106 455680 211354 458044
rect 223022 455682 225270 458046
rect 236862 455680 239110 458044
rect 250792 455682 253040 458046
rect 264708 455684 266956 458048
rect 278542 455692 280790 458056
rect 292472 455694 294720 458058
rect 306388 455696 308636 458060
rect 320222 455692 322470 458056
rect 334152 455694 336400 458058
rect 348068 455696 350316 458060
rect 361678 455682 363926 458046
rect 375608 455684 377856 458048
rect 389524 455686 391772 458050
rect 403364 455684 405612 458048
rect 417294 455686 419542 458050
rect 195136 443954 197384 446318
rect 209066 443956 211314 446320
rect 222982 443958 225230 446322
rect 236822 443956 239070 446320
rect 250752 443958 253000 446322
rect 264668 443960 266916 446324
rect 278502 443968 280750 446332
rect 292432 443970 294680 446334
rect 306348 443972 308596 446336
rect 320182 443968 322430 446332
rect 334112 443970 336360 446334
rect 348028 443972 350276 446336
rect 361638 443958 363886 446322
rect 375568 443960 377816 446324
rect 389484 443962 391732 446326
rect 403324 443960 405572 446324
rect 417254 443962 419502 446326
rect 195216 419828 197464 422192
rect 209146 419830 211394 422194
rect 278582 419842 280830 422206
rect 292512 419844 294760 422208
rect 306428 419846 308676 422210
rect 320262 419842 322510 422206
rect 334192 419844 336440 422208
rect 194668 405568 196916 407932
rect 208598 405570 210846 407934
rect 278034 405582 280282 407946
rect 291964 405584 294212 407948
rect 305880 405586 308128 407950
rect 319714 405582 321962 407946
rect 333644 405584 335892 407948
rect 194884 392742 197132 395106
rect 208814 392744 211062 395108
rect 278250 392756 280498 395120
rect 292180 392758 294428 395122
rect 306096 392760 308344 395124
rect 319930 392756 322178 395120
rect 333860 392758 336108 395122
rect 195190 384042 197438 386406
rect 209120 384044 211368 386408
rect 278556 384056 280804 386420
rect 292486 384058 294734 386422
rect 306402 384060 308650 386424
rect 320236 384056 322484 386420
rect 334166 384058 336414 386422
rect 278008 369796 280256 372160
rect 291938 369798 294186 372162
rect 305854 369800 308102 372164
rect 319688 369796 321936 372160
rect 333618 369798 335866 372162
rect 347534 369800 349782 372164
rect 361144 369786 363392 372150
rect 375074 369788 377322 372152
rect 388990 369790 391238 372154
rect 222704 356960 224952 359324
rect 236544 356958 238792 359322
rect 250474 356960 252722 359324
rect 264390 356962 266638 359326
rect 278224 356970 280472 359334
rect 292154 356972 294402 359336
rect 306070 356974 308318 359338
rect 319904 356970 322152 359334
rect 333834 356972 336082 359336
rect 347750 356974 349998 359338
rect 361360 356960 363608 359324
rect 375290 356962 377538 359326
rect 389206 356964 391454 359328
rect 222134 345132 224382 347496
rect 235974 345130 238222 347494
rect 249904 345132 252152 347496
rect 263820 345134 266068 347498
rect 277654 345142 279902 347506
rect 291584 345144 293832 347508
rect 305500 345146 307748 347510
rect 319334 345142 321582 347506
rect 333264 345144 335512 347508
rect 347180 345146 349428 347510
rect 360790 345132 363038 347496
rect 374720 345134 376968 347498
rect 388636 345136 390884 347500
rect 222350 332306 224598 334670
rect 236190 332304 238438 334668
rect 250120 332306 252368 334670
rect 264036 332308 266284 334672
rect 277870 332316 280118 334680
rect 291800 332318 294048 334682
rect 305716 332320 307964 334684
rect 319550 332316 321798 334680
rect 333480 332318 335728 334682
rect 347396 332320 349644 334684
rect 361006 332306 363254 334670
rect 374936 332308 377184 334672
rect 388852 332310 391100 334674
rect 196038 317624 198286 319988
rect 209968 317626 212216 319990
rect 279404 317638 281652 320002
rect 293334 317640 295582 320004
rect 307250 317642 309498 320006
rect 321084 317638 323332 320002
rect 335014 317640 337262 320004
rect 196608 307958 198856 310322
rect 210538 307960 212786 310324
rect 279974 307972 282222 310336
rect 293904 307974 296152 310338
rect 307820 307976 310068 310340
rect 321654 307972 323902 310336
rect 335584 307974 337832 310338
rect 196750 297438 198998 299802
rect 210680 297440 212928 299804
rect 280116 297452 282364 299816
rect 294046 297454 296294 299818
rect 307962 297456 310210 299820
rect 321796 297452 324044 299816
rect 335726 297454 337974 299818
rect 196608 286490 198856 288854
rect 210538 286492 212786 288856
rect 279974 286504 282222 288868
rect 293904 286506 296152 288870
rect 307820 286508 310068 288872
rect 321654 286504 323902 288868
rect 335584 286506 337832 288870
rect 196892 274266 199140 276630
rect 210822 274268 213070 276632
rect 280258 274280 282506 276644
rect 294188 274282 296436 276646
rect 308104 274284 310352 276648
rect 321938 274280 324186 276644
rect 335868 274282 338116 276646
rect 196472 258518 198720 260882
rect 210402 258520 212650 260884
rect 224318 258522 226566 260886
rect 238158 258520 240406 260884
rect 252088 258522 254336 260886
rect 266004 258524 268252 260888
rect 279838 258532 282086 260896
rect 293768 258534 296016 260898
rect 307684 258536 309932 260900
rect 321518 258532 323766 260896
rect 335448 258534 337696 260898
rect 195506 235886 197754 238250
rect 209436 235888 211684 238252
rect 278872 235900 281120 238264
rect 292802 235902 295050 238266
rect 306718 235904 308966 238268
rect 320552 235900 322800 238264
rect 334482 235902 336730 238266
rect 195916 219982 198164 222346
rect 209846 219984 212094 222348
rect 279282 219996 281530 222360
rect 293212 219998 295460 222362
rect 307128 220000 309376 222364
rect 320962 219996 323210 222360
rect 334892 219998 337140 222362
rect 195916 203530 198164 205894
rect 209846 203532 212094 205896
rect 279282 203544 281530 205908
rect 293212 203546 295460 205910
rect 307128 203548 309376 205912
rect 320962 203544 323210 205908
rect 334892 203546 337140 205910
rect 195506 188722 197754 191086
rect 209436 188724 211684 191088
rect 278872 188736 281120 191100
rect 292802 188738 295050 191102
rect 306718 188740 308966 191104
rect 320552 188736 322800 191100
rect 334482 188738 336730 191102
rect 194958 174462 197206 176826
rect 208888 174464 211136 176828
rect 222804 174466 225052 176830
rect 236644 174464 238892 176828
rect 250574 174466 252822 176830
rect 264490 174468 266738 176832
rect 278324 174476 280572 176840
rect 292254 174478 294502 176842
rect 306170 174480 308418 176844
rect 320004 174476 322252 176840
rect 333934 174478 336182 176842
rect 195174 161636 197422 164000
rect 209104 161638 211352 164002
rect 223020 161640 225268 164004
rect 236860 161638 239108 164002
rect 250790 161640 253038 164004
rect 264706 161642 266954 164006
rect 278540 161650 280788 164014
rect 292470 161652 294718 164016
rect 306386 161654 308634 164018
rect 320220 161650 322468 164014
rect 334150 161652 336398 164016
rect 194906 139276 197154 141640
rect 208836 139278 211084 141642
rect 222752 139280 225000 141644
rect 236592 139278 238840 141642
rect 250522 139280 252770 141644
rect 264438 139282 266686 141646
rect 278272 139290 280520 141654
rect 292202 139292 294450 141656
rect 306118 139294 308366 141658
rect 319952 139290 322200 141654
rect 333882 139292 336130 141656
rect 347798 139294 350046 141658
rect 194836 126796 197084 129160
rect 208766 126798 211014 129162
rect 222682 126800 224930 129164
rect 236522 126798 238770 129162
rect 250452 126800 252700 129164
rect 264368 126802 266616 129166
rect 278202 126810 280450 129174
rect 292132 126812 294380 129176
rect 306048 126814 308296 129178
rect 319882 126810 322130 129174
rect 333812 126812 336060 129176
rect 347728 126814 349976 129178
rect 194766 115362 197014 117726
rect 208696 115364 210944 117728
rect 222612 115366 224860 117730
rect 236452 115364 238700 117728
rect 250382 115366 252630 117730
rect 264298 115368 266546 117732
rect 278132 115376 280380 117740
rect 292062 115378 294310 117742
rect 305978 115380 308226 117744
rect 319812 115376 322060 117740
rect 333742 115378 335990 117742
rect 347658 115380 349906 117744
rect 194628 102952 196876 105316
rect 208558 102954 210806 105318
rect 222474 102956 224722 105320
rect 236314 102954 238562 105318
rect 250244 102956 252492 105320
rect 264160 102958 266408 105322
rect 277994 102966 280242 105330
rect 291924 102968 294172 105332
rect 305840 102970 308088 105334
rect 319674 102966 321922 105330
rect 333604 102968 335852 105332
rect 347520 102970 349768 105334
rect 277418 87250 279666 89614
rect 291348 87252 293596 89616
rect 305264 87254 307512 89618
rect 319098 87250 321346 89614
rect 333028 87252 335276 89616
rect 346944 87254 349192 89618
rect 277418 74662 279666 77026
rect 291348 74664 293596 77028
rect 305264 74666 307512 77030
rect 319098 74662 321346 77026
rect 333028 74664 335276 77028
rect 346944 74666 349192 77030
rect 277418 62074 279666 64438
rect 291348 62076 293596 64440
rect 305264 62078 307512 64442
rect 319098 62074 321346 64438
rect 333028 62076 335276 64440
rect 346944 62078 349192 64442
<< locali >>
rect 201278 666800 205076 670524
rect 282776 666800 286574 670524
rect 379924 666800 383722 670524
rect 189734 665796 214212 666800
rect 189734 665794 207956 665796
rect 189734 663430 194026 665794
rect 196274 663432 207956 665794
rect 210204 663432 214212 665796
rect 196274 663430 214212 663432
rect 189734 662586 214212 663430
rect 272354 665812 420906 666800
rect 272354 665810 305238 665812
rect 272354 665808 291322 665810
rect 272354 663444 277392 665808
rect 279640 663446 291322 665808
rect 293570 663448 305238 665810
rect 307486 665810 346918 665812
rect 307486 665808 333002 665810
rect 307486 663448 319072 665808
rect 293570 663446 319072 663448
rect 279640 663444 319072 663446
rect 321320 665726 333002 665808
rect 321320 663444 328962 665726
rect 272354 663376 328962 663444
rect 331494 663446 333002 665726
rect 335250 663448 346918 665810
rect 349166 665802 420906 665812
rect 349166 665800 388374 665802
rect 349166 665798 374458 665800
rect 349166 663448 360528 665798
rect 335250 663446 360528 663448
rect 331494 663434 360528 663446
rect 362776 663436 374458 665798
rect 376706 663438 388374 665800
rect 390622 665800 416144 665802
rect 390622 663438 402214 665800
rect 376706 663436 402214 663438
rect 404462 663438 416144 665800
rect 418392 663438 420906 665802
rect 404462 663436 420906 663438
rect 362776 663434 420906 663436
rect 331494 663376 420906 663434
rect 272354 662586 420906 663376
rect 201186 661298 205288 662586
rect 282776 661298 286844 662586
rect 201186 654144 205242 661298
rect 282788 655438 286844 661298
rect 282776 654144 286844 655438
rect 379772 661298 383842 662586
rect 379772 654144 383828 661298
rect 189734 653140 214212 654144
rect 189734 653138 208504 653140
rect 189734 650774 194574 653138
rect 196822 650776 208504 653138
rect 210752 650776 214212 653140
rect 196822 650774 214212 650776
rect 189734 649930 214212 650774
rect 272354 653156 420906 654144
rect 272354 653154 305786 653156
rect 272354 653152 291870 653154
rect 272354 650788 277940 653152
rect 280188 650790 291870 653152
rect 294118 650792 305786 653154
rect 308034 653154 347466 653156
rect 308034 653152 333550 653154
rect 308034 650792 319620 653152
rect 294118 650790 319620 650792
rect 280188 650788 319620 650790
rect 321868 652982 333550 653152
rect 321868 650788 329000 652982
rect 272354 650632 329000 650788
rect 331532 650790 333550 652982
rect 335798 650792 347466 653154
rect 349714 653146 420906 653156
rect 349714 653144 388922 653146
rect 349714 653142 375006 653144
rect 349714 650792 361076 653142
rect 335798 650790 361076 650792
rect 331532 650778 361076 650790
rect 363324 650780 375006 653142
rect 377254 650782 388922 653144
rect 391170 653144 416692 653146
rect 391170 650782 402762 653144
rect 377254 650780 402762 650782
rect 405010 650782 416692 653144
rect 418940 650782 420906 653146
rect 405010 650780 420906 650782
rect 363324 650778 420906 650780
rect 331532 650632 420906 650778
rect 272354 649930 420906 650632
rect 201186 639884 205242 649930
rect 282776 639884 286844 649930
rect 379772 639884 383828 649930
rect 189734 638880 214212 639884
rect 189734 638878 207956 638880
rect 189734 636514 194026 638878
rect 196274 636516 207956 638878
rect 210204 636516 214212 638880
rect 196274 636514 214212 636516
rect 189734 635670 214212 636514
rect 272354 638896 420906 639884
rect 272354 638894 305238 638896
rect 272354 638892 291322 638894
rect 272354 636528 277392 638892
rect 279640 636530 291322 638892
rect 293570 636532 305238 638894
rect 307486 638894 346918 638896
rect 307486 638892 333002 638894
rect 307486 636532 319072 638892
rect 293570 636530 319072 636532
rect 279640 636528 319072 636530
rect 321320 638810 333002 638892
rect 321320 636528 328962 638810
rect 272354 636460 328962 636528
rect 331494 636530 333002 638810
rect 335250 636532 346918 638894
rect 349166 638886 420906 638896
rect 349166 638884 388374 638886
rect 349166 638882 374458 638884
rect 349166 636532 360528 638882
rect 335250 636530 360528 636532
rect 331494 636518 360528 636530
rect 362776 636520 374458 638882
rect 376706 636522 388374 638884
rect 390622 638884 416144 638886
rect 390622 636522 402214 638884
rect 376706 636520 402214 636522
rect 404462 636522 416144 638884
rect 418392 636522 420906 638886
rect 404462 636520 420906 636522
rect 362776 636518 420906 636520
rect 331494 636460 420906 636518
rect 272354 635670 420906 636460
rect 201186 634382 205288 635670
rect 282776 634382 286844 635670
rect 201186 626002 205242 634382
rect 282788 626364 286844 634382
rect 379772 634382 383842 635670
rect 201290 625622 205088 626002
rect 282788 625622 286586 626364
rect 379772 626228 383828 634382
rect 379936 625622 383734 626228
rect 189734 624618 214212 625622
rect 189734 624616 208516 624618
rect 189734 622252 194586 624616
rect 196834 622254 208516 624616
rect 210764 622254 214212 624618
rect 196834 622252 214212 622254
rect 189734 621408 214212 622252
rect 272354 624634 420906 625622
rect 272354 624632 305798 624634
rect 272354 624630 291882 624632
rect 272354 622266 277952 624630
rect 280200 622268 291882 624630
rect 294130 622270 305798 624632
rect 308046 624632 347478 624634
rect 308046 624630 333562 624632
rect 308046 622270 319632 624630
rect 294130 622268 319632 622270
rect 280200 622266 319632 622268
rect 321880 624460 333562 624630
rect 321880 622266 329012 624460
rect 272354 622110 329012 622266
rect 331544 622268 333562 624460
rect 335810 622270 347478 624632
rect 349726 624624 420906 624634
rect 349726 624622 388934 624624
rect 349726 624620 375018 624622
rect 349726 622270 361088 624620
rect 335810 622268 361088 622270
rect 331544 622256 361088 622268
rect 363336 622258 375018 624620
rect 377266 622260 388934 624622
rect 391182 624622 416704 624624
rect 391182 622260 402774 624622
rect 377266 622258 402774 622260
rect 405022 622260 416704 624622
rect 418952 622260 420906 624624
rect 405022 622258 420906 622260
rect 363336 622256 420906 622258
rect 331544 622110 420906 622256
rect 272354 621408 420906 622110
rect 201290 611362 205088 621408
rect 282788 611362 286586 621408
rect 379936 611362 383734 621408
rect 157200 610398 420906 611362
rect 157200 610396 180402 610398
rect 157200 608032 166486 610396
rect 168734 608034 180402 610396
rect 182650 610374 420906 610398
rect 182650 610372 305250 610374
rect 182650 610370 291334 610372
rect 182650 610362 277404 610370
rect 182650 610360 263570 610362
rect 182650 610358 221884 610360
rect 182650 610356 207968 610358
rect 182650 608034 194038 610356
rect 168734 608032 194038 608034
rect 157200 607992 194038 608032
rect 196286 607994 207968 610356
rect 210216 607996 221884 610358
rect 224132 610358 249654 610360
rect 224132 607996 235724 610358
rect 210216 607994 235724 607996
rect 237972 607996 249654 610358
rect 251902 607998 263570 610360
rect 265818 608006 277404 610362
rect 279652 608008 291334 610370
rect 293582 608010 305250 610372
rect 307498 610372 346930 610374
rect 307498 610370 333014 610372
rect 307498 608010 319084 610370
rect 293582 608008 319084 608010
rect 279652 608006 319084 608008
rect 321332 610288 333014 610370
rect 321332 608006 328974 610288
rect 265818 607998 328974 608006
rect 251902 607996 328974 607998
rect 237972 607994 328974 607996
rect 196286 607992 328974 607994
rect 157200 607938 328974 607992
rect 331506 608008 333014 610288
rect 335262 608010 346930 610372
rect 349178 610364 420906 610374
rect 349178 610362 388386 610364
rect 349178 610360 374470 610362
rect 349178 608010 360540 610360
rect 335262 608008 360540 608010
rect 331506 607996 360540 608008
rect 362788 607998 374470 610360
rect 376718 608000 388386 610362
rect 390634 610362 416156 610364
rect 390634 608000 402226 610362
rect 376718 607998 402226 608000
rect 404474 608000 416156 610362
rect 418404 608000 420906 610364
rect 404474 607998 420906 608000
rect 362788 607996 420906 607998
rect 331506 607938 420906 607996
rect 157200 607148 420906 607938
rect 201290 605506 205300 607148
rect 282788 605506 286824 607148
rect 201372 593334 205300 605506
rect 282896 593472 286824 605506
rect 379926 594198 383854 607148
rect 379926 593540 383912 594198
rect 201468 592904 205266 593334
rect 282966 592904 286764 593472
rect 380114 592904 383912 593540
rect 189988 591900 215998 592904
rect 189988 591898 208694 591900
rect 189988 589534 194764 591898
rect 197012 589536 208694 591898
rect 210942 589536 215998 591900
rect 197012 589534 215998 589536
rect 189988 588690 215998 589534
rect 272354 591916 340950 592904
rect 272354 591914 305976 591916
rect 272354 591912 292060 591914
rect 272354 589548 278130 591912
rect 280378 589550 292060 591912
rect 294308 589552 305976 591914
rect 308224 591914 340950 591916
rect 308224 591912 333740 591914
rect 308224 589552 319810 591912
rect 294308 589550 319810 589552
rect 280378 589548 319810 589550
rect 322058 591742 333740 591912
rect 322058 589548 329190 591742
rect 272354 589392 329190 589548
rect 331722 589550 333740 591742
rect 335988 589550 340950 591914
rect 331722 589392 340950 589550
rect 272354 588690 340950 589392
rect 366450 591906 395520 592904
rect 366450 591904 389112 591906
rect 366450 589540 375196 591904
rect 377444 589542 389112 591904
rect 391360 589542 395520 591906
rect 377444 589540 395520 589542
rect 366450 588690 395520 589540
rect 201468 578644 205266 588690
rect 282966 578644 286764 588690
rect 380114 578644 383912 588690
rect 189988 577640 215998 578644
rect 189988 577638 208146 577640
rect 189988 575274 194216 577638
rect 196464 575276 208146 577638
rect 210394 575276 215998 577640
rect 196464 575274 215998 575276
rect 189988 574430 215998 575274
rect 272354 577656 340950 578644
rect 272354 577654 305428 577656
rect 272354 577652 291512 577654
rect 272354 575288 277582 577652
rect 279830 575290 291512 577652
rect 293760 575292 305428 577654
rect 307676 577654 340950 577656
rect 307676 577652 333192 577654
rect 307676 575292 319262 577652
rect 293760 575290 319262 575292
rect 279830 575288 319262 575290
rect 321510 577570 333192 577652
rect 321510 575288 329152 577570
rect 272354 575220 329152 575288
rect 331684 575290 333192 577570
rect 335440 575290 340950 577654
rect 331684 575220 340950 575290
rect 272354 574430 340950 575220
rect 366450 577646 395520 578644
rect 366450 577644 388564 577646
rect 366450 575280 374648 577644
rect 376896 575282 388564 577644
rect 390812 575282 395520 577646
rect 376896 575280 395520 575282
rect 366450 574430 395520 575280
rect 201468 565818 205266 574430
rect 282966 565818 286764 574430
rect 380114 565818 383912 574430
rect 189988 564814 215998 565818
rect 189988 564812 208362 564814
rect 189988 562448 194432 564812
rect 196680 562450 208362 564812
rect 210610 562450 215998 564814
rect 196680 562448 215998 562450
rect 189988 561604 215998 562448
rect 272354 564830 340950 565818
rect 272354 564828 305644 564830
rect 272354 564826 291728 564828
rect 272354 562462 277798 564826
rect 280046 562464 291728 564826
rect 293976 562466 305644 564828
rect 307892 564828 340950 564830
rect 307892 564826 333408 564828
rect 307892 562466 319478 564826
rect 293976 562464 319478 562466
rect 280046 562462 319478 562464
rect 321726 564766 333408 564826
rect 321726 562462 329078 564766
rect 272354 562416 329078 562462
rect 331610 562464 333408 564766
rect 335656 562464 340950 564828
rect 331610 562416 340950 562464
rect 272354 561604 340950 562416
rect 366450 564820 395520 565818
rect 366450 564818 388780 564820
rect 366450 562454 374864 564818
rect 377112 562456 388780 564818
rect 391028 562456 395520 564820
rect 377112 562454 395520 562456
rect 366450 561604 395520 562454
rect 200654 548088 205408 561604
rect 282178 548088 286932 561604
rect 378922 549382 383676 561604
rect 378922 548088 384014 549382
rect 188536 547100 420906 548088
rect 188536 547098 306078 547100
rect 188536 547096 292162 547098
rect 188536 547088 278232 547096
rect 188536 547086 264398 547088
rect 188536 547084 222712 547086
rect 188536 547082 208796 547084
rect 188536 544718 194866 547082
rect 197114 544720 208796 547082
rect 211044 544722 222712 547084
rect 224960 547084 250482 547086
rect 224960 544722 236552 547084
rect 211044 544720 236552 544722
rect 238800 544722 250482 547084
rect 252730 544724 264398 547086
rect 266646 544732 278232 547088
rect 280480 544734 292162 547096
rect 294410 544736 306078 547098
rect 308326 547098 347758 547100
rect 308326 547096 333842 547098
rect 308326 544736 319912 547096
rect 294410 544734 319912 544736
rect 280480 544732 319912 544734
rect 322160 546926 333842 547096
rect 322160 544732 329292 546926
rect 266646 544724 329292 544732
rect 252730 544722 329292 544724
rect 238800 544720 329292 544722
rect 197114 544718 329292 544720
rect 188536 544576 329292 544718
rect 331824 544734 333842 546926
rect 336090 544736 347758 547098
rect 350006 547090 420906 547100
rect 350006 547088 389214 547090
rect 350006 547086 375298 547088
rect 350006 544736 361368 547086
rect 336090 544734 361368 544736
rect 331824 544722 361368 544734
rect 363616 544724 375298 547086
rect 377546 544726 389214 547088
rect 391462 547088 416984 547090
rect 391462 544726 403054 547088
rect 377546 544724 403054 544726
rect 405302 544726 416984 547088
rect 419232 544726 420906 547090
rect 405302 544724 420906 544726
rect 363616 544722 420906 544724
rect 331824 544576 420906 544722
rect 188536 543874 420906 544576
rect 201570 533828 205368 543874
rect 283068 533828 286866 543874
rect 380216 533828 384014 543874
rect 188536 532840 420906 533828
rect 188536 532838 305530 532840
rect 188536 532836 291614 532838
rect 188536 532828 277684 532836
rect 188536 532826 263850 532828
rect 188536 532824 222164 532826
rect 188536 532822 208248 532824
rect 188536 530458 194318 532822
rect 196566 530460 208248 532822
rect 210496 530462 222164 532824
rect 224412 532824 249934 532826
rect 224412 530462 236004 532824
rect 210496 530460 236004 530462
rect 238252 530462 249934 532824
rect 252182 530464 263850 532826
rect 266098 530472 277684 532828
rect 279932 530474 291614 532836
rect 293862 530476 305530 532838
rect 307778 532838 347210 532840
rect 307778 532836 333294 532838
rect 307778 530476 319364 532836
rect 293862 530474 319364 530476
rect 279932 530472 319364 530474
rect 321612 532754 333294 532836
rect 321612 530472 329254 532754
rect 266098 530464 329254 530472
rect 252182 530462 329254 530464
rect 238252 530460 329254 530462
rect 196566 530458 329254 530460
rect 188536 530404 329254 530458
rect 331786 530474 333294 532754
rect 335542 530476 347210 532838
rect 349458 532830 420906 532840
rect 349458 532828 388666 532830
rect 349458 532826 374750 532828
rect 349458 530476 360820 532826
rect 335542 530474 360820 530476
rect 331786 530462 360820 530474
rect 363068 530464 374750 532826
rect 376998 530466 388666 532828
rect 390914 532828 416436 532830
rect 390914 530466 402506 532828
rect 376998 530464 402506 530466
rect 404754 530466 416436 532828
rect 418684 530466 420906 532830
rect 404754 530464 420906 530466
rect 363068 530462 420906 530464
rect 331786 530404 420906 530462
rect 188536 529614 420906 530404
rect 201570 521002 205368 529614
rect 283068 521002 286866 529614
rect 380216 521002 384014 529614
rect 188536 520014 420906 521002
rect 188536 520012 305746 520014
rect 188536 520010 291830 520012
rect 188536 520002 277900 520010
rect 188536 520000 264066 520002
rect 188536 519998 222380 520000
rect 188536 519996 208464 519998
rect 188536 517632 194534 519996
rect 196782 517634 208464 519996
rect 210712 517636 222380 519998
rect 224628 519998 250150 520000
rect 224628 517636 236220 519998
rect 210712 517634 236220 517636
rect 238468 517636 250150 519998
rect 252398 517638 264066 520000
rect 266314 517646 277900 520002
rect 280148 517648 291830 520010
rect 294078 517650 305746 520012
rect 307994 520012 347426 520014
rect 307994 520010 333510 520012
rect 307994 517650 319580 520010
rect 294078 517648 319580 517650
rect 280148 517646 319580 517648
rect 321828 519950 333510 520010
rect 321828 517646 329180 519950
rect 266314 517638 329180 517646
rect 252398 517636 329180 517638
rect 238468 517634 329180 517636
rect 196782 517632 329180 517634
rect 188536 517600 329180 517632
rect 331712 517648 333510 519950
rect 335758 517650 347426 520012
rect 349674 520004 420906 520014
rect 349674 520002 388882 520004
rect 349674 520000 374966 520002
rect 349674 517650 361036 520000
rect 335758 517648 361036 517650
rect 331712 517636 361036 517648
rect 363284 517638 374966 520000
rect 377214 517640 388882 520002
rect 391130 520002 416652 520004
rect 391130 517640 402722 520002
rect 377214 517638 402722 517640
rect 404970 517640 416652 520002
rect 418900 517640 420906 520004
rect 404970 517638 420906 517640
rect 363284 517636 420906 517638
rect 331712 517600 420906 517636
rect 188536 516788 420906 517600
rect 200894 515642 205602 516788
rect 282636 515642 287026 516788
rect 201496 500154 205602 515642
rect 282920 500192 287026 515642
rect 379184 500874 383956 516788
rect 201632 499580 205430 500154
rect 283130 499580 286928 500192
rect 379184 499580 384076 500874
rect 190616 498592 420906 499580
rect 190616 498590 306140 498592
rect 190616 498588 292224 498590
rect 190616 498580 278294 498588
rect 190616 498578 264460 498580
rect 190616 498576 222774 498578
rect 190616 498574 208858 498576
rect 190616 496210 194928 498574
rect 197176 496212 208858 498574
rect 211106 496214 222774 498576
rect 225022 498576 250544 498578
rect 225022 496214 236614 498576
rect 211106 496212 236614 496214
rect 238862 496214 250544 498576
rect 252792 496216 264460 498578
rect 266708 496224 278294 498580
rect 280542 496226 292224 498588
rect 294472 496228 306140 498590
rect 308388 498590 347820 498592
rect 308388 498588 333904 498590
rect 308388 496228 319974 498588
rect 294472 496226 319974 496228
rect 280542 496224 319974 496226
rect 322222 498418 333904 498588
rect 322222 496224 329354 498418
rect 266708 496216 329354 496224
rect 252792 496214 329354 496216
rect 238862 496212 329354 496214
rect 197176 496210 329354 496212
rect 190616 496068 329354 496210
rect 331886 496226 333904 498418
rect 336152 496228 347820 498590
rect 350068 498582 420906 498592
rect 350068 498580 389276 498582
rect 350068 498578 375360 498580
rect 350068 496228 361430 498578
rect 336152 496226 361430 496228
rect 331886 496214 361430 496226
rect 363678 496216 375360 498578
rect 377608 496218 389276 498580
rect 391524 498580 417046 498582
rect 391524 496218 403116 498580
rect 377608 496216 403116 496218
rect 405364 496218 417046 498580
rect 419294 496218 420906 498582
rect 405364 496216 420906 496218
rect 363678 496214 420906 496216
rect 331886 496068 420906 496214
rect 190616 495366 420906 496068
rect 201632 485320 205430 495366
rect 283130 485320 286928 495366
rect 380278 485320 384076 495366
rect 190234 484332 420906 485320
rect 190234 484330 305592 484332
rect 190234 484328 291676 484330
rect 190234 484320 277746 484328
rect 190234 484318 263912 484320
rect 190234 484316 222226 484318
rect 190234 484314 208310 484316
rect 190234 481950 194380 484314
rect 196628 481952 208310 484314
rect 210558 481954 222226 484316
rect 224474 484316 249996 484318
rect 224474 481954 236066 484316
rect 210558 481952 236066 481954
rect 238314 481954 249996 484316
rect 252244 481956 263912 484318
rect 266160 481964 277746 484320
rect 279994 481966 291676 484328
rect 293924 481968 305592 484330
rect 307840 484330 347272 484332
rect 307840 484328 333356 484330
rect 307840 481968 319426 484328
rect 293924 481966 319426 481968
rect 279994 481964 319426 481966
rect 321674 484246 333356 484328
rect 321674 481964 329316 484246
rect 266160 481956 329316 481964
rect 252244 481954 329316 481956
rect 238314 481952 329316 481954
rect 196628 481950 329316 481952
rect 190234 481896 329316 481950
rect 331848 481966 333356 484246
rect 335604 481968 347272 484330
rect 349520 484322 420906 484332
rect 349520 484320 388728 484322
rect 349520 484318 374812 484320
rect 349520 481968 360882 484318
rect 335604 481966 360882 481968
rect 331848 481954 360882 481966
rect 363130 481956 374812 484318
rect 377060 481958 388728 484320
rect 390976 484320 416498 484322
rect 390976 481958 402568 484320
rect 377060 481956 402568 481958
rect 404816 481958 416498 484320
rect 418746 481958 420906 484322
rect 404816 481956 420906 481958
rect 363130 481954 420906 481956
rect 331848 481896 420906 481954
rect 190234 481106 420906 481896
rect 201632 472494 205430 481106
rect 283130 472494 286928 481106
rect 380278 472494 384076 481106
rect 190234 471506 420906 472494
rect 190234 471504 305808 471506
rect 190234 471502 291892 471504
rect 190234 471494 277962 471502
rect 190234 471492 264128 471494
rect 190234 471490 222442 471492
rect 190234 471488 208526 471490
rect 190234 469124 194596 471488
rect 196844 469126 208526 471488
rect 210774 469128 222442 471490
rect 224690 471490 250212 471492
rect 224690 469128 236282 471490
rect 210774 469126 236282 469128
rect 238530 469128 250212 471490
rect 252460 469130 264128 471492
rect 266376 469138 277962 471494
rect 280210 469140 291892 471502
rect 294140 469142 305808 471504
rect 308056 471504 347488 471506
rect 308056 471502 333572 471504
rect 308056 469142 319642 471502
rect 294140 469140 319642 469142
rect 280210 469138 319642 469140
rect 321890 471442 333572 471502
rect 321890 469138 329242 471442
rect 266376 469130 329242 469138
rect 252460 469128 329242 469130
rect 238530 469126 329242 469128
rect 196844 469124 329242 469126
rect 190234 469092 329242 469124
rect 331774 469140 333572 471442
rect 335820 469142 347488 471504
rect 349736 471496 420906 471506
rect 349736 471494 388944 471496
rect 349736 471492 375028 471494
rect 349736 469142 361098 471492
rect 335820 469140 361098 469142
rect 331774 469128 361098 469140
rect 363346 469130 375028 471492
rect 377276 469132 388944 471494
rect 391192 471494 416714 471496
rect 391192 469132 402784 471494
rect 377276 469130 402784 469132
rect 405032 469132 416714 471494
rect 418962 469132 420906 471496
rect 405032 469130 420906 469132
rect 363346 469128 420906 469130
rect 331774 469092 420906 469128
rect 190234 468280 420906 469092
rect 200956 467134 205700 468280
rect 282698 467134 286972 468280
rect 201866 460380 205700 467134
rect 201880 459048 205678 460380
rect 282826 459090 286972 467134
rect 379234 467134 383548 468280
rect 282826 459048 287176 459090
rect 379234 459048 383380 467134
rect 190234 459006 383380 459048
rect 384550 459006 420906 459048
rect 190234 458060 420906 459006
rect 190234 458058 306388 458060
rect 190234 458056 292472 458058
rect 190234 458048 278542 458056
rect 190234 458046 264708 458048
rect 190234 458044 223022 458046
rect 190234 458042 209106 458044
rect 190234 455678 195176 458042
rect 197424 455680 209106 458042
rect 211354 455682 223022 458044
rect 225270 458044 250792 458046
rect 225270 455682 236862 458044
rect 211354 455680 236862 455682
rect 239110 455682 250792 458044
rect 253040 455684 264708 458046
rect 266956 455692 278542 458048
rect 280790 455694 292472 458056
rect 294720 455696 306388 458058
rect 308636 458058 348068 458060
rect 308636 458056 334152 458058
rect 308636 455696 320222 458056
rect 294720 455694 320222 455696
rect 280790 455692 320222 455694
rect 322470 457886 334152 458056
rect 322470 455692 329602 457886
rect 266956 455684 329602 455692
rect 253040 455682 329602 455684
rect 239110 455680 329602 455682
rect 197424 455678 329602 455680
rect 190234 455536 329602 455678
rect 332134 455694 334152 457886
rect 336400 455696 348068 458058
rect 350316 458050 420906 458060
rect 350316 458048 389524 458050
rect 350316 458046 375608 458048
rect 350316 455696 361678 458046
rect 336400 455694 361678 455696
rect 332134 455682 361678 455694
rect 363926 455684 375608 458046
rect 377856 455686 389524 458048
rect 391772 458048 417294 458050
rect 391772 455686 403364 458048
rect 377856 455684 403364 455686
rect 405612 455686 417294 458048
rect 419542 455686 420906 458050
rect 405612 455684 420906 455686
rect 363926 455682 420906 455684
rect 332134 455536 420906 455682
rect 190234 454834 420906 455536
rect 201768 453774 205678 454834
rect 283378 453774 287308 454834
rect 201768 447324 205672 453774
rect 283404 449552 287308 453774
rect 283338 447324 287308 449552
rect 380358 453774 384324 454834
rect 380358 449552 384262 453774
rect 380358 447324 384284 449552
rect 190234 446336 420906 447324
rect 190234 446334 306348 446336
rect 190234 446332 292432 446334
rect 190234 446324 278502 446332
rect 190234 446322 264668 446324
rect 190234 446320 222982 446322
rect 190234 446318 209066 446320
rect 190234 443954 195136 446318
rect 197384 443956 209066 446318
rect 211314 443958 222982 446320
rect 225230 446320 250752 446322
rect 225230 443958 236822 446320
rect 211314 443956 236822 443958
rect 239070 443958 250752 446320
rect 253000 443960 264668 446322
rect 266916 443968 278502 446324
rect 280750 443970 292432 446332
rect 294680 443972 306348 446334
rect 308596 446334 348028 446336
rect 308596 446332 334112 446334
rect 308596 443972 320182 446332
rect 294680 443970 320182 443972
rect 280750 443968 320182 443970
rect 322430 446162 334112 446332
rect 322430 443968 329562 446162
rect 266916 443960 329562 443968
rect 253000 443958 329562 443960
rect 239070 443956 329562 443958
rect 197384 443954 329562 443956
rect 190234 443812 329562 443954
rect 332094 443970 334112 446162
rect 336360 443972 348028 446334
rect 350276 446326 420906 446336
rect 350276 446324 389484 446326
rect 350276 446322 375568 446324
rect 350276 443972 361638 446322
rect 336360 443970 361638 443972
rect 332094 443958 361638 443970
rect 363886 443960 375568 446322
rect 377816 443962 389484 446324
rect 391732 446324 417254 446326
rect 391732 443962 403324 446324
rect 377816 443960 403324 443962
rect 405572 443962 417254 446324
rect 419502 443962 420906 446326
rect 405572 443960 420906 443962
rect 363886 443958 420906 443960
rect 332094 443812 420906 443958
rect 190234 443110 420906 443812
rect 201768 426590 205672 443110
rect 283338 442050 287308 443110
rect 201768 425338 205718 426590
rect 188884 423198 193354 423314
rect 201920 423198 205718 425338
rect 283404 424954 287308 442050
rect 380358 442050 384284 443110
rect 380358 433602 384262 442050
rect 283418 423198 287216 424954
rect 188884 422194 217042 423198
rect 188884 422192 209146 422194
rect 188884 419828 195216 422192
rect 197464 419830 209146 422192
rect 211394 419830 217042 422194
rect 197464 419828 217042 419830
rect 188884 419116 217042 419828
rect 189818 418984 217042 419116
rect 272496 422210 341056 423198
rect 272496 422208 306428 422210
rect 272496 422206 292512 422208
rect 272496 419842 278582 422206
rect 280830 419844 292512 422206
rect 294760 419846 306428 422208
rect 308676 422208 341056 422210
rect 308676 422206 334192 422208
rect 308676 419846 320262 422206
rect 294760 419844 320262 419846
rect 280830 419842 320262 419844
rect 322510 422036 334192 422206
rect 322510 419842 329642 422036
rect 272496 419686 329642 419842
rect 332174 419844 334192 422036
rect 336440 419844 341056 422208
rect 332174 419686 341056 419844
rect 272496 418984 341056 419686
rect 201920 408938 205718 418984
rect 283418 408938 287216 418984
rect 189818 407934 217042 408938
rect 189818 407932 208598 407934
rect 189818 405568 194668 407932
rect 196916 405570 208598 407932
rect 210846 405570 217042 407934
rect 196916 405568 217042 405570
rect 189818 404724 217042 405568
rect 272496 407950 341056 408938
rect 272496 407948 305880 407950
rect 272496 407946 291964 407948
rect 272496 405582 278034 407946
rect 280282 405584 291964 407946
rect 294212 405586 305880 407948
rect 308128 407948 341056 407950
rect 308128 407946 333644 407948
rect 308128 405586 319714 407946
rect 294212 405584 319714 405586
rect 280282 405582 319714 405584
rect 321962 407864 333644 407946
rect 321962 405582 329604 407864
rect 272496 405514 329604 405582
rect 332136 405584 333644 407864
rect 335892 405584 341056 407948
rect 332136 405514 341056 405584
rect 272496 404724 341056 405514
rect 201920 396112 205718 404724
rect 283418 396112 287216 404724
rect 189818 395108 217042 396112
rect 189818 395106 208814 395108
rect 189818 392742 194884 395106
rect 197132 392744 208814 395106
rect 211062 392744 217042 395108
rect 197132 392742 217042 392744
rect 189818 391898 217042 392742
rect 272496 395124 341056 396112
rect 272496 395122 306096 395124
rect 272496 395120 292180 395122
rect 272496 392756 278250 395120
rect 280498 392758 292180 395120
rect 294428 392760 306096 395122
rect 308344 395122 341056 395124
rect 308344 395120 333860 395122
rect 308344 392760 319930 395120
rect 294428 392758 319930 392760
rect 280498 392756 319930 392758
rect 322178 395060 333860 395120
rect 322178 392756 329530 395060
rect 272496 392710 329530 392756
rect 332062 392758 333860 395060
rect 336108 392758 341056 395122
rect 332062 392710 341056 392758
rect 272496 391898 341056 392710
rect 201244 389352 205424 391898
rect 282986 389352 287166 391898
rect 201244 387412 205692 389352
rect 282986 387412 287190 389352
rect 189818 386408 217042 387412
rect 189818 386406 209120 386408
rect 189818 384042 195190 386406
rect 197438 384044 209120 386406
rect 211368 384044 217042 386408
rect 197438 384042 217042 384044
rect 189818 383198 217042 384042
rect 272496 386424 341056 387412
rect 272496 386422 306402 386424
rect 272496 386420 292486 386422
rect 272496 384056 278556 386420
rect 280804 384058 292486 386420
rect 294734 384060 306402 386422
rect 308650 386422 341056 386424
rect 308650 386420 334166 386422
rect 308650 384060 320236 386420
rect 294734 384058 320236 384060
rect 280804 384056 320236 384058
rect 322484 386250 334166 386420
rect 322484 384056 329616 386250
rect 272496 383900 329616 384056
rect 332148 384058 334166 386250
rect 336414 384058 341056 386422
rect 332148 383900 341056 384058
rect 272496 383198 341056 383900
rect 201894 377648 205692 383198
rect 283392 373152 287190 383198
rect 380240 379726 384302 433602
rect 380240 377816 384338 379726
rect 380540 373152 384338 377816
rect 272496 372164 394636 373152
rect 272496 372162 305854 372164
rect 272496 372160 291938 372162
rect 272496 369796 278008 372160
rect 280256 369798 291938 372160
rect 294186 369800 305854 372162
rect 308102 372162 347534 372164
rect 308102 372160 333618 372162
rect 308102 369800 319688 372160
rect 294186 369798 319688 369800
rect 280256 369796 319688 369798
rect 321936 372078 333618 372160
rect 321936 369796 329578 372078
rect 272496 369728 329578 369796
rect 332110 369798 333618 372078
rect 335866 369800 347534 372162
rect 349782 372154 394636 372164
rect 349782 372152 388990 372154
rect 349782 372150 375074 372152
rect 349782 369800 361144 372150
rect 335866 369798 361144 369800
rect 332110 369786 361144 369798
rect 363392 369788 375074 372150
rect 377322 369790 388990 372152
rect 391238 369790 394636 372154
rect 377322 369788 394636 369790
rect 363392 369786 394636 369788
rect 332110 369728 394636 369786
rect 272496 368938 394636 369728
rect 283392 360326 287190 368938
rect 380540 360326 384338 368938
rect 218664 359338 394636 360326
rect 218664 359336 306070 359338
rect 218664 359334 292154 359336
rect 218664 359326 278224 359334
rect 218664 359324 264390 359326
rect 218664 356960 222704 359324
rect 224952 359322 250474 359324
rect 224952 356960 236544 359322
rect 218664 356958 236544 356960
rect 238792 356960 250474 359322
rect 252722 356962 264390 359324
rect 266638 356970 278224 359326
rect 280472 356972 292154 359334
rect 294402 356974 306070 359336
rect 308318 359336 347750 359338
rect 308318 359334 333834 359336
rect 308318 356974 319904 359334
rect 294402 356972 319904 356974
rect 280472 356970 319904 356972
rect 322152 359274 333834 359334
rect 322152 356970 329504 359274
rect 266638 356962 329504 356970
rect 252722 356960 329504 356962
rect 238792 356958 329504 356960
rect 218664 356924 329504 356958
rect 332036 356972 333834 359274
rect 336082 356974 347750 359336
rect 349998 359328 394636 359338
rect 349998 359326 389206 359328
rect 349998 359324 375290 359326
rect 349998 356974 361360 359324
rect 336082 356972 361360 356974
rect 332036 356960 361360 356972
rect 363608 356962 375290 359324
rect 377538 356964 389206 359326
rect 391454 356964 394636 359328
rect 377538 356962 394636 356964
rect 363608 356960 394636 356962
rect 332036 356924 394636 356960
rect 218664 356112 394636 356924
rect 282924 348498 287236 356112
rect 379630 352716 384084 356112
rect 379772 348498 384084 352716
rect 216570 347510 394636 348498
rect 216570 347508 305500 347510
rect 216570 347506 291584 347508
rect 216570 347498 277654 347506
rect 216570 347496 263820 347498
rect 216570 345132 222134 347496
rect 224382 347494 249904 347496
rect 224382 345132 235974 347494
rect 216570 345130 235974 345132
rect 238222 345132 249904 347494
rect 252152 345134 263820 347496
rect 266068 345142 277654 347498
rect 279902 345144 291584 347506
rect 293832 345146 305500 347508
rect 307748 347508 347180 347510
rect 307748 347506 333264 347508
rect 307748 345146 319334 347506
rect 293832 345144 319334 345146
rect 279902 345142 319334 345144
rect 321582 347424 333264 347506
rect 321582 345142 329224 347424
rect 266068 345134 329224 345142
rect 252152 345132 329224 345134
rect 238222 345130 329224 345132
rect 216570 345074 329224 345130
rect 331756 345144 333264 347424
rect 335512 345146 347180 347508
rect 349428 347500 394636 347510
rect 349428 347498 388636 347500
rect 349428 347496 374720 347498
rect 349428 345146 360790 347496
rect 335512 345144 360790 345146
rect 331756 345132 360790 345144
rect 363038 345134 374720 347496
rect 376968 345136 388636 347498
rect 390884 345136 394636 347500
rect 376968 345134 394636 345136
rect 363038 345132 394636 345134
rect 331756 345074 394636 345132
rect 216570 344284 394636 345074
rect 282924 335672 287236 344284
rect 379772 335672 384084 344284
rect 216570 334684 394636 335672
rect 216570 334682 305716 334684
rect 216570 334680 291800 334682
rect 216570 334672 277870 334680
rect 216570 334670 264036 334672
rect 216570 332306 222350 334670
rect 224598 334668 250120 334670
rect 224598 332306 236190 334668
rect 216570 332304 236190 332306
rect 238438 332306 250120 334668
rect 252368 332308 264036 334670
rect 266284 332316 277870 334672
rect 280118 332318 291800 334680
rect 294048 332320 305716 334682
rect 307964 334682 347396 334684
rect 307964 334680 333480 334682
rect 307964 332320 319550 334680
rect 294048 332318 319550 332320
rect 280118 332316 319550 332318
rect 321798 334620 333480 334680
rect 321798 332316 329150 334620
rect 266284 332308 329150 332316
rect 252368 332306 329150 332308
rect 238438 332304 329150 332306
rect 216570 332270 329150 332304
rect 331682 332318 333480 334620
rect 335728 332320 347396 334682
rect 349644 334674 394636 334684
rect 349644 334672 388852 334674
rect 349644 334670 374936 334672
rect 349644 332320 361006 334670
rect 335728 332318 361006 332320
rect 331682 332306 361006 332318
rect 363254 332308 374936 334670
rect 377184 332310 388852 334672
rect 391100 332310 394636 334674
rect 377184 332308 394636 332310
rect 363254 332306 394636 332308
rect 331682 332270 394636 332306
rect 216570 331458 394636 332270
rect 200864 329970 205660 330792
rect 282606 329970 287236 331458
rect 379276 329970 384084 331458
rect 201348 320994 205660 329970
rect 282924 320994 287236 329970
rect 379772 322536 384084 329970
rect 190322 319990 217042 320994
rect 190322 319988 209968 319990
rect 190322 317624 196038 319988
rect 198286 317626 209968 319988
rect 212216 317626 217042 319990
rect 198286 317624 217042 317626
rect 190322 316780 217042 317624
rect 273502 320976 287236 320994
rect 288504 320976 343072 320994
rect 273502 320098 343072 320976
rect 273502 320006 329682 320098
rect 273502 320004 307250 320006
rect 273502 320002 293334 320004
rect 273502 317638 279404 320002
rect 281652 317640 293334 320002
rect 295582 317642 307250 320004
rect 309498 320002 329682 320006
rect 309498 317642 321084 320002
rect 295582 317640 321084 317642
rect 281652 317638 321084 317640
rect 323332 317748 329682 320002
rect 332214 320004 343072 320098
rect 332214 317748 335014 320004
rect 323332 317640 335014 317748
rect 337262 317640 343072 320004
rect 323332 317638 343072 317640
rect 273502 316780 343072 317638
rect 202180 316650 206540 316780
rect 282924 316752 288038 316780
rect 283526 316650 288038 316752
rect 202180 311328 206206 316650
rect 283526 311328 287552 316650
rect 190322 310324 217042 311328
rect 190322 310322 210538 310324
rect 190322 307958 196608 310322
rect 198856 307960 210538 310322
rect 212786 307960 217042 310324
rect 198856 307958 217042 307960
rect 190322 307114 217042 307958
rect 273502 310418 343072 311328
rect 273502 310340 329644 310418
rect 273502 310338 307820 310340
rect 273502 310336 293904 310338
rect 273502 307972 279974 310336
rect 282222 307974 293904 310336
rect 296152 307976 307820 310338
rect 310068 310336 329644 310340
rect 310068 307976 321654 310336
rect 296152 307974 321654 307976
rect 282222 307972 321654 307974
rect 323902 308068 329644 310336
rect 332176 310338 343072 310418
rect 332176 308068 335584 310338
rect 323902 307974 335584 308068
rect 337832 307974 343072 310338
rect 323902 307972 343072 307974
rect 273502 307114 343072 307972
rect 202180 306984 207110 307114
rect 283526 306984 288608 307114
rect 202180 300808 206206 306984
rect 283526 300808 287552 306984
rect 190322 299804 217042 300808
rect 190322 299802 210680 299804
rect 190322 297438 196750 299802
rect 198998 297440 210680 299802
rect 212928 297440 217042 299804
rect 198998 297438 217042 297440
rect 190322 296594 217042 297438
rect 273502 299878 343072 300808
rect 273502 299820 329606 299878
rect 273502 299818 307962 299820
rect 273502 299816 294046 299818
rect 273502 297452 280116 299816
rect 282364 297454 294046 299816
rect 296294 297456 307962 299818
rect 310210 299816 329606 299820
rect 310210 297456 321796 299816
rect 296294 297454 321796 297456
rect 282364 297452 321796 297454
rect 324044 297528 329606 299816
rect 332138 299818 343072 299878
rect 332138 297528 335726 299818
rect 324044 297454 335726 297528
rect 337974 297454 343072 299818
rect 324044 297452 343072 297454
rect 273502 296594 343072 297452
rect 202180 296464 207252 296594
rect 283526 296464 288750 296594
rect 202180 289860 206206 296464
rect 283526 289860 287552 296464
rect 190322 288856 217042 289860
rect 190322 288854 210538 288856
rect 190322 286490 196608 288854
rect 198856 286492 210538 288854
rect 212786 286492 217042 288856
rect 198856 286490 217042 286492
rect 190322 285646 217042 286490
rect 273502 288872 343072 289860
rect 273502 288870 307820 288872
rect 273502 288868 293904 288870
rect 273502 286504 279974 288868
rect 282222 286506 293904 288868
rect 296152 286508 307820 288870
rect 310068 288870 343072 288872
rect 310068 288868 335584 288870
rect 310068 286508 321654 288868
rect 296152 286506 321654 286508
rect 282222 286504 321654 286506
rect 323902 288774 335584 288868
rect 323902 286504 329570 288774
rect 273502 286424 329570 286504
rect 332102 286506 335584 288774
rect 337832 286506 343072 288870
rect 332102 286424 343072 286506
rect 273502 285646 343072 286424
rect 202180 285516 207110 285646
rect 283526 285516 288608 285646
rect 202180 277636 206206 285516
rect 283526 277636 287552 285516
rect 190322 276632 217042 277636
rect 190322 276630 210822 276632
rect 190322 274266 196892 276630
rect 199140 274268 210822 276630
rect 213070 274268 217042 276632
rect 199140 274266 217042 274268
rect 190322 273422 217042 274266
rect 273502 276648 343072 277636
rect 273502 276646 308104 276648
rect 273502 276644 294188 276646
rect 273502 274280 280258 276644
rect 282506 274282 294188 276644
rect 296436 274284 308104 276646
rect 310352 276646 343072 276648
rect 310352 276644 335868 276646
rect 310352 274284 321938 276644
rect 296436 274282 321938 274284
rect 282506 274280 321938 274282
rect 324186 276394 335868 276644
rect 324186 274280 329570 276394
rect 273502 274044 329570 274280
rect 332102 274282 335868 276394
rect 338116 274282 343072 276646
rect 332102 274044 343072 274282
rect 273502 273422 343072 274044
rect 202180 273292 207394 273422
rect 283526 273292 288892 273422
rect 202180 261888 206206 273292
rect 283526 261888 287552 273292
rect 189722 260900 341180 261888
rect 189722 260898 307684 260900
rect 189722 260896 293768 260898
rect 189722 260888 279838 260896
rect 189722 260886 266004 260888
rect 189722 260884 224318 260886
rect 189722 260882 210402 260884
rect 189722 258518 196472 260882
rect 198720 258520 210402 260882
rect 212650 258522 224318 260884
rect 226566 260884 252088 260886
rect 226566 258522 238158 260884
rect 212650 258520 238158 258522
rect 240406 258522 252088 260884
rect 254336 258524 266004 260886
rect 268252 258532 279838 260888
rect 282086 258534 293768 260896
rect 296016 258536 307684 260898
rect 309932 260898 341180 260900
rect 309932 260896 335448 260898
rect 309932 258536 321518 260896
rect 296016 258534 321518 258536
rect 282086 258532 321518 258534
rect 323766 258534 335448 260896
rect 337696 258534 341180 260898
rect 323766 258532 341180 258534
rect 268252 258524 341180 258532
rect 254336 258522 341180 258524
rect 240406 258520 341180 258522
rect 198720 258518 341180 258520
rect 189722 257674 341180 258518
rect 202180 257544 206974 257674
rect 283526 257544 288472 257674
rect 202180 239256 206206 257544
rect 283526 239256 287552 257544
rect 192302 238252 215530 239256
rect 192302 238250 209436 238252
rect 192302 235886 195506 238250
rect 197754 235888 209436 238250
rect 211684 235888 215530 238252
rect 197754 235886 215530 235888
rect 192302 235042 215530 235886
rect 276024 238268 342908 239256
rect 276024 238266 306718 238268
rect 276024 238264 292802 238266
rect 276024 235900 278872 238264
rect 281120 235902 292802 238264
rect 295050 235904 306718 238266
rect 308966 238266 342908 238268
rect 308966 238264 334482 238266
rect 308966 235904 320552 238264
rect 295050 235902 320552 235904
rect 281120 235900 320552 235902
rect 322800 238186 334482 238264
rect 322800 235900 329586 238186
rect 276024 235836 329586 235900
rect 332118 235902 334482 238186
rect 336730 235902 342908 238266
rect 332118 235836 342908 235902
rect 276024 235042 342908 235836
rect 202180 233278 206206 235042
rect 283526 234140 287552 235042
rect 202210 223352 206008 233278
rect 283708 223352 287506 234140
rect 192302 222348 215530 223352
rect 192302 222346 209846 222348
rect 192302 219982 195916 222346
rect 198164 219984 209846 222346
rect 212094 219984 215530 222348
rect 198164 219982 215530 219984
rect 192302 219138 215530 219982
rect 276024 222364 342908 223352
rect 276024 222362 307128 222364
rect 276024 222360 293212 222362
rect 276024 219996 279282 222360
rect 281530 219998 293212 222360
rect 295460 220000 307128 222362
rect 309376 222362 342908 222364
rect 309376 222360 334892 222362
rect 309376 220000 320962 222360
rect 295460 219998 320962 220000
rect 281530 219996 320962 219998
rect 323210 222332 334892 222360
rect 323210 219996 329804 222332
rect 276024 219982 329804 219996
rect 332336 219998 334892 222332
rect 337140 219998 342908 222362
rect 332336 219982 342908 219998
rect 276024 219138 342908 219982
rect 202210 206900 206008 219138
rect 283708 206900 287506 219138
rect 192302 205896 215530 206900
rect 192302 205894 209846 205896
rect 100842 204960 101190 204980
rect 97392 204940 101190 204960
rect 97392 204656 100876 204940
rect 101156 204656 101190 204940
rect 97392 204642 101190 204656
rect 100842 204622 101190 204642
rect 192302 203530 195916 205894
rect 198164 203532 209846 205894
rect 212094 203532 215530 205896
rect 198164 203530 215530 203532
rect 192302 202686 215530 203530
rect 276024 205928 342908 206900
rect 276024 205912 330006 205928
rect 276024 205910 307128 205912
rect 276024 205908 293212 205910
rect 276024 203544 279282 205908
rect 281530 203546 293212 205908
rect 295460 203548 307128 205910
rect 309376 205908 330006 205912
rect 309376 203548 320962 205908
rect 295460 203546 320962 203548
rect 281530 203544 320962 203546
rect 323210 203578 330006 205908
rect 332538 205910 342908 205928
rect 332538 203578 334892 205910
rect 323210 203546 334892 203578
rect 337140 203546 342908 205910
rect 323210 203544 342908 203546
rect 276024 202686 342908 203544
rect 202210 192092 206008 202686
rect 283708 192092 287506 202686
rect 192302 191088 215530 192092
rect 192302 191086 209436 191088
rect 192302 188722 195506 191086
rect 197754 188724 209436 191086
rect 211684 188724 215530 191088
rect 197754 188722 215530 188724
rect 192302 187878 215530 188722
rect 276024 191104 342908 192092
rect 276024 191102 306718 191104
rect 276024 191100 292802 191102
rect 276024 188736 278872 191100
rect 281120 188738 292802 191100
rect 295050 188740 306718 191102
rect 308966 191102 342908 191104
rect 308966 191100 334482 191102
rect 308966 188740 320552 191100
rect 295050 188738 320552 188740
rect 281120 188736 320552 188738
rect 322800 190930 334482 191100
rect 322800 188736 329932 190930
rect 276024 188580 329932 188736
rect 332464 188738 334482 190930
rect 336730 188738 342908 191102
rect 332464 188580 342908 188738
rect 276024 187878 342908 188580
rect 202210 177832 206008 187878
rect 283708 177832 287506 187878
rect 192302 176844 342908 177832
rect 192302 176842 306170 176844
rect 192302 176840 292254 176842
rect 192302 176832 278324 176840
rect 192302 176830 264490 176832
rect 192302 176828 222804 176830
rect 192302 176826 208888 176828
rect 192302 174462 194958 176826
rect 197206 174464 208888 176826
rect 211136 174466 222804 176828
rect 225052 176828 250574 176830
rect 225052 174466 236644 176828
rect 211136 174464 236644 174466
rect 238892 174466 250574 176828
rect 252822 174468 264490 176830
rect 266738 174476 278324 176832
rect 280572 174478 292254 176840
rect 294502 174480 306170 176842
rect 308418 176842 342908 176844
rect 308418 176840 333934 176842
rect 308418 174480 320004 176840
rect 294502 174478 320004 174480
rect 280572 174476 320004 174478
rect 322252 176758 333934 176840
rect 322252 174476 329894 176758
rect 266738 174468 329894 174476
rect 252822 174466 329894 174468
rect 238892 174464 329894 174466
rect 197206 174462 329894 174464
rect 192302 174408 329894 174462
rect 332426 174478 333934 176758
rect 336182 174478 342908 176842
rect 332426 174408 342908 174478
rect 192302 173618 342908 174408
rect 202210 165006 206008 173618
rect 283708 165006 287506 173618
rect 192302 164018 342908 165006
rect 192302 164016 306386 164018
rect 192302 164014 292470 164016
rect 192302 164006 278540 164014
rect 192302 164004 264706 164006
rect 192302 164002 223020 164004
rect 192302 164000 209104 164002
rect 192302 161636 195174 164000
rect 197422 161638 209104 164000
rect 211352 161640 223020 164002
rect 225268 164002 250790 164004
rect 225268 161640 236860 164002
rect 211352 161638 236860 161640
rect 239108 161640 250790 164002
rect 253038 161642 264706 164004
rect 266954 161650 278540 164006
rect 280788 161652 292470 164014
rect 294718 161654 306386 164016
rect 308634 164016 342908 164018
rect 308634 164014 334150 164016
rect 308634 161654 320220 164014
rect 294718 161652 320220 161654
rect 280788 161650 320220 161652
rect 322468 163954 334150 164014
rect 322468 161650 329820 163954
rect 266954 161642 329820 161650
rect 253038 161640 329820 161642
rect 239108 161638 329820 161640
rect 197422 161636 329820 161638
rect 192302 161604 329820 161636
rect 332352 161652 334150 163954
rect 336398 161652 342908 164016
rect 332352 161604 342908 161652
rect 192302 160792 342908 161604
rect 201534 143168 205714 160792
rect 201534 142646 205740 143168
rect 283276 142646 287456 160792
rect 187654 141658 352454 142646
rect 187654 141656 306118 141658
rect 187654 141654 292202 141656
rect 187654 141646 278272 141654
rect 187654 141644 264438 141646
rect 187654 141642 222752 141644
rect 187654 141640 208836 141642
rect 187654 139276 194906 141640
rect 197154 139278 208836 141640
rect 211084 139280 222752 141642
rect 225000 141642 250522 141644
rect 225000 139280 236592 141642
rect 211084 139278 236592 139280
rect 238840 139280 250522 141642
rect 252770 139282 264438 141644
rect 266686 139290 278272 141646
rect 280520 139292 292202 141654
rect 294450 139294 306118 141656
rect 308366 141656 347798 141658
rect 308366 141654 333882 141656
rect 308366 139294 319952 141654
rect 294450 139292 319952 139294
rect 280520 139290 319952 139292
rect 322200 141454 333882 141654
rect 322200 139290 329784 141454
rect 266686 139282 329784 139290
rect 252770 139280 329784 139282
rect 238840 139278 329784 139280
rect 197154 139276 329784 139278
rect 187654 139104 329784 139276
rect 332316 139292 333882 141454
rect 336130 139294 347798 141656
rect 350046 139294 352454 141658
rect 336130 139292 352454 139294
rect 332316 139104 352454 139292
rect 187654 138432 352454 139104
rect 201534 130166 205714 138432
rect 283276 130166 287456 138432
rect 187654 129464 352454 130166
rect 187654 129178 329636 129464
rect 187654 129176 306048 129178
rect 187654 129174 292132 129176
rect 187654 129166 278202 129174
rect 187654 129164 264368 129166
rect 187654 129162 222682 129164
rect 187654 129160 208766 129162
rect 187654 126796 194836 129160
rect 197084 126798 208766 129160
rect 211014 126800 222682 129162
rect 224930 129162 250452 129164
rect 224930 126800 236522 129162
rect 211014 126798 236522 126800
rect 238770 126800 250452 129162
rect 252700 126802 264368 129164
rect 266616 126810 278202 129166
rect 280450 126812 292132 129174
rect 294380 126814 306048 129176
rect 308296 129174 329636 129178
rect 308296 126814 319882 129174
rect 294380 126812 319882 126814
rect 280450 126810 319882 126812
rect 322130 127114 329636 129174
rect 332168 129178 352454 129464
rect 332168 129176 347728 129178
rect 332168 127114 333812 129176
rect 322130 126812 333812 127114
rect 336060 126814 347728 129176
rect 349976 126814 352454 129178
rect 336060 126812 352454 126814
rect 322130 126810 352454 126812
rect 266616 126802 352454 126810
rect 252700 126800 352454 126802
rect 238770 126798 352454 126800
rect 197084 126796 352454 126798
rect 187654 125952 352454 126796
rect 201534 118732 205714 125952
rect 283276 118732 287456 125952
rect 187654 117808 352454 118732
rect 187654 117744 329710 117808
rect 187654 117742 305978 117744
rect 187654 117740 292062 117742
rect 187654 117732 278132 117740
rect 187654 117730 264298 117732
rect 187654 117728 222612 117730
rect 187654 117726 208696 117728
rect 187654 115362 194766 117726
rect 197014 115364 208696 117726
rect 210944 115366 222612 117728
rect 224860 117728 250382 117730
rect 224860 115366 236452 117728
rect 210944 115364 236452 115366
rect 238700 115366 250382 117728
rect 252630 115368 264298 117730
rect 266546 115376 278132 117732
rect 280380 115378 292062 117740
rect 294310 115380 305978 117742
rect 308226 117740 329710 117744
rect 308226 115380 319812 117740
rect 294310 115378 319812 115380
rect 280380 115376 319812 115378
rect 322060 115458 329710 117740
rect 332242 117744 352454 117808
rect 332242 117742 347658 117744
rect 332242 115458 333742 117742
rect 322060 115378 333742 115458
rect 335990 115380 347658 117742
rect 349906 115380 352454 117744
rect 335990 115378 352454 115380
rect 322060 115376 352454 115378
rect 266546 115368 352454 115376
rect 252630 115366 352454 115368
rect 238700 115364 352454 115366
rect 197014 115362 352454 115364
rect 187654 114518 352454 115362
rect 201534 106322 205714 114518
rect 283276 106844 287456 114518
rect 283162 106322 287456 106844
rect 187654 105634 352454 106322
rect 187654 105334 329858 105634
rect 187654 105332 305840 105334
rect 187654 105330 291924 105332
rect 187654 105322 277994 105330
rect 187654 105320 264160 105322
rect 187654 105318 222474 105320
rect 187654 105316 208558 105318
rect 187654 102952 194628 105316
rect 196876 102954 208558 105316
rect 210806 102956 222474 105318
rect 224722 105318 250244 105320
rect 224722 102956 236314 105318
rect 210806 102954 236314 102956
rect 238562 102956 250244 105318
rect 252492 102958 264160 105320
rect 266408 102966 277994 105322
rect 280242 102968 291924 105330
rect 294172 102970 305840 105332
rect 308088 105330 329858 105334
rect 308088 102970 319674 105330
rect 294172 102968 319674 102970
rect 280242 102966 319674 102968
rect 321922 103284 329858 105330
rect 332390 105334 352454 105634
rect 332390 105332 347520 105334
rect 332390 103284 333604 105332
rect 321922 102968 333604 103284
rect 335852 102970 347520 105332
rect 349768 102970 352454 105334
rect 335852 102968 352454 102970
rect 321922 102966 352454 102968
rect 266408 102958 352454 102966
rect 252492 102956 352454 102958
rect 238562 102954 352454 102956
rect 196876 102952 352454 102954
rect 187654 102108 352454 102952
rect 200624 94788 205196 102108
rect 282436 90606 287008 102108
rect 270820 89918 352454 90606
rect 270820 89618 329282 89918
rect 270820 89616 305264 89618
rect 270820 89614 291348 89616
rect 270820 87250 277418 89614
rect 279666 87252 291348 89614
rect 293596 87254 305264 89616
rect 307512 89614 329282 89618
rect 307512 87254 319098 89614
rect 293596 87252 319098 87254
rect 279666 87250 319098 87252
rect 321346 87568 329282 89614
rect 331814 89618 352454 89918
rect 331814 89616 346944 89618
rect 331814 87568 333028 89616
rect 321346 87252 333028 87568
rect 335276 87254 346944 89616
rect 349192 87254 352454 89618
rect 335276 87252 352454 87254
rect 321346 87250 352454 87252
rect 270820 86392 352454 87250
rect 282436 78018 287008 86392
rect 270820 77330 352454 78018
rect 270820 77030 329282 77330
rect 270820 77028 305264 77030
rect 270820 77026 291348 77028
rect 270820 74662 277418 77026
rect 279666 74664 291348 77026
rect 293596 74666 305264 77028
rect 307512 77026 329282 77030
rect 307512 74666 319098 77026
rect 293596 74664 319098 74666
rect 279666 74662 319098 74664
rect 321346 74980 329282 77026
rect 331814 77030 352454 77330
rect 331814 77028 346944 77030
rect 331814 74980 333028 77028
rect 321346 74664 333028 74980
rect 335276 74666 346944 77028
rect 349192 74666 352454 77030
rect 335276 74664 352454 74666
rect 321346 74662 352454 74664
rect 270820 73804 352454 74662
rect 282436 65430 287008 73804
rect 270820 64742 352454 65430
rect 270820 64442 329282 64742
rect 270820 64440 305264 64442
rect 270820 64438 291348 64440
rect 270820 62074 277418 64438
rect 279666 62076 291348 64438
rect 293596 62078 305264 64440
rect 307512 64438 329282 64442
rect 307512 62078 319098 64438
rect 293596 62076 319098 62078
rect 279666 62074 319098 62076
rect 321346 62392 329282 64438
rect 331814 64442 352454 64742
rect 331814 64440 346944 64442
rect 331814 62392 333028 64440
rect 321346 62076 333028 62392
rect 335276 62078 346944 64440
rect 349192 62078 352454 64442
rect 335276 62076 352454 62078
rect 321346 62074 352454 62076
rect 270820 61216 352454 62074
rect 282436 47510 287008 61216
<< viali >>
rect 328962 663376 331494 665726
rect 329000 650632 331532 652982
rect 328962 636460 331494 638810
rect 329012 622110 331544 624460
rect 328974 607938 331506 610288
rect 329190 589392 331722 591742
rect 329152 575220 331684 577570
rect 329078 562416 331610 564766
rect 329292 544576 331824 546926
rect 329254 530404 331786 532754
rect 329180 517600 331712 519950
rect 329354 496068 331886 498418
rect 329316 481896 331848 484246
rect 329242 469092 331774 471442
rect 329602 455536 332134 457886
rect 329562 443812 332094 446162
rect 329642 419686 332174 422036
rect 329604 405514 332136 407864
rect 329530 392710 332062 395060
rect 329616 383900 332148 386250
rect 329578 369728 332110 372078
rect 329504 356924 332036 359274
rect 329224 345074 331756 347424
rect 329150 332270 331682 334620
rect 329682 317748 332214 320098
rect 329644 308068 332176 310418
rect 329606 297528 332138 299878
rect 329570 286424 332102 288774
rect 329570 274044 332102 276394
rect 329586 235836 332118 238186
rect 329804 219982 332336 222332
rect 97038 204634 97392 204968
rect 100876 204656 101156 204940
rect 330006 203578 332538 205928
rect 329932 188580 332464 190930
rect 329894 174408 332426 176758
rect 329820 161604 332352 163954
rect 329784 139104 332316 141454
rect 329636 127114 332168 129464
rect 329710 115458 332242 117808
rect 329858 103284 332390 105634
rect 329282 87568 331814 89918
rect 329282 74980 331814 77330
rect 329282 62392 331814 64742
<< metal1 >>
rect 16824 689368 20304 690522
rect 16824 688204 17538 689368
rect 18770 688204 20304 689368
rect 16824 686872 20304 688204
rect 16734 686270 20304 686872
rect 16734 685364 20294 686270
rect 16750 680872 20294 685364
rect 16768 679086 20294 680872
rect 16768 678024 20304 679086
rect 16824 670474 20304 678024
rect 31538 670552 84670 670818
rect 87172 670552 89064 670640
rect 23060 670474 89064 670552
rect 16824 669246 89064 670474
rect 16824 668490 89024 669246
rect 16860 668318 89024 668490
rect 16860 668246 38000 668318
rect 23060 668242 38000 668246
rect 82020 668242 89024 668318
rect 87136 490636 88744 668242
rect 328816 665726 331658 665892
rect 328816 663376 328962 665726
rect 331494 663376 331658 665726
rect 328816 663194 331658 663376
rect 328854 652982 331696 653148
rect 328854 650632 329000 652982
rect 331532 650632 331696 652982
rect 328854 650450 331696 650632
rect 328816 638810 331658 638976
rect 328816 636460 328962 638810
rect 331494 636460 331658 638810
rect 328816 636278 331658 636460
rect 430266 625150 432170 625254
rect 430266 625112 431906 625150
rect 430266 624914 430332 625112
rect 430530 624952 431906 625112
rect 432104 624952 432170 625150
rect 430530 624914 432170 624952
rect 430266 624830 432170 624914
rect 328866 624460 331708 624626
rect 328866 622110 329012 624460
rect 331544 622110 331708 624460
rect 328866 621928 331708 622110
rect 429390 621880 431990 621994
rect 429390 621852 431726 621880
rect 429390 621636 429474 621852
rect 429690 621664 431726 621852
rect 431942 621664 431990 621880
rect 429690 621636 431990 621664
rect 429390 621570 431990 621636
rect 428524 618572 431934 618668
rect 428524 618450 431688 618572
rect 428524 618244 428628 618450
rect 428836 618366 431688 618450
rect 431896 618366 431934 618572
rect 428836 618244 431934 618366
rect 428524 618188 431934 618244
rect 427656 615042 431972 615136
rect 427656 615014 431698 615042
rect 427656 614806 427750 615014
rect 427966 614834 431698 615014
rect 431914 614834 431972 615042
rect 427966 614806 431972 614834
rect 427656 614722 431972 614806
rect 426706 611764 432000 611878
rect 426706 611680 431708 611764
rect 426706 611472 426790 611680
rect 427024 611556 431708 611680
rect 431942 611556 432000 611764
rect 427024 611472 432000 611556
rect 426706 611406 432000 611472
rect 328828 610288 331670 610454
rect 328828 607938 328974 610288
rect 331506 607938 331670 610288
rect 328828 607756 331670 607938
rect 329044 591742 331886 591908
rect 329044 589392 329190 591742
rect 331722 589392 331886 591742
rect 329044 589210 331886 589392
rect 329006 577570 331848 577736
rect 329006 575220 329152 577570
rect 331684 575220 331848 577570
rect 329006 575038 331848 575220
rect 328932 564766 331774 564932
rect 328932 562416 329078 564766
rect 331610 562416 331774 564766
rect 328932 562234 331774 562416
rect 329146 546926 331988 547092
rect 329146 544576 329292 546926
rect 331824 544576 331988 546926
rect 329146 544394 331988 544576
rect 329108 532754 331950 532920
rect 329108 530404 329254 532754
rect 331786 530404 331950 532754
rect 329108 530222 331950 530404
rect 329034 519950 331876 520116
rect 329034 517600 329180 519950
rect 331712 517600 331876 519950
rect 329034 517418 331876 517600
rect 329208 498418 332050 498584
rect 329208 496068 329354 498418
rect 331886 496068 332050 498418
rect 329208 495886 332050 496068
rect 87136 485928 88752 490636
rect 87136 460628 88744 485928
rect 329170 484246 332012 484412
rect 329170 481896 329316 484246
rect 331848 481896 332012 484246
rect 329170 481714 332012 481896
rect 329096 471442 331938 471608
rect 329096 469092 329242 471442
rect 331774 469092 331938 471442
rect 329096 468910 331938 469092
rect 87132 459416 88760 460628
rect 90846 460076 94928 460088
rect 90846 460040 97140 460076
rect 90846 459996 96844 460040
rect 90846 459752 90886 459996
rect 91154 459752 96844 459996
rect 97108 459752 97140 460040
rect 90846 459706 97140 459752
rect 90846 459700 94928 459706
rect 87136 353226 88744 459416
rect 329456 457886 332298 458052
rect 329456 455536 329602 457886
rect 332134 455536 332298 457886
rect 329456 455354 332298 455536
rect 329416 446162 332258 446328
rect 329416 443812 329562 446162
rect 332094 443812 332258 446162
rect 329416 443630 332258 443812
rect 329496 422036 332338 422202
rect 329496 419686 329642 422036
rect 332174 419686 332338 422036
rect 329496 419504 332338 419686
rect 329458 407864 332300 408030
rect 329458 405514 329604 407864
rect 332136 405514 332300 407864
rect 329458 405332 332300 405514
rect 329384 395060 332226 395226
rect 329384 392710 329530 395060
rect 332062 392710 332226 395060
rect 329384 392528 332226 392710
rect 329470 386250 332312 386416
rect 329470 383900 329616 386250
rect 332148 383900 332312 386250
rect 329470 383718 332312 383900
rect 329432 372078 332274 372244
rect 329432 369728 329578 372078
rect 332110 369728 332274 372078
rect 329432 369546 332274 369728
rect 329358 359274 332200 359440
rect 329358 356924 329504 359274
rect 332036 356924 332200 359274
rect 329358 356742 332200 356924
rect 87136 353180 103126 353226
rect 87136 352910 102720 353180
rect 103036 352910 103126 353180
rect 87136 352836 103126 352910
rect 87136 351938 88744 352836
rect 87136 351392 88100 351938
rect 88682 351392 88744 351938
rect 87136 351320 88744 351392
rect 87058 350454 100280 350462
rect 87058 350410 103084 350454
rect 87058 350102 87154 350410
rect 87454 350378 103084 350410
rect 87454 350140 102826 350378
rect 103048 350140 103084 350378
rect 87454 350102 103084 350140
rect 87058 350088 103084 350102
rect 87058 350060 100280 350088
rect 88070 349558 88910 349728
rect 88070 348956 88146 349558
rect 88720 348956 88910 349558
rect 88070 203784 88910 348956
rect 329078 347424 331920 347590
rect 329078 345074 329224 347424
rect 331756 345074 331920 347424
rect 329078 344892 331920 345074
rect 329004 334620 331846 334786
rect 329004 332270 329150 334620
rect 331682 332270 331846 334620
rect 329004 332088 331846 332270
rect 329536 320098 332378 320264
rect 329536 317748 329682 320098
rect 332214 317748 332378 320098
rect 329536 317566 332378 317748
rect 329498 310418 332340 310584
rect 329498 308068 329644 310418
rect 332176 308068 332340 310418
rect 329498 307886 332340 308068
rect 329460 299878 332302 300044
rect 329460 297528 329606 299878
rect 332138 297528 332302 299878
rect 329460 297346 332302 297528
rect 329424 288774 332266 288940
rect 329424 286424 329570 288774
rect 332102 286424 332266 288774
rect 329424 286242 332266 286424
rect 329424 276394 332266 276560
rect 329424 274044 329570 276394
rect 332102 274044 332266 276394
rect 329424 273862 332266 274044
rect 329440 238186 332282 238352
rect 329440 235836 329586 238186
rect 332118 235836 332282 238186
rect 329440 235654 332282 235836
rect 329658 222332 332500 222498
rect 329658 219982 329804 222332
rect 332336 219982 332500 222332
rect 329658 219800 332500 219982
rect 329860 205928 332702 206094
rect 97004 204968 97418 205008
rect 97004 204634 97038 204968
rect 97392 204634 97418 204968
rect 97004 204592 97418 204634
rect 100842 204940 101190 204980
rect 100842 204656 100876 204940
rect 101156 204656 101190 204940
rect 100842 204622 101190 204656
rect 88070 203112 88932 203784
rect 329860 203578 330006 205928
rect 332538 203578 332702 205928
rect 329860 203396 332702 203578
rect 88070 202818 88440 203112
rect 88706 202818 88932 203112
rect 88070 202610 88932 202818
rect 329786 190930 332628 191096
rect 329786 188580 329932 190930
rect 332464 188580 332628 190930
rect 329786 188398 332628 188580
rect 329748 176758 332590 176924
rect 329748 174408 329894 176758
rect 332426 174408 332590 176758
rect 329748 174226 332590 174408
rect 329674 163954 332516 164120
rect 329674 161604 329820 163954
rect 332352 161604 332516 163954
rect 329674 161422 332516 161604
rect 329638 141454 332480 141620
rect 329638 139104 329784 141454
rect 332316 139104 332480 141454
rect 329638 138922 332480 139104
rect 329490 129464 332332 129630
rect 329490 127114 329636 129464
rect 332168 127114 332332 129464
rect 329490 126932 332332 127114
rect 329564 117808 332406 117974
rect 329564 115458 329710 117808
rect 332242 115458 332406 117808
rect 329564 115276 332406 115458
rect 329712 105634 332554 105800
rect 329712 103284 329858 105634
rect 332390 103284 332554 105634
rect 329712 103102 332554 103284
rect 329136 89918 331978 90084
rect 329136 87568 329282 89918
rect 331814 87568 331978 89918
rect 329136 87386 331978 87568
rect 329136 77330 331978 77496
rect 329136 74980 329282 77330
rect 331814 74980 331978 77330
rect 329136 74798 331978 74980
rect 329136 64742 331978 64908
rect 329136 62392 329282 64742
rect 331814 62392 331978 64742
rect 329136 62210 331978 62392
<< via1 >>
rect 17538 688204 18770 689368
rect 328962 663376 331494 665726
rect 329000 650632 331532 652982
rect 328962 636460 331494 638810
rect 430332 624914 430530 625112
rect 431906 624952 432104 625150
rect 329012 622110 331544 624460
rect 429474 621636 429690 621852
rect 431726 621664 431942 621880
rect 428628 618244 428836 618450
rect 431688 618366 431896 618572
rect 427750 614806 427966 615014
rect 431698 614834 431914 615042
rect 426790 611472 427024 611680
rect 431708 611556 431942 611764
rect 328974 607938 331506 610288
rect 329190 589392 331722 591742
rect 329152 575220 331684 577570
rect 329078 562416 331610 564766
rect 329292 544576 331824 546926
rect 329254 530404 331786 532754
rect 329180 517600 331712 519950
rect 329354 496068 331886 498418
rect 329316 481896 331848 484246
rect 329242 469092 331774 471442
rect 90886 459752 91154 459996
rect 96844 459752 97108 460040
rect 329602 455536 332134 457886
rect 329562 443812 332094 446162
rect 329642 419686 332174 422036
rect 329604 405514 332136 407864
rect 329530 392710 332062 395060
rect 329616 383900 332148 386250
rect 329578 369728 332110 372078
rect 329504 356924 332036 359274
rect 102720 352910 103036 353180
rect 88100 351392 88682 351938
rect 87154 350102 87454 350410
rect 102826 350140 103048 350378
rect 88146 348956 88720 349558
rect 329224 345074 331756 347424
rect 329150 332270 331682 334620
rect 329682 317748 332214 320098
rect 329644 308068 332176 310418
rect 329606 297528 332138 299878
rect 329570 286424 332102 288774
rect 329570 274044 332102 276394
rect 329586 235836 332118 238186
rect 329804 219982 332336 222332
rect 97038 204634 97392 204968
rect 100876 204656 101156 204940
rect 330006 203578 332538 205928
rect 88440 202818 88706 203112
rect 329932 188580 332464 190930
rect 329894 174408 332426 176758
rect 329820 161604 332352 163954
rect 329784 139104 332316 141454
rect 329636 127114 332168 129464
rect 329710 115458 332242 117808
rect 329858 103284 332390 105634
rect 329282 87568 331814 89918
rect 329282 74980 331814 77330
rect 329282 62392 331814 64742
<< metal2 >>
rect 122144 699706 123216 699854
rect 69920 699460 70992 699660
rect 69920 698760 70052 699460
rect 70838 698760 70992 699460
rect 17196 689368 18976 689848
rect 17196 688204 17538 689368
rect 18770 688204 18976 689368
rect 17196 687656 18976 688204
rect 2428 683482 11996 683870
rect 2428 683404 10560 683482
rect 2428 682162 2972 683404
rect 4020 682240 10560 683404
rect 11608 682240 11996 683482
rect 4020 682162 11996 682240
rect 2428 681774 11996 682162
rect 69920 677082 70992 698760
rect 69872 675376 70992 677082
rect 122144 699006 122298 699706
rect 123084 699006 123216 699706
rect 122144 676610 123216 699006
rect 177172 699236 178322 699460
rect 330362 699404 331528 699648
rect 177172 698572 177430 699236
rect 178044 698572 178322 699236
rect 177172 678160 178322 698572
rect 228072 699186 229166 699330
rect 228072 698440 228208 699186
rect 228956 698440 229166 699186
rect 228072 679556 229166 698440
rect 330362 698704 330570 699404
rect 331356 698704 331528 699404
rect 330362 680982 331528 698704
rect 415130 699050 415606 699200
rect 415130 698768 415200 699050
rect 415504 698768 415606 699050
rect 415130 682442 415606 698768
rect 415130 681972 431438 682442
rect 330362 680954 414596 680982
rect 330362 680484 430624 680954
rect 330362 680366 414596 680484
rect 289562 679556 413646 679562
rect 228072 679286 413646 679556
rect 228072 679026 429724 679286
rect 228072 678816 429758 679026
rect 228072 678764 413646 678816
rect 228072 678758 293008 678764
rect 228072 678694 229166 678758
rect 177172 678086 293100 678160
rect 177172 677972 413664 678086
rect 177172 677502 428996 677972
rect 177172 677362 413664 677502
rect 177172 677332 178322 677362
rect 289580 677288 413664 677362
rect 122144 676578 171188 676610
rect 289510 676578 413594 676656
rect 122144 676484 413594 676578
rect 122144 676246 428052 676484
rect 122144 676014 428072 676246
rect 122144 675858 413594 676014
rect 122144 675780 293008 675858
rect 122144 675692 171188 675780
rect 122144 675668 123216 675692
rect 69872 675288 73284 675376
rect 69872 675274 169620 675288
rect 69872 675266 292914 675274
rect 69872 675114 413594 675266
rect 69872 674644 427110 675114
rect 69872 674476 413594 674644
rect 69872 674352 169620 674476
rect 289510 674468 413594 674476
rect 72376 674338 169620 674352
rect 328816 665726 331658 665892
rect 328816 663376 328962 665726
rect 331494 663376 331658 665726
rect 328816 663194 331658 663376
rect 87552 655878 91224 656038
rect 87552 655814 91232 655878
rect 87552 655802 93892 655814
rect 87552 655614 90648 655802
rect 90854 655614 93892 655802
rect 87552 655608 93892 655614
rect 87552 655548 91232 655608
rect 87552 655484 91224 655548
rect 87552 653022 88048 655484
rect 87168 652084 88368 653022
rect 86242 651744 88368 652084
rect 328854 652982 331696 653148
rect 86242 650678 88350 651744
rect 86242 491262 87772 650678
rect 328854 650632 329000 652982
rect 331532 650632 331696 652982
rect 328854 650450 331696 650632
rect 328816 638810 331658 638976
rect 328816 636460 328962 638810
rect 331494 636460 331658 638810
rect 328816 636278 331658 636460
rect 328866 624460 331708 624626
rect 328866 622110 329012 624460
rect 331544 622110 331708 624460
rect 328866 621928 331708 622110
rect 426744 611724 427080 674644
rect 427736 615068 428072 676014
rect 428620 618536 428956 677502
rect 429422 621938 429758 678816
rect 430280 625178 430616 680484
rect 431064 628408 431400 681972
rect 431062 628176 438690 628408
rect 431062 628158 431792 628176
rect 431064 627724 431404 628158
rect 430220 625112 430690 625178
rect 430220 624914 430332 625112
rect 430530 624914 430690 625112
rect 430220 624886 430690 624914
rect 429362 621852 429824 621938
rect 429362 621636 429474 621852
rect 429690 621636 429832 621852
rect 429362 621560 429832 621636
rect 428524 618450 428966 618536
rect 428524 618394 428628 618450
rect 428516 618244 428628 618394
rect 428836 618244 428966 618450
rect 427656 615014 428106 615068
rect 427656 614806 427750 615014
rect 427966 614806 428106 615014
rect 426684 611680 427132 611724
rect 426684 611472 426790 611680
rect 427024 611472 427132 611680
rect 328828 610288 331670 610454
rect 328828 607938 328974 610288
rect 331506 607938 331670 610288
rect 328828 607756 331670 607938
rect 426684 609482 427132 611472
rect 329044 591742 331886 591908
rect 329044 589392 329190 591742
rect 331722 589392 331886 591742
rect 329044 589210 331886 589392
rect 329006 577570 331848 577736
rect 329006 575220 329152 577570
rect 331684 575220 331848 577570
rect 329006 575038 331848 575220
rect 328932 564766 331774 564932
rect 328932 562416 329078 564766
rect 331610 562416 331774 564766
rect 328932 562234 331774 562416
rect 329146 546926 331988 547092
rect 329146 544576 329292 546926
rect 331824 544576 331988 546926
rect 329146 544394 331988 544576
rect 92722 536310 97020 536366
rect 92722 536054 92812 536310
rect 93082 536054 97020 536310
rect 92722 536030 97020 536054
rect 329108 532754 331950 532920
rect 329108 530404 329254 532754
rect 331786 530404 331950 532754
rect 329108 530222 331950 530404
rect 92928 520794 93212 520804
rect 92928 520542 96916 520794
rect 92928 511724 93212 520542
rect 329034 519950 331876 520116
rect 329034 517600 329180 519950
rect 331712 517600 331876 519950
rect 329034 517418 331876 517600
rect 92910 511328 93212 511724
rect 92910 509840 93230 511328
rect 92928 509680 93230 509840
rect 92590 509454 93412 509680
rect 92590 509058 92798 509454
rect 93262 509058 93412 509454
rect 92590 508850 93412 509058
rect 329208 498418 332050 498584
rect 329208 496068 329354 498418
rect 331886 496068 332050 498418
rect 329208 495886 332050 496068
rect 86242 485836 87796 491262
rect 86242 460964 87772 485836
rect 329170 484246 332012 484412
rect 329170 481896 329316 484246
rect 331848 481896 332012 484246
rect 329170 481714 332012 481896
rect 329096 471442 331938 471608
rect 329096 469092 329242 471442
rect 331774 469092 331938 471442
rect 329096 468910 331938 469092
rect 86120 460850 87840 460964
rect 86120 460262 87850 460850
rect 86120 459996 91194 460262
rect 86120 459752 90886 459996
rect 91154 459752 91194 459996
rect 86120 459618 91194 459752
rect 96818 460040 97136 460052
rect 96818 459752 96844 460040
rect 97108 459752 97136 460040
rect 96818 459732 97136 459752
rect 86120 459416 87850 459618
rect 86120 421152 87840 459416
rect 329456 457886 332298 458052
rect 329456 455536 329602 457886
rect 332134 455536 332298 457886
rect 329456 455354 332298 455536
rect 426684 448408 427152 609482
rect 427656 609444 428106 614806
rect 428516 612972 428966 618244
rect 429374 616222 429824 621560
rect 429374 616002 429832 616222
rect 428516 612696 428994 612972
rect 427648 609370 428106 609444
rect 427648 451688 428094 609370
rect 428548 455216 428994 612696
rect 429386 458466 429832 616002
rect 430226 467228 430672 624886
rect 430226 467022 430692 467228
rect 430264 461790 430692 467022
rect 431092 465002 431404 627724
rect 431842 625150 438776 625210
rect 431842 624952 431906 625150
rect 432104 624952 438776 625150
rect 431842 624910 438776 624952
rect 431674 621880 438608 621922
rect 431674 621664 431726 621880
rect 431942 621664 438608 621880
rect 431674 621622 438608 621664
rect 431654 618572 438588 618634
rect 431654 618366 431688 618572
rect 431896 618366 438588 618572
rect 431654 618334 438588 618366
rect 431654 615042 438588 615084
rect 431654 614834 431698 615042
rect 431914 614834 438588 615042
rect 431654 614784 438588 614834
rect 431654 611764 438588 611814
rect 431654 611556 431708 611764
rect 431942 611556 438588 611764
rect 431654 611514 438588 611556
rect 431092 464726 436300 465002
rect 430226 461512 436300 461790
rect 430264 461498 430692 461512
rect 429386 458206 436096 458466
rect 429386 458184 429832 458206
rect 428548 454956 436134 455216
rect 428548 454934 429882 454956
rect 427648 451652 429112 451688
rect 427648 451406 435950 451652
rect 427668 451356 435950 451406
rect 427668 451332 429112 451356
rect 426684 448402 428464 448408
rect 426684 448124 436024 448402
rect 426684 448052 428464 448124
rect 329416 446162 332258 446328
rect 329416 443812 329562 446162
rect 332094 443812 332258 446162
rect 329416 443630 332258 443812
rect 86038 420824 87840 421152
rect 329496 422036 332338 422202
rect 86038 350410 87758 420824
rect 329496 419686 329642 422036
rect 332174 419686 332338 422036
rect 329496 419504 332338 419686
rect 329458 407864 332300 408030
rect 329458 405514 329604 407864
rect 332136 405514 332300 407864
rect 329458 405332 332300 405514
rect 329384 395060 332226 395226
rect 329384 392710 329530 395060
rect 332062 392710 332226 395060
rect 329384 392528 332226 392710
rect 329470 386250 332312 386416
rect 329470 383900 329616 386250
rect 332148 383900 332312 386250
rect 329470 383718 332312 383900
rect 329432 372078 332274 372244
rect 329432 369728 329578 372078
rect 332110 369728 332274 372078
rect 329432 369546 332274 369728
rect 329358 359274 332200 359440
rect 329358 356924 329504 359274
rect 332036 356924 332200 359274
rect 329358 356742 332200 356924
rect 102684 353180 103082 353226
rect 102684 352910 102720 353180
rect 103036 352910 103082 353180
rect 102684 352864 103082 352910
rect 88054 351938 88730 352030
rect 88054 351392 88100 351938
rect 88682 351392 88730 351938
rect 88054 351346 88730 351392
rect 86038 350102 87154 350410
rect 87454 350102 87758 350410
rect 86038 349784 87758 350102
rect 85810 349636 87758 349784
rect 88174 349678 88720 351346
rect 102794 350378 103078 350434
rect 102794 350140 102826 350378
rect 103048 350140 103078 350378
rect 102794 350098 103078 350140
rect 85810 200510 87738 349636
rect 88090 349558 88776 349678
rect 88090 348956 88146 349558
rect 88720 348956 88776 349558
rect 88090 348882 88776 348956
rect 329078 347424 331920 347590
rect 329078 345074 329224 347424
rect 331756 345074 331920 347424
rect 329078 344892 331920 345074
rect 329004 334620 331846 334786
rect 329004 332270 329150 334620
rect 331682 332270 331846 334620
rect 329004 332088 331846 332270
rect 329536 320098 332378 320264
rect 329536 317748 329682 320098
rect 332214 317748 332378 320098
rect 329536 317566 332378 317748
rect 329498 310418 332340 310584
rect 329498 308068 329644 310418
rect 332176 308068 332340 310418
rect 329498 307886 332340 308068
rect 329460 299878 332302 300044
rect 329460 297528 329606 299878
rect 332138 297528 332302 299878
rect 329460 297346 332302 297528
rect 329424 288774 332266 288940
rect 329424 286424 329570 288774
rect 332102 286424 332266 288774
rect 329424 286242 332266 286424
rect 329424 276394 332266 276560
rect 329424 274044 329570 276394
rect 332102 274044 332266 276394
rect 329424 273862 332266 274044
rect 407356 259014 410032 259304
rect 329440 238186 332282 238352
rect 329440 235836 329586 238186
rect 332118 235836 332282 238186
rect 329440 235654 332282 235836
rect 329658 222332 332500 222498
rect 329658 219982 329804 222332
rect 332336 219982 332500 222332
rect 329658 219800 332500 219982
rect 329860 205928 332702 206094
rect 97004 204968 97418 205008
rect 97004 204634 97038 204968
rect 97392 204634 97418 204968
rect 97004 204592 97418 204634
rect 100842 204940 101190 204980
rect 100842 204656 100876 204940
rect 101156 204656 101190 204940
rect 100842 204622 101190 204656
rect 329860 203578 330006 205928
rect 332538 203578 332702 205928
rect 329860 203396 332702 203578
rect 88358 203112 101172 203150
rect 88358 202818 88440 203112
rect 88706 202818 101172 203112
rect 88358 202754 101172 202818
rect 85810 200162 97234 200510
rect 85810 199920 101132 200162
rect 85810 199712 97234 199920
rect 329786 190930 332628 191096
rect 329786 188580 329932 190930
rect 332464 188580 332628 190930
rect 329786 188398 332628 188580
rect 329748 176758 332590 176924
rect 329748 174408 329894 176758
rect 332426 174408 332590 176758
rect 329748 174226 332590 174408
rect 329674 163954 332516 164120
rect 329674 161604 329820 163954
rect 332352 161604 332516 163954
rect 329674 161422 332516 161604
rect 329638 141454 332480 141620
rect 329638 139104 329784 141454
rect 332316 139104 332480 141454
rect 329638 138922 332480 139104
rect 329490 129464 332332 129630
rect 329490 127114 329636 129464
rect 332168 127114 332332 129464
rect 329490 126932 332332 127114
rect 329564 117808 332406 117974
rect 329564 115458 329710 117808
rect 332242 115458 332406 117808
rect 329564 115276 332406 115458
rect 329712 105634 332554 105800
rect 329712 103284 329858 105634
rect 332390 103284 332554 105634
rect 329712 103102 332554 103284
rect 329136 89918 331978 90084
rect 329136 87568 329282 89918
rect 331814 87568 331978 89918
rect 329136 87386 331978 87568
rect 329136 77330 331978 77496
rect 329136 74980 329282 77330
rect 331814 74980 331978 77330
rect 329136 74798 331978 74980
rect 329136 64742 331978 64908
rect 329136 62392 329282 64742
rect 331814 62392 331978 64742
rect 329136 62210 331978 62392
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 70052 698760 70838 699460
rect 17538 688204 18770 689368
rect 2972 682162 4020 683404
rect 10560 682240 11608 683482
rect 122298 699006 123084 699706
rect 177430 698572 178044 699236
rect 228208 698440 228956 699186
rect 330570 698704 331356 699404
rect 415200 698768 415504 699050
rect 328962 663376 331494 665726
rect 90648 655614 90854 655802
rect 329000 650632 331532 652982
rect 328962 636460 331494 638810
rect 329012 622110 331544 624460
rect 328974 607938 331506 610288
rect 329190 589392 331722 591742
rect 329152 575220 331684 577570
rect 329078 562416 331610 564766
rect 329292 544576 331824 546926
rect 92812 536054 93082 536310
rect 329254 530404 331786 532754
rect 329180 517600 331712 519950
rect 92798 509058 93262 509454
rect 329354 496068 331886 498418
rect 329316 481896 331848 484246
rect 329242 469092 331774 471442
rect 329602 455536 332134 457886
rect 329562 443812 332094 446162
rect 329642 419686 332174 422036
rect 329604 405514 332136 407864
rect 329530 392710 332062 395060
rect 329616 383900 332148 386250
rect 329578 369728 332110 372078
rect 329504 356924 332036 359274
rect 329224 345074 331756 347424
rect 329150 332270 331682 334620
rect 329682 317748 332214 320098
rect 329644 308068 332176 310418
rect 329606 297528 332138 299878
rect 329570 286424 332102 288774
rect 329570 274044 332102 276394
rect 329586 235836 332118 238186
rect 329804 219982 332336 222332
rect 97038 204634 97392 204968
rect 100876 204656 101156 204940
rect 330006 203578 332538 205928
rect 329932 188580 332464 190930
rect 329894 174408 332426 176758
rect 329820 161604 332352 163954
rect 329784 139104 332316 141454
rect 329636 127114 332168 129464
rect 329710 115458 332242 117808
rect 329858 103284 332390 105634
rect 329282 87568 331814 89918
rect 329282 74980 331814 77330
rect 329282 62392 331814 64742
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 16752 698466 20824 702300
rect 68662 699460 72734 702300
rect 68662 698760 70052 699460
rect 70838 698760 72734 699460
rect 68662 698466 72734 698760
rect 120678 699706 124750 702300
rect 120678 699006 122298 699706
rect 123084 699006 124750 699706
rect 120678 698676 124750 699006
rect 165926 698488 169998 702300
rect 176336 699236 180408 702300
rect 176336 698572 177430 699236
rect 178044 698572 180408 699236
rect 16990 690532 20688 698466
rect 176336 698416 180408 698572
rect 217628 698310 221700 702300
rect 228108 699186 232180 702300
rect 228108 698440 228208 699186
rect 228956 698440 232180 699186
rect 228108 698310 232180 698440
rect 319336 698382 323408 702300
rect 329748 699404 333820 702300
rect 329748 698704 330570 699404
rect 331356 698704 333820 699404
rect 329748 698310 333820 698704
rect 413780 699050 417852 702300
rect 413780 698768 415200 699050
rect 415504 698768 417852 699050
rect 465732 698778 469804 702300
rect 413780 698622 417852 698768
rect 510880 698640 514952 702340
rect 520902 698606 524974 702340
rect 566594 702300 571594 704800
rect 567176 698412 571248 702300
rect 16442 689368 20688 690532
rect 16442 688204 17538 689368
rect 18770 688342 20688 689368
rect 18770 688204 20552 688342
rect 16442 687452 20552 688204
rect -800 684728 1700 685242
rect 11666 684804 18750 684860
rect 11666 684744 20294 684804
rect -800 683404 4602 684728
rect -800 682162 2972 683404
rect 4020 682162 4602 683404
rect -800 680942 4602 682162
rect 10036 683482 20294 684744
rect 10036 682240 10560 683482
rect 11608 682240 20294 683482
rect 582300 682418 584800 682984
rect -800 680242 1700 680942
rect 10036 680936 20294 682240
rect 11666 680900 20294 680936
rect 16750 680872 20294 680900
rect 16768 678024 20294 680872
rect 574234 678344 584800 682418
rect 16860 670474 20166 678024
rect 582300 677984 584800 678344
rect 31538 670552 84670 670818
rect 87172 670552 89064 670640
rect 23060 670474 89064 670552
rect 16860 669246 89064 670474
rect 16860 668318 89024 669246
rect 16860 668246 38000 668318
rect 23060 668242 38000 668246
rect 82020 668242 89024 668318
rect 87422 656140 88852 668242
rect 328816 665726 331658 665892
rect 328816 663376 328962 665726
rect 331494 663376 331658 665726
rect 328816 663194 331658 663376
rect 87394 655802 90980 656140
rect 87394 655614 90648 655802
rect 90854 655614 90980 655802
rect 87394 655386 90980 655614
rect 328854 652982 331696 653148
rect 328854 650632 329000 652982
rect 331532 650632 331696 652982
rect 328854 650450 331696 650632
rect -800 648098 1660 648642
rect -800 644312 20156 648098
rect -800 643842 1660 644312
rect 582340 644184 584800 644584
rect 574030 640110 584800 644184
rect 582340 639784 584800 640110
rect 328816 638810 331658 638976
rect -800 638250 1660 638642
rect -800 634464 20016 638250
rect 328816 636460 328962 638810
rect 331494 636460 331658 638810
rect 328816 636278 331658 636460
rect -800 633842 1660 634464
rect 582340 634254 584800 634584
rect 574228 630180 584800 634254
rect 582340 629784 584800 630180
rect 328866 624460 331708 624626
rect 328866 622110 329012 624460
rect 331544 622110 331708 624460
rect 328866 621928 331708 622110
rect 328828 610288 331670 610454
rect 328828 607938 328974 610288
rect 331506 607938 331670 610288
rect 328828 607756 331670 607938
rect 329044 591742 331886 591908
rect 329044 589392 329190 591742
rect 331722 589392 331886 591742
rect 583520 589472 584800 589584
rect 329044 589210 331886 589392
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 575062 584856 583716 585090
rect 575062 584744 584800 584856
rect 575062 584534 583716 584744
rect 575046 583674 583700 583954
rect 575046 583562 584800 583674
rect 575046 583398 583700 583562
rect 329006 577570 331848 577736
rect 329006 575220 329152 577570
rect 331684 575220 331848 577570
rect 329006 575038 331848 575220
rect 328932 564766 331774 564932
rect -800 563786 1660 564242
rect -800 560000 20086 563786
rect 328932 562416 329078 564766
rect 331610 562416 331774 564766
rect 328932 562234 331774 562416
rect -800 559442 1660 560000
rect -800 553726 1660 554242
rect 512570 553978 529414 554950
rect -800 549940 20016 553726
rect 512570 551694 513626 553978
rect 516246 551694 529414 553978
rect 512570 551006 529414 551694
rect 563414 554848 574574 554950
rect 582340 554848 584800 555362
rect 563414 551062 584800 554848
rect 563414 551006 574574 551062
rect 582340 550562 584800 551062
rect -800 549442 1660 549940
rect 329146 546926 331988 547092
rect 329146 544576 329292 546926
rect 331824 544576 331988 546926
rect 582340 544860 584800 545362
rect 329146 544394 331988 544576
rect 573994 541074 584800 544860
rect 582340 540562 584800 541074
rect 85038 536310 93230 536436
rect 85038 536214 92812 536310
rect 85034 536054 92812 536214
rect 93082 536054 93230 536310
rect 85034 535978 93230 536054
rect 85034 513008 85588 535978
rect 329108 532754 331950 532920
rect 329108 530404 329254 532754
rect 331786 530404 331950 532754
rect 329108 530222 331950 530404
rect 89420 522896 96624 522966
rect 89420 522660 96286 522896
rect 96516 522660 96624 522896
rect 89420 522580 96624 522660
rect 89430 522402 90308 522580
rect 89430 521982 90312 522402
rect 352 511806 3128 511836
rect 85034 511822 85610 513008
rect 82018 511806 85626 511822
rect 352 511788 34802 511806
rect 50488 511788 85626 511806
rect 352 511642 85626 511788
rect -800 511530 85626 511642
rect 352 511334 85626 511530
rect 352 511326 82750 511334
rect 2800 511318 82750 511326
rect 85034 511318 85610 511334
rect 34452 511300 50662 511318
rect 35026 510702 83476 510766
rect 85062 510702 85630 510802
rect 2684 510672 85630 510702
rect 380 510460 85630 510672
rect -800 510348 85630 510460
rect 380 510168 85630 510348
rect 380 510162 38000 510168
rect 82020 510162 85630 510168
rect -800 509166 480 509278
rect 82982 509238 83642 509388
rect 82982 508786 83114 509238
rect 83528 508786 83642 509238
rect 82982 508726 83642 508786
rect 82982 508352 83648 508726
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 11854 468606 28154 468640
rect 11854 468594 51140 468606
rect 82998 468596 83648 508352
rect 85062 500204 85630 510162
rect 2540 468584 51140 468594
rect 306 468574 51140 468584
rect 73058 468574 83648 468596
rect 306 468420 83648 468574
rect -800 468308 83648 468420
rect 306 468074 83648 468308
rect 2540 468068 83648 468074
rect 84488 499444 85630 500204
rect 2540 468052 83532 468068
rect 50782 468038 83532 468052
rect 50782 468020 73912 468038
rect 2628 467470 81170 467472
rect 2628 467468 83538 467470
rect 352 467238 83538 467468
rect -800 467126 83538 467238
rect 352 466970 83538 467126
rect 352 466966 81170 466970
rect 352 466958 3128 466966
rect -800 465944 480 466056
rect 81504 465706 82272 465860
rect 81504 465148 81630 465706
rect 82086 465148 82272 465706
rect 82946 465682 83538 466970
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 342 425198 3118 425454
rect -800 425086 3118 425198
rect 342 424944 3118 425086
rect 81504 424254 82272 465148
rect 39676 424236 82272 424254
rect 3082 424224 8420 424226
rect 350 424202 8420 424224
rect 18682 424202 82272 424236
rect 350 424016 82272 424202
rect -800 423904 82272 424016
rect 350 423738 82272 423904
rect 82926 465444 83538 465682
rect 350 423722 18786 423738
rect 350 423714 3126 423722
rect 39676 423702 81954 423738
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 370 381976 3146 382194
rect -800 381864 3146 381976
rect 370 381684 3146 381864
rect 408 380794 3184 381050
rect -800 380682 3184 380794
rect 408 380540 3184 380682
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 362 338754 3138 339018
rect -800 338642 3138 338754
rect 362 338508 3138 338642
rect 398 337572 3174 337772
rect -800 337460 3174 337572
rect 398 337262 3174 337460
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 380 295532 3156 295794
rect -800 295420 3156 295532
rect 380 295284 3156 295420
rect 436 294350 3212 294640
rect -800 294238 3212 294350
rect 436 294130 3212 294238
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 390 252510 3166 252784
rect -800 252398 3166 252510
rect 390 252274 3166 252398
rect 408 251328 3184 251648
rect -800 251216 3184 251328
rect 408 251138 3184 251216
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect -800 219064 1660 219688
rect -800 215278 20036 219064
rect -800 214888 1660 215278
rect -800 209150 1660 209688
rect -800 205364 20036 209150
rect -800 204888 1660 205364
rect 82926 205028 83476 465444
rect 84488 433756 85554 499444
rect 89446 465708 90312 521982
rect 329034 519950 331876 520116
rect 329034 517600 329180 519950
rect 331712 517600 331876 519950
rect 329034 517418 331876 517600
rect 92742 509454 93346 509540
rect 92742 509058 92798 509454
rect 93262 509058 93346 509454
rect 92742 508992 93346 509058
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 329208 498418 332050 498584
rect 329208 496068 329354 498418
rect 331886 496068 332050 498418
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 329208 495886 332050 496068
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 329170 484246 332012 484412
rect 329170 481896 329316 484246
rect 331848 481896 332012 484246
rect 329170 481714 332012 481896
rect 329096 471442 331938 471608
rect 329096 469092 329242 471442
rect 331774 469092 331938 471442
rect 329096 468910 331938 469092
rect 89446 465182 89586 465708
rect 90146 465182 90312 465708
rect 89446 464920 90312 465182
rect 329456 457886 332298 458052
rect 329456 455536 329602 457886
rect 332134 455536 332298 457886
rect 583520 455628 584800 455740
rect 329456 455354 332298 455536
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 329416 446162 332258 446328
rect 329416 443812 329562 446162
rect 332094 443812 332258 446162
rect 329416 443630 332258 443812
rect 84336 431474 85554 433756
rect 84336 358032 85400 431474
rect 329496 422036 332338 422202
rect 329496 419686 329642 422036
rect 332174 419686 332338 422036
rect 329496 419504 332338 419686
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 329458 407864 332300 408030
rect 329458 405514 329604 407864
rect 332136 405514 332300 407864
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 329458 405332 332300 405514
rect 583520 405296 584800 405408
rect 329384 395060 332226 395226
rect 329384 392710 329530 395060
rect 332062 392710 332226 395060
rect 329384 392528 332226 392710
rect 329470 386250 332312 386416
rect 329470 383900 329616 386250
rect 332148 383900 332312 386250
rect 329470 383718 332312 383900
rect 329432 372078 332274 372244
rect 329432 369728 329578 372078
rect 332110 369728 332274 372078
rect 329432 369546 332274 369728
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 84184 354534 85400 358032
rect 329358 359274 332200 359440
rect 329358 356924 329504 359274
rect 332036 356924 332200 359274
rect 583520 358874 584800 358986
rect 329358 356742 332200 356924
rect 84184 214158 85248 354534
rect 329078 347424 331920 347590
rect 329078 345074 329224 347424
rect 331756 345074 331920 347424
rect 329078 344892 331920 345074
rect 329004 334620 331846 334786
rect 329004 332270 329150 334620
rect 331682 332270 331846 334620
rect 329004 332088 331846 332270
rect 329536 320098 332378 320264
rect 329536 317748 329682 320098
rect 332214 317748 332378 320098
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 329536 317566 332378 317748
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect 329498 310418 332340 310584
rect 329498 308068 329644 310418
rect 332176 308068 332340 310418
rect 329498 307886 332340 308068
rect 329460 299878 332302 300044
rect 329460 297528 329606 299878
rect 332138 297528 332302 299878
rect 329460 297346 332302 297528
rect 329424 288774 332266 288940
rect 329424 286424 329570 288774
rect 332102 286424 332266 288774
rect 329424 286242 332266 286424
rect 329424 276394 332266 276560
rect 329424 274044 329570 276394
rect 332102 274044 332266 276394
rect 583520 275140 584800 275252
rect 329424 273862 332266 274044
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect 329440 238186 332282 238352
rect 329440 235836 329586 238186
rect 332118 235836 332282 238186
rect 329440 235654 332282 235836
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 329658 222332 332500 222498
rect 329658 219982 329804 222332
rect 332336 219982 332500 222332
rect 329658 219800 332500 219982
rect 84184 213874 95042 214158
rect 98844 213874 99504 213904
rect 84184 213672 99504 213874
rect 84184 213302 99000 213672
rect 99330 213302 99504 213672
rect 84184 213206 99504 213302
rect 85388 213202 99504 213206
rect 94702 213176 99504 213202
rect 98844 213128 99504 213176
rect 329860 205928 332702 206094
rect 82926 205012 85170 205028
rect 82926 205008 97410 205012
rect 82926 204968 97418 205008
rect 82926 204634 97038 204968
rect 97392 204634 97418 204968
rect 82926 204592 97418 204634
rect 100842 204940 101190 204980
rect 100842 204656 100876 204940
rect 101156 204656 101190 204940
rect 100842 204622 101190 204656
rect 82926 204578 97410 204592
rect 82926 204558 83476 204578
rect 84700 204566 97410 204578
rect 329860 203578 330006 205928
rect 332538 203578 332702 205928
rect 329860 203396 332702 203578
rect 582340 191430 584800 196230
rect 329786 190930 332628 191096
rect 329786 188580 329932 190930
rect 332464 188580 332628 190930
rect 329786 188398 332628 188580
rect 582340 181430 584800 186230
rect -800 177066 1660 177688
rect -800 173280 20044 177066
rect 329748 176758 332590 176924
rect 329748 174408 329894 176758
rect 332426 174408 332590 176758
rect 329748 174226 332590 174408
rect -800 172888 1660 173280
rect -800 167178 1660 167688
rect -800 163392 20184 167178
rect 329674 163954 332516 164120
rect -800 162888 1660 163392
rect 329674 161604 329820 163954
rect 332352 161604 332516 163954
rect 329674 161422 332516 161604
rect 561626 151098 575864 151442
rect 582340 151098 584800 151630
rect 561626 150902 584800 151098
rect 561626 147496 562246 150902
rect 565960 147496 584800 150902
rect 561626 147312 584800 147496
rect 561626 147054 577510 147312
rect 561626 147032 573062 147054
rect 582340 146830 584800 147312
rect 329638 141454 332480 141620
rect 329638 139104 329784 141454
rect 332316 139104 332480 141454
rect 329638 138922 332480 139104
rect 574134 141070 577510 141090
rect 582340 141070 584800 141630
rect 574134 137968 584800 141070
rect 574190 137284 584800 137968
rect 582340 136830 584800 137284
rect 329490 129464 332332 129630
rect 329490 127114 329636 129464
rect 332168 127114 332332 129464
rect 329490 126932 332332 127114
rect 362 124888 3138 125174
rect -800 124776 3138 124888
rect 362 124664 3138 124776
rect 398 123706 3174 124002
rect -800 123594 3174 123706
rect 398 123492 3174 123594
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 329564 117808 332406 117974
rect 329564 115458 329710 117808
rect 332242 115458 332406 117808
rect 329564 115276 332406 115458
rect 329712 105634 332554 105800
rect 329712 103284 329858 105634
rect 332390 103284 332554 105634
rect 329712 103102 332554 103284
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect 329136 89918 331978 90084
rect 329136 87568 329282 89918
rect 331814 87568 331978 89918
rect 329136 87386 331978 87568
rect 390 81666 3166 82006
rect -800 81554 3166 81666
rect 390 81496 3166 81554
rect 408 80484 3184 80798
rect -800 80372 3184 80484
rect 408 80288 3184 80372
rect -800 79190 480 79302
rect -800 78008 480 78120
rect 329136 77330 331978 77496
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 329136 74980 329282 77330
rect 331814 74980 331978 77330
rect 329136 74798 331978 74980
rect 329136 64742 331978 64908
rect 329136 62392 329282 64742
rect 331814 62392 331978 64742
rect 329136 62210 331978 62392
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect 398 38444 3174 38718
rect -800 38332 3174 38444
rect 398 38208 3174 38332
rect 390 37262 3166 37492
rect -800 37150 3166 37262
rect 390 36982 3166 37150
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect 390 17022 3166 17302
rect -800 16910 3166 17022
rect 583520 16910 584800 17022
rect 390 16792 3166 16910
rect 426 15840 3202 16082
rect -800 15728 3202 15840
rect 583520 15728 584800 15840
rect 426 15572 3202 15728
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 177430 698572 178044 699236
rect 228208 698440 228956 699186
rect 330570 698704 331356 699404
rect 328962 663376 331494 665726
rect 329000 650632 331532 652982
rect 328962 636460 331494 638810
rect 329012 622110 331544 624460
rect 328974 607938 331506 610288
rect 329190 589392 331722 591742
rect 329152 575220 331684 577570
rect 329078 562416 331610 564766
rect 513626 551694 516246 553978
rect 329292 544576 331824 546926
rect 329254 530404 331786 532754
rect 96286 522660 96516 522896
rect 83114 508786 83528 509238
rect 81630 465148 82086 465706
rect 329180 517600 331712 519950
rect 92798 509058 93262 509454
rect 329354 496068 331886 498418
rect 329316 481896 331848 484246
rect 329242 469092 331774 471442
rect 89586 465182 90146 465708
rect 329602 455536 332134 457886
rect 329562 443812 332094 446162
rect 329642 419686 332174 422036
rect 329604 405514 332136 407864
rect 329530 392710 332062 395060
rect 329616 383900 332148 386250
rect 329578 369728 332110 372078
rect 329504 356924 332036 359274
rect 329224 345074 331756 347424
rect 329150 332270 331682 334620
rect 329682 317748 332214 320098
rect 329644 308068 332176 310418
rect 329606 297528 332138 299878
rect 329570 286424 332102 288774
rect 329570 274044 332102 276394
rect 329586 235836 332118 238186
rect 329804 219982 332336 222332
rect 99000 213302 99330 213672
rect 97038 204634 97392 204968
rect 100876 204656 101156 204940
rect 330006 203578 332538 205928
rect 329932 188580 332464 190930
rect 329894 174408 332426 176758
rect 329820 161604 332352 163954
rect 562246 147496 565960 150902
rect 329784 139104 332316 141454
rect 329636 127114 332168 129464
rect 329710 115458 332242 117808
rect 329858 103284 332390 105634
rect 329282 87568 331814 89918
rect 329282 74980 331814 77330
rect 329282 62392 331814 64742
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 165926 698488 169998 702300
rect 176336 699236 180408 702300
rect 176336 698572 177430 699236
rect 178044 698572 180408 699236
rect 176336 698416 180408 698572
rect 217628 698310 221700 702300
rect 228108 699186 232180 702300
rect 228108 698440 228208 699186
rect 228956 698440 232180 699186
rect 228108 698310 232180 698440
rect 319336 698382 323408 702300
rect 329748 699404 333820 702300
rect 329748 698704 330570 699404
rect 331356 698704 333820 699404
rect 329748 698310 333820 698704
rect 327798 667938 333330 670524
rect 327582 665726 333330 667938
rect 327582 663376 328962 665726
rect 331494 663376 333330 665726
rect 327582 663094 333330 663376
rect 327578 661298 333330 663094
rect 328730 657432 333330 661298
rect 328718 656698 333330 657432
rect 328540 655438 333330 656698
rect 327798 652982 333330 655438
rect 327798 650632 329000 652982
rect 331532 650632 333330 652982
rect 327798 641022 333330 650632
rect 327582 638810 333330 641022
rect 90870 636852 92534 637056
rect 90870 602698 92548 636852
rect 327582 636460 328962 638810
rect 331494 636460 333330 638810
rect 327582 636178 333330 636460
rect 327578 634382 333330 636178
rect 328730 628176 333330 634382
rect 328552 626916 333330 628176
rect 327810 624460 333330 626916
rect 327810 622110 329012 624460
rect 331544 622110 333330 624460
rect 327810 612500 333330 622110
rect 327594 610288 333330 612500
rect 327594 607938 328974 610288
rect 331506 607938 333330 610288
rect 327594 607656 333330 607938
rect 327590 605842 333330 607656
rect 327810 605506 333330 605842
rect 88606 602608 107508 602698
rect 88606 602000 189802 602608
rect 328730 602000 333330 605506
rect 433664 602000 434934 612998
rect 448264 602000 448396 602122
rect 88606 598000 448396 602000
rect 88606 597946 189802 598000
rect 88606 597734 107508 597946
rect 328730 594198 333330 598000
rect 327988 591742 333330 594198
rect 327988 589392 329190 591742
rect 331722 589392 333330 591742
rect 327988 579782 333330 589392
rect 327772 577570 333330 579782
rect 327772 575220 329152 577570
rect 331684 575220 333330 577570
rect 327772 574938 333330 575220
rect 327768 573124 333330 574938
rect 327988 564766 333330 573124
rect 327988 562416 329078 564766
rect 331610 564032 333330 564766
rect 331610 562416 333518 564032
rect 327988 562112 333518 562416
rect 327984 560458 333518 562112
rect 328712 549382 333518 560458
rect 512990 553978 516846 554688
rect 512990 551694 513626 553978
rect 516246 551694 516846 553978
rect 512990 551096 516846 551694
rect 328090 546926 333518 549382
rect 328090 544576 329292 546926
rect 331824 545094 333518 546926
rect 331824 545048 333470 545094
rect 331824 544576 333432 545048
rect 328090 534966 333432 544576
rect 327874 532754 333432 534966
rect 327874 530404 329254 532754
rect 331786 530404 333432 532754
rect 327874 530122 333432 530404
rect 327870 528308 333432 530122
rect 96262 522896 96866 522992
rect 96262 522660 96286 522896
rect 96516 522660 96866 522896
rect 96262 522564 96866 522660
rect 93838 514000 94574 521360
rect 328090 519950 333432 528308
rect 328090 517600 329180 519950
rect 331712 519216 333432 519950
rect 331712 517600 333620 519216
rect 328090 517296 333620 517600
rect 328086 515642 333620 517296
rect 328730 514000 333620 515642
rect 499320 514000 501292 518462
rect 93738 513996 104744 514000
rect 128082 513996 516000 514000
rect 93738 510000 516000 513996
rect 92590 509520 93412 509680
rect 89550 509502 93412 509520
rect 83024 509454 93412 509502
rect 83024 509238 92798 509454
rect 83024 508786 83114 509238
rect 83528 509058 92798 509238
rect 93262 509058 93412 509454
rect 83528 508850 93412 509058
rect 83528 508786 93224 508850
rect 83024 508718 93224 508786
rect 89550 508698 93224 508718
rect 328730 500898 333330 510000
rect 328730 500874 333580 500898
rect 328152 498418 333580 500874
rect 328152 496068 329354 498418
rect 331886 496586 333580 498418
rect 331886 496540 333532 496586
rect 331886 496068 333494 496540
rect 328152 486458 333494 496068
rect 327936 484246 333494 486458
rect 327936 481896 329316 484246
rect 331848 481896 333494 484246
rect 327936 481614 333494 481896
rect 327932 479800 333494 481614
rect 328152 471442 333494 479800
rect 328152 469092 329242 471442
rect 331774 470708 333494 471442
rect 331774 469092 333682 470708
rect 328152 468788 333682 469092
rect 328148 467134 333682 468788
rect 328730 466804 333682 467134
rect 81438 465708 90250 465934
rect 81438 465706 89586 465708
rect 81438 465148 81630 465706
rect 82086 465182 89586 465706
rect 90146 465182 90250 465708
rect 82086 465148 90250 465182
rect 81438 464990 90250 465148
rect 328730 464000 333330 466804
rect 419392 464000 432120 464052
rect 190234 462730 432120 464000
rect 190234 461438 426126 462730
rect 431518 461438 432120 462730
rect 190234 460976 426162 461438
rect 431480 460976 432120 461438
rect 190234 460000 432120 460976
rect 282314 459978 289018 460000
rect 328400 457886 333332 460000
rect 419392 459956 432120 460000
rect 328400 455536 329602 457886
rect 332134 455536 333332 457886
rect 328400 455342 333332 455536
rect 328400 453774 333434 455342
rect 328730 449552 333330 453774
rect 328360 446162 333330 449552
rect 328360 443812 329562 446162
rect 332094 443812 333330 446162
rect 328360 443618 333330 443812
rect 328360 442050 333394 443618
rect 328730 440000 333330 442050
rect 89704 439832 96878 440000
rect 153712 439832 420906 440000
rect 89704 436000 420906 439832
rect 328730 426590 333330 436000
rect 328440 424336 333330 426590
rect 328440 422036 333372 424336
rect 328440 419686 329642 422036
rect 332174 419686 333372 422036
rect 328440 419492 333372 419686
rect 328440 417678 333474 419492
rect 328440 410076 333330 417678
rect 328224 407864 333330 410076
rect 328224 405514 329604 407864
rect 332136 405514 333330 407864
rect 328224 405232 333330 405514
rect 328220 403418 333330 405232
rect 328440 395060 333330 403418
rect 328440 392710 329530 395060
rect 332062 392710 333330 395060
rect 328440 392406 333330 392710
rect 328436 389352 333330 392406
rect 328414 388550 333330 389352
rect 328414 386250 333346 388550
rect 328414 383900 329616 386250
rect 332148 383900 333346 386250
rect 328414 383706 333346 383900
rect 328414 381892 333448 383706
rect 328414 374290 333330 381892
rect 328198 372078 333330 374290
rect 328198 369728 329578 372078
rect 332110 369728 333330 372078
rect 328198 369446 333330 369728
rect 328194 367632 333330 369446
rect 328414 359274 333330 367632
rect 328414 356924 329504 359274
rect 332036 356924 333330 359274
rect 328414 356620 333330 356924
rect 328410 352716 333330 356620
rect 328730 350022 333330 352716
rect 328060 349636 333330 350022
rect 327844 347424 333330 349636
rect 327844 345074 329224 347424
rect 331756 345074 333330 347424
rect 327844 344792 333330 345074
rect 327840 342978 333330 344792
rect 100846 330134 101740 337076
rect 328060 334620 333330 342978
rect 328060 332270 329150 334620
rect 331682 332270 333330 334620
rect 328060 331966 333330 332270
rect 100846 330058 103080 330134
rect 100188 330000 103928 330058
rect 141012 330000 142394 330434
rect 183398 330000 186480 330466
rect 328056 330000 333330 331966
rect 100188 326000 394636 330000
rect 100188 325786 103928 326000
rect 328730 321652 333330 326000
rect 328296 320098 334194 321652
rect 328296 317748 329682 320098
rect 332214 317748 334194 320098
rect 328296 317288 334194 317748
rect 328296 316140 334296 317288
rect 328730 311986 333330 316140
rect 328730 310418 334764 311986
rect 328730 308068 329644 310418
rect 332176 308068 334764 310418
rect 328730 307622 334764 308068
rect 328730 306474 334866 307622
rect 328730 301466 333330 306474
rect 328730 299878 334906 301466
rect 328730 297528 329606 299878
rect 332138 297528 334906 299878
rect 328730 297102 334906 297528
rect 328730 295954 335008 297102
rect 328730 290518 333330 295954
rect 328730 288774 334764 290518
rect 328730 286424 329570 288774
rect 332102 286424 334764 288774
rect 328730 286154 334764 286424
rect 328730 285006 334866 286154
rect 328730 278294 333330 285006
rect 328730 276394 335048 278294
rect 328730 274044 329570 276394
rect 332102 274044 335048 276394
rect 328730 273930 335048 274044
rect 328730 272782 335150 273930
rect 328730 262902 333330 272782
rect 328730 258182 334628 262902
rect 328730 256376 334730 258182
rect 328730 254000 333330 256376
rect 398104 254000 419348 254030
rect 106530 250000 419348 254000
rect 328730 240394 333330 250000
rect 398104 249936 419348 250000
rect 328730 238186 333662 240394
rect 328730 235836 329586 238186
rect 332118 235836 333662 238186
rect 328730 235550 333662 235836
rect 328730 233736 333764 235550
rect 328730 224490 333330 233736
rect 328730 222332 334072 224490
rect 328730 219982 329804 222332
rect 332336 219982 334072 222332
rect 328730 219646 334072 219982
rect 328730 217832 334174 219646
rect 98932 213904 101202 213914
rect 98844 213672 101202 213904
rect 98844 213302 99000 213672
rect 99330 213444 101202 213672
rect 99330 213302 99504 213444
rect 98844 213128 99504 213302
rect 328730 208038 333330 217832
rect 328730 205928 334072 208038
rect 97004 204968 97418 205008
rect 97004 204634 97038 204968
rect 97392 204634 97418 204968
rect 97004 204592 97418 204634
rect 100842 204940 101190 204980
rect 100842 204656 100876 204940
rect 101156 204656 101190 204940
rect 100842 204622 101190 204656
rect 328730 203578 330006 205928
rect 332538 203578 334072 205928
rect 328730 203194 334072 203578
rect 328730 201380 334174 203194
rect 328730 193230 333330 201380
rect 328730 190930 333662 193230
rect 328730 188580 329932 190930
rect 332464 188580 333662 190930
rect 328730 188386 333662 188580
rect 328730 186572 333764 188386
rect 96588 151746 98388 181984
rect 328730 178970 333330 186572
rect 328514 176758 333330 178970
rect 328514 174408 329894 176758
rect 332426 174408 333330 176758
rect 328514 174126 333330 174408
rect 328510 172312 333330 174126
rect 328730 163954 333330 172312
rect 328730 161604 329820 163954
rect 332352 161604 333330 163954
rect 328730 161300 333330 161604
rect 104406 151746 106512 156612
rect 328726 151746 333432 161300
rect 83990 151604 379272 151746
rect 544358 151604 558746 151646
rect 83990 151578 558746 151604
rect 83990 150902 566372 151578
rect 83990 147496 562246 150902
rect 565960 147496 566372 150902
rect 83990 146826 566372 147496
rect 83990 146758 549092 146826
rect 557004 146816 566372 146826
rect 328726 143168 333432 146758
rect 375160 146620 549092 146758
rect 328462 141454 333432 143168
rect 328462 139104 329784 141454
rect 332316 139104 333432 141454
rect 328462 138940 333432 139104
rect 328458 138744 333432 138940
rect 328458 137816 333330 138744
rect 328730 130688 333330 137816
rect 328392 129464 333330 130688
rect 328392 127114 329636 129464
rect 332168 127114 333330 129464
rect 328392 126460 333330 127114
rect 328388 125336 333330 126460
rect 328730 119254 333330 125336
rect 328322 117808 333330 119254
rect 328322 115458 329710 117808
rect 332242 115458 333330 117808
rect 328322 115026 333330 115458
rect 328318 113902 333330 115026
rect 328730 106844 333330 113902
rect 328184 105634 333330 106844
rect 328184 103284 329858 105634
rect 332390 103284 333330 105634
rect 328184 102616 333330 103284
rect 328180 101492 333330 102616
rect 328730 91454 333330 101492
rect 328698 90952 333330 91454
rect 327608 89918 333954 90952
rect 327608 87568 329282 89918
rect 331814 87568 333954 89918
rect 327608 86900 333954 87568
rect 327604 86098 333954 86900
rect 328698 85802 333330 86098
rect 328730 78866 333330 85802
rect 328698 78364 333330 78866
rect 327608 77330 333954 78364
rect 327608 74980 329282 77330
rect 331814 74980 333954 77330
rect 327608 74312 333954 74980
rect 327604 73510 333954 74312
rect 328698 73214 333330 73510
rect 328730 66278 333330 73214
rect 328698 65776 333330 66278
rect 327608 64742 333954 65776
rect 327608 62392 329282 64742
rect 331814 62392 333954 64742
rect 327608 61724 333954 62392
rect 327604 60922 333954 61724
rect 328698 60626 333330 60922
rect 91704 55990 108052 56000
rect 122568 55990 124316 59938
rect 328730 56000 333330 60626
rect 173296 55990 199070 56000
rect 91704 55958 199070 55990
rect 208362 55958 352454 56000
rect 91704 52000 352454 55958
rect 191940 51646 215346 52000
rect 328730 48958 333330 52000
<< via4 >>
rect 177430 698572 178044 699236
rect 228208 698440 228956 699186
rect 330570 698704 331356 699404
rect 513626 551694 516246 553978
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 165926 698488 169998 702300
rect 176336 699236 180408 702300
rect 176336 698572 177430 699236
rect 178044 698572 180408 699236
rect 176336 698416 180408 698572
rect 217628 698310 221700 702300
rect 228108 699186 232180 702300
rect 228108 698440 228208 699186
rect 228956 698440 232180 699186
rect 228108 698310 232180 698440
rect 319336 698382 323408 702300
rect 329748 699404 333820 702300
rect 329748 698704 330570 699404
rect 331356 698704 333820 699404
rect 329748 698310 333820 698704
rect 313114 667938 318892 670524
rect 128554 667272 189802 667342
rect 312956 667272 318892 667938
rect 128554 667264 318892 667272
rect 90404 667262 92700 667264
rect 97670 667262 318892 667264
rect 90404 666950 318892 667262
rect 439498 666950 440926 667024
rect 90404 663988 444066 666950
rect 93964 662112 94586 663988
rect 128554 663910 444066 663988
rect 185186 663882 444066 663910
rect 312838 663560 444066 663882
rect 312838 661298 318892 663560
rect 314104 657432 318786 661298
rect 314092 656698 318786 657432
rect 313914 655438 318786 656698
rect 313172 654454 318786 655438
rect 313114 647632 318786 654454
rect 439498 651952 440926 663560
rect 313114 641022 318892 647632
rect 312956 637156 318892 641022
rect 312838 634382 318892 637156
rect 314104 628176 318786 634382
rect 313926 626916 318786 628176
rect 313184 625932 318786 626916
rect 313126 619110 318786 625932
rect 313126 612500 318904 619110
rect 312968 608634 318904 612500
rect 312850 605842 318904 608634
rect 313184 605506 318904 605842
rect 314104 594198 318786 605506
rect 313362 593214 318786 594198
rect 313304 586392 318786 593214
rect 313304 579782 319082 586392
rect 313146 575916 319082 579782
rect 313028 573124 319082 575916
rect 313362 572216 319082 573124
rect 313362 563090 318786 572216
rect 313244 562112 318786 563090
rect 313244 560458 318778 562112
rect 314020 555780 318778 560458
rect 477472 555824 486468 555836
rect 477472 555812 511988 555824
rect 477472 555780 516884 555812
rect 91370 553978 516884 555780
rect 91370 551694 513626 553978
rect 516246 551694 516884 553978
rect 91370 550272 516884 551694
rect 91370 550218 511988 550272
rect 91370 549956 486468 550218
rect 91370 549882 104744 549956
rect 128082 549952 486468 549956
rect 91370 549874 99162 549882
rect 128082 549874 478382 549952
rect 97016 536726 97834 549874
rect 314020 549382 318888 549874
rect 313464 548398 318888 549382
rect 313406 541576 318888 548398
rect 313406 534966 319184 541576
rect 424412 537880 428146 549874
rect 313248 531100 319184 534966
rect 313130 528308 319184 531100
rect 313464 527400 319184 528308
rect 313464 518274 318888 527400
rect 313346 517296 318888 518274
rect 313346 515642 318880 517296
rect 314104 512772 318880 515642
rect 314104 507240 318786 512772
rect 313774 500898 318848 507240
rect 313774 500874 318950 500898
rect 313526 499890 318950 500874
rect 313468 493068 318950 499890
rect 245920 490000 261942 490022
rect 313468 490000 319246 493068
rect 420318 490000 422470 490086
rect 91216 486000 422470 490000
rect 103556 485518 104170 486000
rect 122018 485518 124932 486000
rect 245920 485980 261942 486000
rect 313310 482592 319246 486000
rect 313192 479800 319246 482592
rect 313526 478892 319246 479800
rect 420318 479534 422470 486000
rect 313526 469766 318950 478892
rect 420318 477172 435174 479534
rect 313408 468788 318950 469766
rect 313408 467134 318942 468788
rect 314104 466804 318942 467134
rect 314104 461276 318786 466804
rect 313774 460186 318786 461276
rect 313774 459358 318788 460186
rect 313716 454000 318890 459358
rect 190234 450000 420906 454000
rect 314104 449552 318786 450000
rect 313734 447634 318786 449552
rect 313676 442050 318850 447634
rect 314104 426590 318786 442050
rect 313814 424336 318786 426590
rect 313814 423508 318828 424336
rect 313756 410076 318930 423508
rect 313598 406210 318930 410076
rect 313480 405686 318930 406210
rect 313480 403418 318786 405686
rect 313814 393384 318786 403418
rect 313696 388550 318786 393384
rect 313696 387722 318802 388550
rect 313696 387062 318904 387722
rect 313730 374290 318904 387062
rect 313572 370424 318904 374290
rect 313454 369900 318904 370424
rect 313454 367632 318786 369900
rect 100014 363284 181806 363300
rect 100014 359160 207024 363284
rect 103176 356330 103886 359160
rect 179692 358604 207024 359160
rect 202192 354000 207024 358604
rect 313788 357598 318786 367632
rect 313670 354000 318786 357598
rect 202192 350000 394636 354000
rect 202192 349694 207024 350000
rect 313376 349636 318786 350000
rect 313218 345770 318786 349636
rect 313100 342978 318786 345770
rect 313434 332944 318786 342978
rect 313316 329970 318786 332944
rect 314104 321652 318786 329970
rect 313670 316140 319650 321652
rect 314104 311986 318786 316140
rect 314104 306474 320220 311986
rect 314104 301466 318786 306474
rect 314104 295954 320362 301466
rect 314104 290518 318786 295954
rect 314104 285006 320220 290518
rect 314104 278294 318786 285006
rect 314104 272782 320504 278294
rect 314104 270000 318786 272782
rect 396756 270000 419348 270076
rect 106530 266000 419348 270000
rect 112040 264924 114408 266000
rect 111810 262996 114408 264924
rect 111810 256572 114380 262996
rect 314104 262902 318786 266000
rect 396756 265968 419348 266000
rect 111810 255126 114408 256572
rect 112040 241032 114408 255126
rect 314104 256418 320084 262902
rect 410120 262496 410612 265968
rect 314104 256376 320080 256418
rect 111818 235962 114548 241032
rect 101184 233482 114548 235962
rect 101184 215264 102000 233482
rect 111818 233410 114548 233482
rect 314104 240394 318786 256376
rect 314104 233786 319118 240394
rect 314104 233736 319114 233786
rect 314104 224490 318786 233736
rect 314104 217882 319528 224490
rect 314104 217832 319524 217882
rect 314104 208038 318786 217832
rect 314104 201430 319528 208038
rect 314104 201380 319524 201430
rect 314104 193230 318786 201380
rect 314104 186622 319118 193230
rect 314104 186572 319114 186622
rect 314104 178970 318786 186572
rect 313888 175104 318786 178970
rect 313770 172312 318786 175104
rect 314104 162278 318786 172312
rect 313986 159536 318786 162278
rect 313986 143168 318782 159536
rect 313836 140422 318782 143168
rect 313836 139918 318786 140422
rect 313718 137816 318786 139918
rect 314104 130688 318786 137816
rect 313766 127438 318786 130688
rect 313648 125336 318786 127438
rect 314104 119254 318786 125336
rect 313696 116004 318786 119254
rect 313578 113902 318786 116004
rect 314104 106844 318786 113902
rect 313558 103594 318786 106844
rect 313440 101492 318786 103594
rect 314104 100000 318786 101492
rect 91704 96000 352454 100000
rect 114910 95926 121448 96000
rect 314104 91454 318786 96000
rect 314072 90952 318786 91454
rect 312982 87878 319410 90952
rect 312864 86098 319410 87878
rect 314072 85802 318786 86098
rect 314104 78866 318786 85802
rect 314072 78364 318786 78866
rect 312982 75290 319410 78364
rect 312864 73510 319410 75290
rect 314072 73214 318786 73510
rect 314104 66278 318786 73214
rect 314072 65776 318786 66278
rect 312982 62702 319410 65776
rect 312864 60922 319410 62702
rect 314072 60626 318786 60922
rect 314104 48958 318786 60626
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use pll_full_buffered2  pll_full_buffered2_0
timestamp 1647910864
transform 1 0 100982 0 1 174612
box -3258 0 88322 40874
use filter_buffered  filter_buffered_0
timestamp 1647903160
transform 1 0 115808 0 1 59356
box -2 0 89610 28900
use ashish  ashish_0
timestamp 1647888148
transform 1 0 406076 0 1 64768
box -2100 -2540 8350 2594
use div_pd_buffered  div_pd_buffered_0
timestamp 1647910864
transform 1 0 102890 0 1 341826
box -1894 -6452 88296 14680
use divider_buffered  divider_buffered_0
timestamp 1647903160
transform 1 0 409804 0 1 252392
box -1492 -3136 88296 10326
use pd_buffered  pd_buffered_0
timestamp 1647912062
transform 1 0 96910 0 1 454596
box -1894 -6512 88296 8906
use cp_buffered  cp_buffered_0
timestamp 1647912062
transform 1 0 96826 0 1 525962
box -2796 -7196 88288 10904
use ro_divider_buffered  ro_divider_buffered_0
timestamp 1647903160
transform 1 0 437678 0 1 468106
box -5944 -21716 87550 24552
use pll_full_buffered1  pll_full_buffered1_1
timestamp 1647909110
transform 1 0 93658 0 1 630304
box -2122 0 88316 32243
use ro_complete_buffered  ro_complete_buffered_0
timestamp 1647903160
transform 1 0 440094 0 1 631512
box -5924 -21716 87550 20899
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
