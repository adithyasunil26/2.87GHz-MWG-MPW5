magic
tech sky130A
timestamp 1640770827
<< nwell >>
rect -145 -20 875 200
<< nmos >>
rect -85 -240 -70 -150
rect 40 -240 55 -150
rect 165 -240 180 -150
rect 290 -240 305 -150
rect 415 -240 430 -150
rect 540 -240 555 -150
rect 665 -240 680 -150
rect 790 -240 805 -150
<< pmos >>
rect -85 0 -70 180
rect 90 0 105 180
rect 265 0 280 180
rect 440 0 455 180
rect 615 0 630 180
rect 790 0 805 180
<< ndiff >>
rect -125 -160 -85 -150
rect -125 -185 -120 -160
rect -95 -185 -85 -160
rect -125 -205 -85 -185
rect -125 -230 -120 -205
rect -95 -230 -85 -205
rect -125 -240 -85 -230
rect -70 -160 -30 -150
rect -70 -185 -60 -160
rect -35 -185 -30 -160
rect -70 -205 -30 -185
rect -70 -230 -60 -205
rect -35 -230 -30 -205
rect -70 -240 -30 -230
rect 0 -160 40 -150
rect 0 -185 5 -160
rect 30 -185 40 -160
rect 0 -205 40 -185
rect 0 -230 5 -205
rect 30 -230 40 -205
rect 0 -240 40 -230
rect 55 -160 95 -150
rect 55 -185 65 -160
rect 90 -185 95 -160
rect 55 -205 95 -185
rect 55 -230 65 -205
rect 90 -230 95 -205
rect 55 -240 95 -230
rect 125 -160 165 -150
rect 125 -185 130 -160
rect 155 -185 165 -160
rect 125 -205 165 -185
rect 125 -230 130 -205
rect 155 -230 165 -205
rect 125 -240 165 -230
rect 180 -160 220 -150
rect 180 -185 190 -160
rect 215 -185 220 -160
rect 180 -205 220 -185
rect 180 -230 190 -205
rect 215 -230 220 -205
rect 180 -240 220 -230
rect 250 -160 290 -150
rect 250 -185 255 -160
rect 280 -185 290 -160
rect 250 -205 290 -185
rect 250 -230 255 -205
rect 280 -230 290 -205
rect 250 -240 290 -230
rect 305 -160 345 -150
rect 305 -185 315 -160
rect 340 -185 345 -160
rect 305 -205 345 -185
rect 305 -230 315 -205
rect 340 -230 345 -205
rect 305 -240 345 -230
rect 375 -160 415 -150
rect 375 -185 380 -160
rect 405 -185 415 -160
rect 375 -205 415 -185
rect 375 -230 380 -205
rect 405 -230 415 -205
rect 375 -240 415 -230
rect 430 -160 470 -150
rect 430 -185 440 -160
rect 465 -185 470 -160
rect 430 -205 470 -185
rect 430 -230 440 -205
rect 465 -230 470 -205
rect 430 -240 470 -230
rect 500 -160 540 -150
rect 500 -185 505 -160
rect 530 -185 540 -160
rect 500 -205 540 -185
rect 500 -230 505 -205
rect 530 -230 540 -205
rect 500 -240 540 -230
rect 555 -160 595 -150
rect 555 -185 565 -160
rect 590 -185 595 -160
rect 555 -205 595 -185
rect 555 -230 565 -205
rect 590 -230 595 -205
rect 555 -240 595 -230
rect 625 -160 665 -150
rect 625 -185 630 -160
rect 655 -185 665 -160
rect 625 -205 665 -185
rect 625 -230 630 -205
rect 655 -230 665 -205
rect 625 -240 665 -230
rect 680 -160 720 -150
rect 680 -185 690 -160
rect 715 -185 720 -160
rect 680 -205 720 -185
rect 680 -230 690 -205
rect 715 -230 720 -205
rect 680 -240 720 -230
rect 750 -160 790 -150
rect 750 -185 755 -160
rect 780 -185 790 -160
rect 750 -205 790 -185
rect 750 -230 755 -205
rect 780 -230 790 -205
rect 750 -240 790 -230
rect 805 -160 845 -150
rect 805 -185 815 -160
rect 840 -185 845 -160
rect 805 -205 845 -185
rect 805 -230 815 -205
rect 840 -230 845 -205
rect 805 -240 845 -230
<< pdiff >>
rect -125 170 -85 180
rect -125 145 -120 170
rect -95 145 -85 170
rect -125 125 -85 145
rect -125 100 -120 125
rect -95 100 -85 125
rect -125 80 -85 100
rect -125 55 -120 80
rect -95 55 -85 80
rect -125 35 -85 55
rect -125 10 -120 35
rect -95 10 -85 35
rect -125 0 -85 10
rect -70 170 -30 180
rect -70 145 -60 170
rect -35 145 -30 170
rect -70 125 -30 145
rect -70 100 -60 125
rect -35 100 -30 125
rect -70 80 -30 100
rect -70 55 -60 80
rect -35 55 -30 80
rect -70 35 -30 55
rect -70 10 -60 35
rect -35 10 -30 35
rect -70 0 -30 10
rect 50 170 90 180
rect 50 145 55 170
rect 80 145 90 170
rect 50 125 90 145
rect 50 100 55 125
rect 80 100 90 125
rect 50 80 90 100
rect 50 55 55 80
rect 80 55 90 80
rect 50 35 90 55
rect 50 10 55 35
rect 80 10 90 35
rect 50 0 90 10
rect 105 170 145 180
rect 105 145 115 170
rect 140 145 145 170
rect 105 125 145 145
rect 105 100 115 125
rect 140 100 145 125
rect 105 80 145 100
rect 105 55 115 80
rect 140 55 145 80
rect 105 35 145 55
rect 105 10 115 35
rect 140 10 145 35
rect 105 0 145 10
rect 225 170 265 180
rect 225 145 230 170
rect 255 145 265 170
rect 225 125 265 145
rect 225 100 230 125
rect 255 100 265 125
rect 225 80 265 100
rect 225 55 230 80
rect 255 55 265 80
rect 225 35 265 55
rect 225 10 230 35
rect 255 10 265 35
rect 225 0 265 10
rect 280 170 320 180
rect 280 145 290 170
rect 315 145 320 170
rect 280 125 320 145
rect 280 100 290 125
rect 315 100 320 125
rect 280 80 320 100
rect 280 55 290 80
rect 315 55 320 80
rect 280 35 320 55
rect 280 10 290 35
rect 315 10 320 35
rect 280 0 320 10
rect 400 170 440 180
rect 400 145 405 170
rect 430 145 440 170
rect 400 125 440 145
rect 400 100 405 125
rect 430 100 440 125
rect 400 80 440 100
rect 400 55 405 80
rect 430 55 440 80
rect 400 35 440 55
rect 400 10 405 35
rect 430 10 440 35
rect 400 0 440 10
rect 455 170 495 180
rect 455 145 465 170
rect 490 145 495 170
rect 455 125 495 145
rect 455 100 465 125
rect 490 100 495 125
rect 455 80 495 100
rect 455 55 465 80
rect 490 55 495 80
rect 455 35 495 55
rect 455 10 465 35
rect 490 10 495 35
rect 455 0 495 10
rect 575 170 615 180
rect 575 145 580 170
rect 605 145 615 170
rect 575 125 615 145
rect 575 100 580 125
rect 605 100 615 125
rect 575 80 615 100
rect 575 55 580 80
rect 605 55 615 80
rect 575 35 615 55
rect 575 10 580 35
rect 605 10 615 35
rect 575 0 615 10
rect 630 170 670 180
rect 630 145 640 170
rect 665 145 670 170
rect 630 125 670 145
rect 630 100 640 125
rect 665 100 670 125
rect 630 80 670 100
rect 630 55 640 80
rect 665 55 670 80
rect 630 35 670 55
rect 630 10 640 35
rect 665 10 670 35
rect 630 0 670 10
rect 750 170 790 180
rect 750 145 755 170
rect 780 145 790 170
rect 750 125 790 145
rect 750 100 755 125
rect 780 100 790 125
rect 750 80 790 100
rect 750 55 755 80
rect 780 55 790 80
rect 750 35 790 55
rect 750 10 755 35
rect 780 10 790 35
rect 750 0 790 10
rect 805 170 845 180
rect 805 145 815 170
rect 840 145 845 170
rect 805 125 845 145
rect 805 100 815 125
rect 840 100 845 125
rect 805 80 845 100
rect 805 55 815 80
rect 840 55 845 80
rect 805 35 845 55
rect 805 10 815 35
rect 840 10 845 35
rect 805 0 845 10
<< ndiffc >>
rect -120 -185 -95 -160
rect -120 -230 -95 -205
rect -60 -185 -35 -160
rect -60 -230 -35 -205
rect 5 -185 30 -160
rect 5 -230 30 -205
rect 65 -185 90 -160
rect 65 -230 90 -205
rect 130 -185 155 -160
rect 130 -230 155 -205
rect 190 -185 215 -160
rect 190 -230 215 -205
rect 255 -185 280 -160
rect 255 -230 280 -205
rect 315 -185 340 -160
rect 315 -230 340 -205
rect 380 -185 405 -160
rect 380 -230 405 -205
rect 440 -185 465 -160
rect 440 -230 465 -205
rect 505 -185 530 -160
rect 505 -230 530 -205
rect 565 -185 590 -160
rect 565 -230 590 -205
rect 630 -185 655 -160
rect 630 -230 655 -205
rect 690 -185 715 -160
rect 690 -230 715 -205
rect 755 -185 780 -160
rect 755 -230 780 -205
rect 815 -185 840 -160
rect 815 -230 840 -205
<< pdiffc >>
rect -120 145 -95 170
rect -120 100 -95 125
rect -120 55 -95 80
rect -120 10 -95 35
rect -60 145 -35 170
rect -60 100 -35 125
rect -60 55 -35 80
rect -60 10 -35 35
rect 55 145 80 170
rect 55 100 80 125
rect 55 55 80 80
rect 55 10 80 35
rect 115 145 140 170
rect 115 100 140 125
rect 115 55 140 80
rect 115 10 140 35
rect 230 145 255 170
rect 230 100 255 125
rect 230 55 255 80
rect 230 10 255 35
rect 290 145 315 170
rect 290 100 315 125
rect 290 55 315 80
rect 290 10 315 35
rect 405 145 430 170
rect 405 100 430 125
rect 405 55 430 80
rect 405 10 430 35
rect 465 145 490 170
rect 465 100 490 125
rect 465 55 490 80
rect 465 10 490 35
rect 580 145 605 170
rect 580 100 605 125
rect 580 55 605 80
rect 580 10 605 35
rect 640 145 665 170
rect 640 100 665 125
rect 640 55 665 80
rect 640 10 665 35
rect 755 145 780 170
rect 755 100 780 125
rect 755 55 780 80
rect 755 10 780 35
rect 815 145 840 170
rect 815 100 840 125
rect 815 55 840 80
rect 815 10 840 35
<< poly >>
rect -85 180 -70 200
rect 90 180 105 200
rect 265 180 280 200
rect 440 180 455 200
rect 615 180 630 200
rect 790 180 805 200
rect -85 -30 -70 0
rect 90 -20 105 0
rect 265 -20 280 0
rect 440 -20 455 0
rect -125 -40 -70 -30
rect -125 -60 -115 -40
rect -95 -60 -70 -40
rect 70 -30 110 -20
rect 70 -50 80 -30
rect 100 -50 110 -30
rect 70 -60 110 -50
rect 250 -30 290 -20
rect 250 -50 260 -30
rect 280 -50 290 -30
rect 250 -60 290 -50
rect 425 -30 465 -20
rect 425 -50 435 -30
rect 455 -50 465 -30
rect 425 -60 465 -50
rect -125 -70 -70 -60
rect -85 -150 -70 -70
rect 615 -85 630 0
rect 790 -50 805 0
rect 750 -60 805 -50
rect 750 -80 760 -60
rect 780 -80 805 -60
rect 20 -95 60 -85
rect 20 -115 30 -95
rect 50 -115 60 -95
rect 20 -125 60 -115
rect 150 -95 190 -85
rect 150 -115 160 -95
rect 180 -115 190 -95
rect 150 -125 190 -115
rect 265 -95 305 -85
rect 265 -115 275 -95
rect 295 -115 305 -95
rect 265 -125 305 -115
rect 390 -95 430 -85
rect 390 -115 400 -95
rect 420 -115 430 -95
rect 390 -125 430 -115
rect 520 -95 560 -85
rect 520 -115 530 -95
rect 550 -115 560 -95
rect 520 -125 560 -115
rect 600 -95 640 -85
rect 750 -90 805 -80
rect 600 -115 610 -95
rect 630 -110 640 -95
rect 630 -115 680 -110
rect 600 -125 680 -115
rect 40 -150 55 -125
rect 165 -150 180 -125
rect 280 -130 305 -125
rect 290 -150 305 -130
rect 415 -150 430 -125
rect 540 -150 555 -125
rect 665 -150 680 -125
rect 790 -150 805 -90
rect -85 -270 -70 -240
rect 40 -270 55 -240
rect 165 -270 180 -240
rect 290 -270 305 -240
rect 415 -270 430 -240
rect 540 -270 555 -240
rect 665 -270 680 -240
rect 790 -270 805 -240
<< polycont >>
rect -115 -60 -95 -40
rect 80 -50 100 -30
rect 260 -50 280 -30
rect 435 -50 455 -30
rect 760 -80 780 -60
rect 30 -115 50 -95
rect 160 -115 180 -95
rect 275 -115 295 -95
rect 400 -115 420 -95
rect 530 -115 550 -95
rect 610 -115 630 -95
<< locali >>
rect -120 180 -100 265
rect 115 180 135 220
rect 230 180 250 265
rect 405 180 425 265
rect 580 180 600 265
rect 755 180 775 265
rect -125 170 -90 180
rect -125 145 -120 170
rect -95 145 -90 170
rect -125 125 -90 145
rect -125 100 -120 125
rect -95 100 -90 125
rect -125 80 -90 100
rect -125 55 -120 80
rect -95 55 -90 80
rect -125 35 -90 55
rect -125 10 -120 35
rect -95 10 -90 35
rect -125 0 -90 10
rect -65 170 -30 180
rect -65 145 -60 170
rect -35 145 -30 170
rect -65 125 -30 145
rect -65 100 -60 125
rect -35 100 -30 125
rect -65 80 -30 100
rect 50 170 85 180
rect 50 145 55 170
rect 80 145 85 170
rect 50 125 85 145
rect 50 100 55 125
rect 80 100 85 125
rect 50 80 85 100
rect -65 55 -60 80
rect -35 55 55 80
rect 80 55 85 80
rect -65 35 -30 55
rect -65 10 -60 35
rect -35 10 -30 35
rect -65 0 -30 10
rect 50 35 85 55
rect 50 10 55 35
rect 80 10 85 35
rect 50 0 85 10
rect 110 170 145 180
rect 110 145 115 170
rect 140 145 145 170
rect 110 125 145 145
rect 110 100 115 125
rect 140 100 145 125
rect 110 80 145 100
rect 110 55 115 80
rect 140 55 145 80
rect 110 35 145 55
rect 110 10 115 35
rect 140 10 145 35
rect 110 0 145 10
rect 225 170 260 180
rect 225 145 230 170
rect 255 145 260 170
rect 225 125 260 145
rect 225 100 230 125
rect 255 100 260 125
rect 225 80 260 100
rect 225 55 230 80
rect 255 55 260 80
rect 225 35 260 55
rect 225 10 230 35
rect 255 10 260 35
rect 225 0 260 10
rect 285 170 320 180
rect 285 145 290 170
rect 315 145 320 170
rect 285 125 320 145
rect 285 100 290 125
rect 315 100 320 125
rect 285 80 320 100
rect 285 55 290 80
rect 315 55 320 80
rect 400 170 435 180
rect 400 145 405 170
rect 430 145 435 170
rect 400 125 435 145
rect 400 100 405 125
rect 430 100 435 125
rect 400 80 435 100
rect 400 55 405 80
rect 430 55 435 80
rect 285 35 300 55
rect 320 35 365 55
rect 285 10 290 35
rect 315 10 320 35
rect 285 0 320 10
rect 70 -30 110 -20
rect 250 -30 290 -20
rect 345 -25 365 35
rect 400 35 435 55
rect 400 10 405 35
rect 430 10 435 35
rect 400 0 435 10
rect 460 170 495 180
rect 460 145 465 170
rect 490 145 495 170
rect 460 125 495 145
rect 460 100 465 125
rect 490 100 495 125
rect 460 80 495 100
rect 460 55 465 80
rect 490 55 495 80
rect 460 35 495 55
rect 460 10 465 35
rect 490 30 495 35
rect 460 0 495 10
rect 575 170 610 180
rect 575 145 580 170
rect 605 145 610 170
rect 575 125 610 145
rect 575 100 580 125
rect 605 100 610 125
rect 575 80 610 100
rect 575 55 580 80
rect 605 55 610 80
rect 575 35 610 55
rect 575 10 580 35
rect 605 10 610 35
rect 575 0 610 10
rect 635 170 670 180
rect 635 145 640 170
rect 665 145 670 170
rect 635 125 670 145
rect 635 100 640 125
rect 665 100 670 125
rect 635 80 670 100
rect 635 55 640 80
rect 665 55 670 80
rect 635 35 670 55
rect 635 10 640 35
rect 665 10 670 35
rect 635 0 670 10
rect 750 170 785 180
rect 750 145 755 170
rect 780 145 785 170
rect 750 125 785 145
rect 750 100 755 125
rect 780 100 785 125
rect 750 80 785 100
rect 750 55 755 80
rect 780 55 785 80
rect 750 35 785 55
rect 750 10 755 35
rect 780 10 785 35
rect 750 0 785 10
rect 810 170 845 180
rect 810 145 815 170
rect 840 145 845 170
rect 810 125 845 145
rect 810 100 815 125
rect 840 100 845 125
rect 810 80 845 100
rect 810 55 815 80
rect 840 55 845 80
rect 810 35 845 55
rect 810 10 815 35
rect 840 10 845 35
rect 810 0 845 10
rect 640 -20 665 0
rect 425 -25 465 -20
rect -125 -40 -85 -30
rect -145 -60 -115 -40
rect -95 -60 -85 -40
rect 70 -50 80 -30
rect 100 -50 165 -30
rect 185 -50 260 -30
rect 280 -50 290 -30
rect 70 -60 110 -50
rect -125 -70 -85 -60
rect 160 -85 180 -50
rect 250 -60 290 -50
rect 325 -30 550 -25
rect 325 -45 435 -30
rect 20 -95 60 -85
rect -40 -115 30 -95
rect 50 -115 60 -95
rect -60 -150 -35 -115
rect 20 -125 60 -115
rect 150 -95 190 -85
rect 150 -115 160 -95
rect 180 -115 190 -95
rect 150 -125 190 -115
rect 265 -95 305 -85
rect 265 -115 275 -95
rect 295 -115 305 -95
rect 265 -125 305 -115
rect 325 -150 345 -45
rect 425 -50 435 -45
rect 455 -45 550 -30
rect 640 -40 715 -20
rect 455 -50 465 -45
rect 425 -60 465 -50
rect 530 -85 550 -45
rect 690 -60 715 -40
rect 750 -60 790 -50
rect 690 -80 760 -60
rect 780 -80 790 -60
rect 390 -95 430 -85
rect 390 -115 400 -95
rect 420 -115 430 -95
rect 390 -125 430 -115
rect 520 -95 560 -85
rect 520 -115 530 -95
rect 550 -115 560 -95
rect 520 -125 560 -115
rect 600 -95 640 -85
rect 600 -115 610 -95
rect 630 -115 640 -95
rect 600 -125 640 -115
rect 690 -150 715 -80
rect 750 -90 790 -80
rect 815 -150 840 0
rect -125 -160 -90 -150
rect -125 -185 -120 -160
rect -95 -185 -90 -160
rect -125 -205 -90 -185
rect -125 -230 -120 -205
rect -95 -230 -90 -205
rect -125 -240 -90 -230
rect -65 -160 -30 -150
rect -65 -185 -60 -160
rect -35 -185 -30 -160
rect -65 -205 -30 -185
rect -65 -230 -60 -205
rect -35 -230 -30 -205
rect -65 -240 -30 -230
rect 0 -160 35 -150
rect 0 -185 5 -160
rect 30 -185 35 -160
rect 0 -205 35 -185
rect 0 -230 5 -205
rect 30 -230 35 -205
rect 0 -240 35 -230
rect 60 -160 75 -150
rect 60 -185 65 -160
rect 90 -185 95 -170
rect 60 -205 95 -185
rect 60 -230 65 -205
rect 90 -230 95 -205
rect 60 -240 95 -230
rect 125 -160 160 -150
rect 125 -185 130 -160
rect 155 -185 160 -160
rect 125 -205 160 -185
rect 125 -230 130 -205
rect 155 -230 160 -205
rect 125 -240 160 -230
rect 185 -160 220 -150
rect 185 -185 190 -160
rect 215 -185 220 -160
rect 185 -205 220 -185
rect 185 -230 190 -205
rect 215 -230 220 -205
rect 185 -240 220 -230
rect 250 -160 285 -150
rect 250 -185 255 -160
rect 280 -185 285 -160
rect 250 -205 285 -185
rect 250 -230 255 -205
rect 280 -230 285 -205
rect 250 -240 285 -230
rect 310 -160 345 -150
rect 310 -185 315 -160
rect 340 -185 345 -160
rect 310 -205 345 -185
rect 310 -230 315 -205
rect 340 -230 345 -205
rect 310 -240 345 -230
rect 375 -160 410 -150
rect 375 -185 380 -160
rect 405 -185 410 -160
rect 375 -205 410 -185
rect 375 -230 380 -205
rect 405 -230 410 -205
rect 375 -240 410 -230
rect 435 -160 450 -150
rect 435 -185 440 -160
rect 465 -185 470 -170
rect 435 -205 470 -185
rect 435 -230 440 -205
rect 465 -230 470 -205
rect 435 -240 470 -230
rect 500 -160 535 -150
rect 500 -185 505 -160
rect 530 -185 535 -160
rect 500 -205 535 -185
rect 500 -230 505 -205
rect 530 -230 535 -205
rect 500 -240 535 -230
rect 560 -160 595 -150
rect 560 -185 565 -160
rect 590 -185 595 -160
rect 560 -205 595 -185
rect 560 -230 565 -205
rect 590 -230 595 -205
rect 560 -240 595 -230
rect 625 -160 660 -150
rect 625 -185 630 -160
rect 655 -185 660 -160
rect 625 -205 660 -185
rect 625 -230 630 -205
rect 655 -230 660 -205
rect 625 -240 660 -230
rect 685 -160 720 -150
rect 685 -185 690 -160
rect 715 -185 720 -160
rect 685 -205 720 -185
rect 685 -230 690 -205
rect 715 -230 720 -205
rect 685 -240 720 -230
rect 750 -160 785 -150
rect 750 -185 755 -160
rect 780 -185 785 -160
rect 750 -205 785 -185
rect 750 -230 755 -205
rect 780 -230 785 -205
rect 750 -240 785 -230
rect 810 -160 845 -150
rect 810 -185 815 -160
rect 840 -185 845 -160
rect 810 -205 845 -185
rect 810 -230 815 -205
rect 840 -230 845 -205
rect 810 -240 845 -230
rect -120 -340 -95 -240
rect 5 -280 25 -240
rect -120 -345 -115 -340
rect 130 -340 155 -240
rect 190 -280 210 -240
rect 130 -345 135 -340
rect 255 -340 280 -240
rect 385 -280 405 -240
rect 255 -345 260 -340
rect 505 -340 530 -240
rect 565 -280 585 -240
rect 505 -345 510 -340
rect 630 -340 655 -240
rect 630 -345 635 -340
rect 755 -340 780 -240
rect 755 -345 760 -340
<< viali >>
rect -120 265 -100 285
rect 230 265 250 285
rect 115 220 135 240
rect 405 265 425 285
rect 580 265 600 285
rect 755 265 775 285
rect 300 35 320 55
rect 475 10 490 30
rect 490 10 495 30
rect 165 -50 185 -30
rect 260 -50 280 -30
rect -60 -115 -40 -95
rect 275 -115 295 -95
rect 760 -80 780 -60
rect 400 -115 420 -95
rect 610 -115 630 -95
rect 75 -160 95 -150
rect 75 -170 90 -160
rect 90 -170 95 -160
rect 450 -160 470 -150
rect 450 -170 465 -160
rect 465 -170 470 -160
rect 5 -300 25 -280
rect -115 -360 -95 -340
rect 190 -300 210 -280
rect 135 -360 155 -340
rect 385 -300 405 -280
rect 260 -360 280 -340
rect 565 -300 585 -280
rect 510 -360 530 -340
rect 635 -360 655 -340
rect 760 -360 780 -340
<< metal1 >>
rect -130 290 -90 295
rect -130 260 -125 290
rect -95 260 -90 290
rect -130 255 -90 260
rect 220 290 260 295
rect 220 260 225 290
rect 255 260 260 290
rect 220 255 260 260
rect 395 290 435 295
rect 395 260 400 290
rect 430 260 435 290
rect 395 255 435 260
rect 570 290 610 295
rect 570 260 575 290
rect 605 260 610 290
rect 570 255 610 260
rect 745 290 785 295
rect 745 260 750 290
rect 780 260 785 290
rect 745 255 785 260
rect 105 240 145 250
rect 105 235 115 240
rect -60 220 115 235
rect 135 220 145 240
rect -60 -85 -45 220
rect 105 210 145 220
rect 290 55 330 65
rect 290 50 300 55
rect 80 35 300 50
rect 320 35 330 55
rect -70 -95 -30 -85
rect -70 -115 -60 -95
rect -40 -115 -30 -95
rect -70 -125 -30 -115
rect 80 -140 95 35
rect 290 25 330 35
rect 465 30 505 40
rect 465 10 475 30
rect 495 10 505 30
rect 465 0 505 10
rect 155 -25 195 -20
rect 155 -55 160 -25
rect 190 -55 195 -25
rect 155 -60 195 -55
rect 250 -30 290 -20
rect 250 -50 260 -30
rect 280 -35 290 -30
rect 280 -50 420 -35
rect 250 -60 290 -50
rect 405 -85 420 -50
rect 265 -90 305 -85
rect 265 -120 270 -90
rect 300 -120 305 -90
rect 265 -125 305 -120
rect 390 -95 430 -85
rect 390 -115 400 -95
rect 420 -115 430 -95
rect 480 -100 495 0
rect 750 -60 790 -50
rect 750 -80 760 -60
rect 780 -65 790 -60
rect 780 -80 875 -65
rect 600 -95 640 -85
rect 750 -90 790 -80
rect 600 -100 610 -95
rect 390 -125 430 -115
rect 455 -115 610 -100
rect 630 -115 640 -95
rect 455 -140 470 -115
rect 600 -125 640 -115
rect 65 -150 105 -140
rect 65 -170 75 -150
rect 95 -170 105 -150
rect 65 -180 105 -170
rect 440 -150 480 -140
rect 440 -170 450 -150
rect 470 -170 480 -150
rect 440 -180 480 -170
rect -5 -280 35 -270
rect -5 -300 5 -280
rect 25 -285 35 -280
rect 180 -280 220 -270
rect 180 -285 190 -280
rect 25 -300 190 -285
rect 210 -300 220 -280
rect -5 -310 35 -300
rect 180 -310 220 -300
rect 375 -280 415 -270
rect 375 -300 385 -280
rect 405 -285 415 -280
rect 555 -280 595 -270
rect 555 -285 565 -280
rect 405 -300 565 -285
rect 585 -300 595 -280
rect 375 -310 415 -300
rect 555 -310 595 -300
rect -125 -335 -85 -330
rect -125 -365 -120 -335
rect -90 -365 -85 -335
rect -125 -370 -85 -365
rect 125 -335 165 -330
rect 125 -365 130 -335
rect 160 -365 165 -335
rect 125 -370 165 -365
rect 250 -335 290 -330
rect 250 -365 255 -335
rect 285 -365 290 -335
rect 250 -370 290 -365
rect 500 -335 540 -330
rect 500 -365 505 -335
rect 535 -365 540 -335
rect 500 -370 540 -365
rect 625 -335 665 -330
rect 625 -365 630 -335
rect 660 -365 665 -335
rect 625 -370 665 -365
rect 750 -335 790 -330
rect 750 -365 755 -335
rect 785 -365 790 -335
rect 750 -370 790 -365
<< via1 >>
rect -125 285 -95 290
rect -125 265 -120 285
rect -120 265 -100 285
rect -100 265 -95 285
rect -125 260 -95 265
rect 225 285 255 290
rect 225 265 230 285
rect 230 265 250 285
rect 250 265 255 285
rect 225 260 255 265
rect 400 285 430 290
rect 400 265 405 285
rect 405 265 425 285
rect 425 265 430 285
rect 400 260 430 265
rect 575 285 605 290
rect 575 265 580 285
rect 580 265 600 285
rect 600 265 605 285
rect 575 260 605 265
rect 750 285 780 290
rect 750 265 755 285
rect 755 265 775 285
rect 775 265 780 285
rect 750 260 780 265
rect 160 -30 190 -25
rect 160 -50 165 -30
rect 165 -50 185 -30
rect 185 -50 190 -30
rect 160 -55 190 -50
rect 270 -95 300 -90
rect 270 -115 275 -95
rect 275 -115 295 -95
rect 295 -115 300 -95
rect 270 -120 300 -115
rect -120 -340 -90 -335
rect -120 -360 -115 -340
rect -115 -360 -95 -340
rect -95 -360 -90 -340
rect -120 -365 -90 -360
rect 130 -340 160 -335
rect 130 -360 135 -340
rect 135 -360 155 -340
rect 155 -360 160 -340
rect 130 -365 160 -360
rect 255 -340 285 -335
rect 255 -360 260 -340
rect 260 -360 280 -340
rect 280 -360 285 -340
rect 255 -365 285 -360
rect 505 -340 535 -335
rect 505 -360 510 -340
rect 510 -360 530 -340
rect 530 -360 535 -340
rect 505 -365 535 -360
rect 630 -340 660 -335
rect 630 -360 635 -340
rect 635 -360 655 -340
rect 655 -360 660 -340
rect 630 -365 660 -360
rect 755 -340 785 -335
rect 755 -360 760 -340
rect 760 -360 780 -340
rect 780 -360 785 -340
rect 755 -365 785 -360
<< metal2 >>
rect -135 290 -85 300
rect -135 260 -125 290
rect -95 260 -85 290
rect -135 250 -85 260
rect 215 290 265 300
rect 215 260 225 290
rect 255 260 265 290
rect 215 250 265 260
rect 390 290 440 300
rect 390 260 400 290
rect 430 260 440 290
rect 390 250 440 260
rect 565 290 615 300
rect 565 260 575 290
rect 605 260 615 290
rect 565 250 615 260
rect 740 290 790 300
rect 740 260 750 290
rect 780 260 790 290
rect 740 250 790 260
rect -145 15 180 30
rect 165 -15 180 15
rect 150 -25 200 -15
rect 150 -55 160 -25
rect 190 -55 200 -25
rect 150 -65 200 -55
rect 260 -90 310 -80
rect 260 -100 270 -90
rect -145 -115 270 -100
rect 260 -120 270 -115
rect 300 -120 310 -90
rect 260 -130 310 -120
rect -130 -330 -80 -325
rect -130 -370 -125 -330
rect -85 -370 -80 -330
rect -130 -375 -80 -370
rect 120 -330 170 -325
rect 120 -370 125 -330
rect 165 -370 170 -330
rect 120 -375 170 -370
rect 245 -330 295 -325
rect 245 -370 250 -330
rect 290 -370 295 -330
rect 245 -375 295 -370
rect 495 -330 545 -325
rect 495 -370 500 -330
rect 540 -370 545 -330
rect 495 -375 545 -370
rect 620 -330 670 -325
rect 620 -370 625 -330
rect 665 -370 670 -330
rect 620 -375 670 -370
rect 745 -330 795 -325
rect 745 -370 750 -330
rect 790 -370 795 -330
rect 745 -375 795 -370
<< via2 >>
rect -125 260 -95 290
rect 225 260 255 290
rect 400 260 430 290
rect 575 260 605 290
rect 750 260 780 290
rect -125 -335 -85 -330
rect -125 -365 -120 -335
rect -120 -365 -90 -335
rect -90 -365 -85 -335
rect -125 -370 -85 -365
rect 125 -335 165 -330
rect 125 -365 130 -335
rect 130 -365 160 -335
rect 160 -365 165 -335
rect 125 -370 165 -365
rect 250 -335 290 -330
rect 250 -365 255 -335
rect 255 -365 285 -335
rect 285 -365 290 -335
rect 250 -370 290 -365
rect 500 -335 540 -330
rect 500 -365 505 -335
rect 505 -365 535 -335
rect 535 -365 540 -335
rect 500 -370 540 -365
rect 625 -335 665 -330
rect 625 -365 630 -335
rect 630 -365 660 -335
rect 660 -365 665 -335
rect 625 -370 665 -365
rect 750 -335 790 -330
rect 750 -365 755 -335
rect 755 -365 785 -335
rect 785 -365 790 -335
rect 750 -370 790 -365
<< metal3 >>
rect -135 295 -85 300
rect -135 255 -130 295
rect -90 255 -85 295
rect -135 250 -85 255
rect 215 295 265 300
rect 215 255 220 295
rect 260 255 265 295
rect 215 250 265 255
rect 390 295 440 300
rect 390 255 395 295
rect 435 255 440 295
rect 390 250 440 255
rect 565 295 615 300
rect 565 255 570 295
rect 610 255 615 295
rect 565 250 615 255
rect 740 295 790 300
rect 740 255 745 295
rect 785 255 790 295
rect 740 250 790 255
rect -130 -330 -80 -325
rect -130 -370 -125 -330
rect -85 -370 -80 -330
rect -130 -375 -80 -370
rect 120 -330 170 -325
rect 120 -370 125 -330
rect 165 -370 170 -330
rect 120 -375 170 -370
rect 245 -330 295 -325
rect 245 -370 250 -330
rect 290 -370 295 -330
rect 245 -375 295 -370
rect 495 -330 545 -325
rect 495 -370 500 -330
rect 540 -370 545 -330
rect 495 -375 545 -370
rect 620 -330 670 -325
rect 620 -370 625 -330
rect 665 -370 670 -330
rect 620 -375 670 -370
rect 745 -330 795 -325
rect 745 -370 750 -330
rect 790 -370 795 -330
rect 745 -375 795 -370
<< via3 >>
rect -130 290 -90 295
rect -130 260 -125 290
rect -125 260 -95 290
rect -95 260 -90 290
rect -130 255 -90 260
rect 220 290 260 295
rect 220 260 225 290
rect 225 260 255 290
rect 255 260 260 290
rect 220 255 260 260
rect 395 290 435 295
rect 395 260 400 290
rect 400 260 430 290
rect 430 260 435 290
rect 395 255 435 260
rect 570 290 610 295
rect 570 260 575 290
rect 575 260 605 290
rect 605 260 610 290
rect 570 255 610 260
rect 745 290 785 295
rect 745 260 750 290
rect 750 260 780 290
rect 780 260 785 290
rect 745 255 785 260
rect -125 -370 -85 -330
rect 125 -370 165 -330
rect 250 -370 290 -330
rect 500 -370 540 -330
rect 625 -370 665 -330
rect 750 -370 790 -330
<< metal4 >>
rect -140 295 -80 305
rect -140 255 -130 295
rect -90 290 -80 295
rect 210 295 270 305
rect 210 290 220 295
rect -90 260 220 290
rect -90 255 -80 260
rect -140 245 -80 255
rect 210 255 220 260
rect 260 290 270 295
rect 385 295 445 305
rect 385 290 395 295
rect 260 260 395 290
rect 260 255 270 260
rect 210 245 270 255
rect 385 255 395 260
rect 435 290 445 295
rect 560 295 620 305
rect 560 290 570 295
rect 435 260 570 290
rect 435 255 445 260
rect 385 245 445 255
rect 560 255 570 260
rect 610 290 620 295
rect 735 295 795 305
rect 735 290 745 295
rect 610 260 745 290
rect 610 255 620 260
rect 560 245 620 255
rect 735 255 745 260
rect 785 290 795 295
rect 785 260 875 290
rect 785 255 795 260
rect 735 245 795 255
rect -135 -330 -75 -320
rect 115 -330 175 -320
rect 240 -330 300 -320
rect 490 -330 550 -320
rect 615 -330 675 -320
rect 740 -330 800 -320
rect -135 -370 -125 -330
rect -85 -360 125 -330
rect -85 -370 -75 -360
rect -135 -380 -75 -370
rect 115 -370 125 -360
rect 165 -360 250 -330
rect 165 -370 175 -360
rect 115 -380 175 -370
rect 240 -370 250 -360
rect 290 -360 500 -330
rect 290 -370 300 -360
rect 240 -380 300 -370
rect 490 -370 500 -360
rect 540 -360 625 -330
rect 540 -370 550 -360
rect 490 -380 550 -370
rect 615 -370 625 -360
rect 665 -360 750 -330
rect 665 -370 675 -360
rect 615 -380 675 -370
rect 740 -370 750 -360
rect 790 -360 875 -330
rect 790 -370 800 -360
rect 740 -380 800 -370
<< labels >>
rlabel metal4 -125 260 875 290 1 VDD
rlabel locali 815 -150 840 -105 1 Qbar
rlabel metal1 760 -80 875 -65 1 Q
rlabel metal1 385 -300 585 -285 1 z5
rlabel metal1 455 -115 495 -100 1 Qbar1
rlabel metal1 560 -115 600 -100 1 Qbar1
rlabel metal1 405 -85 420 -45 1 clk
rlabel metal1 260 -50 325 -35 1 clk
rlabel metal2 -145 15 -130 30 1 clk
rlabel locali 110 -50 250 -30 1 clk
rlabel locali -145 -60 -85 -40 1 D
rlabel metal2 -145 -115 -90 -100 1 R
rlabel locali -60 -150 -40 -115 1 Z2
rlabel metal1 -60 -85 -45 0 1 Z2
rlabel locali -30 55 50 80 1 Z1
rlabel metal1 5 -300 210 -285 1 Z4
rlabel locali 325 -150 345 -85 1 Z3
rlabel locali 530 -125 550 -25 1 Z3
rlabel locali 435 -45 475 -25 1 Z3
rlabel metal4 -120 -360 875 -330 1 GND
<< end >>
