magic
tech sky130A
timestamp 1640012992
<< nwell >>
rect -60 160 500 505
<< nmos >>
rect 10 -10 40 90
rect 205 -10 235 90
rect 400 -10 430 90
<< pmos >>
rect 10 180 40 380
rect 205 180 235 380
rect 400 180 430 380
<< ndiff >>
rect -40 75 10 90
rect -40 5 -25 75
rect -5 5 10 75
rect -40 -10 10 5
rect 40 75 90 90
rect 40 5 55 75
rect 75 5 90 75
rect 40 -10 90 5
rect 155 75 205 90
rect 155 5 170 75
rect 190 5 205 75
rect 155 -10 205 5
rect 235 75 285 90
rect 235 5 250 75
rect 270 5 285 75
rect 235 -10 285 5
rect 350 75 400 90
rect 350 5 365 75
rect 385 5 400 75
rect 350 -10 400 5
rect 430 75 480 90
rect 430 5 445 75
rect 465 5 480 75
rect 430 -10 480 5
<< pdiff >>
rect -40 365 10 380
rect -40 195 -25 365
rect -5 195 10 365
rect -40 180 10 195
rect 40 365 90 380
rect 40 195 55 365
rect 75 195 90 365
rect 40 180 90 195
rect 155 365 205 380
rect 155 195 170 365
rect 190 195 205 365
rect 155 180 205 195
rect 235 365 285 380
rect 235 195 250 365
rect 270 195 285 365
rect 235 180 285 195
rect 350 365 400 380
rect 350 195 365 365
rect 385 195 400 365
rect 350 180 400 195
rect 430 365 480 380
rect 430 195 445 365
rect 465 195 480 365
rect 430 180 480 195
<< ndiffc >>
rect -25 5 -5 75
rect 55 5 75 75
rect 170 5 190 75
rect 250 5 270 75
rect 365 5 385 75
rect 445 5 465 75
<< pdiffc >>
rect -25 195 -5 365
rect 55 195 75 365
rect 170 195 190 365
rect 250 195 270 365
rect 365 195 385 365
rect 445 195 465 365
<< psubdiff >>
rect 100 -60 325 -45
rect 100 -90 115 -60
rect 310 -90 325 -60
rect 100 -100 325 -90
<< nsubdiff >>
rect 120 475 350 485
rect 120 440 135 475
rect 330 440 350 475
rect 120 430 350 440
<< psubdiffcont >>
rect 115 -90 310 -60
<< nsubdiffcont >>
rect 135 440 330 475
<< poly >>
rect 10 380 40 395
rect 205 380 235 395
rect 400 380 430 395
rect 10 150 40 180
rect 205 150 235 180
rect 400 150 430 180
rect -30 140 40 150
rect -30 120 -20 140
rect 0 120 40 140
rect -30 110 40 120
rect 165 140 235 150
rect 165 120 175 140
rect 195 120 235 140
rect 165 110 235 120
rect 360 140 430 150
rect 360 120 370 140
rect 390 120 430 140
rect 360 110 430 120
rect 10 90 40 110
rect 205 90 235 110
rect 400 90 430 110
rect 10 -25 40 -10
rect 205 -25 235 -10
rect 400 -25 430 -10
<< polycont >>
rect -20 120 0 140
rect 175 120 195 140
rect 370 120 390 140
<< locali >>
rect -60 475 500 505
rect -60 440 135 475
rect 330 440 500 475
rect -60 415 500 440
rect -35 365 5 415
rect -35 195 -25 365
rect -5 195 5 365
rect -35 185 5 195
rect 45 365 85 375
rect 45 195 55 365
rect 75 195 85 365
rect -30 145 10 150
rect -30 115 -25 145
rect 5 115 10 145
rect -30 110 10 115
rect 45 145 85 195
rect 160 365 200 415
rect 160 195 170 365
rect 190 195 200 365
rect 160 185 200 195
rect 240 365 280 375
rect 240 195 250 365
rect 270 195 280 365
rect 165 145 205 150
rect 45 140 205 145
rect 45 120 175 140
rect 195 120 205 140
rect 45 115 205 120
rect -35 75 5 85
rect -35 5 -25 75
rect -5 5 5 75
rect -35 -40 5 5
rect 45 75 85 115
rect 165 110 205 115
rect 240 145 280 195
rect 355 365 395 415
rect 355 195 365 365
rect 385 195 395 365
rect 355 185 395 195
rect 435 365 475 375
rect 435 195 445 365
rect 465 195 475 365
rect 360 145 400 150
rect 240 140 400 145
rect 240 120 370 140
rect 390 120 400 140
rect 240 115 400 120
rect 45 5 55 75
rect 75 5 85 75
rect 45 -5 85 5
rect 160 75 200 85
rect 160 5 170 75
rect 190 5 200 75
rect 160 -40 200 5
rect 240 75 280 115
rect 360 110 400 115
rect 240 5 250 75
rect 270 5 280 75
rect 240 -5 280 5
rect 355 75 395 85
rect 355 5 365 75
rect 385 5 395 75
rect 355 -40 395 5
rect 435 75 475 195
rect 435 5 445 75
rect 465 5 475 75
rect 435 -5 475 5
rect -50 -60 500 -40
rect -50 -90 115 -60
rect 310 -90 500 -60
rect -50 -110 500 -90
<< viali >>
rect -25 140 5 145
rect -25 120 -20 140
rect -20 120 0 140
rect 0 120 5 140
rect -25 115 5 120
rect 475 115 505 145
<< metal1 >>
rect -35 150 10 155
rect 470 150 515 155
rect -35 145 515 150
rect -35 115 -25 145
rect 5 115 475 145
rect 505 115 515 145
rect -35 110 515 115
rect -35 105 10 110
rect 470 105 515 110
<< labels >>
rlabel locali 400 450 400 450 1 vdd
rlabel locali 380 -80 380 -80 1 gnd
rlabel viali 490 130 490 130 1 out3
<< end >>
