magic
tech sky130A
magscale 1 2
timestamp 1647891597
<< psubdiff >>
rect 166784 680094 169514 680314
rect 166784 677730 167022 680094
rect 169270 677730 169514 680094
rect 166784 677524 169514 677730
rect 180700 680096 183430 680316
rect 180700 677732 180938 680096
rect 183186 677732 183430 680096
rect 180700 677526 183430 677732
rect 194336 680054 197066 680274
rect 194336 677690 194574 680054
rect 196822 677690 197066 680054
rect 194336 677484 197066 677690
rect 208266 680056 210996 680276
rect 208266 677692 208504 680056
rect 210752 677692 210996 680056
rect 208266 677486 210996 677692
rect 222182 680058 224912 680278
rect 222182 677694 222420 680058
rect 224668 677694 224912 680058
rect 222182 677488 224912 677694
rect 236022 680056 238752 680276
rect 236022 677692 236260 680056
rect 238508 677692 238752 680056
rect 236022 677486 238752 677692
rect 249952 680058 252682 680278
rect 249952 677694 250190 680058
rect 252438 677694 252682 680058
rect 249952 677488 252682 677694
rect 263868 680060 266598 680280
rect 263868 677696 264106 680060
rect 266354 677696 266598 680060
rect 263868 677490 266598 677696
rect 277702 680068 280432 680288
rect 277702 677704 277940 680068
rect 280188 677704 280432 680068
rect 277702 677498 280432 677704
rect 291632 680070 294362 680290
rect 291632 677706 291870 680070
rect 294118 677706 294362 680070
rect 291632 677500 294362 677706
rect 305548 680072 308278 680292
rect 305548 677708 305786 680072
rect 308034 677708 308278 680072
rect 305548 677502 308278 677708
rect 319382 680068 322112 680288
rect 319382 677704 319620 680068
rect 321868 677704 322112 680068
rect 319382 677498 322112 677704
rect 333312 680070 336042 680290
rect 333312 677706 333550 680070
rect 335798 677706 336042 680070
rect 333312 677500 336042 677706
rect 347228 680072 349958 680292
rect 347228 677708 347466 680072
rect 349714 677708 349958 680072
rect 347228 677502 349958 677708
rect 360838 680058 363568 680278
rect 360838 677694 361076 680058
rect 363324 677694 363568 680058
rect 360838 677488 363568 677694
rect 374768 680060 377498 680280
rect 374768 677696 375006 680060
rect 377254 677696 377498 680060
rect 374768 677490 377498 677696
rect 388684 680062 391414 680282
rect 388684 677698 388922 680062
rect 391170 677698 391414 680062
rect 388684 677492 391414 677698
rect 402524 680060 405254 680280
rect 402524 677696 402762 680060
rect 405010 677696 405254 680060
rect 402524 677490 405254 677696
rect 416454 680062 419184 680282
rect 416454 677698 416692 680062
rect 418940 677698 419184 680062
rect 416454 677492 419184 677698
rect 430370 680064 433100 680284
rect 430370 677700 430608 680064
rect 432856 677700 433100 680064
rect 430370 677494 433100 677700
rect 193788 665794 196518 666014
rect 193788 663430 194026 665794
rect 196274 663430 196518 665794
rect 193788 663224 196518 663430
rect 207718 665796 210448 666016
rect 207718 663432 207956 665796
rect 210204 663432 210448 665796
rect 207718 663226 210448 663432
rect 277154 665808 279884 666028
rect 277154 663444 277392 665808
rect 279640 663444 279884 665808
rect 277154 663238 279884 663444
rect 291084 665810 293814 666030
rect 291084 663446 291322 665810
rect 293570 663446 293814 665810
rect 291084 663240 293814 663446
rect 305000 665812 307730 666032
rect 305000 663448 305238 665812
rect 307486 663448 307730 665812
rect 305000 663242 307730 663448
rect 318834 665808 321564 666028
rect 318834 663444 319072 665808
rect 321320 663444 321564 665808
rect 318834 663238 321564 663444
rect 332764 665810 335494 666030
rect 332764 663446 333002 665810
rect 335250 663446 335494 665810
rect 332764 663240 335494 663446
rect 346680 665812 349410 666032
rect 346680 663448 346918 665812
rect 349166 663448 349410 665812
rect 346680 663242 349410 663448
rect 360290 665798 363020 666018
rect 360290 663434 360528 665798
rect 362776 663434 363020 665798
rect 360290 663228 363020 663434
rect 374220 665800 376950 666020
rect 374220 663436 374458 665800
rect 376706 663436 376950 665800
rect 374220 663230 376950 663436
rect 388136 665802 390866 666022
rect 388136 663438 388374 665802
rect 390622 663438 390866 665802
rect 388136 663232 390866 663438
rect 401976 665800 404706 666020
rect 401976 663436 402214 665800
rect 404462 663436 404706 665800
rect 401976 663230 404706 663436
rect 415906 665802 418636 666022
rect 415906 663438 416144 665802
rect 418392 663438 418636 665802
rect 415906 663232 418636 663438
rect 429822 665804 432552 666024
rect 429822 663440 430060 665804
rect 432308 663440 432552 665804
rect 429822 663234 432552 663440
rect 194336 653138 197066 653358
rect 194336 650774 194574 653138
rect 196822 650774 197066 653138
rect 194336 650568 197066 650774
rect 208266 653140 210996 653360
rect 208266 650776 208504 653140
rect 210752 650776 210996 653140
rect 208266 650570 210996 650776
rect 277702 653152 280432 653372
rect 277702 650788 277940 653152
rect 280188 650788 280432 653152
rect 277702 650582 280432 650788
rect 291632 653154 294362 653374
rect 291632 650790 291870 653154
rect 294118 650790 294362 653154
rect 291632 650584 294362 650790
rect 305548 653156 308278 653376
rect 305548 650792 305786 653156
rect 308034 650792 308278 653156
rect 305548 650586 308278 650792
rect 319382 653152 322112 653372
rect 319382 650788 319620 653152
rect 321868 650788 322112 653152
rect 319382 650582 322112 650788
rect 333312 653154 336042 653374
rect 333312 650790 333550 653154
rect 335798 650790 336042 653154
rect 333312 650584 336042 650790
rect 347228 653156 349958 653376
rect 347228 650792 347466 653156
rect 349714 650792 349958 653156
rect 347228 650586 349958 650792
rect 360838 653142 363568 653362
rect 360838 650778 361076 653142
rect 363324 650778 363568 653142
rect 360838 650572 363568 650778
rect 374768 653144 377498 653364
rect 374768 650780 375006 653144
rect 377254 650780 377498 653144
rect 374768 650574 377498 650780
rect 388684 653146 391414 653366
rect 388684 650782 388922 653146
rect 391170 650782 391414 653146
rect 388684 650576 391414 650782
rect 402524 653144 405254 653364
rect 402524 650780 402762 653144
rect 405010 650780 405254 653144
rect 402524 650574 405254 650780
rect 416454 653146 419184 653366
rect 416454 650782 416692 653146
rect 418940 650782 419184 653146
rect 416454 650576 419184 650782
rect 430370 653148 433100 653368
rect 430370 650784 430608 653148
rect 432856 650784 433100 653148
rect 430370 650578 433100 650784
rect 193788 638878 196518 639098
rect 193788 636514 194026 638878
rect 196274 636514 196518 638878
rect 193788 636308 196518 636514
rect 207718 638880 210448 639100
rect 207718 636516 207956 638880
rect 210204 636516 210448 638880
rect 207718 636310 210448 636516
rect 277154 638892 279884 639112
rect 277154 636528 277392 638892
rect 279640 636528 279884 638892
rect 277154 636322 279884 636528
rect 291084 638894 293814 639114
rect 291084 636530 291322 638894
rect 293570 636530 293814 638894
rect 291084 636324 293814 636530
rect 305000 638896 307730 639116
rect 305000 636532 305238 638896
rect 307486 636532 307730 638896
rect 305000 636326 307730 636532
rect 318834 638892 321564 639112
rect 318834 636528 319072 638892
rect 321320 636528 321564 638892
rect 318834 636322 321564 636528
rect 332764 638894 335494 639114
rect 332764 636530 333002 638894
rect 335250 636530 335494 638894
rect 332764 636324 335494 636530
rect 346680 638896 349410 639116
rect 346680 636532 346918 638896
rect 349166 636532 349410 638896
rect 346680 636326 349410 636532
rect 360290 638882 363020 639102
rect 360290 636518 360528 638882
rect 362776 636518 363020 638882
rect 360290 636312 363020 636518
rect 374220 638884 376950 639104
rect 374220 636520 374458 638884
rect 376706 636520 376950 638884
rect 374220 636314 376950 636520
rect 388136 638886 390866 639106
rect 388136 636522 388374 638886
rect 390622 636522 390866 638886
rect 388136 636316 390866 636522
rect 401976 638884 404706 639104
rect 401976 636520 402214 638884
rect 404462 636520 404706 638884
rect 401976 636314 404706 636520
rect 415906 638886 418636 639106
rect 415906 636522 416144 638886
rect 418392 636522 418636 638886
rect 415906 636316 418636 636522
rect 429822 638888 432552 639108
rect 429822 636524 430060 638888
rect 432308 636524 432552 638888
rect 429822 636318 432552 636524
rect 194348 624616 197078 624836
rect 194348 622252 194586 624616
rect 196834 622252 197078 624616
rect 194348 622046 197078 622252
rect 208278 624618 211008 624838
rect 208278 622254 208516 624618
rect 210764 622254 211008 624618
rect 208278 622048 211008 622254
rect 277714 624630 280444 624850
rect 277714 622266 277952 624630
rect 280200 622266 280444 624630
rect 277714 622060 280444 622266
rect 291644 624632 294374 624852
rect 291644 622268 291882 624632
rect 294130 622268 294374 624632
rect 291644 622062 294374 622268
rect 305560 624634 308290 624854
rect 305560 622270 305798 624634
rect 308046 622270 308290 624634
rect 305560 622064 308290 622270
rect 319394 624630 322124 624850
rect 319394 622266 319632 624630
rect 321880 622266 322124 624630
rect 319394 622060 322124 622266
rect 333324 624632 336054 624852
rect 333324 622268 333562 624632
rect 335810 622268 336054 624632
rect 333324 622062 336054 622268
rect 347240 624634 349970 624854
rect 347240 622270 347478 624634
rect 349726 622270 349970 624634
rect 347240 622064 349970 622270
rect 360850 624620 363580 624840
rect 360850 622256 361088 624620
rect 363336 622256 363580 624620
rect 360850 622050 363580 622256
rect 374780 624622 377510 624842
rect 374780 622258 375018 624622
rect 377266 622258 377510 624622
rect 374780 622052 377510 622258
rect 388696 624624 391426 624844
rect 388696 622260 388934 624624
rect 391182 622260 391426 624624
rect 388696 622054 391426 622260
rect 402536 624622 405266 624842
rect 402536 622258 402774 624622
rect 405022 622258 405266 624622
rect 402536 622052 405266 622258
rect 416466 624624 419196 624844
rect 416466 622260 416704 624624
rect 418952 622260 419196 624624
rect 416466 622054 419196 622260
rect 430382 624626 433112 624846
rect 430382 622262 430620 624626
rect 432868 622262 433112 624626
rect 430382 622056 433112 622262
rect 166248 610396 168978 610616
rect 166248 608032 166486 610396
rect 168734 608032 168978 610396
rect 166248 607826 168978 608032
rect 180164 610398 182894 610618
rect 180164 608034 180402 610398
rect 182650 608034 182894 610398
rect 180164 607828 182894 608034
rect 193800 610356 196530 610576
rect 193800 607992 194038 610356
rect 196286 607992 196530 610356
rect 193800 607786 196530 607992
rect 207730 610358 210460 610578
rect 207730 607994 207968 610358
rect 210216 607994 210460 610358
rect 207730 607788 210460 607994
rect 221646 610360 224376 610580
rect 221646 607996 221884 610360
rect 224132 607996 224376 610360
rect 221646 607790 224376 607996
rect 235486 610358 238216 610578
rect 235486 607994 235724 610358
rect 237972 607994 238216 610358
rect 235486 607788 238216 607994
rect 249416 610360 252146 610580
rect 249416 607996 249654 610360
rect 251902 607996 252146 610360
rect 249416 607790 252146 607996
rect 263332 610362 266062 610582
rect 263332 607998 263570 610362
rect 265818 607998 266062 610362
rect 263332 607792 266062 607998
rect 277166 610370 279896 610590
rect 277166 608006 277404 610370
rect 279652 608006 279896 610370
rect 277166 607800 279896 608006
rect 291096 610372 293826 610592
rect 291096 608008 291334 610372
rect 293582 608008 293826 610372
rect 291096 607802 293826 608008
rect 305012 610374 307742 610594
rect 305012 608010 305250 610374
rect 307498 608010 307742 610374
rect 305012 607804 307742 608010
rect 318846 610370 321576 610590
rect 318846 608006 319084 610370
rect 321332 608006 321576 610370
rect 318846 607800 321576 608006
rect 332776 610372 335506 610592
rect 332776 608008 333014 610372
rect 335262 608008 335506 610372
rect 332776 607802 335506 608008
rect 346692 610374 349422 610594
rect 346692 608010 346930 610374
rect 349178 608010 349422 610374
rect 346692 607804 349422 608010
rect 360302 610360 363032 610580
rect 360302 607996 360540 610360
rect 362788 607996 363032 610360
rect 360302 607790 363032 607996
rect 374232 610362 376962 610582
rect 374232 607998 374470 610362
rect 376718 607998 376962 610362
rect 374232 607792 376962 607998
rect 388148 610364 390878 610584
rect 388148 608000 388386 610364
rect 390634 608000 390878 610364
rect 388148 607794 390878 608000
rect 401988 610362 404718 610582
rect 401988 607998 402226 610362
rect 404474 607998 404718 610362
rect 401988 607792 404718 607998
rect 415918 610364 418648 610584
rect 415918 608000 416156 610364
rect 418404 608000 418648 610364
rect 415918 607794 418648 608000
rect 429834 610366 432564 610586
rect 429834 608002 430072 610366
rect 432320 608002 432564 610366
rect 429834 607796 432564 608002
rect 194526 591898 197256 592118
rect 194526 589534 194764 591898
rect 197012 589534 197256 591898
rect 194526 589328 197256 589534
rect 208456 591900 211186 592120
rect 208456 589536 208694 591900
rect 210942 589536 211186 591900
rect 208456 589330 211186 589536
rect 277892 591912 280622 592132
rect 277892 589548 278130 591912
rect 280378 589548 280622 591912
rect 277892 589342 280622 589548
rect 291822 591914 294552 592134
rect 291822 589550 292060 591914
rect 294308 589550 294552 591914
rect 291822 589344 294552 589550
rect 305738 591916 308468 592136
rect 305738 589552 305976 591916
rect 308224 589552 308468 591916
rect 305738 589346 308468 589552
rect 319572 591912 322302 592132
rect 319572 589548 319810 591912
rect 322058 589548 322302 591912
rect 319572 589342 322302 589548
rect 333502 591914 336232 592134
rect 333502 589550 333740 591914
rect 335988 589550 336232 591914
rect 333502 589344 336232 589550
rect 374958 591904 377688 592124
rect 374958 589540 375196 591904
rect 377444 589540 377688 591904
rect 374958 589334 377688 589540
rect 388874 591906 391604 592126
rect 388874 589542 389112 591906
rect 391360 589542 391604 591906
rect 388874 589336 391604 589542
rect 193978 577638 196708 577858
rect 193978 575274 194216 577638
rect 196464 575274 196708 577638
rect 193978 575068 196708 575274
rect 207908 577640 210638 577860
rect 207908 575276 208146 577640
rect 210394 575276 210638 577640
rect 207908 575070 210638 575276
rect 277344 577652 280074 577872
rect 277344 575288 277582 577652
rect 279830 575288 280074 577652
rect 277344 575082 280074 575288
rect 291274 577654 294004 577874
rect 291274 575290 291512 577654
rect 293760 575290 294004 577654
rect 291274 575084 294004 575290
rect 305190 577656 307920 577876
rect 305190 575292 305428 577656
rect 307676 575292 307920 577656
rect 305190 575086 307920 575292
rect 319024 577652 321754 577872
rect 319024 575288 319262 577652
rect 321510 575288 321754 577652
rect 319024 575082 321754 575288
rect 332954 577654 335684 577874
rect 332954 575290 333192 577654
rect 335440 575290 335684 577654
rect 332954 575084 335684 575290
rect 374410 577644 377140 577864
rect 374410 575280 374648 577644
rect 376896 575280 377140 577644
rect 374410 575074 377140 575280
rect 388326 577646 391056 577866
rect 388326 575282 388564 577646
rect 390812 575282 391056 577646
rect 388326 575076 391056 575282
rect 194194 564812 196924 565032
rect 194194 562448 194432 564812
rect 196680 562448 196924 564812
rect 194194 562242 196924 562448
rect 208124 564814 210854 565034
rect 208124 562450 208362 564814
rect 210610 562450 210854 564814
rect 208124 562244 210854 562450
rect 277560 564826 280290 565046
rect 277560 562462 277798 564826
rect 280046 562462 280290 564826
rect 277560 562256 280290 562462
rect 291490 564828 294220 565048
rect 291490 562464 291728 564828
rect 293976 562464 294220 564828
rect 291490 562258 294220 562464
rect 305406 564830 308136 565050
rect 305406 562466 305644 564830
rect 307892 562466 308136 564830
rect 305406 562260 308136 562466
rect 319240 564826 321970 565046
rect 319240 562462 319478 564826
rect 321726 562462 321970 564826
rect 319240 562256 321970 562462
rect 333170 564828 335900 565048
rect 333170 562464 333408 564828
rect 335656 562464 335900 564828
rect 333170 562258 335900 562464
rect 374626 564818 377356 565038
rect 374626 562454 374864 564818
rect 377112 562454 377356 564818
rect 374626 562248 377356 562454
rect 388542 564820 391272 565040
rect 388542 562456 388780 564820
rect 391028 562456 391272 564820
rect 388542 562250 391272 562456
rect 139312 547124 142042 547344
rect 139312 544760 139550 547124
rect 141798 544760 142042 547124
rect 139312 544554 142042 544760
rect 153146 547120 155876 547340
rect 153146 544756 153384 547120
rect 155632 544756 155876 547120
rect 153146 544550 155876 544756
rect 167076 547122 169806 547342
rect 167076 544758 167314 547122
rect 169562 544758 169806 547122
rect 167076 544552 169806 544758
rect 180992 547124 183722 547344
rect 180992 544760 181230 547124
rect 183478 544760 183722 547124
rect 180992 544554 183722 544760
rect 194628 547082 197358 547302
rect 194628 544718 194866 547082
rect 197114 544718 197358 547082
rect 194628 544512 197358 544718
rect 208558 547084 211288 547304
rect 208558 544720 208796 547084
rect 211044 544720 211288 547084
rect 208558 544514 211288 544720
rect 222474 547086 225204 547306
rect 222474 544722 222712 547086
rect 224960 544722 225204 547086
rect 222474 544516 225204 544722
rect 236314 547084 239044 547304
rect 236314 544720 236552 547084
rect 238800 544720 239044 547084
rect 236314 544514 239044 544720
rect 250244 547086 252974 547306
rect 250244 544722 250482 547086
rect 252730 544722 252974 547086
rect 250244 544516 252974 544722
rect 264160 547088 266890 547308
rect 264160 544724 264398 547088
rect 266646 544724 266890 547088
rect 264160 544518 266890 544724
rect 277994 547096 280724 547316
rect 277994 544732 278232 547096
rect 280480 544732 280724 547096
rect 277994 544526 280724 544732
rect 291924 547098 294654 547318
rect 291924 544734 292162 547098
rect 294410 544734 294654 547098
rect 291924 544528 294654 544734
rect 305840 547100 308570 547320
rect 305840 544736 306078 547100
rect 308326 544736 308570 547100
rect 305840 544530 308570 544736
rect 319674 547096 322404 547316
rect 319674 544732 319912 547096
rect 322160 544732 322404 547096
rect 319674 544526 322404 544732
rect 333604 547098 336334 547318
rect 333604 544734 333842 547098
rect 336090 544734 336334 547098
rect 333604 544528 336334 544734
rect 347520 547100 350250 547320
rect 347520 544736 347758 547100
rect 350006 544736 350250 547100
rect 347520 544530 350250 544736
rect 361130 547086 363860 547306
rect 361130 544722 361368 547086
rect 363616 544722 363860 547086
rect 361130 544516 363860 544722
rect 375060 547088 377790 547308
rect 375060 544724 375298 547088
rect 377546 544724 377790 547088
rect 375060 544518 377790 544724
rect 388976 547090 391706 547310
rect 388976 544726 389214 547090
rect 391462 544726 391706 547090
rect 388976 544520 391706 544726
rect 402816 547088 405546 547308
rect 402816 544724 403054 547088
rect 405302 544724 405546 547088
rect 402816 544518 405546 544724
rect 416746 547090 419476 547310
rect 416746 544726 416984 547090
rect 419232 544726 419476 547090
rect 416746 544520 419476 544726
rect 430662 547092 433392 547312
rect 430662 544728 430900 547092
rect 433148 544728 433392 547092
rect 430662 544522 433392 544728
rect 444496 547100 447226 547320
rect 444496 544736 444734 547100
rect 446982 544736 447226 547100
rect 444496 544530 447226 544736
rect 138764 532864 141494 533084
rect 138764 530500 139002 532864
rect 141250 530500 141494 532864
rect 138764 530294 141494 530500
rect 152598 532860 155328 533080
rect 152598 530496 152836 532860
rect 155084 530496 155328 532860
rect 152598 530290 155328 530496
rect 166528 532862 169258 533082
rect 166528 530498 166766 532862
rect 169014 530498 169258 532862
rect 166528 530292 169258 530498
rect 180444 532864 183174 533084
rect 180444 530500 180682 532864
rect 182930 530500 183174 532864
rect 180444 530294 183174 530500
rect 194080 532822 196810 533042
rect 194080 530458 194318 532822
rect 196566 530458 196810 532822
rect 194080 530252 196810 530458
rect 208010 532824 210740 533044
rect 208010 530460 208248 532824
rect 210496 530460 210740 532824
rect 208010 530254 210740 530460
rect 221926 532826 224656 533046
rect 221926 530462 222164 532826
rect 224412 530462 224656 532826
rect 221926 530256 224656 530462
rect 235766 532824 238496 533044
rect 235766 530460 236004 532824
rect 238252 530460 238496 532824
rect 235766 530254 238496 530460
rect 249696 532826 252426 533046
rect 249696 530462 249934 532826
rect 252182 530462 252426 532826
rect 249696 530256 252426 530462
rect 263612 532828 266342 533048
rect 263612 530464 263850 532828
rect 266098 530464 266342 532828
rect 263612 530258 266342 530464
rect 277446 532836 280176 533056
rect 277446 530472 277684 532836
rect 279932 530472 280176 532836
rect 277446 530266 280176 530472
rect 291376 532838 294106 533058
rect 291376 530474 291614 532838
rect 293862 530474 294106 532838
rect 291376 530268 294106 530474
rect 305292 532840 308022 533060
rect 305292 530476 305530 532840
rect 307778 530476 308022 532840
rect 305292 530270 308022 530476
rect 319126 532836 321856 533056
rect 319126 530472 319364 532836
rect 321612 530472 321856 532836
rect 319126 530266 321856 530472
rect 333056 532838 335786 533058
rect 333056 530474 333294 532838
rect 335542 530474 335786 532838
rect 333056 530268 335786 530474
rect 346972 532840 349702 533060
rect 346972 530476 347210 532840
rect 349458 530476 349702 532840
rect 346972 530270 349702 530476
rect 360582 532826 363312 533046
rect 360582 530462 360820 532826
rect 363068 530462 363312 532826
rect 360582 530256 363312 530462
rect 374512 532828 377242 533048
rect 374512 530464 374750 532828
rect 376998 530464 377242 532828
rect 374512 530258 377242 530464
rect 388428 532830 391158 533050
rect 388428 530466 388666 532830
rect 390914 530466 391158 532830
rect 388428 530260 391158 530466
rect 402268 532828 404998 533048
rect 402268 530464 402506 532828
rect 404754 530464 404998 532828
rect 402268 530258 404998 530464
rect 416198 532830 418928 533050
rect 416198 530466 416436 532830
rect 418684 530466 418928 532830
rect 416198 530260 418928 530466
rect 430114 532832 432844 533052
rect 430114 530468 430352 532832
rect 432600 530468 432844 532832
rect 430114 530262 432844 530468
rect 443948 532840 446678 533060
rect 443948 530476 444186 532840
rect 446434 530476 446678 532840
rect 443948 530270 446678 530476
rect 138980 520038 141710 520258
rect 138980 517674 139218 520038
rect 141466 517674 141710 520038
rect 138980 517468 141710 517674
rect 152814 520034 155544 520254
rect 152814 517670 153052 520034
rect 155300 517670 155544 520034
rect 152814 517464 155544 517670
rect 166744 520036 169474 520256
rect 166744 517672 166982 520036
rect 169230 517672 169474 520036
rect 166744 517466 169474 517672
rect 180660 520038 183390 520258
rect 180660 517674 180898 520038
rect 183146 517674 183390 520038
rect 180660 517468 183390 517674
rect 194296 519996 197026 520216
rect 194296 517632 194534 519996
rect 196782 517632 197026 519996
rect 194296 517426 197026 517632
rect 208226 519998 210956 520218
rect 208226 517634 208464 519998
rect 210712 517634 210956 519998
rect 208226 517428 210956 517634
rect 222142 520000 224872 520220
rect 222142 517636 222380 520000
rect 224628 517636 224872 520000
rect 222142 517430 224872 517636
rect 235982 519998 238712 520218
rect 235982 517634 236220 519998
rect 238468 517634 238712 519998
rect 235982 517428 238712 517634
rect 249912 520000 252642 520220
rect 249912 517636 250150 520000
rect 252398 517636 252642 520000
rect 249912 517430 252642 517636
rect 263828 520002 266558 520222
rect 263828 517638 264066 520002
rect 266314 517638 266558 520002
rect 263828 517432 266558 517638
rect 277662 520010 280392 520230
rect 277662 517646 277900 520010
rect 280148 517646 280392 520010
rect 277662 517440 280392 517646
rect 291592 520012 294322 520232
rect 291592 517648 291830 520012
rect 294078 517648 294322 520012
rect 291592 517442 294322 517648
rect 305508 520014 308238 520234
rect 305508 517650 305746 520014
rect 307994 517650 308238 520014
rect 305508 517444 308238 517650
rect 319342 520010 322072 520230
rect 319342 517646 319580 520010
rect 321828 517646 322072 520010
rect 319342 517440 322072 517646
rect 333272 520012 336002 520232
rect 333272 517648 333510 520012
rect 335758 517648 336002 520012
rect 333272 517442 336002 517648
rect 347188 520014 349918 520234
rect 347188 517650 347426 520014
rect 349674 517650 349918 520014
rect 347188 517444 349918 517650
rect 360798 520000 363528 520220
rect 360798 517636 361036 520000
rect 363284 517636 363528 520000
rect 360798 517430 363528 517636
rect 374728 520002 377458 520222
rect 374728 517638 374966 520002
rect 377214 517638 377458 520002
rect 374728 517432 377458 517638
rect 388644 520004 391374 520224
rect 388644 517640 388882 520004
rect 391130 517640 391374 520004
rect 388644 517434 391374 517640
rect 402484 520002 405214 520222
rect 402484 517638 402722 520002
rect 404970 517638 405214 520002
rect 402484 517432 405214 517638
rect 416414 520004 419144 520224
rect 416414 517640 416652 520004
rect 418900 517640 419144 520004
rect 416414 517434 419144 517640
rect 430330 520006 433060 520226
rect 430330 517642 430568 520006
rect 432816 517642 433060 520006
rect 430330 517436 433060 517642
rect 444164 520014 446894 520234
rect 444164 517650 444402 520014
rect 446650 517650 446894 520014
rect 444164 517444 446894 517650
rect 167138 498614 169868 498834
rect 167138 496250 167376 498614
rect 169624 496250 169868 498614
rect 167138 496044 169868 496250
rect 181054 498616 183784 498836
rect 181054 496252 181292 498616
rect 183540 496252 183784 498616
rect 181054 496046 183784 496252
rect 194690 498574 197420 498794
rect 194690 496210 194928 498574
rect 197176 496210 197420 498574
rect 194690 496004 197420 496210
rect 208620 498576 211350 498796
rect 208620 496212 208858 498576
rect 211106 496212 211350 498576
rect 208620 496006 211350 496212
rect 222536 498578 225266 498798
rect 222536 496214 222774 498578
rect 225022 496214 225266 498578
rect 222536 496008 225266 496214
rect 236376 498576 239106 498796
rect 236376 496212 236614 498576
rect 238862 496212 239106 498576
rect 236376 496006 239106 496212
rect 250306 498578 253036 498798
rect 250306 496214 250544 498578
rect 252792 496214 253036 498578
rect 250306 496008 253036 496214
rect 264222 498580 266952 498800
rect 264222 496216 264460 498580
rect 266708 496216 266952 498580
rect 264222 496010 266952 496216
rect 278056 498588 280786 498808
rect 278056 496224 278294 498588
rect 280542 496224 280786 498588
rect 278056 496018 280786 496224
rect 291986 498590 294716 498810
rect 291986 496226 292224 498590
rect 294472 496226 294716 498590
rect 291986 496020 294716 496226
rect 305902 498592 308632 498812
rect 305902 496228 306140 498592
rect 308388 496228 308632 498592
rect 305902 496022 308632 496228
rect 319736 498588 322466 498808
rect 319736 496224 319974 498588
rect 322222 496224 322466 498588
rect 319736 496018 322466 496224
rect 333666 498590 336396 498810
rect 333666 496226 333904 498590
rect 336152 496226 336396 498590
rect 333666 496020 336396 496226
rect 347582 498592 350312 498812
rect 347582 496228 347820 498592
rect 350068 496228 350312 498592
rect 347582 496022 350312 496228
rect 361192 498578 363922 498798
rect 361192 496214 361430 498578
rect 363678 496214 363922 498578
rect 361192 496008 363922 496214
rect 375122 498580 377852 498800
rect 375122 496216 375360 498580
rect 377608 496216 377852 498580
rect 375122 496010 377852 496216
rect 389038 498582 391768 498802
rect 389038 496218 389276 498582
rect 391524 496218 391768 498582
rect 389038 496012 391768 496218
rect 402878 498580 405608 498800
rect 402878 496216 403116 498580
rect 405364 496216 405608 498580
rect 402878 496010 405608 496216
rect 416808 498582 419538 498802
rect 416808 496218 417046 498582
rect 419294 496218 419538 498582
rect 416808 496012 419538 496218
rect 430724 498584 433454 498804
rect 430724 496220 430962 498584
rect 433210 496220 433454 498584
rect 430724 496014 433454 496220
rect 444558 498592 447288 498812
rect 444558 496228 444796 498592
rect 447044 496228 447288 498592
rect 444558 496022 447288 496228
rect 166590 484354 169320 484574
rect 166590 481990 166828 484354
rect 169076 481990 169320 484354
rect 166590 481784 169320 481990
rect 180506 484356 183236 484576
rect 180506 481992 180744 484356
rect 182992 481992 183236 484356
rect 180506 481786 183236 481992
rect 194142 484314 196872 484534
rect 194142 481950 194380 484314
rect 196628 481950 196872 484314
rect 194142 481744 196872 481950
rect 208072 484316 210802 484536
rect 208072 481952 208310 484316
rect 210558 481952 210802 484316
rect 208072 481746 210802 481952
rect 221988 484318 224718 484538
rect 221988 481954 222226 484318
rect 224474 481954 224718 484318
rect 221988 481748 224718 481954
rect 235828 484316 238558 484536
rect 235828 481952 236066 484316
rect 238314 481952 238558 484316
rect 235828 481746 238558 481952
rect 249758 484318 252488 484538
rect 249758 481954 249996 484318
rect 252244 481954 252488 484318
rect 249758 481748 252488 481954
rect 263674 484320 266404 484540
rect 263674 481956 263912 484320
rect 266160 481956 266404 484320
rect 263674 481750 266404 481956
rect 277508 484328 280238 484548
rect 277508 481964 277746 484328
rect 279994 481964 280238 484328
rect 277508 481758 280238 481964
rect 291438 484330 294168 484550
rect 291438 481966 291676 484330
rect 293924 481966 294168 484330
rect 291438 481760 294168 481966
rect 305354 484332 308084 484552
rect 305354 481968 305592 484332
rect 307840 481968 308084 484332
rect 305354 481762 308084 481968
rect 319188 484328 321918 484548
rect 319188 481964 319426 484328
rect 321674 481964 321918 484328
rect 319188 481758 321918 481964
rect 333118 484330 335848 484550
rect 333118 481966 333356 484330
rect 335604 481966 335848 484330
rect 333118 481760 335848 481966
rect 347034 484332 349764 484552
rect 347034 481968 347272 484332
rect 349520 481968 349764 484332
rect 347034 481762 349764 481968
rect 360644 484318 363374 484538
rect 360644 481954 360882 484318
rect 363130 481954 363374 484318
rect 360644 481748 363374 481954
rect 374574 484320 377304 484540
rect 374574 481956 374812 484320
rect 377060 481956 377304 484320
rect 374574 481750 377304 481956
rect 388490 484322 391220 484542
rect 388490 481958 388728 484322
rect 390976 481958 391220 484322
rect 388490 481752 391220 481958
rect 402330 484320 405060 484540
rect 402330 481956 402568 484320
rect 404816 481956 405060 484320
rect 402330 481750 405060 481956
rect 416260 484322 418990 484542
rect 416260 481958 416498 484322
rect 418746 481958 418990 484322
rect 416260 481752 418990 481958
rect 430176 484324 432906 484544
rect 430176 481960 430414 484324
rect 432662 481960 432906 484324
rect 430176 481754 432906 481960
rect 444010 484332 446740 484552
rect 444010 481968 444248 484332
rect 446496 481968 446740 484332
rect 444010 481762 446740 481968
rect 166806 471528 169536 471748
rect 166806 469164 167044 471528
rect 169292 469164 169536 471528
rect 166806 468958 169536 469164
rect 180722 471530 183452 471750
rect 180722 469166 180960 471530
rect 183208 469166 183452 471530
rect 180722 468960 183452 469166
rect 194358 471488 197088 471708
rect 194358 469124 194596 471488
rect 196844 469124 197088 471488
rect 194358 468918 197088 469124
rect 208288 471490 211018 471710
rect 208288 469126 208526 471490
rect 210774 469126 211018 471490
rect 208288 468920 211018 469126
rect 222204 471492 224934 471712
rect 222204 469128 222442 471492
rect 224690 469128 224934 471492
rect 222204 468922 224934 469128
rect 236044 471490 238774 471710
rect 236044 469126 236282 471490
rect 238530 469126 238774 471490
rect 236044 468920 238774 469126
rect 249974 471492 252704 471712
rect 249974 469128 250212 471492
rect 252460 469128 252704 471492
rect 249974 468922 252704 469128
rect 263890 471494 266620 471714
rect 263890 469130 264128 471494
rect 266376 469130 266620 471494
rect 263890 468924 266620 469130
rect 277724 471502 280454 471722
rect 277724 469138 277962 471502
rect 280210 469138 280454 471502
rect 277724 468932 280454 469138
rect 291654 471504 294384 471724
rect 291654 469140 291892 471504
rect 294140 469140 294384 471504
rect 291654 468934 294384 469140
rect 305570 471506 308300 471726
rect 305570 469142 305808 471506
rect 308056 469142 308300 471506
rect 305570 468936 308300 469142
rect 319404 471502 322134 471722
rect 319404 469138 319642 471502
rect 321890 469138 322134 471502
rect 319404 468932 322134 469138
rect 333334 471504 336064 471724
rect 333334 469140 333572 471504
rect 335820 469140 336064 471504
rect 333334 468934 336064 469140
rect 347250 471506 349980 471726
rect 347250 469142 347488 471506
rect 349736 469142 349980 471506
rect 347250 468936 349980 469142
rect 360860 471492 363590 471712
rect 360860 469128 361098 471492
rect 363346 469128 363590 471492
rect 360860 468922 363590 469128
rect 374790 471494 377520 471714
rect 374790 469130 375028 471494
rect 377276 469130 377520 471494
rect 374790 468924 377520 469130
rect 388706 471496 391436 471716
rect 388706 469132 388944 471496
rect 391192 469132 391436 471496
rect 388706 468926 391436 469132
rect 402546 471494 405276 471714
rect 402546 469130 402784 471494
rect 405032 469130 405276 471494
rect 402546 468924 405276 469130
rect 416476 471496 419206 471716
rect 416476 469132 416714 471496
rect 418962 469132 419206 471496
rect 416476 468926 419206 469132
rect 430392 471498 433122 471718
rect 430392 469134 430630 471498
rect 432878 469134 433122 471498
rect 430392 468928 433122 469134
rect 444226 471506 446956 471726
rect 444226 469142 444464 471506
rect 446712 469142 446956 471506
rect 444226 468936 446956 469142
rect 139622 458084 142352 458304
rect 139622 455720 139860 458084
rect 142108 455720 142352 458084
rect 139622 455514 142352 455720
rect 153456 458080 156186 458300
rect 153456 455716 153694 458080
rect 155942 455716 156186 458080
rect 153456 455510 156186 455716
rect 167386 458082 170116 458302
rect 167386 455718 167624 458082
rect 169872 455718 170116 458082
rect 167386 455512 170116 455718
rect 181302 458084 184032 458304
rect 181302 455720 181540 458084
rect 183788 455720 184032 458084
rect 181302 455514 184032 455720
rect 194938 458042 197668 458262
rect 194938 455678 195176 458042
rect 197424 455678 197668 458042
rect 194938 455472 197668 455678
rect 208868 458044 211598 458264
rect 208868 455680 209106 458044
rect 211354 455680 211598 458044
rect 208868 455474 211598 455680
rect 222784 458046 225514 458266
rect 222784 455682 223022 458046
rect 225270 455682 225514 458046
rect 222784 455476 225514 455682
rect 236624 458044 239354 458264
rect 236624 455680 236862 458044
rect 239110 455680 239354 458044
rect 236624 455474 239354 455680
rect 250554 458046 253284 458266
rect 250554 455682 250792 458046
rect 253040 455682 253284 458046
rect 250554 455476 253284 455682
rect 264470 458048 267200 458268
rect 264470 455684 264708 458048
rect 266956 455684 267200 458048
rect 264470 455478 267200 455684
rect 278304 458056 281034 458276
rect 278304 455692 278542 458056
rect 280790 455692 281034 458056
rect 278304 455486 281034 455692
rect 292234 458058 294964 458278
rect 292234 455694 292472 458058
rect 294720 455694 294964 458058
rect 292234 455488 294964 455694
rect 306150 458060 308880 458280
rect 306150 455696 306388 458060
rect 308636 455696 308880 458060
rect 306150 455490 308880 455696
rect 319984 458056 322714 458276
rect 319984 455692 320222 458056
rect 322470 455692 322714 458056
rect 319984 455486 322714 455692
rect 333914 458058 336644 458278
rect 333914 455694 334152 458058
rect 336400 455694 336644 458058
rect 333914 455488 336644 455694
rect 347830 458060 350560 458280
rect 347830 455696 348068 458060
rect 350316 455696 350560 458060
rect 347830 455490 350560 455696
rect 361440 458046 364170 458266
rect 361440 455682 361678 458046
rect 363926 455682 364170 458046
rect 361440 455476 364170 455682
rect 375370 458048 378100 458268
rect 375370 455684 375608 458048
rect 377856 455684 378100 458048
rect 375370 455478 378100 455684
rect 389286 458050 392016 458270
rect 389286 455686 389524 458050
rect 391772 455686 392016 458050
rect 389286 455480 392016 455686
rect 403126 458048 405856 458268
rect 403126 455684 403364 458048
rect 405612 455684 405856 458048
rect 403126 455478 405856 455684
rect 417056 458050 419786 458270
rect 417056 455686 417294 458050
rect 419542 455686 419786 458050
rect 417056 455480 419786 455686
rect 430972 458052 433702 458272
rect 430972 455688 431210 458052
rect 433458 455688 433702 458052
rect 430972 455482 433702 455688
rect 444806 458060 447536 458280
rect 444806 455696 445044 458060
rect 447292 455696 447536 458060
rect 444806 455490 447536 455696
rect 139582 446360 142312 446580
rect 139582 443996 139820 446360
rect 142068 443996 142312 446360
rect 139582 443790 142312 443996
rect 153416 446356 156146 446576
rect 153416 443992 153654 446356
rect 155902 443992 156146 446356
rect 153416 443786 156146 443992
rect 167346 446358 170076 446578
rect 167346 443994 167584 446358
rect 169832 443994 170076 446358
rect 167346 443788 170076 443994
rect 181262 446360 183992 446580
rect 181262 443996 181500 446360
rect 183748 443996 183992 446360
rect 181262 443790 183992 443996
rect 194898 446318 197628 446538
rect 194898 443954 195136 446318
rect 197384 443954 197628 446318
rect 194898 443748 197628 443954
rect 208828 446320 211558 446540
rect 208828 443956 209066 446320
rect 211314 443956 211558 446320
rect 208828 443750 211558 443956
rect 222744 446322 225474 446542
rect 222744 443958 222982 446322
rect 225230 443958 225474 446322
rect 222744 443752 225474 443958
rect 236584 446320 239314 446540
rect 236584 443956 236822 446320
rect 239070 443956 239314 446320
rect 236584 443750 239314 443956
rect 250514 446322 253244 446542
rect 250514 443958 250752 446322
rect 253000 443958 253244 446322
rect 250514 443752 253244 443958
rect 264430 446324 267160 446544
rect 264430 443960 264668 446324
rect 266916 443960 267160 446324
rect 264430 443754 267160 443960
rect 278264 446332 280994 446552
rect 278264 443968 278502 446332
rect 280750 443968 280994 446332
rect 278264 443762 280994 443968
rect 292194 446334 294924 446554
rect 292194 443970 292432 446334
rect 294680 443970 294924 446334
rect 292194 443764 294924 443970
rect 306110 446336 308840 446556
rect 306110 443972 306348 446336
rect 308596 443972 308840 446336
rect 306110 443766 308840 443972
rect 319944 446332 322674 446552
rect 319944 443968 320182 446332
rect 322430 443968 322674 446332
rect 319944 443762 322674 443968
rect 333874 446334 336604 446554
rect 333874 443970 334112 446334
rect 336360 443970 336604 446334
rect 333874 443764 336604 443970
rect 347790 446336 350520 446556
rect 347790 443972 348028 446336
rect 350276 443972 350520 446336
rect 347790 443766 350520 443972
rect 361400 446322 364130 446542
rect 361400 443958 361638 446322
rect 363886 443958 364130 446322
rect 361400 443752 364130 443958
rect 375330 446324 378060 446544
rect 375330 443960 375568 446324
rect 377816 443960 378060 446324
rect 375330 443754 378060 443960
rect 389246 446326 391976 446546
rect 389246 443962 389484 446326
rect 391732 443962 391976 446326
rect 389246 443756 391976 443962
rect 403086 446324 405816 446544
rect 403086 443960 403324 446324
rect 405572 443960 405816 446324
rect 403086 443754 405816 443960
rect 417016 446326 419746 446546
rect 417016 443962 417254 446326
rect 419502 443962 419746 446326
rect 417016 443756 419746 443962
rect 430932 446328 433662 446548
rect 430932 443964 431170 446328
rect 433418 443964 433662 446328
rect 430932 443758 433662 443964
rect 444766 446336 447496 446556
rect 444766 443972 445004 446336
rect 447252 443972 447496 446336
rect 444766 443766 447496 443972
rect 42380 422218 45110 422438
rect 42380 419854 42618 422218
rect 44866 419854 45110 422218
rect 42380 419648 45110 419854
rect 56296 422220 59026 422440
rect 56296 419856 56534 422220
rect 58782 419856 59026 422220
rect 56296 419650 59026 419856
rect 70136 422218 72866 422438
rect 70136 419854 70374 422218
rect 72622 419854 72866 422218
rect 70136 419648 72866 419854
rect 84066 422220 86796 422440
rect 84066 419856 84304 422220
rect 86552 419856 86796 422220
rect 84066 419650 86796 419856
rect 97982 422222 100712 422442
rect 97982 419858 98220 422222
rect 100468 419858 100712 422222
rect 97982 419652 100712 419858
rect 111816 422230 114546 422450
rect 111816 419866 112054 422230
rect 114302 419866 114546 422230
rect 111816 419660 114546 419866
rect 125746 422232 128476 422452
rect 125746 419868 125984 422232
rect 128232 419868 128476 422232
rect 125746 419662 128476 419868
rect 194978 422192 197708 422412
rect 194978 419828 195216 422192
rect 197464 419828 197708 422192
rect 194978 419622 197708 419828
rect 208908 422194 211638 422414
rect 208908 419830 209146 422194
rect 211394 419830 211638 422194
rect 208908 419624 211638 419830
rect 278344 422206 281074 422426
rect 278344 419842 278582 422206
rect 280830 419842 281074 422206
rect 278344 419636 281074 419842
rect 292274 422208 295004 422428
rect 292274 419844 292512 422208
rect 294760 419844 295004 422208
rect 292274 419638 295004 419844
rect 306190 422210 308920 422430
rect 306190 419846 306428 422210
rect 308676 419846 308920 422210
rect 306190 419640 308920 419846
rect 320024 422206 322754 422426
rect 320024 419842 320262 422206
rect 322510 419842 322754 422206
rect 320024 419636 322754 419842
rect 333954 422208 336684 422428
rect 333954 419844 334192 422208
rect 336440 419844 336684 422208
rect 333954 419638 336684 419844
rect 528652 422214 531382 422434
rect 528652 419850 528890 422214
rect 531138 419850 531382 422214
rect 528652 419644 531382 419850
rect 542568 422216 545298 422436
rect 542568 419852 542806 422216
rect 545054 419852 545298 422216
rect 542568 419646 545298 419852
rect 41832 407958 44562 408178
rect 41832 405594 42070 407958
rect 44318 405594 44562 407958
rect 41832 405388 44562 405594
rect 55748 407960 58478 408180
rect 55748 405596 55986 407960
rect 58234 405596 58478 407960
rect 55748 405390 58478 405596
rect 69588 407958 72318 408178
rect 69588 405594 69826 407958
rect 72074 405594 72318 407958
rect 69588 405388 72318 405594
rect 83518 407960 86248 408180
rect 83518 405596 83756 407960
rect 86004 405596 86248 407960
rect 83518 405390 86248 405596
rect 97434 407962 100164 408182
rect 97434 405598 97672 407962
rect 99920 405598 100164 407962
rect 97434 405392 100164 405598
rect 111268 407970 113998 408190
rect 111268 405606 111506 407970
rect 113754 405606 113998 407970
rect 111268 405400 113998 405606
rect 125198 407972 127928 408192
rect 125198 405608 125436 407972
rect 127684 405608 127928 407972
rect 125198 405402 127928 405608
rect 194430 407932 197160 408152
rect 194430 405568 194668 407932
rect 196916 405568 197160 407932
rect 194430 405362 197160 405568
rect 208360 407934 211090 408154
rect 208360 405570 208598 407934
rect 210846 405570 211090 407934
rect 208360 405364 211090 405570
rect 277796 407946 280526 408166
rect 277796 405582 278034 407946
rect 280282 405582 280526 407946
rect 277796 405376 280526 405582
rect 291726 407948 294456 408168
rect 291726 405584 291964 407948
rect 294212 405584 294456 407948
rect 291726 405378 294456 405584
rect 305642 407950 308372 408170
rect 305642 405586 305880 407950
rect 308128 405586 308372 407950
rect 305642 405380 308372 405586
rect 319476 407946 322206 408166
rect 319476 405582 319714 407946
rect 321962 405582 322206 407946
rect 319476 405376 322206 405582
rect 333406 407948 336136 408168
rect 333406 405584 333644 407948
rect 335892 405584 336136 407948
rect 333406 405378 336136 405584
rect 528104 407954 530834 408174
rect 528104 405590 528342 407954
rect 530590 405590 530834 407954
rect 528104 405384 530834 405590
rect 542020 407956 544750 408176
rect 542020 405592 542258 407956
rect 544506 405592 544750 407956
rect 542020 405386 544750 405592
rect 42048 395132 44778 395352
rect 42048 392768 42286 395132
rect 44534 392768 44778 395132
rect 42048 392562 44778 392768
rect 55964 395134 58694 395354
rect 55964 392770 56202 395134
rect 58450 392770 58694 395134
rect 55964 392564 58694 392770
rect 69804 395132 72534 395352
rect 69804 392768 70042 395132
rect 72290 392768 72534 395132
rect 69804 392562 72534 392768
rect 83734 395134 86464 395354
rect 83734 392770 83972 395134
rect 86220 392770 86464 395134
rect 83734 392564 86464 392770
rect 97650 395136 100380 395356
rect 97650 392772 97888 395136
rect 100136 392772 100380 395136
rect 97650 392566 100380 392772
rect 111484 395144 114214 395364
rect 111484 392780 111722 395144
rect 113970 392780 114214 395144
rect 111484 392574 114214 392780
rect 125414 395146 128144 395366
rect 125414 392782 125652 395146
rect 127900 392782 128144 395146
rect 125414 392576 128144 392782
rect 194646 395106 197376 395326
rect 194646 392742 194884 395106
rect 197132 392742 197376 395106
rect 194646 392536 197376 392742
rect 208576 395108 211306 395328
rect 208576 392744 208814 395108
rect 211062 392744 211306 395108
rect 208576 392538 211306 392744
rect 278012 395120 280742 395340
rect 278012 392756 278250 395120
rect 280498 392756 280742 395120
rect 278012 392550 280742 392756
rect 291942 395122 294672 395342
rect 291942 392758 292180 395122
rect 294428 392758 294672 395122
rect 291942 392552 294672 392758
rect 305858 395124 308588 395344
rect 305858 392760 306096 395124
rect 308344 392760 308588 395124
rect 305858 392554 308588 392760
rect 319692 395120 322422 395340
rect 319692 392756 319930 395120
rect 322178 392756 322422 395120
rect 319692 392550 322422 392756
rect 333622 395122 336352 395342
rect 333622 392758 333860 395122
rect 336108 392758 336352 395122
rect 333622 392552 336352 392758
rect 528320 395128 531050 395348
rect 528320 392764 528558 395128
rect 530806 392764 531050 395128
rect 528320 392558 531050 392764
rect 542236 395130 544966 395350
rect 542236 392766 542474 395130
rect 544722 392766 544966 395130
rect 542236 392560 544966 392766
rect 194952 386406 197682 386626
rect 194952 384042 195190 386406
rect 197438 384042 197682 386406
rect 194952 383836 197682 384042
rect 208882 386408 211612 386628
rect 208882 384044 209120 386408
rect 211368 384044 211612 386408
rect 208882 383838 211612 384044
rect 278318 386420 281048 386640
rect 278318 384056 278556 386420
rect 280804 384056 281048 386420
rect 278318 383850 281048 384056
rect 292248 386422 294978 386642
rect 292248 384058 292486 386422
rect 294734 384058 294978 386422
rect 292248 383852 294978 384058
rect 306164 386424 308894 386644
rect 306164 384060 306402 386424
rect 308650 384060 308894 386424
rect 306164 383854 308894 384060
rect 319998 386420 322728 386640
rect 319998 384056 320236 386420
rect 322484 384056 322728 386420
rect 319998 383850 322728 384056
rect 333928 386422 336658 386642
rect 333928 384058 334166 386422
rect 336414 384058 336658 386422
rect 333928 383852 336658 384058
rect 528626 386428 531356 386648
rect 528626 384064 528864 386428
rect 531112 384064 531356 386428
rect 528626 383858 531356 384064
rect 542542 386430 545272 386650
rect 542542 384066 542780 386430
rect 545028 384066 545272 386430
rect 542542 383860 545272 384066
rect 152922 372184 155652 372404
rect 152922 369820 153160 372184
rect 155408 369820 155652 372184
rect 152922 369614 155652 369820
rect 166852 372186 169582 372406
rect 166852 369822 167090 372186
rect 169338 369822 169582 372186
rect 166852 369616 169582 369822
rect 180768 372188 183498 372408
rect 180768 369824 181006 372188
rect 183254 369824 183498 372188
rect 180768 369618 183498 369824
rect 194404 372146 197134 372366
rect 194404 369782 194642 372146
rect 196890 369782 197134 372146
rect 194404 369576 197134 369782
rect 208334 372148 211064 372368
rect 208334 369784 208572 372148
rect 210820 369784 211064 372148
rect 208334 369578 211064 369784
rect 277770 372160 280500 372380
rect 277770 369796 278008 372160
rect 280256 369796 280500 372160
rect 277770 369590 280500 369796
rect 291700 372162 294430 372382
rect 291700 369798 291938 372162
rect 294186 369798 294430 372162
rect 291700 369592 294430 369798
rect 305616 372164 308346 372384
rect 305616 369800 305854 372164
rect 308102 369800 308346 372164
rect 305616 369594 308346 369800
rect 319450 372160 322180 372380
rect 319450 369796 319688 372160
rect 321936 369796 322180 372160
rect 319450 369590 322180 369796
rect 333380 372162 336110 372382
rect 333380 369798 333618 372162
rect 335866 369798 336110 372162
rect 333380 369592 336110 369798
rect 347296 372164 350026 372384
rect 347296 369800 347534 372164
rect 349782 369800 350026 372164
rect 347296 369594 350026 369800
rect 360906 372150 363636 372370
rect 360906 369786 361144 372150
rect 363392 369786 363636 372150
rect 360906 369580 363636 369786
rect 374836 372152 377566 372372
rect 374836 369788 375074 372152
rect 377322 369788 377566 372152
rect 374836 369582 377566 369788
rect 388752 372154 391482 372374
rect 388752 369790 388990 372154
rect 391238 369790 391482 372154
rect 388752 369584 391482 369790
rect 402592 372152 405322 372372
rect 402592 369788 402830 372152
rect 405078 369788 405322 372152
rect 402592 369582 405322 369788
rect 416522 372154 419252 372374
rect 416522 369790 416760 372154
rect 419008 369790 419252 372154
rect 416522 369584 419252 369790
rect 430438 372156 433168 372376
rect 430438 369792 430676 372156
rect 432924 369792 433168 372156
rect 430438 369586 433168 369792
rect 444272 372164 447002 372384
rect 444272 369800 444510 372164
rect 446758 369800 447002 372164
rect 444272 369594 447002 369800
rect 458202 372166 460932 372386
rect 458202 369802 458440 372166
rect 460688 369802 460932 372166
rect 458202 369596 460932 369802
rect 472118 372168 474848 372388
rect 472118 369804 472356 372168
rect 474604 369804 474848 372168
rect 472118 369598 474848 369804
rect 485952 372164 488682 372384
rect 485952 369800 486190 372164
rect 488438 369800 488682 372164
rect 485952 369594 488682 369800
rect 499882 372166 502612 372386
rect 499882 369802 500120 372166
rect 502368 369802 502612 372166
rect 499882 369596 502612 369802
rect 513798 372168 516528 372388
rect 513798 369804 514036 372168
rect 516284 369804 516528 372168
rect 513798 369598 516528 369804
rect 528078 372168 530808 372388
rect 528078 369804 528316 372168
rect 530564 369804 530808 372168
rect 528078 369598 530808 369804
rect 541994 372170 544724 372390
rect 541994 369806 542232 372170
rect 544480 369806 544724 372170
rect 541994 369600 544724 369806
rect 556266 372150 558996 372370
rect 556266 369786 556504 372150
rect 558752 369786 558996 372150
rect 556266 369580 558996 369786
rect 153138 359358 155868 359578
rect 153138 356994 153376 359358
rect 155624 356994 155868 359358
rect 153138 356788 155868 356994
rect 167068 359360 169798 359580
rect 167068 356996 167306 359360
rect 169554 356996 169798 359360
rect 167068 356790 169798 356996
rect 180984 359362 183714 359582
rect 180984 356998 181222 359362
rect 183470 356998 183714 359362
rect 180984 356792 183714 356998
rect 194620 359320 197350 359540
rect 194620 356956 194858 359320
rect 197106 356956 197350 359320
rect 194620 356750 197350 356956
rect 208550 359322 211280 359542
rect 208550 356958 208788 359322
rect 211036 356958 211280 359322
rect 208550 356752 211280 356958
rect 222466 359324 225196 359544
rect 222466 356960 222704 359324
rect 224952 356960 225196 359324
rect 222466 356754 225196 356960
rect 236306 359322 239036 359542
rect 236306 356958 236544 359322
rect 238792 356958 239036 359322
rect 236306 356752 239036 356958
rect 250236 359324 252966 359544
rect 250236 356960 250474 359324
rect 252722 356960 252966 359324
rect 250236 356754 252966 356960
rect 264152 359326 266882 359546
rect 264152 356962 264390 359326
rect 266638 356962 266882 359326
rect 264152 356756 266882 356962
rect 277986 359334 280716 359554
rect 277986 356970 278224 359334
rect 280472 356970 280716 359334
rect 277986 356764 280716 356970
rect 291916 359336 294646 359556
rect 291916 356972 292154 359336
rect 294402 356972 294646 359336
rect 291916 356766 294646 356972
rect 305832 359338 308562 359558
rect 305832 356974 306070 359338
rect 308318 356974 308562 359338
rect 305832 356768 308562 356974
rect 319666 359334 322396 359554
rect 319666 356970 319904 359334
rect 322152 356970 322396 359334
rect 319666 356764 322396 356970
rect 333596 359336 336326 359556
rect 333596 356972 333834 359336
rect 336082 356972 336326 359336
rect 333596 356766 336326 356972
rect 347512 359338 350242 359558
rect 347512 356974 347750 359338
rect 349998 356974 350242 359338
rect 347512 356768 350242 356974
rect 361122 359324 363852 359544
rect 361122 356960 361360 359324
rect 363608 356960 363852 359324
rect 361122 356754 363852 356960
rect 375052 359326 377782 359546
rect 375052 356962 375290 359326
rect 377538 356962 377782 359326
rect 375052 356756 377782 356962
rect 388968 359328 391698 359548
rect 388968 356964 389206 359328
rect 391454 356964 391698 359328
rect 388968 356758 391698 356964
rect 402808 359326 405538 359546
rect 402808 356962 403046 359326
rect 405294 356962 405538 359326
rect 402808 356756 405538 356962
rect 416738 359328 419468 359548
rect 416738 356964 416976 359328
rect 419224 356964 419468 359328
rect 416738 356758 419468 356964
rect 430654 359330 433384 359550
rect 430654 356966 430892 359330
rect 433140 356966 433384 359330
rect 430654 356760 433384 356966
rect 444488 359338 447218 359558
rect 444488 356974 444726 359338
rect 446974 356974 447218 359338
rect 444488 356768 447218 356974
rect 458418 359340 461148 359560
rect 458418 356976 458656 359340
rect 460904 356976 461148 359340
rect 458418 356770 461148 356976
rect 472334 359342 475064 359562
rect 472334 356978 472572 359342
rect 474820 356978 475064 359342
rect 472334 356772 475064 356978
rect 486168 359338 488898 359558
rect 486168 356974 486406 359338
rect 488654 356974 488898 359338
rect 486168 356768 488898 356974
rect 500098 359340 502828 359560
rect 500098 356976 500336 359340
rect 502584 356976 502828 359340
rect 500098 356770 502828 356976
rect 514014 359342 516744 359562
rect 514014 356978 514252 359342
rect 516500 356978 516744 359342
rect 514014 356772 516744 356978
rect 528294 359342 531024 359562
rect 528294 356978 528532 359342
rect 530780 356978 531024 359342
rect 528294 356772 531024 356978
rect 542210 359344 544940 359564
rect 542210 356980 542448 359344
rect 544696 356980 544940 359344
rect 542210 356774 544940 356980
rect 556482 359324 559212 359544
rect 556482 356960 556720 359324
rect 558968 356960 559212 359324
rect 556482 356754 559212 356960
rect 138734 347534 141464 347754
rect 138734 345170 138972 347534
rect 141220 345170 141464 347534
rect 138734 344964 141464 345170
rect 152568 347530 155298 347750
rect 152568 345166 152806 347530
rect 155054 345166 155298 347530
rect 152568 344960 155298 345166
rect 166498 347532 169228 347752
rect 166498 345168 166736 347532
rect 168984 345168 169228 347532
rect 166498 344962 169228 345168
rect 180414 347534 183144 347754
rect 180414 345170 180652 347534
rect 182900 345170 183144 347534
rect 180414 344964 183144 345170
rect 194050 347492 196780 347712
rect 194050 345128 194288 347492
rect 196536 345128 196780 347492
rect 194050 344922 196780 345128
rect 207980 347494 210710 347714
rect 207980 345130 208218 347494
rect 210466 345130 210710 347494
rect 207980 344924 210710 345130
rect 221896 347496 224626 347716
rect 221896 345132 222134 347496
rect 224382 345132 224626 347496
rect 221896 344926 224626 345132
rect 235736 347494 238466 347714
rect 235736 345130 235974 347494
rect 238222 345130 238466 347494
rect 235736 344924 238466 345130
rect 249666 347496 252396 347716
rect 249666 345132 249904 347496
rect 252152 345132 252396 347496
rect 249666 344926 252396 345132
rect 263582 347498 266312 347718
rect 263582 345134 263820 347498
rect 266068 345134 266312 347498
rect 263582 344928 266312 345134
rect 277416 347506 280146 347726
rect 277416 345142 277654 347506
rect 279902 345142 280146 347506
rect 277416 344936 280146 345142
rect 291346 347508 294076 347728
rect 291346 345144 291584 347508
rect 293832 345144 294076 347508
rect 291346 344938 294076 345144
rect 305262 347510 307992 347730
rect 305262 345146 305500 347510
rect 307748 345146 307992 347510
rect 305262 344940 307992 345146
rect 319096 347506 321826 347726
rect 319096 345142 319334 347506
rect 321582 345142 321826 347506
rect 319096 344936 321826 345142
rect 333026 347508 335756 347728
rect 333026 345144 333264 347508
rect 335512 345144 335756 347508
rect 333026 344938 335756 345144
rect 346942 347510 349672 347730
rect 346942 345146 347180 347510
rect 349428 345146 349672 347510
rect 346942 344940 349672 345146
rect 360552 347496 363282 347716
rect 360552 345132 360790 347496
rect 363038 345132 363282 347496
rect 360552 344926 363282 345132
rect 374482 347498 377212 347718
rect 374482 345134 374720 347498
rect 376968 345134 377212 347498
rect 374482 344928 377212 345134
rect 388398 347500 391128 347720
rect 388398 345136 388636 347500
rect 390884 345136 391128 347500
rect 388398 344930 391128 345136
rect 402238 347498 404968 347718
rect 402238 345134 402476 347498
rect 404724 345134 404968 347498
rect 402238 344928 404968 345134
rect 416168 347500 418898 347720
rect 416168 345136 416406 347500
rect 418654 345136 418898 347500
rect 416168 344930 418898 345136
rect 430084 347502 432814 347722
rect 430084 345138 430322 347502
rect 432570 345138 432814 347502
rect 430084 344932 432814 345138
rect 443918 347510 446648 347730
rect 443918 345146 444156 347510
rect 446404 345146 446648 347510
rect 443918 344940 446648 345146
rect 457848 347512 460578 347732
rect 457848 345148 458086 347512
rect 460334 345148 460578 347512
rect 457848 344942 460578 345148
rect 471764 347514 474494 347734
rect 471764 345150 472002 347514
rect 474250 345150 474494 347514
rect 471764 344944 474494 345150
rect 485598 347510 488328 347730
rect 485598 345146 485836 347510
rect 488084 345146 488328 347510
rect 485598 344940 488328 345146
rect 499528 347512 502258 347732
rect 499528 345148 499766 347512
rect 502014 345148 502258 347512
rect 499528 344942 502258 345148
rect 513444 347514 516174 347734
rect 513444 345150 513682 347514
rect 515930 345150 516174 347514
rect 513444 344944 516174 345150
rect 527724 347514 530454 347734
rect 527724 345150 527962 347514
rect 530210 345150 530454 347514
rect 527724 344944 530454 345150
rect 541640 347516 544370 347736
rect 541640 345152 541878 347516
rect 544126 345152 544370 347516
rect 541640 344946 544370 345152
rect 555912 347496 558642 347716
rect 555912 345132 556150 347496
rect 558398 345132 558642 347496
rect 555912 344926 558642 345132
rect 138950 334708 141680 334928
rect 138950 332344 139188 334708
rect 141436 332344 141680 334708
rect 138950 332138 141680 332344
rect 152784 334704 155514 334924
rect 152784 332340 153022 334704
rect 155270 332340 155514 334704
rect 152784 332134 155514 332340
rect 166714 334706 169444 334926
rect 166714 332342 166952 334706
rect 169200 332342 169444 334706
rect 166714 332136 169444 332342
rect 180630 334708 183360 334928
rect 180630 332344 180868 334708
rect 183116 332344 183360 334708
rect 180630 332138 183360 332344
rect 194266 334666 196996 334886
rect 194266 332302 194504 334666
rect 196752 332302 196996 334666
rect 194266 332096 196996 332302
rect 208196 334668 210926 334888
rect 208196 332304 208434 334668
rect 210682 332304 210926 334668
rect 208196 332098 210926 332304
rect 222112 334670 224842 334890
rect 222112 332306 222350 334670
rect 224598 332306 224842 334670
rect 222112 332100 224842 332306
rect 235952 334668 238682 334888
rect 235952 332304 236190 334668
rect 238438 332304 238682 334668
rect 235952 332098 238682 332304
rect 249882 334670 252612 334890
rect 249882 332306 250120 334670
rect 252368 332306 252612 334670
rect 249882 332100 252612 332306
rect 263798 334672 266528 334892
rect 263798 332308 264036 334672
rect 266284 332308 266528 334672
rect 263798 332102 266528 332308
rect 277632 334680 280362 334900
rect 277632 332316 277870 334680
rect 280118 332316 280362 334680
rect 277632 332110 280362 332316
rect 291562 334682 294292 334902
rect 291562 332318 291800 334682
rect 294048 332318 294292 334682
rect 291562 332112 294292 332318
rect 305478 334684 308208 334904
rect 305478 332320 305716 334684
rect 307964 332320 308208 334684
rect 305478 332114 308208 332320
rect 319312 334680 322042 334900
rect 319312 332316 319550 334680
rect 321798 332316 322042 334680
rect 319312 332110 322042 332316
rect 333242 334682 335972 334902
rect 333242 332318 333480 334682
rect 335728 332318 335972 334682
rect 333242 332112 335972 332318
rect 347158 334684 349888 334904
rect 347158 332320 347396 334684
rect 349644 332320 349888 334684
rect 347158 332114 349888 332320
rect 360768 334670 363498 334890
rect 360768 332306 361006 334670
rect 363254 332306 363498 334670
rect 360768 332100 363498 332306
rect 374698 334672 377428 334892
rect 374698 332308 374936 334672
rect 377184 332308 377428 334672
rect 374698 332102 377428 332308
rect 388614 334674 391344 334894
rect 388614 332310 388852 334674
rect 391100 332310 391344 334674
rect 388614 332104 391344 332310
rect 402454 334672 405184 334892
rect 402454 332308 402692 334672
rect 404940 332308 405184 334672
rect 402454 332102 405184 332308
rect 416384 334674 419114 334894
rect 416384 332310 416622 334674
rect 418870 332310 419114 334674
rect 416384 332104 419114 332310
rect 430300 334676 433030 334896
rect 430300 332312 430538 334676
rect 432786 332312 433030 334676
rect 430300 332106 433030 332312
rect 444134 334684 446864 334904
rect 444134 332320 444372 334684
rect 446620 332320 446864 334684
rect 444134 332114 446864 332320
rect 458064 334686 460794 334906
rect 458064 332322 458302 334686
rect 460550 332322 460794 334686
rect 458064 332116 460794 332322
rect 471980 334688 474710 334908
rect 471980 332324 472218 334688
rect 474466 332324 474710 334688
rect 471980 332118 474710 332324
rect 485814 334684 488544 334904
rect 485814 332320 486052 334684
rect 488300 332320 488544 334684
rect 485814 332114 488544 332320
rect 499744 334686 502474 334906
rect 499744 332322 499982 334686
rect 502230 332322 502474 334686
rect 499744 332116 502474 332322
rect 513660 334688 516390 334908
rect 513660 332324 513898 334688
rect 516146 332324 516390 334688
rect 513660 332118 516390 332324
rect 527940 334688 530670 334908
rect 527940 332324 528178 334688
rect 530426 332324 530670 334688
rect 527940 332118 530670 332324
rect 541856 334690 544586 334910
rect 541856 332326 542094 334690
rect 544342 332326 544586 334690
rect 541856 332120 544586 332326
rect 556128 334670 558858 334890
rect 556128 332306 556366 334670
rect 558614 332306 558858 334670
rect 556128 332100 558858 332306
rect 43202 320014 45932 320234
rect 43202 317650 43440 320014
rect 45688 317650 45932 320014
rect 43202 317444 45932 317650
rect 57118 320016 59848 320236
rect 57118 317652 57356 320016
rect 59604 317652 59848 320016
rect 57118 317446 59848 317652
rect 70958 320014 73688 320234
rect 70958 317650 71196 320014
rect 73444 317650 73688 320014
rect 70958 317444 73688 317650
rect 112638 320026 115368 320246
rect 112638 317662 112876 320026
rect 115124 317662 115368 320026
rect 112638 317456 115368 317662
rect 126568 320028 129298 320248
rect 126568 317664 126806 320028
rect 129054 317664 129298 320028
rect 126568 317458 129298 317664
rect 195800 319988 198530 320208
rect 195800 317624 196038 319988
rect 198286 317624 198530 319988
rect 195800 317418 198530 317624
rect 209730 319990 212460 320210
rect 209730 317626 209968 319990
rect 212216 317626 212460 319990
rect 209730 317420 212460 317626
rect 279166 320002 281896 320222
rect 279166 317638 279404 320002
rect 281652 317638 281896 320002
rect 279166 317432 281896 317638
rect 293096 320004 295826 320224
rect 293096 317640 293334 320004
rect 295582 317640 295826 320004
rect 293096 317434 295826 317640
rect 307012 320006 309742 320226
rect 307012 317642 307250 320006
rect 309498 317642 309742 320006
rect 307012 317436 309742 317642
rect 320846 320002 323576 320222
rect 320846 317638 321084 320002
rect 323332 317638 323576 320002
rect 320846 317432 323576 317638
rect 334776 320004 337506 320224
rect 334776 317640 335014 320004
rect 337262 317640 337506 320004
rect 334776 317434 337506 317640
rect 376232 319994 378962 320214
rect 376232 317630 376470 319994
rect 378718 317630 378962 319994
rect 376232 317424 378962 317630
rect 390148 319996 392878 320216
rect 390148 317632 390386 319996
rect 392634 317632 392878 319996
rect 390148 317426 392878 317632
rect 459346 319996 462076 320216
rect 459346 317632 459584 319996
rect 461832 317632 462076 319996
rect 459346 317426 462076 317632
rect 473276 319998 476006 320218
rect 473276 317634 473514 319998
rect 475762 317634 476006 319998
rect 473276 317428 476006 317634
rect 487192 320000 489922 320220
rect 487192 317636 487430 320000
rect 489678 317636 489922 320000
rect 487192 317430 489922 317636
rect 501026 320008 503756 320228
rect 501026 317644 501264 320008
rect 503512 317644 503756 320008
rect 501026 317438 503756 317644
rect 514810 319974 517540 320194
rect 514810 317610 515048 319974
rect 517296 317610 517540 319974
rect 514810 317404 517540 317610
rect 528740 319976 531470 320196
rect 528740 317612 528978 319976
rect 531226 317612 531470 319976
rect 528740 317406 531470 317612
rect 542656 319978 545386 320198
rect 542656 317614 542894 319978
rect 545142 317614 545386 319978
rect 542656 317408 545386 317614
rect 556490 319986 559220 320206
rect 556490 317622 556728 319986
rect 558976 317622 559220 319986
rect 556490 317416 559220 317622
rect 43772 310348 46502 310568
rect 43772 307984 44010 310348
rect 46258 307984 46502 310348
rect 43772 307778 46502 307984
rect 57688 310350 60418 310570
rect 57688 307986 57926 310350
rect 60174 307986 60418 310350
rect 57688 307780 60418 307986
rect 71528 310348 74258 310568
rect 71528 307984 71766 310348
rect 74014 307984 74258 310348
rect 71528 307778 74258 307984
rect 113208 310360 115938 310580
rect 113208 307996 113446 310360
rect 115694 307996 115938 310360
rect 113208 307790 115938 307996
rect 127138 310362 129868 310582
rect 127138 307998 127376 310362
rect 129624 307998 129868 310362
rect 127138 307792 129868 307998
rect 196370 310322 199100 310542
rect 196370 307958 196608 310322
rect 198856 307958 199100 310322
rect 196370 307752 199100 307958
rect 210300 310324 213030 310544
rect 210300 307960 210538 310324
rect 212786 307960 213030 310324
rect 210300 307754 213030 307960
rect 279736 310336 282466 310556
rect 279736 307972 279974 310336
rect 282222 307972 282466 310336
rect 279736 307766 282466 307972
rect 293666 310338 296396 310558
rect 293666 307974 293904 310338
rect 296152 307974 296396 310338
rect 293666 307768 296396 307974
rect 307582 310340 310312 310560
rect 307582 307976 307820 310340
rect 310068 307976 310312 310340
rect 307582 307770 310312 307976
rect 321416 310336 324146 310556
rect 321416 307972 321654 310336
rect 323902 307972 324146 310336
rect 321416 307766 324146 307972
rect 335346 310338 338076 310558
rect 335346 307974 335584 310338
rect 337832 307974 338076 310338
rect 335346 307768 338076 307974
rect 376802 310328 379532 310548
rect 376802 307964 377040 310328
rect 379288 307964 379532 310328
rect 376802 307758 379532 307964
rect 390718 310330 393448 310550
rect 390718 307966 390956 310330
rect 393204 307966 393448 310330
rect 390718 307760 393448 307966
rect 459916 310330 462646 310550
rect 459916 307966 460154 310330
rect 462402 307966 462646 310330
rect 459916 307760 462646 307966
rect 473846 310332 476576 310552
rect 473846 307968 474084 310332
rect 476332 307968 476576 310332
rect 473846 307762 476576 307968
rect 487762 310334 490492 310554
rect 487762 307970 488000 310334
rect 490248 307970 490492 310334
rect 487762 307764 490492 307970
rect 501596 310342 504326 310562
rect 501596 307978 501834 310342
rect 504082 307978 504326 310342
rect 501596 307772 504326 307978
rect 515380 310308 518110 310528
rect 515380 307944 515618 310308
rect 517866 307944 518110 310308
rect 515380 307738 518110 307944
rect 529310 310310 532040 310530
rect 529310 307946 529548 310310
rect 531796 307946 532040 310310
rect 529310 307740 532040 307946
rect 543226 310312 545956 310532
rect 543226 307948 543464 310312
rect 545712 307948 545956 310312
rect 543226 307742 545956 307948
rect 557060 310320 559790 310540
rect 557060 307956 557298 310320
rect 559546 307956 559790 310320
rect 557060 307750 559790 307956
rect 43914 299828 46644 300048
rect 43914 297464 44152 299828
rect 46400 297464 46644 299828
rect 43914 297258 46644 297464
rect 57830 299830 60560 300050
rect 57830 297466 58068 299830
rect 60316 297466 60560 299830
rect 57830 297260 60560 297466
rect 71670 299828 74400 300048
rect 71670 297464 71908 299828
rect 74156 297464 74400 299828
rect 71670 297258 74400 297464
rect 113350 299840 116080 300060
rect 113350 297476 113588 299840
rect 115836 297476 116080 299840
rect 113350 297270 116080 297476
rect 127280 299842 130010 300062
rect 127280 297478 127518 299842
rect 129766 297478 130010 299842
rect 127280 297272 130010 297478
rect 196512 299802 199242 300022
rect 196512 297438 196750 299802
rect 198998 297438 199242 299802
rect 196512 297232 199242 297438
rect 210442 299804 213172 300024
rect 210442 297440 210680 299804
rect 212928 297440 213172 299804
rect 210442 297234 213172 297440
rect 279878 299816 282608 300036
rect 279878 297452 280116 299816
rect 282364 297452 282608 299816
rect 279878 297246 282608 297452
rect 293808 299818 296538 300038
rect 293808 297454 294046 299818
rect 296294 297454 296538 299818
rect 293808 297248 296538 297454
rect 307724 299820 310454 300040
rect 307724 297456 307962 299820
rect 310210 297456 310454 299820
rect 307724 297250 310454 297456
rect 321558 299816 324288 300036
rect 321558 297452 321796 299816
rect 324044 297452 324288 299816
rect 321558 297246 324288 297452
rect 335488 299818 338218 300038
rect 335488 297454 335726 299818
rect 337974 297454 338218 299818
rect 335488 297248 338218 297454
rect 376944 299808 379674 300028
rect 376944 297444 377182 299808
rect 379430 297444 379674 299808
rect 376944 297238 379674 297444
rect 390860 299810 393590 300030
rect 390860 297446 391098 299810
rect 393346 297446 393590 299810
rect 390860 297240 393590 297446
rect 460058 299810 462788 300030
rect 460058 297446 460296 299810
rect 462544 297446 462788 299810
rect 460058 297240 462788 297446
rect 473988 299812 476718 300032
rect 473988 297448 474226 299812
rect 476474 297448 476718 299812
rect 473988 297242 476718 297448
rect 487904 299814 490634 300034
rect 487904 297450 488142 299814
rect 490390 297450 490634 299814
rect 487904 297244 490634 297450
rect 501738 299822 504468 300042
rect 501738 297458 501976 299822
rect 504224 297458 504468 299822
rect 501738 297252 504468 297458
rect 515522 299788 518252 300008
rect 515522 297424 515760 299788
rect 518008 297424 518252 299788
rect 515522 297218 518252 297424
rect 529452 299790 532182 300010
rect 529452 297426 529690 299790
rect 531938 297426 532182 299790
rect 529452 297220 532182 297426
rect 543368 299792 546098 300012
rect 543368 297428 543606 299792
rect 545854 297428 546098 299792
rect 543368 297222 546098 297428
rect 557202 299800 559932 300020
rect 557202 297436 557440 299800
rect 559688 297436 559932 299800
rect 557202 297230 559932 297436
rect 43772 288880 46502 289100
rect 43772 286516 44010 288880
rect 46258 286516 46502 288880
rect 43772 286310 46502 286516
rect 57688 288882 60418 289102
rect 57688 286518 57926 288882
rect 60174 286518 60418 288882
rect 57688 286312 60418 286518
rect 71528 288880 74258 289100
rect 71528 286516 71766 288880
rect 74014 286516 74258 288880
rect 71528 286310 74258 286516
rect 113208 288892 115938 289112
rect 113208 286528 113446 288892
rect 115694 286528 115938 288892
rect 113208 286322 115938 286528
rect 127138 288894 129868 289114
rect 127138 286530 127376 288894
rect 129624 286530 129868 288894
rect 127138 286324 129868 286530
rect 196370 288854 199100 289074
rect 196370 286490 196608 288854
rect 198856 286490 199100 288854
rect 196370 286284 199100 286490
rect 210300 288856 213030 289076
rect 210300 286492 210538 288856
rect 212786 286492 213030 288856
rect 210300 286286 213030 286492
rect 279736 288868 282466 289088
rect 279736 286504 279974 288868
rect 282222 286504 282466 288868
rect 279736 286298 282466 286504
rect 293666 288870 296396 289090
rect 293666 286506 293904 288870
rect 296152 286506 296396 288870
rect 293666 286300 296396 286506
rect 307582 288872 310312 289092
rect 307582 286508 307820 288872
rect 310068 286508 310312 288872
rect 307582 286302 310312 286508
rect 321416 288868 324146 289088
rect 321416 286504 321654 288868
rect 323902 286504 324146 288868
rect 321416 286298 324146 286504
rect 335346 288870 338076 289090
rect 335346 286506 335584 288870
rect 337832 286506 338076 288870
rect 335346 286300 338076 286506
rect 376802 288860 379532 289080
rect 376802 286496 377040 288860
rect 379288 286496 379532 288860
rect 376802 286290 379532 286496
rect 390718 288862 393448 289082
rect 390718 286498 390956 288862
rect 393204 286498 393448 288862
rect 390718 286292 393448 286498
rect 44056 276656 46786 276876
rect 44056 274292 44294 276656
rect 46542 274292 46786 276656
rect 44056 274086 46786 274292
rect 57972 276658 60702 276878
rect 57972 274294 58210 276658
rect 60458 274294 60702 276658
rect 57972 274088 60702 274294
rect 71812 276656 74542 276876
rect 71812 274292 72050 276656
rect 74298 274292 74542 276656
rect 71812 274086 74542 274292
rect 113492 276668 116222 276888
rect 113492 274304 113730 276668
rect 115978 274304 116222 276668
rect 113492 274098 116222 274304
rect 127422 276670 130152 276890
rect 127422 274306 127660 276670
rect 129908 274306 130152 276670
rect 127422 274100 130152 274306
rect 196654 276630 199384 276850
rect 196654 274266 196892 276630
rect 199140 274266 199384 276630
rect 196654 274060 199384 274266
rect 210584 276632 213314 276852
rect 210584 274268 210822 276632
rect 213070 274268 213314 276632
rect 210584 274062 213314 274268
rect 280020 276644 282750 276864
rect 280020 274280 280258 276644
rect 282506 274280 282750 276644
rect 280020 274074 282750 274280
rect 293950 276646 296680 276866
rect 293950 274282 294188 276646
rect 296436 274282 296680 276646
rect 293950 274076 296680 274282
rect 307866 276648 310596 276868
rect 307866 274284 308104 276648
rect 310352 274284 310596 276648
rect 307866 274078 310596 274284
rect 321700 276644 324430 276864
rect 321700 274280 321938 276644
rect 324186 274280 324430 276644
rect 321700 274074 324430 274280
rect 335630 276646 338360 276866
rect 335630 274282 335868 276646
rect 338116 274282 338360 276646
rect 335630 274076 338360 274282
rect 377086 276636 379816 276856
rect 377086 274272 377324 276636
rect 379572 274272 379816 276636
rect 377086 274066 379816 274272
rect 391002 276638 393732 276858
rect 391002 274274 391240 276638
rect 393488 274274 393732 276638
rect 391002 274068 393732 274274
rect 43636 260908 46366 261128
rect 43636 258544 43874 260908
rect 46122 258544 46366 260908
rect 43636 258338 46366 258544
rect 57552 260910 60282 261130
rect 57552 258546 57790 260910
rect 60038 258546 60282 260910
rect 57552 258340 60282 258546
rect 71392 260908 74122 261128
rect 71392 258544 71630 260908
rect 73878 258544 74122 260908
rect 71392 258338 74122 258544
rect 85322 260910 88052 261130
rect 85322 258546 85560 260910
rect 87808 258546 88052 260910
rect 85322 258340 88052 258546
rect 99238 260912 101968 261132
rect 99238 258548 99476 260912
rect 101724 258548 101968 260912
rect 99238 258342 101968 258548
rect 113072 260920 115802 261140
rect 113072 258556 113310 260920
rect 115558 258556 115802 260920
rect 113072 258350 115802 258556
rect 127002 260922 129732 261142
rect 127002 258558 127240 260922
rect 129488 258558 129732 260922
rect 127002 258352 129732 258558
rect 140918 260924 143648 261144
rect 140918 258560 141156 260924
rect 143404 258560 143648 260924
rect 140918 258354 143648 258560
rect 154752 260920 157482 261140
rect 154752 258556 154990 260920
rect 157238 258556 157482 260920
rect 154752 258350 157482 258556
rect 168682 260922 171412 261142
rect 168682 258558 168920 260922
rect 171168 258558 171412 260922
rect 168682 258352 171412 258558
rect 182598 260924 185328 261144
rect 182598 258560 182836 260924
rect 185084 258560 185328 260924
rect 182598 258354 185328 258560
rect 196234 260882 198964 261102
rect 196234 258518 196472 260882
rect 198720 258518 198964 260882
rect 196234 258312 198964 258518
rect 210164 260884 212894 261104
rect 210164 258520 210402 260884
rect 212650 258520 212894 260884
rect 210164 258314 212894 258520
rect 224080 260886 226810 261106
rect 224080 258522 224318 260886
rect 226566 258522 226810 260886
rect 224080 258316 226810 258522
rect 237920 260884 240650 261104
rect 237920 258520 238158 260884
rect 240406 258520 240650 260884
rect 237920 258314 240650 258520
rect 251850 260886 254580 261106
rect 251850 258522 252088 260886
rect 254336 258522 254580 260886
rect 251850 258316 254580 258522
rect 265766 260888 268496 261108
rect 265766 258524 266004 260888
rect 268252 258524 268496 260888
rect 265766 258318 268496 258524
rect 279600 260896 282330 261116
rect 279600 258532 279838 260896
rect 282086 258532 282330 260896
rect 279600 258326 282330 258532
rect 293530 260898 296260 261118
rect 293530 258534 293768 260898
rect 296016 258534 296260 260898
rect 293530 258328 296260 258534
rect 307446 260900 310176 261120
rect 307446 258536 307684 260900
rect 309932 258536 310176 260900
rect 307446 258330 310176 258536
rect 321280 260896 324010 261116
rect 321280 258532 321518 260896
rect 323766 258532 324010 260896
rect 321280 258326 324010 258532
rect 335210 260898 337940 261118
rect 335210 258534 335448 260898
rect 337696 258534 337940 260898
rect 335210 258328 337940 258534
rect 349126 260900 351856 261120
rect 349126 258536 349364 260900
rect 351612 258536 351856 260900
rect 349126 258330 351856 258536
rect 362736 260886 365466 261106
rect 362736 258522 362974 260886
rect 365222 258522 365466 260886
rect 362736 258316 365466 258522
rect 376666 260888 379396 261108
rect 376666 258524 376904 260888
rect 379152 258524 379396 260888
rect 376666 258318 379396 258524
rect 390582 260890 393312 261110
rect 390582 258526 390820 260890
rect 393068 258526 393312 260890
rect 390582 258320 393312 258526
rect 195268 238250 197998 238470
rect 195268 235886 195506 238250
rect 197754 235886 197998 238250
rect 195268 235680 197998 235886
rect 209198 238252 211928 238472
rect 209198 235888 209436 238252
rect 211684 235888 211928 238252
rect 209198 235682 211928 235888
rect 278634 238264 281364 238484
rect 278634 235900 278872 238264
rect 281120 235900 281364 238264
rect 278634 235694 281364 235900
rect 292564 238266 295294 238486
rect 292564 235902 292802 238266
rect 295050 235902 295294 238266
rect 292564 235696 295294 235902
rect 306480 238268 309210 238488
rect 306480 235904 306718 238268
rect 308966 235904 309210 238268
rect 306480 235698 309210 235904
rect 320314 238264 323044 238484
rect 320314 235900 320552 238264
rect 322800 235900 323044 238264
rect 320314 235694 323044 235900
rect 334244 238266 336974 238486
rect 334244 235902 334482 238266
rect 336730 235902 336974 238266
rect 334244 235696 336974 235902
rect 195678 222346 198408 222566
rect 195678 219982 195916 222346
rect 198164 219982 198408 222346
rect 195678 219776 198408 219982
rect 209608 222348 212338 222568
rect 209608 219984 209846 222348
rect 212094 219984 212338 222348
rect 209608 219778 212338 219984
rect 279044 222360 281774 222580
rect 279044 219996 279282 222360
rect 281530 219996 281774 222360
rect 279044 219790 281774 219996
rect 292974 222362 295704 222582
rect 292974 219998 293212 222362
rect 295460 219998 295704 222362
rect 292974 219792 295704 219998
rect 306890 222364 309620 222584
rect 306890 220000 307128 222364
rect 309376 220000 309620 222364
rect 306890 219794 309620 220000
rect 320724 222360 323454 222580
rect 320724 219996 320962 222360
rect 323210 219996 323454 222360
rect 320724 219790 323454 219996
rect 334654 222362 337384 222582
rect 334654 219998 334892 222362
rect 337140 219998 337384 222362
rect 334654 219792 337384 219998
rect 195678 205894 198408 206114
rect 195678 203530 195916 205894
rect 198164 203530 198408 205894
rect 195678 203324 198408 203530
rect 209608 205896 212338 206116
rect 209608 203532 209846 205896
rect 212094 203532 212338 205896
rect 209608 203326 212338 203532
rect 279044 205908 281774 206128
rect 279044 203544 279282 205908
rect 281530 203544 281774 205908
rect 279044 203338 281774 203544
rect 292974 205910 295704 206130
rect 292974 203546 293212 205910
rect 295460 203546 295704 205910
rect 292974 203340 295704 203546
rect 306890 205912 309620 206132
rect 306890 203548 307128 205912
rect 309376 203548 309620 205912
rect 306890 203342 309620 203548
rect 320724 205908 323454 206128
rect 320724 203544 320962 205908
rect 323210 203544 323454 205908
rect 320724 203338 323454 203544
rect 334654 205910 337384 206130
rect 334654 203546 334892 205910
rect 337140 203546 337384 205910
rect 334654 203340 337384 203546
rect 195268 191086 197998 191306
rect 195268 188722 195506 191086
rect 197754 188722 197998 191086
rect 195268 188516 197998 188722
rect 209198 191088 211928 191308
rect 209198 188724 209436 191088
rect 211684 188724 211928 191088
rect 209198 188518 211928 188724
rect 278634 191100 281364 191320
rect 278634 188736 278872 191100
rect 281120 188736 281364 191100
rect 278634 188530 281364 188736
rect 292564 191102 295294 191322
rect 292564 188738 292802 191102
rect 295050 188738 295294 191102
rect 292564 188532 295294 188738
rect 306480 191104 309210 191324
rect 306480 188740 306718 191104
rect 308966 188740 309210 191104
rect 306480 188534 309210 188740
rect 320314 191100 323044 191320
rect 320314 188736 320552 191100
rect 322800 188736 323044 191100
rect 320314 188530 323044 188736
rect 334244 191102 336974 191322
rect 334244 188738 334482 191102
rect 336730 188738 336974 191102
rect 334244 188532 336974 188738
rect 194720 176826 197450 177046
rect 194720 174462 194958 176826
rect 197206 174462 197450 176826
rect 194720 174256 197450 174462
rect 208650 176828 211380 177048
rect 208650 174464 208888 176828
rect 211136 174464 211380 176828
rect 208650 174258 211380 174464
rect 222566 176830 225296 177050
rect 222566 174466 222804 176830
rect 225052 174466 225296 176830
rect 222566 174260 225296 174466
rect 236406 176828 239136 177048
rect 236406 174464 236644 176828
rect 238892 174464 239136 176828
rect 236406 174258 239136 174464
rect 250336 176830 253066 177050
rect 250336 174466 250574 176830
rect 252822 174466 253066 176830
rect 250336 174260 253066 174466
rect 264252 176832 266982 177052
rect 264252 174468 264490 176832
rect 266738 174468 266982 176832
rect 264252 174262 266982 174468
rect 278086 176840 280816 177060
rect 278086 174476 278324 176840
rect 280572 174476 280816 176840
rect 278086 174270 280816 174476
rect 292016 176842 294746 177062
rect 292016 174478 292254 176842
rect 294502 174478 294746 176842
rect 292016 174272 294746 174478
rect 305932 176844 308662 177064
rect 305932 174480 306170 176844
rect 308418 174480 308662 176844
rect 305932 174274 308662 174480
rect 319766 176840 322496 177060
rect 319766 174476 320004 176840
rect 322252 174476 322496 176840
rect 319766 174270 322496 174476
rect 333696 176842 336426 177062
rect 333696 174478 333934 176842
rect 336182 174478 336426 176842
rect 333696 174272 336426 174478
rect 194936 164000 197666 164220
rect 194936 161636 195174 164000
rect 197422 161636 197666 164000
rect 194936 161430 197666 161636
rect 208866 164002 211596 164222
rect 208866 161638 209104 164002
rect 211352 161638 211596 164002
rect 208866 161432 211596 161638
rect 222782 164004 225512 164224
rect 222782 161640 223020 164004
rect 225268 161640 225512 164004
rect 222782 161434 225512 161640
rect 236622 164002 239352 164222
rect 236622 161638 236860 164002
rect 239108 161638 239352 164002
rect 236622 161432 239352 161638
rect 250552 164004 253282 164224
rect 250552 161640 250790 164004
rect 253038 161640 253282 164004
rect 250552 161434 253282 161640
rect 264468 164006 267198 164226
rect 264468 161642 264706 164006
rect 266954 161642 267198 164006
rect 264468 161436 267198 161642
rect 278302 164014 281032 164234
rect 278302 161650 278540 164014
rect 280788 161650 281032 164014
rect 278302 161444 281032 161650
rect 292232 164016 294962 164236
rect 292232 161652 292470 164016
rect 294718 161652 294962 164016
rect 292232 161446 294962 161652
rect 306148 164018 308878 164238
rect 306148 161654 306386 164018
rect 308634 161654 308878 164018
rect 306148 161448 308878 161654
rect 319982 164014 322712 164234
rect 319982 161650 320220 164014
rect 322468 161650 322712 164014
rect 319982 161444 322712 161650
rect 333912 164016 336642 164236
rect 333912 161652 334150 164016
rect 336398 161652 336642 164016
rect 333912 161446 336642 161652
rect 42070 141666 44800 141886
rect 42070 139302 42308 141666
rect 44556 139302 44800 141666
rect 42070 139096 44800 139302
rect 55986 141668 58716 141888
rect 55986 139304 56224 141668
rect 58472 139304 58716 141668
rect 55986 139098 58716 139304
rect 69826 141666 72556 141886
rect 69826 139302 70064 141666
rect 72312 139302 72556 141666
rect 69826 139096 72556 139302
rect 83756 141668 86486 141888
rect 83756 139304 83994 141668
rect 86242 139304 86486 141668
rect 83756 139098 86486 139304
rect 97672 141670 100402 141890
rect 97672 139306 97910 141670
rect 100158 139306 100402 141670
rect 97672 139100 100402 139306
rect 111506 141678 114236 141898
rect 111506 139314 111744 141678
rect 113992 139314 114236 141678
rect 111506 139108 114236 139314
rect 125436 141680 128166 141900
rect 125436 139316 125674 141680
rect 127922 139316 128166 141680
rect 125436 139110 128166 139316
rect 139352 141682 142082 141902
rect 139352 139318 139590 141682
rect 141838 139318 142082 141682
rect 139352 139112 142082 139318
rect 153186 141678 155916 141898
rect 153186 139314 153424 141678
rect 155672 139314 155916 141678
rect 153186 139108 155916 139314
rect 167116 141680 169846 141900
rect 167116 139316 167354 141680
rect 169602 139316 169846 141680
rect 167116 139110 169846 139316
rect 181032 141682 183762 141902
rect 181032 139318 181270 141682
rect 183518 139318 183762 141682
rect 181032 139112 183762 139318
rect 194668 141640 197398 141860
rect 194668 139276 194906 141640
rect 197154 139276 197398 141640
rect 194668 139070 197398 139276
rect 208598 141642 211328 141862
rect 208598 139278 208836 141642
rect 211084 139278 211328 141642
rect 208598 139072 211328 139278
rect 222514 141644 225244 141864
rect 222514 139280 222752 141644
rect 225000 139280 225244 141644
rect 222514 139074 225244 139280
rect 236354 141642 239084 141862
rect 236354 139278 236592 141642
rect 238840 139278 239084 141642
rect 236354 139072 239084 139278
rect 250284 141644 253014 141864
rect 250284 139280 250522 141644
rect 252770 139280 253014 141644
rect 250284 139074 253014 139280
rect 264200 141646 266930 141866
rect 264200 139282 264438 141646
rect 266686 139282 266930 141646
rect 264200 139076 266930 139282
rect 278034 141654 280764 141874
rect 278034 139290 278272 141654
rect 280520 139290 280764 141654
rect 278034 139084 280764 139290
rect 291964 141656 294694 141876
rect 291964 139292 292202 141656
rect 294450 139292 294694 141656
rect 291964 139086 294694 139292
rect 305880 141658 308610 141878
rect 305880 139294 306118 141658
rect 308366 139294 308610 141658
rect 305880 139088 308610 139294
rect 319714 141654 322444 141874
rect 319714 139290 319952 141654
rect 322200 139290 322444 141654
rect 319714 139084 322444 139290
rect 333644 141656 336374 141876
rect 333644 139292 333882 141656
rect 336130 139292 336374 141656
rect 333644 139086 336374 139292
rect 347560 141658 350290 141878
rect 347560 139294 347798 141658
rect 350046 139294 350290 141658
rect 347560 139088 350290 139294
rect 42000 129186 44730 129406
rect 42000 126822 42238 129186
rect 44486 126822 44730 129186
rect 42000 126616 44730 126822
rect 55916 129188 58646 129408
rect 55916 126824 56154 129188
rect 58402 126824 58646 129188
rect 55916 126618 58646 126824
rect 69756 129186 72486 129406
rect 69756 126822 69994 129186
rect 72242 126822 72486 129186
rect 69756 126616 72486 126822
rect 83686 129188 86416 129408
rect 83686 126824 83924 129188
rect 86172 126824 86416 129188
rect 83686 126618 86416 126824
rect 97602 129190 100332 129410
rect 97602 126826 97840 129190
rect 100088 126826 100332 129190
rect 97602 126620 100332 126826
rect 111436 129198 114166 129418
rect 111436 126834 111674 129198
rect 113922 126834 114166 129198
rect 111436 126628 114166 126834
rect 125366 129200 128096 129420
rect 125366 126836 125604 129200
rect 127852 126836 128096 129200
rect 125366 126630 128096 126836
rect 139282 129202 142012 129422
rect 139282 126838 139520 129202
rect 141768 126838 142012 129202
rect 139282 126632 142012 126838
rect 153116 129198 155846 129418
rect 153116 126834 153354 129198
rect 155602 126834 155846 129198
rect 153116 126628 155846 126834
rect 167046 129200 169776 129420
rect 167046 126836 167284 129200
rect 169532 126836 169776 129200
rect 167046 126630 169776 126836
rect 180962 129202 183692 129422
rect 180962 126838 181200 129202
rect 183448 126838 183692 129202
rect 180962 126632 183692 126838
rect 194598 129160 197328 129380
rect 194598 126796 194836 129160
rect 197084 126796 197328 129160
rect 194598 126590 197328 126796
rect 208528 129162 211258 129382
rect 208528 126798 208766 129162
rect 211014 126798 211258 129162
rect 208528 126592 211258 126798
rect 222444 129164 225174 129384
rect 222444 126800 222682 129164
rect 224930 126800 225174 129164
rect 222444 126594 225174 126800
rect 236284 129162 239014 129382
rect 236284 126798 236522 129162
rect 238770 126798 239014 129162
rect 236284 126592 239014 126798
rect 250214 129164 252944 129384
rect 250214 126800 250452 129164
rect 252700 126800 252944 129164
rect 250214 126594 252944 126800
rect 264130 129166 266860 129386
rect 264130 126802 264368 129166
rect 266616 126802 266860 129166
rect 264130 126596 266860 126802
rect 277964 129174 280694 129394
rect 277964 126810 278202 129174
rect 280450 126810 280694 129174
rect 277964 126604 280694 126810
rect 291894 129176 294624 129396
rect 291894 126812 292132 129176
rect 294380 126812 294624 129176
rect 291894 126606 294624 126812
rect 305810 129178 308540 129398
rect 305810 126814 306048 129178
rect 308296 126814 308540 129178
rect 305810 126608 308540 126814
rect 319644 129174 322374 129394
rect 319644 126810 319882 129174
rect 322130 126810 322374 129174
rect 319644 126604 322374 126810
rect 333574 129176 336304 129396
rect 333574 126812 333812 129176
rect 336060 126812 336304 129176
rect 333574 126606 336304 126812
rect 347490 129178 350220 129398
rect 347490 126814 347728 129178
rect 349976 126814 350220 129178
rect 347490 126608 350220 126814
rect 41930 117752 44660 117972
rect 41930 115388 42168 117752
rect 44416 115388 44660 117752
rect 41930 115182 44660 115388
rect 55846 117754 58576 117974
rect 55846 115390 56084 117754
rect 58332 115390 58576 117754
rect 55846 115184 58576 115390
rect 69686 117752 72416 117972
rect 69686 115388 69924 117752
rect 72172 115388 72416 117752
rect 69686 115182 72416 115388
rect 83616 117754 86346 117974
rect 83616 115390 83854 117754
rect 86102 115390 86346 117754
rect 83616 115184 86346 115390
rect 97532 117756 100262 117976
rect 97532 115392 97770 117756
rect 100018 115392 100262 117756
rect 97532 115186 100262 115392
rect 111366 117764 114096 117984
rect 111366 115400 111604 117764
rect 113852 115400 114096 117764
rect 111366 115194 114096 115400
rect 125296 117766 128026 117986
rect 125296 115402 125534 117766
rect 127782 115402 128026 117766
rect 125296 115196 128026 115402
rect 139212 117768 141942 117988
rect 139212 115404 139450 117768
rect 141698 115404 141942 117768
rect 139212 115198 141942 115404
rect 153046 117764 155776 117984
rect 153046 115400 153284 117764
rect 155532 115400 155776 117764
rect 153046 115194 155776 115400
rect 166976 117766 169706 117986
rect 166976 115402 167214 117766
rect 169462 115402 169706 117766
rect 166976 115196 169706 115402
rect 180892 117768 183622 117988
rect 180892 115404 181130 117768
rect 183378 115404 183622 117768
rect 180892 115198 183622 115404
rect 194528 117726 197258 117946
rect 194528 115362 194766 117726
rect 197014 115362 197258 117726
rect 194528 115156 197258 115362
rect 208458 117728 211188 117948
rect 208458 115364 208696 117728
rect 210944 115364 211188 117728
rect 208458 115158 211188 115364
rect 222374 117730 225104 117950
rect 222374 115366 222612 117730
rect 224860 115366 225104 117730
rect 222374 115160 225104 115366
rect 236214 117728 238944 117948
rect 236214 115364 236452 117728
rect 238700 115364 238944 117728
rect 236214 115158 238944 115364
rect 250144 117730 252874 117950
rect 250144 115366 250382 117730
rect 252630 115366 252874 117730
rect 250144 115160 252874 115366
rect 264060 117732 266790 117952
rect 264060 115368 264298 117732
rect 266546 115368 266790 117732
rect 264060 115162 266790 115368
rect 277894 117740 280624 117960
rect 277894 115376 278132 117740
rect 280380 115376 280624 117740
rect 277894 115170 280624 115376
rect 291824 117742 294554 117962
rect 291824 115378 292062 117742
rect 294310 115378 294554 117742
rect 291824 115172 294554 115378
rect 305740 117744 308470 117964
rect 305740 115380 305978 117744
rect 308226 115380 308470 117744
rect 305740 115174 308470 115380
rect 319574 117740 322304 117960
rect 319574 115376 319812 117740
rect 322060 115376 322304 117740
rect 319574 115170 322304 115376
rect 333504 117742 336234 117962
rect 333504 115378 333742 117742
rect 335990 115378 336234 117742
rect 333504 115172 336234 115378
rect 347420 117744 350150 117964
rect 347420 115380 347658 117744
rect 349906 115380 350150 117744
rect 347420 115174 350150 115380
rect 41792 105342 44522 105562
rect 41792 102978 42030 105342
rect 44278 102978 44522 105342
rect 41792 102772 44522 102978
rect 55708 105344 58438 105564
rect 55708 102980 55946 105344
rect 58194 102980 58438 105344
rect 55708 102774 58438 102980
rect 69548 105342 72278 105562
rect 69548 102978 69786 105342
rect 72034 102978 72278 105342
rect 69548 102772 72278 102978
rect 83478 105344 86208 105564
rect 83478 102980 83716 105344
rect 85964 102980 86208 105344
rect 83478 102774 86208 102980
rect 97394 105346 100124 105566
rect 97394 102982 97632 105346
rect 99880 102982 100124 105346
rect 97394 102776 100124 102982
rect 111228 105354 113958 105574
rect 111228 102990 111466 105354
rect 113714 102990 113958 105354
rect 111228 102784 113958 102990
rect 125158 105356 127888 105576
rect 125158 102992 125396 105356
rect 127644 102992 127888 105356
rect 125158 102786 127888 102992
rect 139074 105358 141804 105578
rect 139074 102994 139312 105358
rect 141560 102994 141804 105358
rect 139074 102788 141804 102994
rect 152908 105354 155638 105574
rect 152908 102990 153146 105354
rect 155394 102990 155638 105354
rect 152908 102784 155638 102990
rect 166838 105356 169568 105576
rect 166838 102992 167076 105356
rect 169324 102992 169568 105356
rect 166838 102786 169568 102992
rect 180754 105358 183484 105578
rect 180754 102994 180992 105358
rect 183240 102994 183484 105358
rect 180754 102788 183484 102994
rect 194390 105316 197120 105536
rect 194390 102952 194628 105316
rect 196876 102952 197120 105316
rect 194390 102746 197120 102952
rect 208320 105318 211050 105538
rect 208320 102954 208558 105318
rect 210806 102954 211050 105318
rect 208320 102748 211050 102954
rect 222236 105320 224966 105540
rect 222236 102956 222474 105320
rect 224722 102956 224966 105320
rect 222236 102750 224966 102956
rect 236076 105318 238806 105538
rect 236076 102954 236314 105318
rect 238562 102954 238806 105318
rect 236076 102748 238806 102954
rect 250006 105320 252736 105540
rect 250006 102956 250244 105320
rect 252492 102956 252736 105320
rect 250006 102750 252736 102956
rect 263922 105322 266652 105542
rect 263922 102958 264160 105322
rect 266408 102958 266652 105322
rect 263922 102752 266652 102958
rect 277756 105330 280486 105550
rect 277756 102966 277994 105330
rect 280242 102966 280486 105330
rect 277756 102760 280486 102966
rect 291686 105332 294416 105552
rect 291686 102968 291924 105332
rect 294172 102968 294416 105332
rect 291686 102762 294416 102968
rect 305602 105334 308332 105554
rect 305602 102970 305840 105334
rect 308088 102970 308332 105334
rect 305602 102764 308332 102970
rect 319436 105330 322166 105550
rect 319436 102966 319674 105330
rect 321922 102966 322166 105330
rect 319436 102760 322166 102966
rect 333366 105332 336096 105552
rect 333366 102968 333604 105332
rect 335852 102968 336096 105332
rect 333366 102762 336096 102968
rect 347282 105334 350012 105554
rect 347282 102970 347520 105334
rect 349768 102970 350012 105334
rect 347282 102764 350012 102970
rect 277180 89614 279910 89834
rect 277180 87250 277418 89614
rect 279666 87250 279910 89614
rect 277180 87044 279910 87250
rect 291110 89616 293840 89836
rect 291110 87252 291348 89616
rect 293596 87252 293840 89616
rect 291110 87046 293840 87252
rect 305026 89618 307756 89838
rect 305026 87254 305264 89618
rect 307512 87254 307756 89618
rect 305026 87048 307756 87254
rect 318860 89614 321590 89834
rect 318860 87250 319098 89614
rect 321346 87250 321590 89614
rect 318860 87044 321590 87250
rect 332790 89616 335520 89836
rect 332790 87252 333028 89616
rect 335276 87252 335520 89616
rect 332790 87046 335520 87252
rect 346706 89618 349436 89838
rect 346706 87254 346944 89618
rect 349192 87254 349436 89618
rect 346706 87048 349436 87254
rect 277180 77026 279910 77246
rect 277180 74662 277418 77026
rect 279666 74662 279910 77026
rect 277180 74456 279910 74662
rect 291110 77028 293840 77248
rect 291110 74664 291348 77028
rect 293596 74664 293840 77028
rect 291110 74458 293840 74664
rect 305026 77030 307756 77250
rect 305026 74666 305264 77030
rect 307512 74666 307756 77030
rect 305026 74460 307756 74666
rect 318860 77026 321590 77246
rect 318860 74662 319098 77026
rect 321346 74662 321590 77026
rect 318860 74456 321590 74662
rect 332790 77028 335520 77248
rect 332790 74664 333028 77028
rect 335276 74664 335520 77028
rect 332790 74458 335520 74664
rect 346706 77030 349436 77250
rect 346706 74666 346944 77030
rect 349192 74666 349436 77030
rect 346706 74460 349436 74666
rect 277180 64438 279910 64658
rect 277180 62074 277418 64438
rect 279666 62074 279910 64438
rect 277180 61868 279910 62074
rect 291110 64440 293840 64660
rect 291110 62076 291348 64440
rect 293596 62076 293840 64440
rect 291110 61870 293840 62076
rect 305026 64442 307756 64662
rect 305026 62078 305264 64442
rect 307512 62078 307756 64442
rect 305026 61872 307756 62078
rect 318860 64438 321590 64658
rect 318860 62074 319098 64438
rect 321346 62074 321590 64438
rect 318860 61868 321590 62074
rect 332790 64440 335520 64660
rect 332790 62076 333028 64440
rect 335276 62076 335520 64440
rect 332790 61870 335520 62076
rect 346706 64442 349436 64662
rect 346706 62078 346944 64442
rect 349192 62078 349436 64442
rect 346706 61872 349436 62078
<< psubdiffcont >>
rect 167022 677730 169270 680094
rect 180938 677732 183186 680096
rect 194574 677690 196822 680054
rect 208504 677692 210752 680056
rect 222420 677694 224668 680058
rect 236260 677692 238508 680056
rect 250190 677694 252438 680058
rect 264106 677696 266354 680060
rect 277940 677704 280188 680068
rect 291870 677706 294118 680070
rect 305786 677708 308034 680072
rect 319620 677704 321868 680068
rect 333550 677706 335798 680070
rect 347466 677708 349714 680072
rect 361076 677694 363324 680058
rect 375006 677696 377254 680060
rect 388922 677698 391170 680062
rect 402762 677696 405010 680060
rect 416692 677698 418940 680062
rect 430608 677700 432856 680064
rect 194026 663430 196274 665794
rect 207956 663432 210204 665796
rect 277392 663444 279640 665808
rect 291322 663446 293570 665810
rect 305238 663448 307486 665812
rect 319072 663444 321320 665808
rect 333002 663446 335250 665810
rect 346918 663448 349166 665812
rect 360528 663434 362776 665798
rect 374458 663436 376706 665800
rect 388374 663438 390622 665802
rect 402214 663436 404462 665800
rect 416144 663438 418392 665802
rect 430060 663440 432308 665804
rect 194574 650774 196822 653138
rect 208504 650776 210752 653140
rect 277940 650788 280188 653152
rect 291870 650790 294118 653154
rect 305786 650792 308034 653156
rect 319620 650788 321868 653152
rect 333550 650790 335798 653154
rect 347466 650792 349714 653156
rect 361076 650778 363324 653142
rect 375006 650780 377254 653144
rect 388922 650782 391170 653146
rect 402762 650780 405010 653144
rect 416692 650782 418940 653146
rect 430608 650784 432856 653148
rect 194026 636514 196274 638878
rect 207956 636516 210204 638880
rect 277392 636528 279640 638892
rect 291322 636530 293570 638894
rect 305238 636532 307486 638896
rect 319072 636528 321320 638892
rect 333002 636530 335250 638894
rect 346918 636532 349166 638896
rect 360528 636518 362776 638882
rect 374458 636520 376706 638884
rect 388374 636522 390622 638886
rect 402214 636520 404462 638884
rect 416144 636522 418392 638886
rect 430060 636524 432308 638888
rect 194586 622252 196834 624616
rect 208516 622254 210764 624618
rect 277952 622266 280200 624630
rect 291882 622268 294130 624632
rect 305798 622270 308046 624634
rect 319632 622266 321880 624630
rect 333562 622268 335810 624632
rect 347478 622270 349726 624634
rect 361088 622256 363336 624620
rect 375018 622258 377266 624622
rect 388934 622260 391182 624624
rect 402774 622258 405022 624622
rect 416704 622260 418952 624624
rect 430620 622262 432868 624626
rect 166486 608032 168734 610396
rect 180402 608034 182650 610398
rect 194038 607992 196286 610356
rect 207968 607994 210216 610358
rect 221884 607996 224132 610360
rect 235724 607994 237972 610358
rect 249654 607996 251902 610360
rect 263570 607998 265818 610362
rect 277404 608006 279652 610370
rect 291334 608008 293582 610372
rect 305250 608010 307498 610374
rect 319084 608006 321332 610370
rect 333014 608008 335262 610372
rect 346930 608010 349178 610374
rect 360540 607996 362788 610360
rect 374470 607998 376718 610362
rect 388386 608000 390634 610364
rect 402226 607998 404474 610362
rect 416156 608000 418404 610364
rect 430072 608002 432320 610366
rect 194764 589534 197012 591898
rect 208694 589536 210942 591900
rect 278130 589548 280378 591912
rect 292060 589550 294308 591914
rect 305976 589552 308224 591916
rect 319810 589548 322058 591912
rect 333740 589550 335988 591914
rect 375196 589540 377444 591904
rect 389112 589542 391360 591906
rect 194216 575274 196464 577638
rect 208146 575276 210394 577640
rect 277582 575288 279830 577652
rect 291512 575290 293760 577654
rect 305428 575292 307676 577656
rect 319262 575288 321510 577652
rect 333192 575290 335440 577654
rect 374648 575280 376896 577644
rect 388564 575282 390812 577646
rect 194432 562448 196680 564812
rect 208362 562450 210610 564814
rect 277798 562462 280046 564826
rect 291728 562464 293976 564828
rect 305644 562466 307892 564830
rect 319478 562462 321726 564826
rect 333408 562464 335656 564828
rect 374864 562454 377112 564818
rect 388780 562456 391028 564820
rect 139550 544760 141798 547124
rect 153384 544756 155632 547120
rect 167314 544758 169562 547122
rect 181230 544760 183478 547124
rect 194866 544718 197114 547082
rect 208796 544720 211044 547084
rect 222712 544722 224960 547086
rect 236552 544720 238800 547084
rect 250482 544722 252730 547086
rect 264398 544724 266646 547088
rect 278232 544732 280480 547096
rect 292162 544734 294410 547098
rect 306078 544736 308326 547100
rect 319912 544732 322160 547096
rect 333842 544734 336090 547098
rect 347758 544736 350006 547100
rect 361368 544722 363616 547086
rect 375298 544724 377546 547088
rect 389214 544726 391462 547090
rect 403054 544724 405302 547088
rect 416984 544726 419232 547090
rect 430900 544728 433148 547092
rect 444734 544736 446982 547100
rect 139002 530500 141250 532864
rect 152836 530496 155084 532860
rect 166766 530498 169014 532862
rect 180682 530500 182930 532864
rect 194318 530458 196566 532822
rect 208248 530460 210496 532824
rect 222164 530462 224412 532826
rect 236004 530460 238252 532824
rect 249934 530462 252182 532826
rect 263850 530464 266098 532828
rect 277684 530472 279932 532836
rect 291614 530474 293862 532838
rect 305530 530476 307778 532840
rect 319364 530472 321612 532836
rect 333294 530474 335542 532838
rect 347210 530476 349458 532840
rect 360820 530462 363068 532826
rect 374750 530464 376998 532828
rect 388666 530466 390914 532830
rect 402506 530464 404754 532828
rect 416436 530466 418684 532830
rect 430352 530468 432600 532832
rect 444186 530476 446434 532840
rect 139218 517674 141466 520038
rect 153052 517670 155300 520034
rect 166982 517672 169230 520036
rect 180898 517674 183146 520038
rect 194534 517632 196782 519996
rect 208464 517634 210712 519998
rect 222380 517636 224628 520000
rect 236220 517634 238468 519998
rect 250150 517636 252398 520000
rect 264066 517638 266314 520002
rect 277900 517646 280148 520010
rect 291830 517648 294078 520012
rect 305746 517650 307994 520014
rect 319580 517646 321828 520010
rect 333510 517648 335758 520012
rect 347426 517650 349674 520014
rect 361036 517636 363284 520000
rect 374966 517638 377214 520002
rect 388882 517640 391130 520004
rect 402722 517638 404970 520002
rect 416652 517640 418900 520004
rect 430568 517642 432816 520006
rect 444402 517650 446650 520014
rect 167376 496250 169624 498614
rect 181292 496252 183540 498616
rect 194928 496210 197176 498574
rect 208858 496212 211106 498576
rect 222774 496214 225022 498578
rect 236614 496212 238862 498576
rect 250544 496214 252792 498578
rect 264460 496216 266708 498580
rect 278294 496224 280542 498588
rect 292224 496226 294472 498590
rect 306140 496228 308388 498592
rect 319974 496224 322222 498588
rect 333904 496226 336152 498590
rect 347820 496228 350068 498592
rect 361430 496214 363678 498578
rect 375360 496216 377608 498580
rect 389276 496218 391524 498582
rect 403116 496216 405364 498580
rect 417046 496218 419294 498582
rect 430962 496220 433210 498584
rect 444796 496228 447044 498592
rect 166828 481990 169076 484354
rect 180744 481992 182992 484356
rect 194380 481950 196628 484314
rect 208310 481952 210558 484316
rect 222226 481954 224474 484318
rect 236066 481952 238314 484316
rect 249996 481954 252244 484318
rect 263912 481956 266160 484320
rect 277746 481964 279994 484328
rect 291676 481966 293924 484330
rect 305592 481968 307840 484332
rect 319426 481964 321674 484328
rect 333356 481966 335604 484330
rect 347272 481968 349520 484332
rect 360882 481954 363130 484318
rect 374812 481956 377060 484320
rect 388728 481958 390976 484322
rect 402568 481956 404816 484320
rect 416498 481958 418746 484322
rect 430414 481960 432662 484324
rect 444248 481968 446496 484332
rect 167044 469164 169292 471528
rect 180960 469166 183208 471530
rect 194596 469124 196844 471488
rect 208526 469126 210774 471490
rect 222442 469128 224690 471492
rect 236282 469126 238530 471490
rect 250212 469128 252460 471492
rect 264128 469130 266376 471494
rect 277962 469138 280210 471502
rect 291892 469140 294140 471504
rect 305808 469142 308056 471506
rect 319642 469138 321890 471502
rect 333572 469140 335820 471504
rect 347488 469142 349736 471506
rect 361098 469128 363346 471492
rect 375028 469130 377276 471494
rect 388944 469132 391192 471496
rect 402784 469130 405032 471494
rect 416714 469132 418962 471496
rect 430630 469134 432878 471498
rect 444464 469142 446712 471506
rect 139860 455720 142108 458084
rect 153694 455716 155942 458080
rect 167624 455718 169872 458082
rect 181540 455720 183788 458084
rect 195176 455678 197424 458042
rect 209106 455680 211354 458044
rect 223022 455682 225270 458046
rect 236862 455680 239110 458044
rect 250792 455682 253040 458046
rect 264708 455684 266956 458048
rect 278542 455692 280790 458056
rect 292472 455694 294720 458058
rect 306388 455696 308636 458060
rect 320222 455692 322470 458056
rect 334152 455694 336400 458058
rect 348068 455696 350316 458060
rect 361678 455682 363926 458046
rect 375608 455684 377856 458048
rect 389524 455686 391772 458050
rect 403364 455684 405612 458048
rect 417294 455686 419542 458050
rect 431210 455688 433458 458052
rect 445044 455696 447292 458060
rect 139820 443996 142068 446360
rect 153654 443992 155902 446356
rect 167584 443994 169832 446358
rect 181500 443996 183748 446360
rect 195136 443954 197384 446318
rect 209066 443956 211314 446320
rect 222982 443958 225230 446322
rect 236822 443956 239070 446320
rect 250752 443958 253000 446322
rect 264668 443960 266916 446324
rect 278502 443968 280750 446332
rect 292432 443970 294680 446334
rect 306348 443972 308596 446336
rect 320182 443968 322430 446332
rect 334112 443970 336360 446334
rect 348028 443972 350276 446336
rect 361638 443958 363886 446322
rect 375568 443960 377816 446324
rect 389484 443962 391732 446326
rect 403324 443960 405572 446324
rect 417254 443962 419502 446326
rect 431170 443964 433418 446328
rect 445004 443972 447252 446336
rect 42618 419854 44866 422218
rect 56534 419856 58782 422220
rect 70374 419854 72622 422218
rect 84304 419856 86552 422220
rect 98220 419858 100468 422222
rect 112054 419866 114302 422230
rect 125984 419868 128232 422232
rect 195216 419828 197464 422192
rect 209146 419830 211394 422194
rect 278582 419842 280830 422206
rect 292512 419844 294760 422208
rect 306428 419846 308676 422210
rect 320262 419842 322510 422206
rect 334192 419844 336440 422208
rect 528890 419850 531138 422214
rect 542806 419852 545054 422216
rect 42070 405594 44318 407958
rect 55986 405596 58234 407960
rect 69826 405594 72074 407958
rect 83756 405596 86004 407960
rect 97672 405598 99920 407962
rect 111506 405606 113754 407970
rect 125436 405608 127684 407972
rect 194668 405568 196916 407932
rect 208598 405570 210846 407934
rect 278034 405582 280282 407946
rect 291964 405584 294212 407948
rect 305880 405586 308128 407950
rect 319714 405582 321962 407946
rect 333644 405584 335892 407948
rect 528342 405590 530590 407954
rect 542258 405592 544506 407956
rect 42286 392768 44534 395132
rect 56202 392770 58450 395134
rect 70042 392768 72290 395132
rect 83972 392770 86220 395134
rect 97888 392772 100136 395136
rect 111722 392780 113970 395144
rect 125652 392782 127900 395146
rect 194884 392742 197132 395106
rect 208814 392744 211062 395108
rect 278250 392756 280498 395120
rect 292180 392758 294428 395122
rect 306096 392760 308344 395124
rect 319930 392756 322178 395120
rect 333860 392758 336108 395122
rect 528558 392764 530806 395128
rect 542474 392766 544722 395130
rect 195190 384042 197438 386406
rect 209120 384044 211368 386408
rect 278556 384056 280804 386420
rect 292486 384058 294734 386422
rect 306402 384060 308650 386424
rect 320236 384056 322484 386420
rect 334166 384058 336414 386422
rect 528864 384064 531112 386428
rect 542780 384066 545028 386430
rect 153160 369820 155408 372184
rect 167090 369822 169338 372186
rect 181006 369824 183254 372188
rect 194642 369782 196890 372146
rect 208572 369784 210820 372148
rect 278008 369796 280256 372160
rect 291938 369798 294186 372162
rect 305854 369800 308102 372164
rect 319688 369796 321936 372160
rect 333618 369798 335866 372162
rect 347534 369800 349782 372164
rect 361144 369786 363392 372150
rect 375074 369788 377322 372152
rect 388990 369790 391238 372154
rect 402830 369788 405078 372152
rect 416760 369790 419008 372154
rect 430676 369792 432924 372156
rect 444510 369800 446758 372164
rect 458440 369802 460688 372166
rect 472356 369804 474604 372168
rect 486190 369800 488438 372164
rect 500120 369802 502368 372166
rect 514036 369804 516284 372168
rect 528316 369804 530564 372168
rect 542232 369806 544480 372170
rect 556504 369786 558752 372150
rect 153376 356994 155624 359358
rect 167306 356996 169554 359360
rect 181222 356998 183470 359362
rect 194858 356956 197106 359320
rect 208788 356958 211036 359322
rect 222704 356960 224952 359324
rect 236544 356958 238792 359322
rect 250474 356960 252722 359324
rect 264390 356962 266638 359326
rect 278224 356970 280472 359334
rect 292154 356972 294402 359336
rect 306070 356974 308318 359338
rect 319904 356970 322152 359334
rect 333834 356972 336082 359336
rect 347750 356974 349998 359338
rect 361360 356960 363608 359324
rect 375290 356962 377538 359326
rect 389206 356964 391454 359328
rect 403046 356962 405294 359326
rect 416976 356964 419224 359328
rect 430892 356966 433140 359330
rect 444726 356974 446974 359338
rect 458656 356976 460904 359340
rect 472572 356978 474820 359342
rect 486406 356974 488654 359338
rect 500336 356976 502584 359340
rect 514252 356978 516500 359342
rect 528532 356978 530780 359342
rect 542448 356980 544696 359344
rect 556720 356960 558968 359324
rect 138972 345170 141220 347534
rect 152806 345166 155054 347530
rect 166736 345168 168984 347532
rect 180652 345170 182900 347534
rect 194288 345128 196536 347492
rect 208218 345130 210466 347494
rect 222134 345132 224382 347496
rect 235974 345130 238222 347494
rect 249904 345132 252152 347496
rect 263820 345134 266068 347498
rect 277654 345142 279902 347506
rect 291584 345144 293832 347508
rect 305500 345146 307748 347510
rect 319334 345142 321582 347506
rect 333264 345144 335512 347508
rect 347180 345146 349428 347510
rect 360790 345132 363038 347496
rect 374720 345134 376968 347498
rect 388636 345136 390884 347500
rect 402476 345134 404724 347498
rect 416406 345136 418654 347500
rect 430322 345138 432570 347502
rect 444156 345146 446404 347510
rect 458086 345148 460334 347512
rect 472002 345150 474250 347514
rect 485836 345146 488084 347510
rect 499766 345148 502014 347512
rect 513682 345150 515930 347514
rect 527962 345150 530210 347514
rect 541878 345152 544126 347516
rect 556150 345132 558398 347496
rect 139188 332344 141436 334708
rect 153022 332340 155270 334704
rect 166952 332342 169200 334706
rect 180868 332344 183116 334708
rect 194504 332302 196752 334666
rect 208434 332304 210682 334668
rect 222350 332306 224598 334670
rect 236190 332304 238438 334668
rect 250120 332306 252368 334670
rect 264036 332308 266284 334672
rect 277870 332316 280118 334680
rect 291800 332318 294048 334682
rect 305716 332320 307964 334684
rect 319550 332316 321798 334680
rect 333480 332318 335728 334682
rect 347396 332320 349644 334684
rect 361006 332306 363254 334670
rect 374936 332308 377184 334672
rect 388852 332310 391100 334674
rect 402692 332308 404940 334672
rect 416622 332310 418870 334674
rect 430538 332312 432786 334676
rect 444372 332320 446620 334684
rect 458302 332322 460550 334686
rect 472218 332324 474466 334688
rect 486052 332320 488300 334684
rect 499982 332322 502230 334686
rect 513898 332324 516146 334688
rect 528178 332324 530426 334688
rect 542094 332326 544342 334690
rect 556366 332306 558614 334670
rect 43440 317650 45688 320014
rect 57356 317652 59604 320016
rect 71196 317650 73444 320014
rect 112876 317662 115124 320026
rect 126806 317664 129054 320028
rect 196038 317624 198286 319988
rect 209968 317626 212216 319990
rect 279404 317638 281652 320002
rect 293334 317640 295582 320004
rect 307250 317642 309498 320006
rect 321084 317638 323332 320002
rect 335014 317640 337262 320004
rect 376470 317630 378718 319994
rect 390386 317632 392634 319996
rect 459584 317632 461832 319996
rect 473514 317634 475762 319998
rect 487430 317636 489678 320000
rect 501264 317644 503512 320008
rect 515048 317610 517296 319974
rect 528978 317612 531226 319976
rect 542894 317614 545142 319978
rect 556728 317622 558976 319986
rect 44010 307984 46258 310348
rect 57926 307986 60174 310350
rect 71766 307984 74014 310348
rect 113446 307996 115694 310360
rect 127376 307998 129624 310362
rect 196608 307958 198856 310322
rect 210538 307960 212786 310324
rect 279974 307972 282222 310336
rect 293904 307974 296152 310338
rect 307820 307976 310068 310340
rect 321654 307972 323902 310336
rect 335584 307974 337832 310338
rect 377040 307964 379288 310328
rect 390956 307966 393204 310330
rect 460154 307966 462402 310330
rect 474084 307968 476332 310332
rect 488000 307970 490248 310334
rect 501834 307978 504082 310342
rect 515618 307944 517866 310308
rect 529548 307946 531796 310310
rect 543464 307948 545712 310312
rect 557298 307956 559546 310320
rect 44152 297464 46400 299828
rect 58068 297466 60316 299830
rect 71908 297464 74156 299828
rect 113588 297476 115836 299840
rect 127518 297478 129766 299842
rect 196750 297438 198998 299802
rect 210680 297440 212928 299804
rect 280116 297452 282364 299816
rect 294046 297454 296294 299818
rect 307962 297456 310210 299820
rect 321796 297452 324044 299816
rect 335726 297454 337974 299818
rect 377182 297444 379430 299808
rect 391098 297446 393346 299810
rect 460296 297446 462544 299810
rect 474226 297448 476474 299812
rect 488142 297450 490390 299814
rect 501976 297458 504224 299822
rect 515760 297424 518008 299788
rect 529690 297426 531938 299790
rect 543606 297428 545854 299792
rect 557440 297436 559688 299800
rect 44010 286516 46258 288880
rect 57926 286518 60174 288882
rect 71766 286516 74014 288880
rect 113446 286528 115694 288892
rect 127376 286530 129624 288894
rect 196608 286490 198856 288854
rect 210538 286492 212786 288856
rect 279974 286504 282222 288868
rect 293904 286506 296152 288870
rect 307820 286508 310068 288872
rect 321654 286504 323902 288868
rect 335584 286506 337832 288870
rect 377040 286496 379288 288860
rect 390956 286498 393204 288862
rect 44294 274292 46542 276656
rect 58210 274294 60458 276658
rect 72050 274292 74298 276656
rect 113730 274304 115978 276668
rect 127660 274306 129908 276670
rect 196892 274266 199140 276630
rect 210822 274268 213070 276632
rect 280258 274280 282506 276644
rect 294188 274282 296436 276646
rect 308104 274284 310352 276648
rect 321938 274280 324186 276644
rect 335868 274282 338116 276646
rect 377324 274272 379572 276636
rect 391240 274274 393488 276638
rect 43874 258544 46122 260908
rect 57790 258546 60038 260910
rect 71630 258544 73878 260908
rect 85560 258546 87808 260910
rect 99476 258548 101724 260912
rect 113310 258556 115558 260920
rect 127240 258558 129488 260922
rect 141156 258560 143404 260924
rect 154990 258556 157238 260920
rect 168920 258558 171168 260922
rect 182836 258560 185084 260924
rect 196472 258518 198720 260882
rect 210402 258520 212650 260884
rect 224318 258522 226566 260886
rect 238158 258520 240406 260884
rect 252088 258522 254336 260886
rect 266004 258524 268252 260888
rect 279838 258532 282086 260896
rect 293768 258534 296016 260898
rect 307684 258536 309932 260900
rect 321518 258532 323766 260896
rect 335448 258534 337696 260898
rect 349364 258536 351612 260900
rect 362974 258522 365222 260886
rect 376904 258524 379152 260888
rect 390820 258526 393068 260890
rect 195506 235886 197754 238250
rect 209436 235888 211684 238252
rect 278872 235900 281120 238264
rect 292802 235902 295050 238266
rect 306718 235904 308966 238268
rect 320552 235900 322800 238264
rect 334482 235902 336730 238266
rect 195916 219982 198164 222346
rect 209846 219984 212094 222348
rect 279282 219996 281530 222360
rect 293212 219998 295460 222362
rect 307128 220000 309376 222364
rect 320962 219996 323210 222360
rect 334892 219998 337140 222362
rect 195916 203530 198164 205894
rect 209846 203532 212094 205896
rect 279282 203544 281530 205908
rect 293212 203546 295460 205910
rect 307128 203548 309376 205912
rect 320962 203544 323210 205908
rect 334892 203546 337140 205910
rect 195506 188722 197754 191086
rect 209436 188724 211684 191088
rect 278872 188736 281120 191100
rect 292802 188738 295050 191102
rect 306718 188740 308966 191104
rect 320552 188736 322800 191100
rect 334482 188738 336730 191102
rect 194958 174462 197206 176826
rect 208888 174464 211136 176828
rect 222804 174466 225052 176830
rect 236644 174464 238892 176828
rect 250574 174466 252822 176830
rect 264490 174468 266738 176832
rect 278324 174476 280572 176840
rect 292254 174478 294502 176842
rect 306170 174480 308418 176844
rect 320004 174476 322252 176840
rect 333934 174478 336182 176842
rect 195174 161636 197422 164000
rect 209104 161638 211352 164002
rect 223020 161640 225268 164004
rect 236860 161638 239108 164002
rect 250790 161640 253038 164004
rect 264706 161642 266954 164006
rect 278540 161650 280788 164014
rect 292470 161652 294718 164016
rect 306386 161654 308634 164018
rect 320220 161650 322468 164014
rect 334150 161652 336398 164016
rect 42308 139302 44556 141666
rect 56224 139304 58472 141668
rect 70064 139302 72312 141666
rect 83994 139304 86242 141668
rect 97910 139306 100158 141670
rect 111744 139314 113992 141678
rect 125674 139316 127922 141680
rect 139590 139318 141838 141682
rect 153424 139314 155672 141678
rect 167354 139316 169602 141680
rect 181270 139318 183518 141682
rect 194906 139276 197154 141640
rect 208836 139278 211084 141642
rect 222752 139280 225000 141644
rect 236592 139278 238840 141642
rect 250522 139280 252770 141644
rect 264438 139282 266686 141646
rect 278272 139290 280520 141654
rect 292202 139292 294450 141656
rect 306118 139294 308366 141658
rect 319952 139290 322200 141654
rect 333882 139292 336130 141656
rect 347798 139294 350046 141658
rect 42238 126822 44486 129186
rect 56154 126824 58402 129188
rect 69994 126822 72242 129186
rect 83924 126824 86172 129188
rect 97840 126826 100088 129190
rect 111674 126834 113922 129198
rect 125604 126836 127852 129200
rect 139520 126838 141768 129202
rect 153354 126834 155602 129198
rect 167284 126836 169532 129200
rect 181200 126838 183448 129202
rect 194836 126796 197084 129160
rect 208766 126798 211014 129162
rect 222682 126800 224930 129164
rect 236522 126798 238770 129162
rect 250452 126800 252700 129164
rect 264368 126802 266616 129166
rect 278202 126810 280450 129174
rect 292132 126812 294380 129176
rect 306048 126814 308296 129178
rect 319882 126810 322130 129174
rect 333812 126812 336060 129176
rect 347728 126814 349976 129178
rect 42168 115388 44416 117752
rect 56084 115390 58332 117754
rect 69924 115388 72172 117752
rect 83854 115390 86102 117754
rect 97770 115392 100018 117756
rect 111604 115400 113852 117764
rect 125534 115402 127782 117766
rect 139450 115404 141698 117768
rect 153284 115400 155532 117764
rect 167214 115402 169462 117766
rect 181130 115404 183378 117768
rect 194766 115362 197014 117726
rect 208696 115364 210944 117728
rect 222612 115366 224860 117730
rect 236452 115364 238700 117728
rect 250382 115366 252630 117730
rect 264298 115368 266546 117732
rect 278132 115376 280380 117740
rect 292062 115378 294310 117742
rect 305978 115380 308226 117744
rect 319812 115376 322060 117740
rect 333742 115378 335990 117742
rect 347658 115380 349906 117744
rect 42030 102978 44278 105342
rect 55946 102980 58194 105344
rect 69786 102978 72034 105342
rect 83716 102980 85964 105344
rect 97632 102982 99880 105346
rect 111466 102990 113714 105354
rect 125396 102992 127644 105356
rect 139312 102994 141560 105358
rect 153146 102990 155394 105354
rect 167076 102992 169324 105356
rect 180992 102994 183240 105358
rect 194628 102952 196876 105316
rect 208558 102954 210806 105318
rect 222474 102956 224722 105320
rect 236314 102954 238562 105318
rect 250244 102956 252492 105320
rect 264160 102958 266408 105322
rect 277994 102966 280242 105330
rect 291924 102968 294172 105332
rect 305840 102970 308088 105334
rect 319674 102966 321922 105330
rect 333604 102968 335852 105332
rect 347520 102970 349768 105334
rect 277418 87250 279666 89614
rect 291348 87252 293596 89616
rect 305264 87254 307512 89618
rect 319098 87250 321346 89614
rect 333028 87252 335276 89616
rect 346944 87254 349192 89618
rect 277418 74662 279666 77026
rect 291348 74664 293596 77028
rect 305264 74666 307512 77030
rect 319098 74662 321346 77026
rect 333028 74664 335276 77028
rect 346944 74666 349192 77030
rect 277418 62074 279666 64438
rect 291348 62076 293596 64440
rect 305264 62078 307512 64442
rect 319098 62074 321346 64438
rect 333028 62076 335276 64440
rect 346944 62078 349192 64442
<< locali >>
rect 159392 680984 200972 681060
rect 205506 681034 282128 681060
rect 287026 681034 379306 681060
rect 205506 680990 379306 681034
rect 384006 680990 440060 681060
rect 205506 680984 440060 680990
rect 159392 680096 440060 680984
rect 159392 680094 180938 680096
rect 159392 677730 167022 680094
rect 169270 677732 180938 680094
rect 183186 680072 440060 680096
rect 183186 680070 305786 680072
rect 183186 680068 291870 680070
rect 183186 680060 277940 680068
rect 183186 680058 264106 680060
rect 183186 680056 222420 680058
rect 183186 680054 208504 680056
rect 183186 677732 194574 680054
rect 169270 677730 194574 677732
rect 159392 677690 194574 677730
rect 196822 677692 208504 680054
rect 210752 677694 222420 680056
rect 224668 680056 250190 680058
rect 224668 677694 236260 680056
rect 210752 677692 236260 677694
rect 238508 677694 250190 680056
rect 252438 677696 264106 680058
rect 266354 677704 277940 680060
rect 280188 677706 291870 680068
rect 294118 677708 305786 680070
rect 308034 680070 347466 680072
rect 308034 680068 333550 680070
rect 308034 677708 319620 680068
rect 294118 677706 319620 677708
rect 280188 677704 319620 677706
rect 321868 679898 333550 680068
rect 321868 677704 329000 679898
rect 266354 677696 329000 677704
rect 252438 677694 329000 677696
rect 238508 677692 329000 677694
rect 196822 677690 329000 677692
rect 159392 677548 329000 677690
rect 331532 677706 333550 679898
rect 335798 677708 347466 680070
rect 349714 680064 440060 680072
rect 349714 680062 430608 680064
rect 349714 680060 388922 680062
rect 349714 680058 375006 680060
rect 349714 677708 361076 680058
rect 335798 677706 361076 677708
rect 331532 677694 361076 677706
rect 363324 677696 375006 680058
rect 377254 677698 388922 680060
rect 391170 680060 416692 680062
rect 391170 677698 402762 680060
rect 377254 677696 402762 677698
rect 405010 677698 416692 680060
rect 418940 677700 430608 680062
rect 432856 677700 440060 680064
rect 418940 677698 440060 677700
rect 405010 677696 440060 677698
rect 363324 677694 440060 677696
rect 331532 677548 440060 677694
rect 159392 676846 440060 677548
rect 201278 666800 205076 676846
rect 282776 666800 286574 676846
rect 379924 666800 383722 676846
rect 189734 665796 214212 666800
rect 189734 665794 207956 665796
rect 189734 663430 194026 665794
rect 196274 663432 207956 665794
rect 210204 663432 214212 665796
rect 196274 663430 214212 663432
rect 189734 662586 214212 663430
rect 272354 665812 440060 666800
rect 272354 665810 305238 665812
rect 272354 665808 291322 665810
rect 272354 663444 277392 665808
rect 279640 663446 291322 665808
rect 293570 663448 305238 665810
rect 307486 665810 346918 665812
rect 307486 665808 333002 665810
rect 307486 663448 319072 665808
rect 293570 663446 319072 663448
rect 279640 663444 319072 663446
rect 321320 665726 333002 665808
rect 321320 663444 328962 665726
rect 272354 663376 328962 663444
rect 331494 663446 333002 665726
rect 335250 663448 346918 665810
rect 349166 665804 440060 665812
rect 349166 665802 430060 665804
rect 349166 665800 388374 665802
rect 349166 665798 374458 665800
rect 349166 663448 360528 665798
rect 335250 663446 360528 663448
rect 331494 663434 360528 663446
rect 362776 663436 374458 665798
rect 376706 663438 388374 665800
rect 390622 665800 416144 665802
rect 390622 663438 402214 665800
rect 376706 663436 402214 663438
rect 404462 663438 416144 665800
rect 418392 663440 430060 665802
rect 432308 663440 440060 665804
rect 418392 663438 440060 663440
rect 404462 663436 440060 663438
rect 362776 663434 440060 663436
rect 331494 663376 440060 663434
rect 272354 662586 440060 663376
rect 201186 661298 205288 662586
rect 282776 661298 286844 662586
rect 201186 654144 205242 661298
rect 282788 655438 286844 661298
rect 282776 654144 286844 655438
rect 379772 661298 383842 662586
rect 379772 654144 383828 661298
rect 189734 653140 214212 654144
rect 189734 653138 208504 653140
rect 189734 650774 194574 653138
rect 196822 650776 208504 653138
rect 210752 650776 214212 653140
rect 196822 650774 214212 650776
rect 189734 649930 214212 650774
rect 272354 653156 440060 654144
rect 272354 653154 305786 653156
rect 272354 653152 291870 653154
rect 272354 650788 277940 653152
rect 280188 650790 291870 653152
rect 294118 650792 305786 653154
rect 308034 653154 347466 653156
rect 308034 653152 333550 653154
rect 308034 650792 319620 653152
rect 294118 650790 319620 650792
rect 280188 650788 319620 650790
rect 321868 652982 333550 653152
rect 321868 650788 329000 652982
rect 272354 650632 329000 650788
rect 331532 650790 333550 652982
rect 335798 650792 347466 653154
rect 349714 653148 440060 653156
rect 349714 653146 430608 653148
rect 349714 653144 388922 653146
rect 349714 653142 375006 653144
rect 349714 650792 361076 653142
rect 335798 650790 361076 650792
rect 331532 650778 361076 650790
rect 363324 650780 375006 653142
rect 377254 650782 388922 653144
rect 391170 653144 416692 653146
rect 391170 650782 402762 653144
rect 377254 650780 402762 650782
rect 405010 650782 416692 653144
rect 418940 650784 430608 653146
rect 432856 650784 440060 653148
rect 418940 650782 440060 650784
rect 405010 650780 440060 650782
rect 363324 650778 440060 650780
rect 331532 650632 440060 650778
rect 272354 649930 440060 650632
rect 201186 639884 205242 649930
rect 282776 639884 286844 649930
rect 379772 639884 383828 649930
rect 189734 638880 214212 639884
rect 189734 638878 207956 638880
rect 189734 636514 194026 638878
rect 196274 636516 207956 638878
rect 210204 636516 214212 638880
rect 196274 636514 214212 636516
rect 189734 635670 214212 636514
rect 272354 638896 440060 639884
rect 272354 638894 305238 638896
rect 272354 638892 291322 638894
rect 272354 636528 277392 638892
rect 279640 636530 291322 638892
rect 293570 636532 305238 638894
rect 307486 638894 346918 638896
rect 307486 638892 333002 638894
rect 307486 636532 319072 638892
rect 293570 636530 319072 636532
rect 279640 636528 319072 636530
rect 321320 638810 333002 638892
rect 321320 636528 328962 638810
rect 272354 636460 328962 636528
rect 331494 636530 333002 638810
rect 335250 636532 346918 638894
rect 349166 638888 440060 638896
rect 349166 638886 430060 638888
rect 349166 638884 388374 638886
rect 349166 638882 374458 638884
rect 349166 636532 360528 638882
rect 335250 636530 360528 636532
rect 331494 636518 360528 636530
rect 362776 636520 374458 638882
rect 376706 636522 388374 638884
rect 390622 638884 416144 638886
rect 390622 636522 402214 638884
rect 376706 636520 402214 636522
rect 404462 636522 416144 638884
rect 418392 636524 430060 638886
rect 432308 636524 440060 638888
rect 418392 636522 440060 636524
rect 404462 636520 440060 636522
rect 362776 636518 440060 636520
rect 331494 636460 440060 636518
rect 272354 635670 440060 636460
rect 201186 634382 205288 635670
rect 282776 634382 286844 635670
rect 201186 626002 205242 634382
rect 282788 626364 286844 634382
rect 379772 634382 383842 635670
rect 201290 625622 205088 626002
rect 282788 625622 286586 626364
rect 379772 626228 383828 634382
rect 379936 625622 383734 626228
rect 189734 624618 214212 625622
rect 189734 624616 208516 624618
rect 189734 622252 194586 624616
rect 196834 622254 208516 624616
rect 210764 622254 214212 624618
rect 196834 622252 214212 622254
rect 189734 621408 214212 622252
rect 272354 624634 440072 625622
rect 272354 624632 305798 624634
rect 272354 624630 291882 624632
rect 272354 622266 277952 624630
rect 280200 622268 291882 624630
rect 294130 622270 305798 624632
rect 308046 624632 347478 624634
rect 308046 624630 333562 624632
rect 308046 622270 319632 624630
rect 294130 622268 319632 622270
rect 280200 622266 319632 622268
rect 321880 624460 333562 624630
rect 321880 622266 329012 624460
rect 272354 622110 329012 622266
rect 331544 622268 333562 624460
rect 335810 622270 347478 624632
rect 349726 624626 440072 624634
rect 349726 624624 430620 624626
rect 349726 624622 388934 624624
rect 349726 624620 375018 624622
rect 349726 622270 361088 624620
rect 335810 622268 361088 622270
rect 331544 622256 361088 622268
rect 363336 622258 375018 624620
rect 377266 622260 388934 624622
rect 391182 624622 416704 624624
rect 391182 622260 402774 624622
rect 377266 622258 402774 622260
rect 405022 622260 416704 624622
rect 418952 622262 430620 624624
rect 432868 622262 440072 624626
rect 418952 622260 440072 622262
rect 405022 622258 440072 622260
rect 363336 622256 440072 622258
rect 331544 622110 440072 622256
rect 272354 621408 440072 622110
rect 201290 611362 205088 621408
rect 282788 611362 286586 621408
rect 379936 611362 383734 621408
rect 157200 610398 440072 611362
rect 157200 610396 180402 610398
rect 157200 608032 166486 610396
rect 168734 608034 180402 610396
rect 182650 610374 440072 610398
rect 182650 610372 305250 610374
rect 182650 610370 291334 610372
rect 182650 610362 277404 610370
rect 182650 610360 263570 610362
rect 182650 610358 221884 610360
rect 182650 610356 207968 610358
rect 182650 608034 194038 610356
rect 168734 608032 194038 608034
rect 157200 607992 194038 608032
rect 196286 607994 207968 610356
rect 210216 607996 221884 610358
rect 224132 610358 249654 610360
rect 224132 607996 235724 610358
rect 210216 607994 235724 607996
rect 237972 607996 249654 610358
rect 251902 607998 263570 610360
rect 265818 608006 277404 610362
rect 279652 608008 291334 610370
rect 293582 608010 305250 610372
rect 307498 610372 346930 610374
rect 307498 610370 333014 610372
rect 307498 608010 319084 610370
rect 293582 608008 319084 608010
rect 279652 608006 319084 608008
rect 321332 610288 333014 610370
rect 321332 608006 328974 610288
rect 265818 607998 328974 608006
rect 251902 607996 328974 607998
rect 237972 607994 328974 607996
rect 196286 607992 328974 607994
rect 157200 607938 328974 607992
rect 331506 608008 333014 610288
rect 335262 608010 346930 610372
rect 349178 610366 440072 610374
rect 349178 610364 430072 610366
rect 349178 610362 388386 610364
rect 349178 610360 374470 610362
rect 349178 608010 360540 610360
rect 335262 608008 360540 608010
rect 331506 607996 360540 608008
rect 362788 607998 374470 610360
rect 376718 608000 388386 610362
rect 390634 610362 416156 610364
rect 390634 608000 402226 610362
rect 376718 607998 402226 608000
rect 404474 608000 416156 610362
rect 418404 608002 430072 610364
rect 432320 608002 440072 610366
rect 418404 608000 440072 608002
rect 404474 607998 440072 608000
rect 362788 607996 440072 607998
rect 331506 607938 440072 607996
rect 157200 607148 440072 607938
rect 201290 605506 205300 607148
rect 282788 605506 286824 607148
rect 201372 593334 205300 605506
rect 282896 593472 286824 605506
rect 379926 594198 383854 607148
rect 379926 593540 383912 594198
rect 201468 592904 205266 593334
rect 282966 592904 286764 593472
rect 380114 592904 383912 593540
rect 189988 591900 215998 592904
rect 189988 591898 208694 591900
rect 189988 589534 194764 591898
rect 197012 589536 208694 591898
rect 210942 589536 215998 591900
rect 197012 589534 215998 589536
rect 189988 588690 215998 589534
rect 272354 591916 340950 592904
rect 272354 591914 305976 591916
rect 272354 591912 292060 591914
rect 272354 589548 278130 591912
rect 280378 589550 292060 591912
rect 294308 589552 305976 591914
rect 308224 591914 340950 591916
rect 308224 591912 333740 591914
rect 308224 589552 319810 591912
rect 294308 589550 319810 589552
rect 280378 589548 319810 589550
rect 322058 591742 333740 591912
rect 322058 589548 329190 591742
rect 272354 589392 329190 589548
rect 331722 589550 333740 591742
rect 335988 589550 340950 591914
rect 331722 589392 340950 589550
rect 272354 588690 340950 589392
rect 366450 591906 395520 592904
rect 366450 591904 389112 591906
rect 366450 589540 375196 591904
rect 377444 589542 389112 591904
rect 391360 589542 395520 591906
rect 377444 589540 395520 589542
rect 366450 588690 395520 589540
rect 201468 578644 205266 588690
rect 282966 578644 286764 588690
rect 380114 578644 383912 588690
rect 189988 577640 215998 578644
rect 189988 577638 208146 577640
rect 189988 575274 194216 577638
rect 196464 575276 208146 577638
rect 210394 575276 215998 577640
rect 196464 575274 215998 575276
rect 189988 574430 215998 575274
rect 272354 577656 340950 578644
rect 272354 577654 305428 577656
rect 272354 577652 291512 577654
rect 272354 575288 277582 577652
rect 279830 575290 291512 577652
rect 293760 575292 305428 577654
rect 307676 577654 340950 577656
rect 307676 577652 333192 577654
rect 307676 575292 319262 577652
rect 293760 575290 319262 575292
rect 279830 575288 319262 575290
rect 321510 577570 333192 577652
rect 321510 575288 329152 577570
rect 272354 575220 329152 575288
rect 331684 575290 333192 577570
rect 335440 575290 340950 577654
rect 331684 575220 340950 575290
rect 272354 574430 340950 575220
rect 366450 577646 395520 578644
rect 366450 577644 388564 577646
rect 366450 575280 374648 577644
rect 376896 575282 388564 577644
rect 390812 575282 395520 577646
rect 376896 575280 395520 575282
rect 366450 574430 395520 575280
rect 201468 565818 205266 574430
rect 282966 565818 286764 574430
rect 380114 565818 383912 574430
rect 189988 564814 215998 565818
rect 189988 564812 208362 564814
rect 189988 562448 194432 564812
rect 196680 562450 208362 564812
rect 210610 562450 215998 564814
rect 196680 562448 215998 562450
rect 189988 561604 215998 562448
rect 272354 564830 340950 565818
rect 272354 564828 305644 564830
rect 272354 564826 291728 564828
rect 272354 562462 277798 564826
rect 280046 562464 291728 564826
rect 293976 562466 305644 564828
rect 307892 564828 340950 564830
rect 307892 564826 333408 564828
rect 307892 562466 319478 564826
rect 293976 562464 319478 562466
rect 280046 562462 319478 562464
rect 321726 564766 333408 564826
rect 321726 562462 329078 564766
rect 272354 562416 329078 562462
rect 331610 562464 333408 564766
rect 335656 562464 340950 564828
rect 331610 562416 340950 562464
rect 272354 561604 340950 562416
rect 366450 564820 395520 565818
rect 366450 564818 388780 564820
rect 366450 562454 374864 564818
rect 377112 562456 388780 564818
rect 391028 562456 395520 564820
rect 377112 562454 395520 562456
rect 366450 561604 395520 562454
rect 200654 548088 205408 561604
rect 282178 548088 286932 561604
rect 378922 549382 383676 561604
rect 378922 548088 384014 549382
rect 132646 547124 452188 548088
rect 132646 544760 139550 547124
rect 141798 547122 181230 547124
rect 141798 547120 167314 547122
rect 141798 544760 153384 547120
rect 132646 544756 153384 544760
rect 155632 544758 167314 547120
rect 169562 544760 181230 547122
rect 183478 547100 452188 547124
rect 183478 547098 306078 547100
rect 183478 547096 292162 547098
rect 183478 547088 278232 547096
rect 183478 547086 264398 547088
rect 183478 547084 222712 547086
rect 183478 547082 208796 547084
rect 183478 544760 194866 547082
rect 169562 544758 194866 544760
rect 155632 544756 194866 544758
rect 132646 544718 194866 544756
rect 197114 544720 208796 547082
rect 211044 544722 222712 547084
rect 224960 547084 250482 547086
rect 224960 544722 236552 547084
rect 211044 544720 236552 544722
rect 238800 544722 250482 547084
rect 252730 544724 264398 547086
rect 266646 544732 278232 547088
rect 280480 544734 292162 547096
rect 294410 544736 306078 547098
rect 308326 547098 347758 547100
rect 308326 547096 333842 547098
rect 308326 544736 319912 547096
rect 294410 544734 319912 544736
rect 280480 544732 319912 544734
rect 322160 546926 333842 547096
rect 322160 544732 329292 546926
rect 266646 544724 329292 544732
rect 252730 544722 329292 544724
rect 238800 544720 329292 544722
rect 197114 544718 329292 544720
rect 132646 544576 329292 544718
rect 331824 544734 333842 546926
rect 336090 544736 347758 547098
rect 350006 547092 444734 547100
rect 350006 547090 430900 547092
rect 350006 547088 389214 547090
rect 350006 547086 375298 547088
rect 350006 544736 361368 547086
rect 336090 544734 361368 544736
rect 331824 544722 361368 544734
rect 363616 544724 375298 547086
rect 377546 544726 389214 547088
rect 391462 547088 416984 547090
rect 391462 544726 403054 547088
rect 377546 544724 403054 544726
rect 405302 544726 416984 547088
rect 419232 544728 430900 547090
rect 433148 544736 444734 547092
rect 446982 544736 452188 547100
rect 433148 544728 452188 544736
rect 419232 544726 452188 544728
rect 405302 544724 452188 544726
rect 363616 544722 452188 544724
rect 331824 544576 452188 544722
rect 132646 543874 452188 544576
rect 201570 533828 205368 543874
rect 283068 533828 286866 543874
rect 380216 533828 384014 543874
rect 132646 532864 452188 533828
rect 132646 530500 139002 532864
rect 141250 532862 180682 532864
rect 141250 532860 166766 532862
rect 141250 530500 152836 532860
rect 132646 530496 152836 530500
rect 155084 530498 166766 532860
rect 169014 530500 180682 532862
rect 182930 532840 452188 532864
rect 182930 532838 305530 532840
rect 182930 532836 291614 532838
rect 182930 532828 277684 532836
rect 182930 532826 263850 532828
rect 182930 532824 222164 532826
rect 182930 532822 208248 532824
rect 182930 530500 194318 532822
rect 169014 530498 194318 530500
rect 155084 530496 194318 530498
rect 132646 530458 194318 530496
rect 196566 530460 208248 532822
rect 210496 530462 222164 532824
rect 224412 532824 249934 532826
rect 224412 530462 236004 532824
rect 210496 530460 236004 530462
rect 238252 530462 249934 532824
rect 252182 530464 263850 532826
rect 266098 530472 277684 532828
rect 279932 530474 291614 532836
rect 293862 530476 305530 532838
rect 307778 532838 347210 532840
rect 307778 532836 333294 532838
rect 307778 530476 319364 532836
rect 293862 530474 319364 530476
rect 279932 530472 319364 530474
rect 321612 532754 333294 532836
rect 321612 530472 329254 532754
rect 266098 530464 329254 530472
rect 252182 530462 329254 530464
rect 238252 530460 329254 530462
rect 196566 530458 329254 530460
rect 132646 530404 329254 530458
rect 331786 530474 333294 532754
rect 335542 530476 347210 532838
rect 349458 532832 444186 532840
rect 349458 532830 430352 532832
rect 349458 532828 388666 532830
rect 349458 532826 374750 532828
rect 349458 530476 360820 532826
rect 335542 530474 360820 530476
rect 331786 530462 360820 530474
rect 363068 530464 374750 532826
rect 376998 530466 388666 532828
rect 390914 532828 416436 532830
rect 390914 530466 402506 532828
rect 376998 530464 402506 530466
rect 404754 530466 416436 532828
rect 418684 530468 430352 532830
rect 432600 530476 444186 532832
rect 446434 530476 452188 532840
rect 432600 530468 452188 530476
rect 418684 530466 452188 530468
rect 404754 530464 452188 530466
rect 363068 530462 452188 530464
rect 331786 530404 452188 530462
rect 132646 529614 452188 530404
rect 201570 521002 205368 529614
rect 283068 521002 286866 529614
rect 380216 521002 384014 529614
rect 132646 520038 452188 521002
rect 132646 517674 139218 520038
rect 141466 520036 180898 520038
rect 141466 520034 166982 520036
rect 141466 517674 153052 520034
rect 132646 517670 153052 517674
rect 155300 517672 166982 520034
rect 169230 517674 180898 520036
rect 183146 520014 452188 520038
rect 183146 520012 305746 520014
rect 183146 520010 291830 520012
rect 183146 520002 277900 520010
rect 183146 520000 264066 520002
rect 183146 519998 222380 520000
rect 183146 519996 208464 519998
rect 183146 517674 194534 519996
rect 169230 517672 194534 517674
rect 155300 517670 194534 517672
rect 132646 517632 194534 517670
rect 196782 517634 208464 519996
rect 210712 517636 222380 519998
rect 224628 519998 250150 520000
rect 224628 517636 236220 519998
rect 210712 517634 236220 517636
rect 238468 517636 250150 519998
rect 252398 517638 264066 520000
rect 266314 517646 277900 520002
rect 280148 517648 291830 520010
rect 294078 517650 305746 520012
rect 307994 520012 347426 520014
rect 307994 520010 333510 520012
rect 307994 517650 319580 520010
rect 294078 517648 319580 517650
rect 280148 517646 319580 517648
rect 321828 519950 333510 520010
rect 321828 517646 329180 519950
rect 266314 517638 329180 517646
rect 252398 517636 329180 517638
rect 238468 517634 329180 517636
rect 196782 517632 329180 517634
rect 132646 517600 329180 517632
rect 331712 517648 333510 519950
rect 335758 517650 347426 520012
rect 349674 520006 444402 520014
rect 349674 520004 430568 520006
rect 349674 520002 388882 520004
rect 349674 520000 374966 520002
rect 349674 517650 361036 520000
rect 335758 517648 361036 517650
rect 331712 517636 361036 517648
rect 363284 517638 374966 520000
rect 377214 517640 388882 520002
rect 391130 520002 416652 520004
rect 391130 517640 402722 520002
rect 377214 517638 402722 517640
rect 404970 517640 416652 520002
rect 418900 517642 430568 520004
rect 432816 517650 444402 520006
rect 446650 517650 452188 520014
rect 432816 517642 452188 517650
rect 418900 517640 452188 517642
rect 404970 517638 452188 517640
rect 363284 517636 452188 517638
rect 331712 517600 452188 517636
rect 132646 516788 452188 517600
rect 200894 515642 205602 516788
rect 282636 515642 287026 516788
rect 201496 500154 205602 515642
rect 282920 500192 287026 515642
rect 379184 500874 383956 516788
rect 201632 499580 205430 500154
rect 283130 499580 286928 500192
rect 379184 499580 384076 500874
rect 161038 498616 452250 499580
rect 161038 498614 181292 498616
rect 161038 496250 167376 498614
rect 169624 496252 181292 498614
rect 183540 498592 452250 498616
rect 183540 498590 306140 498592
rect 183540 498588 292224 498590
rect 183540 498580 278294 498588
rect 183540 498578 264460 498580
rect 183540 498576 222774 498578
rect 183540 498574 208858 498576
rect 183540 496252 194928 498574
rect 169624 496250 194928 496252
rect 161038 496210 194928 496250
rect 197176 496212 208858 498574
rect 211106 496214 222774 498576
rect 225022 498576 250544 498578
rect 225022 496214 236614 498576
rect 211106 496212 236614 496214
rect 238862 496214 250544 498576
rect 252792 496216 264460 498578
rect 266708 496224 278294 498580
rect 280542 496226 292224 498588
rect 294472 496228 306140 498590
rect 308388 498590 347820 498592
rect 308388 498588 333904 498590
rect 308388 496228 319974 498588
rect 294472 496226 319974 496228
rect 280542 496224 319974 496226
rect 322222 498418 333904 498588
rect 322222 496224 329354 498418
rect 266708 496216 329354 496224
rect 252792 496214 329354 496216
rect 238862 496212 329354 496214
rect 197176 496210 329354 496212
rect 161038 496068 329354 496210
rect 331886 496226 333904 498418
rect 336152 496228 347820 498590
rect 350068 498584 444796 498592
rect 350068 498582 430962 498584
rect 350068 498580 389276 498582
rect 350068 498578 375360 498580
rect 350068 496228 361430 498578
rect 336152 496226 361430 496228
rect 331886 496214 361430 496226
rect 363678 496216 375360 498578
rect 377608 496218 389276 498580
rect 391524 498580 417046 498582
rect 391524 496218 403116 498580
rect 377608 496216 403116 496218
rect 405364 496218 417046 498580
rect 419294 496220 430962 498582
rect 433210 496228 444796 498584
rect 447044 496228 452250 498592
rect 433210 496220 452250 496228
rect 419294 496218 452250 496220
rect 405364 496216 452250 496218
rect 363678 496214 452250 496216
rect 331886 496068 452250 496214
rect 161038 495366 452250 496068
rect 201632 485320 205430 495366
rect 283130 485320 286928 495366
rect 380278 485320 384076 495366
rect 161038 484356 452250 485320
rect 161038 484354 180744 484356
rect 161038 481990 166828 484354
rect 169076 481992 180744 484354
rect 182992 484332 452250 484356
rect 182992 484330 305592 484332
rect 182992 484328 291676 484330
rect 182992 484320 277746 484328
rect 182992 484318 263912 484320
rect 182992 484316 222226 484318
rect 182992 484314 208310 484316
rect 182992 481992 194380 484314
rect 169076 481990 194380 481992
rect 161038 481950 194380 481990
rect 196628 481952 208310 484314
rect 210558 481954 222226 484316
rect 224474 484316 249996 484318
rect 224474 481954 236066 484316
rect 210558 481952 236066 481954
rect 238314 481954 249996 484316
rect 252244 481956 263912 484318
rect 266160 481964 277746 484320
rect 279994 481966 291676 484328
rect 293924 481968 305592 484330
rect 307840 484330 347272 484332
rect 307840 484328 333356 484330
rect 307840 481968 319426 484328
rect 293924 481966 319426 481968
rect 279994 481964 319426 481966
rect 321674 484246 333356 484328
rect 321674 481964 329316 484246
rect 266160 481956 329316 481964
rect 252244 481954 329316 481956
rect 238314 481952 329316 481954
rect 196628 481950 329316 481952
rect 161038 481896 329316 481950
rect 331848 481966 333356 484246
rect 335604 481968 347272 484330
rect 349520 484324 444248 484332
rect 349520 484322 430414 484324
rect 349520 484320 388728 484322
rect 349520 484318 374812 484320
rect 349520 481968 360882 484318
rect 335604 481966 360882 481968
rect 331848 481954 360882 481966
rect 363130 481956 374812 484318
rect 377060 481958 388728 484320
rect 390976 484320 416498 484322
rect 390976 481958 402568 484320
rect 377060 481956 402568 481958
rect 404816 481958 416498 484320
rect 418746 481960 430414 484322
rect 432662 481968 444248 484324
rect 446496 481968 452250 484332
rect 432662 481960 452250 481968
rect 418746 481958 452250 481960
rect 404816 481956 452250 481958
rect 363130 481954 452250 481956
rect 331848 481896 452250 481954
rect 161038 481106 452250 481896
rect 201632 472494 205430 481106
rect 283130 472494 286928 481106
rect 380278 472494 384076 481106
rect 161038 471530 452250 472494
rect 161038 471528 180960 471530
rect 161038 469164 167044 471528
rect 169292 469166 180960 471528
rect 183208 471506 452250 471530
rect 183208 471504 305808 471506
rect 183208 471502 291892 471504
rect 183208 471494 277962 471502
rect 183208 471492 264128 471494
rect 183208 471490 222442 471492
rect 183208 471488 208526 471490
rect 183208 469166 194596 471488
rect 169292 469164 194596 469166
rect 161038 469124 194596 469164
rect 196844 469126 208526 471488
rect 210774 469128 222442 471490
rect 224690 471490 250212 471492
rect 224690 469128 236282 471490
rect 210774 469126 236282 469128
rect 238530 469128 250212 471490
rect 252460 469130 264128 471492
rect 266376 469138 277962 471494
rect 280210 469140 291892 471502
rect 294140 469142 305808 471504
rect 308056 471504 347488 471506
rect 308056 471502 333572 471504
rect 308056 469142 319642 471502
rect 294140 469140 319642 469142
rect 280210 469138 319642 469140
rect 321890 471442 333572 471502
rect 321890 469138 329242 471442
rect 266376 469130 329242 469138
rect 252460 469128 329242 469130
rect 238530 469126 329242 469128
rect 196844 469124 329242 469126
rect 161038 469092 329242 469124
rect 331774 469140 333572 471442
rect 335820 469142 347488 471504
rect 349736 471498 444464 471506
rect 349736 471496 430630 471498
rect 349736 471494 388944 471496
rect 349736 471492 375028 471494
rect 349736 469142 361098 471492
rect 335820 469140 361098 469142
rect 331774 469128 361098 469140
rect 363346 469130 375028 471492
rect 377276 469132 388944 471494
rect 391192 471494 416714 471496
rect 391192 469132 402784 471494
rect 377276 469130 402784 469132
rect 405032 469132 416714 471494
rect 418962 469134 430630 471496
rect 432878 469142 444464 471498
rect 446712 469142 452250 471506
rect 432878 469134 452250 469142
rect 418962 469132 452250 469134
rect 405032 469130 452250 469132
rect 363346 469128 452250 469130
rect 331774 469092 452250 469128
rect 161038 468280 452250 469092
rect 200956 467134 205700 468280
rect 282698 467134 286972 468280
rect 201866 460380 205700 467134
rect 201880 459048 205678 460380
rect 282826 459090 286972 467134
rect 379234 467134 383548 468280
rect 282826 459048 287176 459090
rect 379234 459048 383380 467134
rect 139118 459006 383380 459048
rect 384550 459006 453088 459048
rect 139118 458084 453088 459006
rect 139118 455720 139860 458084
rect 142108 458082 181540 458084
rect 142108 458080 167624 458082
rect 142108 455720 153694 458080
rect 139118 455716 153694 455720
rect 155942 455718 167624 458080
rect 169872 455720 181540 458082
rect 183788 458060 453088 458084
rect 183788 458058 306388 458060
rect 183788 458056 292472 458058
rect 183788 458048 278542 458056
rect 183788 458046 264708 458048
rect 183788 458044 223022 458046
rect 183788 458042 209106 458044
rect 183788 455720 195176 458042
rect 169872 455718 195176 455720
rect 155942 455716 195176 455718
rect 139118 455678 195176 455716
rect 197424 455680 209106 458042
rect 211354 455682 223022 458044
rect 225270 458044 250792 458046
rect 225270 455682 236862 458044
rect 211354 455680 236862 455682
rect 239110 455682 250792 458044
rect 253040 455684 264708 458046
rect 266956 455692 278542 458048
rect 280790 455694 292472 458056
rect 294720 455696 306388 458058
rect 308636 458058 348068 458060
rect 308636 458056 334152 458058
rect 308636 455696 320222 458056
rect 294720 455694 320222 455696
rect 280790 455692 320222 455694
rect 322470 457886 334152 458056
rect 322470 455692 329602 457886
rect 266956 455684 329602 455692
rect 253040 455682 329602 455684
rect 239110 455680 329602 455682
rect 197424 455678 329602 455680
rect 139118 455536 329602 455678
rect 332134 455694 334152 457886
rect 336400 455696 348068 458058
rect 350316 458052 445044 458060
rect 350316 458050 431210 458052
rect 350316 458048 389524 458050
rect 350316 458046 375608 458048
rect 350316 455696 361678 458046
rect 336400 455694 361678 455696
rect 332134 455682 361678 455694
rect 363926 455684 375608 458046
rect 377856 455686 389524 458048
rect 391772 458048 417294 458050
rect 391772 455686 403364 458048
rect 377856 455684 403364 455686
rect 405612 455686 417294 458048
rect 419542 455688 431210 458050
rect 433458 455696 445044 458052
rect 447292 455696 453088 458060
rect 433458 455688 453088 455696
rect 419542 455686 453088 455688
rect 405612 455684 453088 455686
rect 363926 455682 453088 455684
rect 332134 455536 453088 455682
rect 139118 454834 453088 455536
rect 201768 453774 205678 454834
rect 283378 453774 287308 454834
rect 201768 447324 205672 453774
rect 283404 449552 287308 453774
rect 283338 447324 287308 449552
rect 380358 453774 384324 454834
rect 380358 449552 384262 453774
rect 380358 447324 384284 449552
rect 139118 446360 453088 447324
rect 139118 443996 139820 446360
rect 142068 446358 181500 446360
rect 142068 446356 167584 446358
rect 142068 443996 153654 446356
rect 139118 443992 153654 443996
rect 155902 443994 167584 446356
rect 169832 443996 181500 446358
rect 183748 446336 453088 446360
rect 183748 446334 306348 446336
rect 183748 446332 292432 446334
rect 183748 446324 278502 446332
rect 183748 446322 264668 446324
rect 183748 446320 222982 446322
rect 183748 446318 209066 446320
rect 183748 443996 195136 446318
rect 169832 443994 195136 443996
rect 155902 443992 195136 443994
rect 139118 443954 195136 443992
rect 197384 443956 209066 446318
rect 211314 443958 222982 446320
rect 225230 446320 250752 446322
rect 225230 443958 236822 446320
rect 211314 443956 236822 443958
rect 239070 443958 250752 446320
rect 253000 443960 264668 446322
rect 266916 443968 278502 446324
rect 280750 443970 292432 446332
rect 294680 443972 306348 446334
rect 308596 446334 348028 446336
rect 308596 446332 334112 446334
rect 308596 443972 320182 446332
rect 294680 443970 320182 443972
rect 280750 443968 320182 443970
rect 322430 446162 334112 446332
rect 322430 443968 329562 446162
rect 266916 443960 329562 443968
rect 253000 443958 329562 443960
rect 239070 443956 329562 443958
rect 197384 443954 329562 443956
rect 139118 443812 329562 443954
rect 332094 443970 334112 446162
rect 336360 443972 348028 446334
rect 350276 446328 445004 446336
rect 350276 446326 431170 446328
rect 350276 446324 389484 446326
rect 350276 446322 375568 446324
rect 350276 443972 361638 446322
rect 336360 443970 361638 443972
rect 332094 443958 361638 443970
rect 363886 443960 375568 446322
rect 377816 443962 389484 446324
rect 391732 446324 417254 446326
rect 391732 443962 403324 446324
rect 377816 443960 403324 443962
rect 405572 443962 417254 446324
rect 419502 443964 431170 446326
rect 433418 443972 445004 446328
rect 447252 443972 453088 446336
rect 433418 443964 453088 443972
rect 419502 443962 453088 443964
rect 405572 443960 453088 443962
rect 363886 443958 453088 443960
rect 332094 443812 453088 443958
rect 139118 443110 453088 443812
rect 118094 424360 121998 441392
rect 201768 426590 205672 443110
rect 283338 442050 287308 443110
rect 201768 425338 205718 426590
rect 118168 423198 121966 424360
rect 132016 423198 193354 423314
rect 201920 423198 205718 425338
rect 283404 424954 287308 442050
rect 380358 442050 384284 443110
rect 380358 433602 384262 442050
rect 283418 423198 287216 424954
rect 36446 423156 62048 423198
rect 67192 423156 217042 423198
rect 36446 422232 217042 423156
rect 36446 422230 125984 422232
rect 36446 422222 112054 422230
rect 36446 422220 98220 422222
rect 36446 422218 56534 422220
rect 36446 419854 42618 422218
rect 44866 419856 56534 422218
rect 58782 422218 84304 422220
rect 58782 419856 70374 422218
rect 44866 419854 70374 419856
rect 72622 419856 84304 422218
rect 86552 419858 98220 422220
rect 100468 419866 112054 422222
rect 114302 419868 125984 422230
rect 128232 422194 217042 422232
rect 128232 422192 209146 422194
rect 128232 419868 195216 422192
rect 114302 419866 195216 419868
rect 100468 419858 195216 419866
rect 86552 419856 195216 419858
rect 72622 419854 195216 419856
rect 36446 419828 195216 419854
rect 197464 419830 209146 422192
rect 211394 419830 217042 422194
rect 197464 419828 217042 419830
rect 36446 419116 217042 419828
rect 36446 418984 134366 419116
rect 189818 418984 217042 419116
rect 272496 422210 341056 423198
rect 272496 422208 306428 422210
rect 272496 422206 292512 422208
rect 272496 419842 278582 422206
rect 280830 419844 292512 422206
rect 294760 419846 306428 422208
rect 308676 422208 341056 422210
rect 308676 422206 334192 422208
rect 308676 419846 320262 422206
rect 294760 419844 320262 419846
rect 280830 419842 320262 419844
rect 322510 422036 334192 422206
rect 322510 419842 329642 422036
rect 272496 419686 329642 419842
rect 332174 419844 334192 422036
rect 336440 419844 341056 422208
rect 332174 419686 341056 419844
rect 272496 418984 341056 419686
rect 62476 408938 66274 418984
rect 118168 408938 121966 418984
rect 201920 408938 205718 418984
rect 283418 408938 287216 418984
rect 36446 407972 134366 408938
rect 36446 407970 125436 407972
rect 36446 407962 111506 407970
rect 36446 407960 97672 407962
rect 36446 407958 55986 407960
rect 36446 405594 42070 407958
rect 44318 405596 55986 407958
rect 58234 407958 83756 407960
rect 58234 405596 69826 407958
rect 44318 405594 69826 405596
rect 72074 405596 83756 407958
rect 86004 405598 97672 407960
rect 99920 405606 111506 407962
rect 113754 405608 125436 407970
rect 127684 405608 134366 407972
rect 113754 405606 134366 405608
rect 99920 405598 134366 405606
rect 86004 405596 134366 405598
rect 72074 405594 134366 405596
rect 36446 404724 134366 405594
rect 189818 407934 217042 408938
rect 189818 407932 208598 407934
rect 189818 405568 194668 407932
rect 196916 405570 208598 407932
rect 210846 405570 217042 407934
rect 196916 405568 217042 405570
rect 189818 404724 217042 405568
rect 272496 407950 341056 408938
rect 272496 407948 305880 407950
rect 272496 407946 291964 407948
rect 272496 405582 278034 407946
rect 280282 405584 291964 407946
rect 294212 405586 305880 407948
rect 308128 407948 341056 407950
rect 308128 407946 333644 407948
rect 308128 405586 319714 407946
rect 294212 405584 319714 405586
rect 280282 405582 319714 405584
rect 321962 407864 333644 407946
rect 321962 405582 329604 407864
rect 272496 405514 329604 405582
rect 332136 405584 333644 407864
rect 335892 405584 341056 407948
rect 332136 405514 341056 405584
rect 272496 404724 341056 405514
rect 62476 396112 66274 404724
rect 118168 396112 121966 404724
rect 201920 396112 205718 404724
rect 283418 396112 287216 404724
rect 36446 395146 134366 396112
rect 36446 395144 125652 395146
rect 36446 395136 111722 395144
rect 36446 395134 97888 395136
rect 36446 395132 56202 395134
rect 36446 392768 42286 395132
rect 44534 392770 56202 395132
rect 58450 395132 83972 395134
rect 58450 392770 70042 395132
rect 44534 392768 70042 392770
rect 72290 392770 83972 395132
rect 86220 392772 97888 395134
rect 100136 392780 111722 395136
rect 113970 392782 125652 395144
rect 127900 392782 134366 395146
rect 113970 392780 134366 392782
rect 100136 392772 134366 392780
rect 86220 392770 134366 392772
rect 72290 392768 134366 392770
rect 36446 391898 134366 392768
rect 189818 395108 217042 396112
rect 189818 395106 208814 395108
rect 189818 392742 194884 395106
rect 197132 392744 208814 395106
rect 211062 392744 217042 395108
rect 197132 392742 217042 392744
rect 189818 391898 217042 392742
rect 272496 395124 341056 396112
rect 272496 395122 306096 395124
rect 272496 395120 292180 395122
rect 272496 392756 278250 395120
rect 280498 392758 292180 395120
rect 294428 392760 306096 395122
rect 308344 395122 341056 395124
rect 308344 395120 333860 395122
rect 308344 392760 319930 395120
rect 294428 392758 319930 392760
rect 280498 392756 319930 392758
rect 322178 395060 333860 395120
rect 322178 392756 329530 395060
rect 272496 392710 329530 392756
rect 332062 392758 333860 395060
rect 336108 392758 341056 395122
rect 332062 392710 341056 392758
rect 272496 391898 341056 392710
rect 61828 391772 66008 391898
rect 117370 391856 121550 391898
rect 201244 389352 205424 391898
rect 282986 389352 287166 391898
rect 201244 387412 205692 389352
rect 282986 387412 287190 389352
rect 189818 386408 217042 387412
rect 189818 386406 209120 386408
rect 189818 384042 195190 386406
rect 197438 384044 209120 386406
rect 211368 384044 217042 386408
rect 197438 384042 217042 384044
rect 189818 383198 217042 384042
rect 272496 386424 341056 387412
rect 272496 386422 306402 386424
rect 272496 386420 292486 386422
rect 272496 384056 278556 386420
rect 280804 384058 292486 386420
rect 294734 384060 306402 386422
rect 308650 386422 341056 386424
rect 308650 386420 334166 386422
rect 308650 384060 320236 386420
rect 294734 384058 320236 384060
rect 280804 384056 320236 384058
rect 322484 386250 334166 386420
rect 322484 384056 329616 386250
rect 272496 383900 329616 384056
rect 332148 384058 334166 386250
rect 336414 384058 341056 386422
rect 332148 383900 341056 384058
rect 272496 383198 341056 383900
rect 201894 373152 205692 383198
rect 283392 373152 287190 383198
rect 380240 379726 384302 433602
rect 534744 424916 538648 430872
rect 534836 423198 538634 424916
rect 521028 422216 550770 423198
rect 521028 422214 542806 422216
rect 521028 419850 528890 422214
rect 531138 419852 542806 422214
rect 545054 419852 550770 422216
rect 531138 419850 550770 419852
rect 521028 418984 550770 419850
rect 534836 408938 538634 418984
rect 521028 407956 550770 408938
rect 521028 407954 542258 407956
rect 521028 405590 528342 407954
rect 530590 405592 542258 407954
rect 544506 405592 550770 407956
rect 530590 405590 550770 405592
rect 521028 404724 550770 405590
rect 534836 396112 538634 404724
rect 521028 395130 550770 396112
rect 521028 395128 542474 395130
rect 521028 392764 528558 395128
rect 530806 392766 542474 395128
rect 544722 392766 550770 395130
rect 530806 392764 550770 392766
rect 521028 391898 550770 392764
rect 534610 387412 538790 391898
rect 521028 386430 550770 387412
rect 521028 386428 542780 386430
rect 521028 384064 528864 386428
rect 531112 384066 542780 386428
rect 545028 384066 550770 386430
rect 531112 384064 550770 384066
rect 521028 383198 550770 384064
rect 380240 377816 384338 379726
rect 380540 373152 384338 377816
rect 465106 373152 468904 379726
rect 534810 373152 538608 383198
rect 147056 372188 217042 373152
rect 147056 372186 181006 372188
rect 147056 372184 167090 372186
rect 147056 369820 153160 372184
rect 155408 369822 167090 372184
rect 169338 369824 181006 372186
rect 183254 372148 217042 372188
rect 183254 372146 208572 372148
rect 183254 369824 194642 372146
rect 169338 369822 194642 369824
rect 155408 369820 194642 369822
rect 147056 369782 194642 369820
rect 196890 369784 208572 372146
rect 210820 369784 217042 372148
rect 196890 369782 217042 369784
rect 147056 368938 217042 369782
rect 272496 373076 559818 373152
rect 272496 372170 561904 373076
rect 272496 372168 542232 372170
rect 272496 372166 472356 372168
rect 272496 372164 458440 372166
rect 272496 372162 305854 372164
rect 272496 372160 291938 372162
rect 272496 369796 278008 372160
rect 280256 369798 291938 372160
rect 294186 369800 305854 372162
rect 308102 372162 347534 372164
rect 308102 372160 333618 372162
rect 308102 369800 319688 372160
rect 294186 369798 319688 369800
rect 280256 369796 319688 369798
rect 321936 372078 333618 372160
rect 321936 369796 329578 372078
rect 272496 369728 329578 369796
rect 332110 369798 333618 372078
rect 335866 369800 347534 372162
rect 349782 372156 444510 372164
rect 349782 372154 430676 372156
rect 349782 372152 388990 372154
rect 349782 372150 375074 372152
rect 349782 369800 361144 372150
rect 335866 369798 361144 369800
rect 332110 369786 361144 369798
rect 363392 369788 375074 372150
rect 377322 369790 388990 372152
rect 391238 372152 416760 372154
rect 391238 369790 402830 372152
rect 377322 369788 402830 369790
rect 405078 369790 416760 372152
rect 419008 369792 430676 372154
rect 432924 369800 444510 372156
rect 446758 369802 458440 372164
rect 460688 369804 472356 372166
rect 474604 372166 514036 372168
rect 474604 372164 500120 372166
rect 474604 369804 486190 372164
rect 460688 369802 486190 369804
rect 446758 369800 486190 369802
rect 488438 369802 500120 372164
rect 502368 369804 514036 372166
rect 516284 369804 528316 372168
rect 530564 369806 542232 372168
rect 544480 372150 561904 372170
rect 544480 369806 556504 372150
rect 530564 369804 556504 369806
rect 502368 369802 556504 369804
rect 488438 369800 556504 369802
rect 432924 369792 556504 369800
rect 419008 369790 556504 369792
rect 405078 369788 556504 369790
rect 363392 369786 556504 369788
rect 558752 369786 561904 372150
rect 332110 369728 561904 369786
rect 272496 368976 561904 369728
rect 272496 368938 559818 368976
rect 201894 360326 205692 368938
rect 283392 360326 287190 368938
rect 380540 360326 384338 368938
rect 465106 360326 468904 368938
rect 534810 360326 538608 368938
rect 147056 360250 560034 360326
rect 147056 359362 562120 360250
rect 147056 359360 181222 359362
rect 147056 359358 167306 359360
rect 147056 356994 153376 359358
rect 155624 356996 167306 359358
rect 169554 356998 181222 359360
rect 183470 359344 562120 359362
rect 183470 359342 542448 359344
rect 183470 359340 472572 359342
rect 183470 359338 458656 359340
rect 183470 359336 306070 359338
rect 183470 359334 292154 359336
rect 183470 359326 278224 359334
rect 183470 359324 264390 359326
rect 183470 359322 222704 359324
rect 183470 359320 208788 359322
rect 183470 356998 194858 359320
rect 169554 356996 194858 356998
rect 155624 356994 194858 356996
rect 147056 356956 194858 356994
rect 197106 356958 208788 359320
rect 211036 356960 222704 359322
rect 224952 359322 250474 359324
rect 224952 356960 236544 359322
rect 211036 356958 236544 356960
rect 238792 356960 250474 359322
rect 252722 356962 264390 359324
rect 266638 356970 278224 359326
rect 280472 356972 292154 359334
rect 294402 356974 306070 359336
rect 308318 359336 347750 359338
rect 308318 359334 333834 359336
rect 308318 356974 319904 359334
rect 294402 356972 319904 356974
rect 280472 356970 319904 356972
rect 322152 359274 333834 359334
rect 322152 356970 329504 359274
rect 266638 356962 329504 356970
rect 252722 356960 329504 356962
rect 238792 356958 329504 356960
rect 197106 356956 329504 356958
rect 147056 356924 329504 356956
rect 332036 356972 333834 359274
rect 336082 356974 347750 359336
rect 349998 359330 444726 359338
rect 349998 359328 430892 359330
rect 349998 359326 389206 359328
rect 349998 359324 375290 359326
rect 349998 356974 361360 359324
rect 336082 356972 361360 356974
rect 332036 356960 361360 356972
rect 363608 356962 375290 359324
rect 377538 356964 389206 359326
rect 391454 359326 416976 359328
rect 391454 356964 403046 359326
rect 377538 356962 403046 356964
rect 405294 356964 416976 359326
rect 419224 356966 430892 359328
rect 433140 356974 444726 359330
rect 446974 356976 458656 359338
rect 460904 356978 472572 359340
rect 474820 359340 514252 359342
rect 474820 359338 500336 359340
rect 474820 356978 486406 359338
rect 460904 356976 486406 356978
rect 446974 356974 486406 356976
rect 488654 356976 500336 359338
rect 502584 356978 514252 359340
rect 516500 356978 528532 359342
rect 530780 356980 542448 359342
rect 544696 359324 562120 359344
rect 544696 356980 556720 359324
rect 530780 356978 556720 356980
rect 502584 356976 556720 356978
rect 488654 356974 556720 356976
rect 433140 356966 556720 356974
rect 419224 356964 556720 356966
rect 405294 356962 556720 356964
rect 363608 356960 556720 356962
rect 558968 356960 562120 359324
rect 332036 356924 562120 356960
rect 147056 356150 562120 356924
rect 147056 356112 560034 356150
rect 201218 352716 205660 356112
rect 201348 348498 205660 352716
rect 282924 348498 287236 356112
rect 379630 352716 384084 356112
rect 379772 348498 384084 352716
rect 464342 352716 468538 356112
rect 534532 352716 538764 356112
rect 464342 350022 468530 352716
rect 534532 350022 538720 352716
rect 464342 348498 468550 350022
rect 534456 348498 538720 350022
rect 130354 348422 559464 348498
rect 130354 347534 561550 348422
rect 130354 345170 138972 347534
rect 141220 347532 180652 347534
rect 141220 347530 166736 347532
rect 141220 345170 152806 347530
rect 130354 345166 152806 345170
rect 155054 345168 166736 347530
rect 168984 345170 180652 347532
rect 182900 347516 561550 347534
rect 182900 347514 541878 347516
rect 182900 347512 472002 347514
rect 182900 347510 458086 347512
rect 182900 347508 305500 347510
rect 182900 347506 291584 347508
rect 182900 347498 277654 347506
rect 182900 347496 263820 347498
rect 182900 347494 222134 347496
rect 182900 347492 208218 347494
rect 182900 345170 194288 347492
rect 168984 345168 194288 345170
rect 155054 345166 194288 345168
rect 130354 345128 194288 345166
rect 196536 345130 208218 347492
rect 210466 345132 222134 347494
rect 224382 347494 249904 347496
rect 224382 345132 235974 347494
rect 210466 345130 235974 345132
rect 238222 345132 249904 347494
rect 252152 345134 263820 347496
rect 266068 345142 277654 347498
rect 279902 345144 291584 347506
rect 293832 345146 305500 347508
rect 307748 347508 347180 347510
rect 307748 347506 333264 347508
rect 307748 345146 319334 347506
rect 293832 345144 319334 345146
rect 279902 345142 319334 345144
rect 321582 347424 333264 347506
rect 321582 345142 329224 347424
rect 266068 345134 329224 345142
rect 252152 345132 329224 345134
rect 238222 345130 329224 345132
rect 196536 345128 329224 345130
rect 130354 345074 329224 345128
rect 331756 345144 333264 347424
rect 335512 345146 347180 347508
rect 349428 347502 444156 347510
rect 349428 347500 430322 347502
rect 349428 347498 388636 347500
rect 349428 347496 374720 347498
rect 349428 345146 360790 347496
rect 335512 345144 360790 345146
rect 331756 345132 360790 345144
rect 363038 345134 374720 347496
rect 376968 345136 388636 347498
rect 390884 347498 416406 347500
rect 390884 345136 402476 347498
rect 376968 345134 402476 345136
rect 404724 345136 416406 347498
rect 418654 345138 430322 347500
rect 432570 345146 444156 347502
rect 446404 345148 458086 347510
rect 460334 345150 472002 347512
rect 474250 347512 513682 347514
rect 474250 347510 499766 347512
rect 474250 345150 485836 347510
rect 460334 345148 485836 345150
rect 446404 345146 485836 345148
rect 488084 345148 499766 347510
rect 502014 345150 513682 347512
rect 515930 345150 527962 347514
rect 530210 345152 541878 347514
rect 544126 347496 561550 347516
rect 544126 345152 556150 347496
rect 530210 345150 556150 345152
rect 502014 345148 556150 345150
rect 488084 345146 556150 345148
rect 432570 345138 556150 345146
rect 418654 345136 556150 345138
rect 404724 345134 556150 345136
rect 363038 345132 556150 345134
rect 558398 345132 561550 347496
rect 331756 345074 561550 345132
rect 130354 344322 561550 345074
rect 130354 344284 559464 344322
rect 201348 335672 205660 344284
rect 282924 335672 287236 344284
rect 379772 335672 384084 344284
rect 464342 335672 468550 344284
rect 534456 335672 538720 344284
rect 130354 335596 559680 335672
rect 130354 334708 561766 335596
rect 130354 332344 139188 334708
rect 141436 334706 180868 334708
rect 141436 334704 166952 334706
rect 141436 332344 153022 334704
rect 130354 332340 153022 332344
rect 155270 332342 166952 334704
rect 169200 332344 180868 334706
rect 183116 334690 561766 334708
rect 183116 334688 542094 334690
rect 183116 334686 472218 334688
rect 183116 334684 458302 334686
rect 183116 334682 305716 334684
rect 183116 334680 291800 334682
rect 183116 334672 277870 334680
rect 183116 334670 264036 334672
rect 183116 334668 222350 334670
rect 183116 334666 208434 334668
rect 183116 332344 194504 334666
rect 169200 332342 194504 332344
rect 155270 332340 194504 332342
rect 130354 332302 194504 332340
rect 196752 332304 208434 334666
rect 210682 332306 222350 334668
rect 224598 334668 250120 334670
rect 224598 332306 236190 334668
rect 210682 332304 236190 332306
rect 238438 332306 250120 334668
rect 252368 332308 264036 334670
rect 266284 332316 277870 334672
rect 280118 332318 291800 334680
rect 294048 332320 305716 334682
rect 307964 334682 347396 334684
rect 307964 334680 333480 334682
rect 307964 332320 319550 334680
rect 294048 332318 319550 332320
rect 280118 332316 319550 332318
rect 321798 334620 333480 334680
rect 321798 332316 329150 334620
rect 266284 332308 329150 332316
rect 252368 332306 329150 332308
rect 238438 332304 329150 332306
rect 196752 332302 329150 332304
rect 130354 332270 329150 332302
rect 331682 332318 333480 334620
rect 335728 332320 347396 334682
rect 349644 334676 444372 334684
rect 349644 334674 430538 334676
rect 349644 334672 388852 334674
rect 349644 334670 374936 334672
rect 349644 332320 361006 334670
rect 335728 332318 361006 332320
rect 331682 332306 361006 332318
rect 363254 332308 374936 334670
rect 377184 332310 388852 334672
rect 391100 334672 416622 334674
rect 391100 332310 402692 334672
rect 377184 332308 402692 332310
rect 404940 332310 416622 334672
rect 418870 332312 430538 334674
rect 432786 332320 444372 334676
rect 446620 332322 458302 334684
rect 460550 332324 472218 334686
rect 474466 334686 513898 334688
rect 474466 334684 499982 334686
rect 474466 332324 486052 334684
rect 460550 332322 486052 332324
rect 446620 332320 486052 332322
rect 488300 332322 499982 334684
rect 502230 332324 513898 334686
rect 516146 332324 528178 334688
rect 530426 332326 542094 334688
rect 544342 334670 561766 334690
rect 544342 332326 556366 334670
rect 530426 332324 556366 332326
rect 502230 332322 556366 332324
rect 488300 332320 556366 332322
rect 432786 332312 556366 332320
rect 418870 332310 556366 332312
rect 404940 332308 556366 332310
rect 363254 332306 556366 332308
rect 558614 332306 561766 334670
rect 331682 332270 561766 332306
rect 130354 331496 561766 332270
rect 130354 331458 559680 331496
rect 200864 329970 205660 331458
rect 282606 329970 287236 331458
rect 379276 329970 384084 331458
rect 464004 329970 468530 331458
rect 534230 329970 538720 331458
rect 201348 320994 205660 329970
rect 282924 320994 287236 329970
rect 379772 320994 384084 329970
rect 464342 320996 468530 329970
rect 37268 320016 76392 320994
rect 37268 320014 57356 320016
rect 37268 317650 43440 320014
rect 45688 317652 57356 320014
rect 59604 320014 76392 320016
rect 59604 317652 71196 320014
rect 45688 317650 71196 317652
rect 73444 317650 76392 320014
rect 37268 316788 76392 317650
rect 37268 316780 62200 316788
rect 62628 311328 66654 316788
rect 68330 316780 76392 316788
rect 108656 320028 133862 320994
rect 108656 320026 126806 320028
rect 108656 317662 112876 320026
rect 115124 317664 126806 320026
rect 129054 317664 133862 320028
rect 115124 317662 133862 317664
rect 108656 316780 133862 317662
rect 190322 319990 217042 320994
rect 190322 319988 209968 319990
rect 190322 317624 196038 319988
rect 198286 317626 209968 319988
rect 212216 317626 217042 319990
rect 198286 317624 217042 317626
rect 190322 316780 217042 317624
rect 273502 320976 287236 320994
rect 288504 320976 343072 320994
rect 273502 320098 343072 320976
rect 273502 320006 329682 320098
rect 273502 320004 307250 320006
rect 273502 320002 293334 320004
rect 273502 317638 279404 320002
rect 281652 317640 293334 320002
rect 295582 317642 307250 320004
rect 309498 320002 329682 320006
rect 309498 317642 321084 320002
rect 295582 317640 321084 317642
rect 281652 317638 321084 317640
rect 323332 317748 329682 320002
rect 332214 320004 343072 320098
rect 332214 317748 335014 320004
rect 323332 317640 335014 317748
rect 337262 317640 343072 320004
rect 323332 317638 343072 317640
rect 273502 316780 343072 317638
rect 370800 319996 395502 320994
rect 370800 319994 390386 319996
rect 370800 317630 376470 319994
rect 378718 317632 390386 319994
rect 392634 317632 395502 319996
rect 378718 317630 395502 317632
rect 370800 316780 395502 317630
rect 454988 320008 507460 320996
rect 534532 320974 538720 329970
rect 454988 320000 501264 320008
rect 454988 319998 487430 320000
rect 454988 319996 473514 319998
rect 454988 317632 459584 319996
rect 461832 317634 473514 319996
rect 475762 317636 487430 319998
rect 489678 317644 501264 320000
rect 503512 317644 507460 320008
rect 489678 317636 507460 317644
rect 475762 317634 507460 317636
rect 461832 317632 507460 317634
rect 454988 316782 507460 317632
rect 507574 319986 562924 320974
rect 507574 319978 556728 319986
rect 507574 319976 542894 319978
rect 507574 319974 528978 319976
rect 507574 317610 515048 319974
rect 517296 317612 528978 319974
rect 531226 317614 542894 319976
rect 545142 317622 556728 319978
rect 558976 317622 562924 319986
rect 545142 317614 562924 317622
rect 531226 317612 562924 317614
rect 517296 317610 562924 317612
rect 118248 316650 122788 316780
rect 202180 316650 206540 316780
rect 282924 316752 288038 316780
rect 283526 316650 288038 316752
rect 380680 316720 385186 316780
rect 118248 311328 122274 316650
rect 202180 311328 206206 316650
rect 283526 311328 287552 316650
rect 380680 311328 384706 316720
rect 464342 311330 468530 316782
rect 507574 316760 562924 317610
rect 37838 310350 76392 311328
rect 37838 310348 57926 310350
rect 37838 307984 44010 310348
rect 46258 307986 57926 310348
rect 60174 310348 76392 310350
rect 60174 307986 71766 310348
rect 46258 307984 71766 307986
rect 74014 307984 76392 310348
rect 37838 307122 76392 307984
rect 37838 307114 66654 307122
rect 68900 307114 76392 307122
rect 108656 310362 133862 311328
rect 108656 310360 127376 310362
rect 108656 307996 113446 310360
rect 115694 307998 127376 310360
rect 129624 307998 133862 310362
rect 115694 307996 133862 307998
rect 108656 307114 133862 307996
rect 190322 310324 217042 311328
rect 190322 310322 210538 310324
rect 190322 307958 196608 310322
rect 198856 307960 210538 310322
rect 212786 307960 217042 310324
rect 198856 307958 217042 307960
rect 190322 307114 217042 307958
rect 273502 310418 343072 311328
rect 273502 310340 329644 310418
rect 273502 310338 307820 310340
rect 273502 310336 293904 310338
rect 273502 307972 279974 310336
rect 282222 307974 293904 310336
rect 296152 307976 307820 310338
rect 310068 310336 329644 310340
rect 310068 307976 321654 310336
rect 296152 307974 321654 307976
rect 282222 307972 321654 307974
rect 323902 308068 329644 310336
rect 332176 310338 343072 310418
rect 332176 308068 335584 310338
rect 323902 307974 335584 308068
rect 337832 307974 343072 310338
rect 323902 307972 343072 307974
rect 273502 307114 343072 307972
rect 370800 310330 395502 311328
rect 370800 310328 390956 310330
rect 370800 307964 377040 310328
rect 379288 307966 390956 310328
rect 393204 307966 395502 310330
rect 379288 307964 395502 307966
rect 370800 307114 395502 307964
rect 454988 311308 508030 311330
rect 534532 311308 538720 316760
rect 454988 310342 563494 311308
rect 454988 310334 501834 310342
rect 454988 310332 488000 310334
rect 454988 310330 474084 310332
rect 454988 307966 460154 310330
rect 462402 307968 474084 310330
rect 476332 307970 488000 310332
rect 490248 307978 501834 310334
rect 504082 310320 563494 310342
rect 504082 310312 557298 310320
rect 504082 310310 543464 310312
rect 504082 310308 529548 310310
rect 504082 307978 515618 310308
rect 490248 307970 515618 307978
rect 476332 307968 515618 307970
rect 462402 307966 515618 307968
rect 454988 307944 515618 307966
rect 517866 307946 529548 310308
rect 531796 307948 543464 310310
rect 545712 307956 557298 310312
rect 559546 307956 563494 310320
rect 545712 307948 563494 307956
rect 531796 307946 563494 307948
rect 517866 307944 563494 307946
rect 454988 307116 563494 307944
rect 62628 300808 66654 307114
rect 118248 306984 123358 307114
rect 202180 306984 207110 307114
rect 283526 306984 288608 307114
rect 380680 307054 385756 307114
rect 118248 300808 122274 306984
rect 202180 300808 206206 306984
rect 283526 300808 287552 306984
rect 380680 300808 384706 307054
rect 464342 300810 468530 307116
rect 507574 307094 563494 307116
rect 37980 299830 76392 300808
rect 37980 299828 58068 299830
rect 37980 297464 44152 299828
rect 46400 297466 58068 299828
rect 60316 299828 76392 299830
rect 60316 297466 71908 299828
rect 46400 297464 71908 297466
rect 74156 297464 76392 299828
rect 37980 296602 76392 297464
rect 37980 296594 66654 296602
rect 69042 296594 76392 296602
rect 108656 299842 133862 300808
rect 108656 299840 127518 299842
rect 108656 297476 113588 299840
rect 115836 297478 127518 299840
rect 129766 297478 133862 299842
rect 115836 297476 133862 297478
rect 108656 296594 133862 297476
rect 190322 299804 217042 300808
rect 190322 299802 210680 299804
rect 190322 297438 196750 299802
rect 198998 297440 210680 299802
rect 212928 297440 217042 299804
rect 198998 297438 217042 297440
rect 190322 296594 217042 297438
rect 273502 299878 343072 300808
rect 273502 299820 329606 299878
rect 273502 299818 307962 299820
rect 273502 299816 294046 299818
rect 273502 297452 280116 299816
rect 282364 297454 294046 299816
rect 296294 297456 307962 299818
rect 310210 299816 329606 299820
rect 310210 297456 321796 299816
rect 296294 297454 321796 297456
rect 282364 297452 321796 297454
rect 324044 297528 329606 299816
rect 332138 299818 343072 299878
rect 332138 297528 335726 299818
rect 324044 297454 335726 297528
rect 337974 297454 343072 299818
rect 324044 297452 343072 297454
rect 273502 296594 343072 297452
rect 370800 299810 395502 300808
rect 370800 299808 391098 299810
rect 370800 297444 377182 299808
rect 379430 297446 391098 299808
rect 393346 297446 395502 299810
rect 379430 297444 395502 297446
rect 370800 296594 395502 297444
rect 454988 300788 508172 300810
rect 534532 300788 538720 307094
rect 454988 299822 563636 300788
rect 454988 299814 501976 299822
rect 454988 299812 488142 299814
rect 454988 299810 474226 299812
rect 454988 297446 460296 299810
rect 462544 297448 474226 299810
rect 476474 297450 488142 299812
rect 490390 297458 501976 299814
rect 504224 299800 563636 299822
rect 504224 299792 557440 299800
rect 504224 299790 543606 299792
rect 504224 299788 529690 299790
rect 504224 297458 515760 299788
rect 490390 297450 515760 297458
rect 476474 297448 515760 297450
rect 462544 297446 515760 297448
rect 454988 297424 515760 297446
rect 518008 297426 529690 299788
rect 531938 297428 543606 299790
rect 545854 297436 557440 299792
rect 559688 297436 563636 299800
rect 545854 297428 563636 297436
rect 531938 297426 563636 297428
rect 518008 297424 563636 297426
rect 454988 296596 563636 297424
rect 62628 289860 66654 296594
rect 118248 296464 123500 296594
rect 202180 296464 207252 296594
rect 283526 296464 288750 296594
rect 380680 296534 385898 296594
rect 507574 296574 563636 296596
rect 118248 289860 122274 296464
rect 202180 289860 206206 296464
rect 283526 289860 287552 296464
rect 380680 289860 384706 296534
rect 37838 288882 76392 289860
rect 37838 288880 57926 288882
rect 37838 286516 44010 288880
rect 46258 286518 57926 288880
rect 60174 288880 76392 288882
rect 60174 286518 71766 288880
rect 46258 286516 71766 286518
rect 74014 286516 76392 288880
rect 37838 285654 76392 286516
rect 37838 285646 66654 285654
rect 68900 285646 76392 285654
rect 108656 288894 133862 289860
rect 108656 288892 127376 288894
rect 108656 286528 113446 288892
rect 115694 286530 127376 288892
rect 129624 286530 133862 288894
rect 115694 286528 133862 286530
rect 108656 285646 133862 286528
rect 190322 288856 217042 289860
rect 190322 288854 210538 288856
rect 190322 286490 196608 288854
rect 198856 286492 210538 288854
rect 212786 286492 217042 288856
rect 198856 286490 217042 286492
rect 190322 285646 217042 286490
rect 273502 288872 343072 289860
rect 273502 288870 307820 288872
rect 273502 288868 293904 288870
rect 273502 286504 279974 288868
rect 282222 286506 293904 288868
rect 296152 286508 307820 288870
rect 310068 288870 343072 288872
rect 310068 288868 335584 288870
rect 310068 286508 321654 288868
rect 296152 286506 321654 286508
rect 282222 286504 321654 286506
rect 323902 288774 335584 288868
rect 323902 286504 329570 288774
rect 273502 286424 329570 286504
rect 332102 286506 335584 288774
rect 337832 286506 343072 288870
rect 332102 286424 343072 286506
rect 273502 285646 343072 286424
rect 370800 288862 395502 289860
rect 370800 288860 390956 288862
rect 370800 286496 377040 288860
rect 379288 286498 390956 288860
rect 393204 286498 395502 288862
rect 379288 286496 395502 286498
rect 370800 285646 395502 286496
rect 62628 277636 66654 285646
rect 118248 285516 123358 285646
rect 202180 285516 207110 285646
rect 283526 285516 288608 285646
rect 380680 285586 385756 285646
rect 118248 277636 122274 285516
rect 202180 277636 206206 285516
rect 283526 277636 287552 285516
rect 380680 277636 384706 285586
rect 38122 276658 76392 277636
rect 38122 276656 58210 276658
rect 38122 274292 44294 276656
rect 46542 274294 58210 276656
rect 60458 276656 76392 276658
rect 60458 274294 72050 276656
rect 46542 274292 72050 274294
rect 74298 274292 76392 276656
rect 38122 273430 76392 274292
rect 38122 273422 66654 273430
rect 69184 273422 76392 273430
rect 108656 276670 133862 277636
rect 108656 276668 127660 276670
rect 108656 274304 113730 276668
rect 115978 274306 127660 276668
rect 129908 274306 133862 276670
rect 115978 274304 133862 274306
rect 108656 273422 133862 274304
rect 190322 276632 217042 277636
rect 190322 276630 210822 276632
rect 190322 274266 196892 276630
rect 199140 274268 210822 276630
rect 213070 274268 217042 276632
rect 199140 274266 217042 274268
rect 190322 273422 217042 274266
rect 273502 276648 343072 277636
rect 273502 276646 308104 276648
rect 273502 276644 294188 276646
rect 273502 274280 280258 276644
rect 282506 274282 294188 276644
rect 296436 274284 308104 276646
rect 310352 276646 343072 276648
rect 310352 276644 335868 276646
rect 310352 274284 321938 276644
rect 296436 274282 321938 274284
rect 282506 274280 321938 274282
rect 324186 276394 335868 276644
rect 324186 274280 329570 276394
rect 273502 274044 329570 274280
rect 332102 274282 335868 276394
rect 338116 274282 343072 276646
rect 332102 274044 343072 274282
rect 273502 273422 343072 274044
rect 370800 276638 395502 277636
rect 370800 276636 391240 276638
rect 370800 274272 377324 276636
rect 379572 274274 391240 276636
rect 393488 274274 395502 276638
rect 379572 274272 395502 274274
rect 370800 273422 395502 274272
rect 62628 261888 66654 273422
rect 118248 273292 123642 273422
rect 202180 273292 207394 273422
rect 283526 273292 288892 273422
rect 380680 273362 386040 273422
rect 118248 261888 122274 273292
rect 202180 261888 206206 273292
rect 283526 261888 287552 273292
rect 380680 261888 384706 273362
rect 37702 260924 400336 261888
rect 37702 260922 141156 260924
rect 37702 260920 127240 260922
rect 37702 260912 113310 260920
rect 37702 260910 99476 260912
rect 37702 260908 57790 260910
rect 37702 258544 43874 260908
rect 46122 258546 57790 260908
rect 60038 260908 85560 260910
rect 60038 258546 71630 260908
rect 46122 258544 71630 258546
rect 73878 258546 85560 260908
rect 87808 258548 99476 260910
rect 101724 258556 113310 260912
rect 115558 258558 127240 260920
rect 129488 258560 141156 260922
rect 143404 260922 182836 260924
rect 143404 260920 168920 260922
rect 143404 258560 154990 260920
rect 129488 258558 154990 258560
rect 115558 258556 154990 258558
rect 157238 258558 168920 260920
rect 171168 258560 182836 260922
rect 185084 260900 400336 260924
rect 185084 260898 307684 260900
rect 185084 260896 293768 260898
rect 185084 260888 279838 260896
rect 185084 260886 266004 260888
rect 185084 260884 224318 260886
rect 185084 260882 210402 260884
rect 185084 258560 196472 260882
rect 171168 258558 196472 258560
rect 157238 258556 196472 258558
rect 101724 258548 196472 258556
rect 87808 258546 196472 258548
rect 73878 258544 196472 258546
rect 37702 258518 196472 258544
rect 198720 258520 210402 260882
rect 212650 258522 224318 260884
rect 226566 260884 252088 260886
rect 226566 258522 238158 260884
rect 212650 258520 238158 258522
rect 240406 258522 252088 260884
rect 254336 258524 266004 260886
rect 268252 258532 279838 260888
rect 282086 258534 293768 260896
rect 296016 258536 307684 260898
rect 309932 260898 349364 260900
rect 309932 260896 335448 260898
rect 309932 258536 321518 260896
rect 296016 258534 321518 258536
rect 282086 258532 321518 258534
rect 323766 258534 335448 260896
rect 337696 258536 349364 260898
rect 351612 260890 400336 260900
rect 351612 260888 390820 260890
rect 351612 260886 376904 260888
rect 351612 258536 362974 260886
rect 337696 258534 362974 258536
rect 323766 258532 362974 258534
rect 268252 258524 362974 258532
rect 254336 258522 362974 258524
rect 365222 258524 376904 260886
rect 379152 258526 390820 260888
rect 393068 258526 400336 260890
rect 379152 258524 400336 258526
rect 365222 258522 400336 258524
rect 240406 258520 400336 258522
rect 198720 258518 400336 258520
rect 37702 257682 400336 258518
rect 37702 257674 66654 257682
rect 68764 257674 400336 257682
rect 62628 243046 66654 257674
rect 118248 257544 123222 257674
rect 202180 257544 206974 257674
rect 283526 257544 288472 257674
rect 380680 257614 385620 257674
rect 118248 243046 122274 257544
rect 202180 239256 206206 257544
rect 283526 239256 287552 257544
rect 380680 243370 384706 257614
rect 189818 238252 215530 239256
rect 189818 238250 209436 238252
rect 189818 235886 195506 238250
rect 197754 235888 209436 238250
rect 211684 235888 215530 238252
rect 197754 235886 215530 235888
rect 189818 235042 215530 235886
rect 276024 238268 342908 239256
rect 276024 238266 306718 238268
rect 276024 238264 292802 238266
rect 276024 235900 278872 238264
rect 281120 235902 292802 238264
rect 295050 235904 306718 238266
rect 308966 238266 342908 238268
rect 308966 238264 334482 238266
rect 308966 235904 320552 238264
rect 295050 235902 320552 235904
rect 281120 235900 320552 235902
rect 322800 238186 334482 238264
rect 322800 235900 329586 238186
rect 276024 235836 329586 235900
rect 332118 235902 334482 238186
rect 336730 235902 342908 238266
rect 332118 235836 342908 235902
rect 276024 235042 342908 235836
rect 202180 233278 206206 235042
rect 283526 234140 287552 235042
rect 202210 223352 206008 233278
rect 283708 223352 287506 234140
rect 189818 222348 215530 223352
rect 189818 222346 209846 222348
rect 189818 219982 195916 222346
rect 198164 219984 209846 222346
rect 212094 219984 215530 222348
rect 198164 219982 215530 219984
rect 189818 219138 215530 219982
rect 276024 222364 342908 223352
rect 276024 222362 307128 222364
rect 276024 222360 293212 222362
rect 276024 219996 279282 222360
rect 281530 219998 293212 222360
rect 295460 220000 307128 222362
rect 309376 222362 342908 222364
rect 309376 222360 334892 222362
rect 309376 220000 320962 222360
rect 295460 219998 320962 220000
rect 281530 219996 320962 219998
rect 323210 222332 334892 222360
rect 323210 219996 329804 222332
rect 276024 219982 329804 219996
rect 332336 219998 334892 222332
rect 337140 219998 342908 222362
rect 332336 219982 342908 219998
rect 276024 219138 342908 219982
rect 202210 206900 206008 219138
rect 283708 206900 287506 219138
rect 189818 205896 215530 206900
rect 189818 205894 209846 205896
rect 189818 203530 195916 205894
rect 198164 203532 209846 205894
rect 212094 203532 215530 205896
rect 198164 203530 215530 203532
rect 189818 202686 215530 203530
rect 276024 205928 342908 206900
rect 276024 205912 330006 205928
rect 276024 205910 307128 205912
rect 276024 205908 293212 205910
rect 276024 203544 279282 205908
rect 281530 203546 293212 205908
rect 295460 203548 307128 205910
rect 309376 205908 330006 205912
rect 309376 203548 320962 205908
rect 295460 203546 320962 203548
rect 281530 203544 320962 203546
rect 323210 203578 330006 205908
rect 332538 205910 342908 205928
rect 332538 203578 334892 205910
rect 323210 203546 334892 203578
rect 337140 203546 342908 205910
rect 323210 203544 342908 203546
rect 276024 202686 342908 203544
rect 202210 192092 206008 202686
rect 283708 192092 287506 202686
rect 189818 191088 215530 192092
rect 189818 191086 209436 191088
rect 189818 188722 195506 191086
rect 197754 188724 209436 191086
rect 211684 188724 215530 191088
rect 197754 188722 215530 188724
rect 189818 187878 215530 188722
rect 276024 191104 342908 192092
rect 276024 191102 306718 191104
rect 276024 191100 292802 191102
rect 276024 188736 278872 191100
rect 281120 188738 292802 191100
rect 295050 188740 306718 191102
rect 308966 191102 342908 191104
rect 308966 191100 334482 191102
rect 308966 188740 320552 191100
rect 295050 188738 320552 188740
rect 281120 188736 320552 188738
rect 322800 190930 334482 191100
rect 322800 188736 329932 190930
rect 276024 188580 329932 188736
rect 332464 188738 334482 190930
rect 336730 188738 342908 191102
rect 332464 188580 342908 188738
rect 276024 187878 342908 188580
rect 202210 177832 206008 187878
rect 283708 177832 287506 187878
rect 188908 176844 342908 177832
rect 188908 176842 306170 176844
rect 188908 176840 292254 176842
rect 188908 176832 278324 176840
rect 188908 176830 264490 176832
rect 188908 176828 222804 176830
rect 188908 176826 208888 176828
rect 188908 174462 194958 176826
rect 197206 174464 208888 176826
rect 211136 174466 222804 176828
rect 225052 176828 250574 176830
rect 225052 174466 236644 176828
rect 211136 174464 236644 174466
rect 238892 174466 250574 176828
rect 252822 174468 264490 176830
rect 266738 174476 278324 176832
rect 280572 174478 292254 176840
rect 294502 174480 306170 176842
rect 308418 176842 342908 176844
rect 308418 176840 333934 176842
rect 308418 174480 320004 176840
rect 294502 174478 320004 174480
rect 280572 174476 320004 174478
rect 322252 176758 333934 176840
rect 322252 174476 329894 176758
rect 266738 174468 329894 174476
rect 252822 174466 329894 174468
rect 238892 174464 329894 174466
rect 197206 174462 329894 174464
rect 188908 174408 329894 174462
rect 332426 174478 333934 176758
rect 336182 174478 342908 176842
rect 332426 174408 342908 174478
rect 188908 173618 342908 174408
rect 202210 165006 206008 173618
rect 283708 165006 287506 173618
rect 188908 164018 342908 165006
rect 188908 164016 306386 164018
rect 188908 164014 292470 164016
rect 188908 164006 278540 164014
rect 188908 164004 264706 164006
rect 188908 164002 223020 164004
rect 188908 164000 209104 164002
rect 188908 161636 195174 164000
rect 197422 161638 209104 164000
rect 211352 161640 223020 164002
rect 225268 164002 250790 164004
rect 225268 161640 236860 164002
rect 211352 161638 236860 161640
rect 239108 161640 250790 164002
rect 253038 161642 264706 164004
rect 266954 161650 278540 164006
rect 280788 161652 292470 164014
rect 294718 161654 306386 164016
rect 308634 164016 342908 164018
rect 308634 164014 334150 164016
rect 308634 161654 320220 164014
rect 294718 161652 320220 161654
rect 280788 161650 320220 161652
rect 322468 163954 334150 164014
rect 322468 161650 329820 163954
rect 266954 161642 329820 161650
rect 253038 161640 329820 161642
rect 239108 161638 329820 161640
rect 197422 161636 329820 161638
rect 188908 161604 329820 161636
rect 332352 161652 334150 163954
rect 336398 161652 342908 164016
rect 332352 161604 342908 161652
rect 188908 160792 342908 161604
rect 201534 143168 205714 160792
rect 62118 142646 67398 143110
rect 121840 142646 121988 143168
rect 201534 142646 205740 143168
rect 283276 142646 287456 160792
rect 36468 142548 117660 142646
rect 121840 142548 352454 142646
rect 36468 141682 352454 142548
rect 36468 141680 139590 141682
rect 36468 141678 125674 141680
rect 36468 141670 111744 141678
rect 36468 141668 97910 141670
rect 36468 141666 56224 141668
rect 36468 139302 42308 141666
rect 44556 139304 56224 141666
rect 58472 141666 83994 141668
rect 58472 139304 70064 141666
rect 44556 139302 70064 139304
rect 72312 139304 83994 141666
rect 86242 139306 97910 141668
rect 100158 139314 111744 141670
rect 113992 139316 125674 141678
rect 127922 139318 139590 141680
rect 141838 141680 181270 141682
rect 141838 141678 167354 141680
rect 141838 139318 153424 141678
rect 127922 139316 153424 139318
rect 113992 139314 153424 139316
rect 155672 139316 167354 141678
rect 169602 139318 181270 141680
rect 183518 141658 352454 141682
rect 183518 141656 306118 141658
rect 183518 141654 292202 141656
rect 183518 141646 278272 141654
rect 183518 141644 264438 141646
rect 183518 141642 222752 141644
rect 183518 141640 208836 141642
rect 183518 139318 194906 141640
rect 169602 139316 194906 139318
rect 155672 139314 194906 139316
rect 100158 139306 194906 139314
rect 86242 139304 194906 139306
rect 72312 139302 194906 139304
rect 36468 139276 194906 139302
rect 197154 139278 208836 141640
rect 211084 139280 222752 141642
rect 225000 141642 250522 141644
rect 225000 139280 236592 141642
rect 211084 139278 236592 139280
rect 238840 139280 250522 141642
rect 252770 139282 264438 141644
rect 266686 139290 278272 141646
rect 280520 139292 292202 141654
rect 294450 139294 306118 141656
rect 308366 141656 347798 141658
rect 308366 141654 333882 141656
rect 308366 139294 319952 141654
rect 294450 139292 319952 139294
rect 280520 139290 319952 139292
rect 322200 141454 333882 141654
rect 322200 139290 329784 141454
rect 266686 139282 329784 139290
rect 252770 139280 329784 139282
rect 238840 139278 329784 139280
rect 197154 139276 329784 139278
rect 36468 139104 329784 139276
rect 332316 139292 333882 141454
rect 336130 139294 347798 141656
rect 350046 139294 352454 141658
rect 336130 139292 352454 139294
rect 332316 139104 352454 139292
rect 36468 138432 352454 139104
rect 62118 130166 67398 138432
rect 117660 130166 122808 138432
rect 201534 130166 205714 138432
rect 283276 130166 287456 138432
rect 36398 129464 352454 130166
rect 36398 129202 329636 129464
rect 36398 129200 139520 129202
rect 36398 129198 125604 129200
rect 36398 129190 111674 129198
rect 36398 129188 97840 129190
rect 36398 129186 56154 129188
rect 36398 126822 42238 129186
rect 44486 126824 56154 129186
rect 58402 129186 83924 129188
rect 58402 126824 69994 129186
rect 44486 126822 69994 126824
rect 72242 126824 83924 129186
rect 86172 126826 97840 129188
rect 100088 126834 111674 129190
rect 113922 126836 125604 129198
rect 127852 126838 139520 129200
rect 141768 129200 181200 129202
rect 141768 129198 167284 129200
rect 141768 126838 153354 129198
rect 127852 126836 153354 126838
rect 113922 126834 153354 126836
rect 155602 126836 167284 129198
rect 169532 126838 181200 129200
rect 183448 129178 329636 129202
rect 183448 129176 306048 129178
rect 183448 129174 292132 129176
rect 183448 129166 278202 129174
rect 183448 129164 264368 129166
rect 183448 129162 222682 129164
rect 183448 129160 208766 129162
rect 183448 126838 194836 129160
rect 169532 126836 194836 126838
rect 155602 126834 194836 126836
rect 100088 126826 194836 126834
rect 86172 126824 194836 126826
rect 72242 126822 194836 126824
rect 36398 126796 194836 126822
rect 197084 126798 208766 129160
rect 211014 126800 222682 129162
rect 224930 129162 250452 129164
rect 224930 126800 236522 129162
rect 211014 126798 236522 126800
rect 238770 126800 250452 129162
rect 252700 126802 264368 129164
rect 266616 126810 278202 129166
rect 280450 126812 292132 129174
rect 294380 126814 306048 129176
rect 308296 129174 329636 129178
rect 308296 126814 319882 129174
rect 294380 126812 319882 126814
rect 280450 126810 319882 126812
rect 322130 127114 329636 129174
rect 332168 129178 352454 129464
rect 332168 129176 347728 129178
rect 332168 127114 333812 129176
rect 322130 126812 333812 127114
rect 336060 126814 347728 129176
rect 349976 126814 352454 129178
rect 336060 126812 352454 126814
rect 322130 126810 352454 126812
rect 266616 126802 352454 126810
rect 252700 126800 352454 126802
rect 238770 126798 352454 126800
rect 197084 126796 352454 126798
rect 36398 125952 352454 126796
rect 62118 118732 67398 125952
rect 117660 118732 122808 125952
rect 201534 118732 205714 125952
rect 283276 118732 287456 125952
rect 36328 117808 352454 118732
rect 36328 117768 329710 117808
rect 36328 117766 139450 117768
rect 36328 117764 125534 117766
rect 36328 117756 111604 117764
rect 36328 117754 97770 117756
rect 36328 117752 56084 117754
rect 36328 115388 42168 117752
rect 44416 115390 56084 117752
rect 58332 117752 83854 117754
rect 58332 115390 69924 117752
rect 44416 115388 69924 115390
rect 72172 115390 83854 117752
rect 86102 115392 97770 117754
rect 100018 115400 111604 117756
rect 113852 115402 125534 117764
rect 127782 115404 139450 117766
rect 141698 117766 181130 117768
rect 141698 117764 167214 117766
rect 141698 115404 153284 117764
rect 127782 115402 153284 115404
rect 113852 115400 153284 115402
rect 155532 115402 167214 117764
rect 169462 115404 181130 117766
rect 183378 117744 329710 117768
rect 183378 117742 305978 117744
rect 183378 117740 292062 117742
rect 183378 117732 278132 117740
rect 183378 117730 264298 117732
rect 183378 117728 222612 117730
rect 183378 117726 208696 117728
rect 183378 115404 194766 117726
rect 169462 115402 194766 115404
rect 155532 115400 194766 115402
rect 100018 115392 194766 115400
rect 86102 115390 194766 115392
rect 72172 115388 194766 115390
rect 36328 115362 194766 115388
rect 197014 115364 208696 117726
rect 210944 115366 222612 117728
rect 224860 117728 250382 117730
rect 224860 115366 236452 117728
rect 210944 115364 236452 115366
rect 238700 115366 250382 117728
rect 252630 115368 264298 117730
rect 266546 115376 278132 117732
rect 280380 115378 292062 117740
rect 294310 115380 305978 117742
rect 308226 117740 329710 117744
rect 308226 115380 319812 117740
rect 294310 115378 319812 115380
rect 280380 115376 319812 115378
rect 322060 115458 329710 117740
rect 332242 117744 352454 117808
rect 332242 117742 347658 117744
rect 332242 115458 333742 117742
rect 322060 115378 333742 115458
rect 335990 115380 347658 117742
rect 349906 115380 352454 117744
rect 335990 115378 352454 115380
rect 322060 115376 352454 115378
rect 266546 115368 352454 115376
rect 252630 115366 352454 115368
rect 238700 115364 352454 115366
rect 197014 115362 352454 115364
rect 36328 114518 352454 115362
rect 62118 106322 67398 114518
rect 117660 106322 122808 114518
rect 201534 106322 205714 114518
rect 283276 106844 287456 114518
rect 283162 106322 287456 106844
rect 36190 105634 352454 106322
rect 36190 105358 329858 105634
rect 36190 105356 139312 105358
rect 36190 105354 125396 105356
rect 36190 105346 111466 105354
rect 36190 105344 97632 105346
rect 36190 105342 55946 105344
rect 36190 102978 42030 105342
rect 44278 102980 55946 105342
rect 58194 105342 83716 105344
rect 58194 102980 69786 105342
rect 44278 102978 69786 102980
rect 72034 102980 83716 105342
rect 85964 102982 97632 105344
rect 99880 102990 111466 105346
rect 113714 102992 125396 105354
rect 127644 102994 139312 105356
rect 141560 105356 180992 105358
rect 141560 105354 167076 105356
rect 141560 102994 153146 105354
rect 127644 102992 153146 102994
rect 113714 102990 153146 102992
rect 155394 102992 167076 105354
rect 169324 102994 180992 105356
rect 183240 105334 329858 105358
rect 183240 105332 305840 105334
rect 183240 105330 291924 105332
rect 183240 105322 277994 105330
rect 183240 105320 264160 105322
rect 183240 105318 222474 105320
rect 183240 105316 208558 105318
rect 183240 102994 194628 105316
rect 169324 102992 194628 102994
rect 155394 102990 194628 102992
rect 99880 102982 194628 102990
rect 85964 102980 194628 102982
rect 72034 102978 194628 102980
rect 36190 102952 194628 102978
rect 196876 102954 208558 105316
rect 210806 102956 222474 105318
rect 224722 105318 250244 105320
rect 224722 102956 236314 105318
rect 210806 102954 236314 102956
rect 238562 102956 250244 105318
rect 252492 102958 264160 105320
rect 266408 102966 277994 105322
rect 280242 102968 291924 105330
rect 294172 102970 305840 105332
rect 308088 105330 329858 105334
rect 308088 102970 319674 105330
rect 294172 102968 319674 102970
rect 280242 102966 319674 102968
rect 321922 103284 329858 105330
rect 332390 105334 352454 105634
rect 332390 105332 347520 105334
rect 332390 103284 333604 105332
rect 321922 102968 333604 103284
rect 335852 102970 347520 105332
rect 349768 102970 352454 105334
rect 335852 102968 352454 102970
rect 321922 102966 352454 102968
rect 266408 102958 352454 102966
rect 252492 102956 352454 102958
rect 238562 102954 352454 102956
rect 196876 102952 352454 102954
rect 36190 102108 352454 102952
rect 200624 94788 205196 102108
rect 282436 90606 287008 102108
rect 270820 89918 352454 90606
rect 270820 89618 329282 89918
rect 270820 89616 305264 89618
rect 270820 89614 291348 89616
rect 270820 87250 277418 89614
rect 279666 87252 291348 89614
rect 293596 87254 305264 89616
rect 307512 89614 329282 89618
rect 307512 87254 319098 89614
rect 293596 87252 319098 87254
rect 279666 87250 319098 87252
rect 321346 87568 329282 89614
rect 331814 89618 352454 89918
rect 331814 89616 346944 89618
rect 331814 87568 333028 89616
rect 321346 87252 333028 87568
rect 335276 87254 346944 89616
rect 349192 87254 352454 89618
rect 335276 87252 352454 87254
rect 321346 87250 352454 87252
rect 270820 86392 352454 87250
rect 282436 78018 287008 86392
rect 270820 77330 352454 78018
rect 270820 77030 329282 77330
rect 270820 77028 305264 77030
rect 270820 77026 291348 77028
rect 270820 74662 277418 77026
rect 279666 74664 291348 77026
rect 293596 74666 305264 77028
rect 307512 77026 329282 77030
rect 307512 74666 319098 77026
rect 293596 74664 319098 74666
rect 279666 74662 319098 74664
rect 321346 74980 329282 77026
rect 331814 77030 352454 77330
rect 331814 77028 346944 77030
rect 331814 74980 333028 77028
rect 321346 74664 333028 74980
rect 335276 74666 346944 77028
rect 349192 74666 352454 77030
rect 335276 74664 352454 74666
rect 321346 74662 352454 74664
rect 270820 73804 352454 74662
rect 282436 65430 287008 73804
rect 270820 64742 352454 65430
rect 270820 64442 329282 64742
rect 270820 64440 305264 64442
rect 270820 64438 291348 64440
rect 270820 62074 277418 64438
rect 279666 62076 291348 64438
rect 293596 62078 305264 64440
rect 307512 64438 329282 64442
rect 307512 62078 319098 64438
rect 293596 62076 319098 62078
rect 279666 62074 319098 62076
rect 321346 62392 329282 64438
rect 331814 64442 352454 64742
rect 331814 64440 346944 64442
rect 331814 62392 333028 64440
rect 321346 62076 333028 62392
rect 335276 62078 346944 64440
rect 349192 62078 352454 64442
rect 335276 62076 352454 62078
rect 321346 62074 352454 62076
rect 270820 61216 352454 62074
rect 282436 47510 287008 61216
<< viali >>
rect 329000 677548 331532 679898
rect 328962 663376 331494 665726
rect 329000 650632 331532 652982
rect 328962 636460 331494 638810
rect 329012 622110 331544 624460
rect 328974 607938 331506 610288
rect 329190 589392 331722 591742
rect 329152 575220 331684 577570
rect 329078 562416 331610 564766
rect 329292 544576 331824 546926
rect 329254 530404 331786 532754
rect 329180 517600 331712 519950
rect 329354 496068 331886 498418
rect 329316 481896 331848 484246
rect 329242 469092 331774 471442
rect 329602 455536 332134 457886
rect 329562 443812 332094 446162
rect 329642 419686 332174 422036
rect 329604 405514 332136 407864
rect 329530 392710 332062 395060
rect 329616 383900 332148 386250
rect 329578 369728 332110 372078
rect 329504 356924 332036 359274
rect 329224 345074 331756 347424
rect 329150 332270 331682 334620
rect 329682 317748 332214 320098
rect 329644 308068 332176 310418
rect 329606 297528 332138 299878
rect 329570 286424 332102 288774
rect 329570 274044 332102 276394
rect 329586 235836 332118 238186
rect 329804 219982 332336 222332
rect 330006 203578 332538 205928
rect 329932 188580 332464 190930
rect 329894 174408 332426 176758
rect 329820 161604 332352 163954
rect 329784 139104 332316 141454
rect 329636 127114 332168 129464
rect 329710 115458 332242 117808
rect 329858 103284 332390 105634
rect 329282 87568 331814 89918
rect 329282 74980 331814 77330
rect 329282 62392 331814 64742
<< metal1 >>
rect 328854 679898 331696 680064
rect 328854 677548 329000 679898
rect 331532 677548 331696 679898
rect 328854 677366 331696 677548
rect 328816 665726 331658 665892
rect 328816 663376 328962 665726
rect 331494 663376 331658 665726
rect 328816 663194 331658 663376
rect 328854 652982 331696 653148
rect 328854 650632 329000 652982
rect 331532 650632 331696 652982
rect 328854 650450 331696 650632
rect 328816 638810 331658 638976
rect 328816 636460 328962 638810
rect 331494 636460 331658 638810
rect 328816 636278 331658 636460
rect 328866 624460 331708 624626
rect 328866 622110 329012 624460
rect 331544 622110 331708 624460
rect 328866 621928 331708 622110
rect 328828 610288 331670 610454
rect 328828 607938 328974 610288
rect 331506 607938 331670 610288
rect 328828 607756 331670 607938
rect 329044 591742 331886 591908
rect 329044 589392 329190 591742
rect 331722 589392 331886 591742
rect 329044 589210 331886 589392
rect 329006 577570 331848 577736
rect 329006 575220 329152 577570
rect 331684 575220 331848 577570
rect 329006 575038 331848 575220
rect 328932 564766 331774 564932
rect 328932 562416 329078 564766
rect 331610 562416 331774 564766
rect 328932 562234 331774 562416
rect 329146 546926 331988 547092
rect 329146 544576 329292 546926
rect 331824 544576 331988 546926
rect 329146 544394 331988 544576
rect 329108 532754 331950 532920
rect 329108 530404 329254 532754
rect 331786 530404 331950 532754
rect 329108 530222 331950 530404
rect 329034 519950 331876 520116
rect 329034 517600 329180 519950
rect 331712 517600 331876 519950
rect 329034 517418 331876 517600
rect 329208 498418 332050 498584
rect 329208 496068 329354 498418
rect 331886 496068 332050 498418
rect 329208 495886 332050 496068
rect 329170 484246 332012 484412
rect 329170 481896 329316 484246
rect 331848 481896 332012 484246
rect 329170 481714 332012 481896
rect 329096 471442 331938 471608
rect 329096 469092 329242 471442
rect 331774 469092 331938 471442
rect 329096 468910 331938 469092
rect 329456 457886 332298 458052
rect 329456 455536 329602 457886
rect 332134 455536 332298 457886
rect 329456 455354 332298 455536
rect 329416 446162 332258 446328
rect 329416 443812 329562 446162
rect 332094 443812 332258 446162
rect 329416 443630 332258 443812
rect 329496 422036 332338 422202
rect 329496 419686 329642 422036
rect 332174 419686 332338 422036
rect 329496 419504 332338 419686
rect 329458 407864 332300 408030
rect 329458 405514 329604 407864
rect 332136 405514 332300 407864
rect 329458 405332 332300 405514
rect 329384 395060 332226 395226
rect 329384 392710 329530 395060
rect 332062 392710 332226 395060
rect 329384 392528 332226 392710
rect 329470 386250 332312 386416
rect 329470 383900 329616 386250
rect 332148 383900 332312 386250
rect 329470 383718 332312 383900
rect 329432 372078 332274 372244
rect 329432 369728 329578 372078
rect 332110 369728 332274 372078
rect 329432 369546 332274 369728
rect 329358 359274 332200 359440
rect 329358 356924 329504 359274
rect 332036 356924 332200 359274
rect 329358 356742 332200 356924
rect 329078 347424 331920 347590
rect 329078 345074 329224 347424
rect 331756 345074 331920 347424
rect 329078 344892 331920 345074
rect 329004 334620 331846 334786
rect 329004 332270 329150 334620
rect 331682 332270 331846 334620
rect 329004 332088 331846 332270
rect 329536 320098 332378 320264
rect 329536 317748 329682 320098
rect 332214 317748 332378 320098
rect 329536 317566 332378 317748
rect 329498 310418 332340 310584
rect 329498 308068 329644 310418
rect 332176 308068 332340 310418
rect 329498 307886 332340 308068
rect 329460 299878 332302 300044
rect 329460 297528 329606 299878
rect 332138 297528 332302 299878
rect 329460 297346 332302 297528
rect 329424 288774 332266 288940
rect 329424 286424 329570 288774
rect 332102 286424 332266 288774
rect 329424 286242 332266 286424
rect 329424 276394 332266 276560
rect 329424 274044 329570 276394
rect 332102 274044 332266 276394
rect 329424 273862 332266 274044
rect 329440 238186 332282 238352
rect 329440 235836 329586 238186
rect 332118 235836 332282 238186
rect 329440 235654 332282 235836
rect 329658 222332 332500 222498
rect 329658 219982 329804 222332
rect 332336 219982 332500 222332
rect 329658 219800 332500 219982
rect 329860 205928 332702 206094
rect 329860 203578 330006 205928
rect 332538 203578 332702 205928
rect 329860 203396 332702 203578
rect 329786 190930 332628 191096
rect 329786 188580 329932 190930
rect 332464 188580 332628 190930
rect 329786 188398 332628 188580
rect 329748 176758 332590 176924
rect 329748 174408 329894 176758
rect 332426 174408 332590 176758
rect 329748 174226 332590 174408
rect 329674 163954 332516 164120
rect 329674 161604 329820 163954
rect 332352 161604 332516 163954
rect 329674 161422 332516 161604
rect 329638 141454 332480 141620
rect 329638 139104 329784 141454
rect 332316 139104 332480 141454
rect 329638 138922 332480 139104
rect 329490 129464 332332 129630
rect 329490 127114 329636 129464
rect 332168 127114 332332 129464
rect 329490 126932 332332 127114
rect 329564 117808 332406 117974
rect 329564 115458 329710 117808
rect 332242 115458 332406 117808
rect 329564 115276 332406 115458
rect 329712 105634 332554 105800
rect 329712 103284 329858 105634
rect 332390 103284 332554 105634
rect 329712 103102 332554 103284
rect 329136 89918 331978 90084
rect 329136 87568 329282 89918
rect 331814 87568 331978 89918
rect 329136 87386 331978 87568
rect 329136 77330 331978 77496
rect 329136 74980 329282 77330
rect 331814 74980 331978 77330
rect 329136 74798 331978 74980
rect 329136 64742 331978 64908
rect 329136 62392 329282 64742
rect 331814 62392 331978 64742
rect 329136 62210 331978 62392
<< via1 >>
rect 329000 677548 331532 679898
rect 328962 663376 331494 665726
rect 329000 650632 331532 652982
rect 328962 636460 331494 638810
rect 329012 622110 331544 624460
rect 328974 607938 331506 610288
rect 329190 589392 331722 591742
rect 329152 575220 331684 577570
rect 329078 562416 331610 564766
rect 329292 544576 331824 546926
rect 329254 530404 331786 532754
rect 329180 517600 331712 519950
rect 329354 496068 331886 498418
rect 329316 481896 331848 484246
rect 329242 469092 331774 471442
rect 329602 455536 332134 457886
rect 329562 443812 332094 446162
rect 329642 419686 332174 422036
rect 329604 405514 332136 407864
rect 329530 392710 332062 395060
rect 329616 383900 332148 386250
rect 329578 369728 332110 372078
rect 329504 356924 332036 359274
rect 329224 345074 331756 347424
rect 329150 332270 331682 334620
rect 329682 317748 332214 320098
rect 329644 308068 332176 310418
rect 329606 297528 332138 299878
rect 329570 286424 332102 288774
rect 329570 274044 332102 276394
rect 329586 235836 332118 238186
rect 329804 219982 332336 222332
rect 330006 203578 332538 205928
rect 329932 188580 332464 190930
rect 329894 174408 332426 176758
rect 329820 161604 332352 163954
rect 329784 139104 332316 141454
rect 329636 127114 332168 129464
rect 329710 115458 332242 117808
rect 329858 103284 332390 105634
rect 329282 87568 331814 89918
rect 329282 74980 331814 77330
rect 329282 62392 331814 64742
<< metal2 >>
rect 328854 679898 331696 680064
rect 328854 677548 329000 679898
rect 331532 677548 331696 679898
rect 328854 677366 331696 677548
rect 328816 665726 331658 665892
rect 328816 663376 328962 665726
rect 331494 663376 331658 665726
rect 328816 663194 331658 663376
rect 328854 652982 331696 653148
rect 328854 650632 329000 652982
rect 331532 650632 331696 652982
rect 328854 650450 331696 650632
rect 328816 638810 331658 638976
rect 328816 636460 328962 638810
rect 331494 636460 331658 638810
rect 328816 636278 331658 636460
rect 328866 624460 331708 624626
rect 328866 622110 329012 624460
rect 331544 622110 331708 624460
rect 328866 621928 331708 622110
rect 328828 610288 331670 610454
rect 328828 607938 328974 610288
rect 331506 607938 331670 610288
rect 328828 607756 331670 607938
rect 329044 591742 331886 591908
rect 329044 589392 329190 591742
rect 331722 589392 331886 591742
rect 329044 589210 331886 589392
rect 329006 577570 331848 577736
rect 329006 575220 329152 577570
rect 331684 575220 331848 577570
rect 329006 575038 331848 575220
rect 328932 564766 331774 564932
rect 328932 562416 329078 564766
rect 331610 562416 331774 564766
rect 328932 562234 331774 562416
rect 329146 546926 331988 547092
rect 329146 544576 329292 546926
rect 331824 544576 331988 546926
rect 329146 544394 331988 544576
rect 329108 532754 331950 532920
rect 329108 530404 329254 532754
rect 331786 530404 331950 532754
rect 329108 530222 331950 530404
rect 329034 519950 331876 520116
rect 329034 517600 329180 519950
rect 331712 517600 331876 519950
rect 329034 517418 331876 517600
rect 329208 498418 332050 498584
rect 329208 496068 329354 498418
rect 331886 496068 332050 498418
rect 329208 495886 332050 496068
rect 329170 484246 332012 484412
rect 329170 481896 329316 484246
rect 331848 481896 332012 484246
rect 329170 481714 332012 481896
rect 329096 471442 331938 471608
rect 329096 469092 329242 471442
rect 331774 469092 331938 471442
rect 329096 468910 331938 469092
rect 329456 457886 332298 458052
rect 329456 455536 329602 457886
rect 332134 455536 332298 457886
rect 329456 455354 332298 455536
rect 329416 446162 332258 446328
rect 329416 443812 329562 446162
rect 332094 443812 332258 446162
rect 329416 443630 332258 443812
rect 329496 422036 332338 422202
rect 329496 419686 329642 422036
rect 332174 419686 332338 422036
rect 329496 419504 332338 419686
rect 329458 407864 332300 408030
rect 329458 405514 329604 407864
rect 332136 405514 332300 407864
rect 329458 405332 332300 405514
rect 329384 395060 332226 395226
rect 329384 392710 329530 395060
rect 332062 392710 332226 395060
rect 329384 392528 332226 392710
rect 329470 386250 332312 386416
rect 329470 383900 329616 386250
rect 332148 383900 332312 386250
rect 329470 383718 332312 383900
rect 329432 372078 332274 372244
rect 329432 369728 329578 372078
rect 332110 369728 332274 372078
rect 329432 369546 332274 369728
rect 329358 359274 332200 359440
rect 329358 356924 329504 359274
rect 332036 356924 332200 359274
rect 329358 356742 332200 356924
rect 329078 347424 331920 347590
rect 329078 345074 329224 347424
rect 331756 345074 331920 347424
rect 329078 344892 331920 345074
rect 329004 334620 331846 334786
rect 329004 332270 329150 334620
rect 331682 332270 331846 334620
rect 329004 332088 331846 332270
rect 329536 320098 332378 320264
rect 329536 317748 329682 320098
rect 332214 317748 332378 320098
rect 329536 317566 332378 317748
rect 329498 310418 332340 310584
rect 329498 308068 329644 310418
rect 332176 308068 332340 310418
rect 329498 307886 332340 308068
rect 329460 299878 332302 300044
rect 329460 297528 329606 299878
rect 332138 297528 332302 299878
rect 329460 297346 332302 297528
rect 329424 288774 332266 288940
rect 329424 286424 329570 288774
rect 332102 286424 332266 288774
rect 329424 286242 332266 286424
rect 329424 276394 332266 276560
rect 329424 274044 329570 276394
rect 332102 274044 332266 276394
rect 329424 273862 332266 274044
rect 329440 238186 332282 238352
rect 329440 235836 329586 238186
rect 332118 235836 332282 238186
rect 329440 235654 332282 235836
rect 329658 222332 332500 222498
rect 329658 219982 329804 222332
rect 332336 219982 332500 222332
rect 329658 219800 332500 219982
rect 329860 205928 332702 206094
rect 329860 203578 330006 205928
rect 332538 203578 332702 205928
rect 329860 203396 332702 203578
rect 329786 190930 332628 191096
rect 329786 188580 329932 190930
rect 332464 188580 332628 190930
rect 329786 188398 332628 188580
rect 329748 176758 332590 176924
rect 329748 174408 329894 176758
rect 332426 174408 332590 176758
rect 329748 174226 332590 174408
rect 329674 163954 332516 164120
rect 329674 161604 329820 163954
rect 332352 161604 332516 163954
rect 329674 161422 332516 161604
rect 329638 141454 332480 141620
rect 329638 139104 329784 141454
rect 332316 139104 332480 141454
rect 329638 138922 332480 139104
rect 329490 129464 332332 129630
rect 329490 127114 329636 129464
rect 332168 127114 332332 129464
rect 329490 126932 332332 127114
rect 329564 117808 332406 117974
rect 329564 115458 329710 117808
rect 332242 115458 332406 117808
rect 329564 115276 332406 115458
rect 329712 105634 332554 105800
rect 329712 103284 329858 105634
rect 332390 103284 332554 105634
rect 329712 103102 332554 103284
rect 329136 89918 331978 90084
rect 329136 87568 329282 89918
rect 331814 87568 331978 89918
rect 329136 87386 331978 87568
rect 329136 77330 331978 77496
rect 329136 74980 329282 77330
rect 331814 74980 331978 77330
rect 329136 74798 331978 74980
rect 329136 64742 331978 64908
rect 329136 62392 329282 64742
rect 331814 62392 331978 64742
rect 329136 62210 331978 62392
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 329000 677548 331532 679898
rect 328962 663376 331494 665726
rect 329000 650632 331532 652982
rect 328962 636460 331494 638810
rect 329012 622110 331544 624460
rect 328974 607938 331506 610288
rect 329190 589392 331722 591742
rect 329152 575220 331684 577570
rect 329078 562416 331610 564766
rect 329292 544576 331824 546926
rect 329254 530404 331786 532754
rect 329180 517600 331712 519950
rect 329354 496068 331886 498418
rect 329316 481896 331848 484246
rect 329242 469092 331774 471442
rect 329602 455536 332134 457886
rect 329562 443812 332094 446162
rect 329642 419686 332174 422036
rect 329604 405514 332136 407864
rect 329530 392710 332062 395060
rect 329616 383900 332148 386250
rect 329578 369728 332110 372078
rect 329504 356924 332036 359274
rect 329224 345074 331756 347424
rect 329150 332270 331682 334620
rect 329682 317748 332214 320098
rect 329644 308068 332176 310418
rect 329606 297528 332138 299878
rect 329570 286424 332102 288774
rect 329570 274044 332102 276394
rect 329586 235836 332118 238186
rect 329804 219982 332336 222332
rect 330006 203578 332538 205928
rect 329932 188580 332464 190930
rect 329894 174408 332426 176758
rect 329820 161604 332352 163954
rect 329784 139104 332316 141454
rect 329636 127114 332168 129464
rect 329710 115458 332242 117808
rect 329858 103284 332390 105634
rect 329282 87568 331814 89918
rect 329282 74980 331814 77330
rect 329282 62392 331814 64742
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 16752 698466 20824 702300
rect 68662 698466 72734 702300
rect 120678 698676 124750 702300
rect 165926 698488 169998 702300
rect 176336 698416 180408 702300
rect 217628 698310 221700 702300
rect 228108 698310 232180 702300
rect 319336 698382 323408 702300
rect 329748 698310 333820 702300
rect 413780 698622 417852 702300
rect 465732 698778 469804 702300
rect 510880 698640 514952 702340
rect 520902 698606 524974 702340
rect 566594 702300 571594 704800
rect 567176 698412 571248 702300
rect -800 684728 1700 685242
rect -800 680942 9812 684728
rect 582300 682418 584800 682984
rect -800 680242 1700 680942
rect 328854 679898 331696 680064
rect 328854 677548 329000 679898
rect 331532 677548 331696 679898
rect 574234 678344 584800 682418
rect 582300 677984 584800 678344
rect 328854 677366 331696 677548
rect 328816 665726 331658 665892
rect 328816 663376 328962 665726
rect 331494 663376 331658 665726
rect 328816 663194 331658 663376
rect 328854 652982 331696 653148
rect 328854 650632 329000 652982
rect 331532 650632 331696 652982
rect 328854 650450 331696 650632
rect -800 648098 1660 648642
rect -800 644312 9952 648098
rect -800 643842 1660 644312
rect 582340 644184 584800 644584
rect 574030 640110 584800 644184
rect 582340 639784 584800 640110
rect 328816 638810 331658 638976
rect -800 638250 1660 638642
rect -800 634464 9812 638250
rect 328816 636460 328962 638810
rect 331494 636460 331658 638810
rect 328816 636278 331658 636460
rect -800 633842 1660 634464
rect 582340 634254 584800 634584
rect 574228 630180 584800 634254
rect 582340 629784 584800 630180
rect 328866 624460 331708 624626
rect 328866 622110 329012 624460
rect 331544 622110 331708 624460
rect 328866 621928 331708 622110
rect 328828 610288 331670 610454
rect 328828 607938 328974 610288
rect 331506 607938 331670 610288
rect 328828 607756 331670 607938
rect 329044 591742 331886 591908
rect 329044 589392 329190 591742
rect 331722 589392 331886 591742
rect 583520 589472 584800 589584
rect 329044 589210 331886 589392
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 575062 584856 583716 585090
rect 575062 584744 584800 584856
rect 575062 584534 583716 584744
rect 575046 583674 583700 583954
rect 575046 583562 584800 583674
rect 575046 583398 583700 583562
rect 329006 577570 331848 577736
rect 329006 575220 329152 577570
rect 331684 575220 331848 577570
rect 329006 575038 331848 575220
rect 328932 564766 331774 564932
rect -800 563786 1660 564242
rect -800 560000 9882 563786
rect 328932 562416 329078 564766
rect 331610 562416 331774 564766
rect 328932 562234 331774 562416
rect -800 559442 1660 560000
rect 546570 554848 574574 554950
rect 582340 554848 584800 555362
rect -800 553726 1660 554242
rect 546570 553978 584800 554848
rect -800 549940 9812 553726
rect 546570 551694 547626 553978
rect 550246 551694 584800 553978
rect 546570 551062 584800 551694
rect 546570 551006 574574 551062
rect 582340 550562 584800 551062
rect -800 549442 1660 549940
rect 329146 546926 331988 547092
rect 329146 544576 329292 546926
rect 331824 544576 331988 546926
rect 582340 544860 584800 545362
rect 329146 544394 331988 544576
rect 573994 541074 584800 544860
rect 582340 540562 584800 541074
rect 329108 532754 331950 532920
rect 329108 530404 329254 532754
rect 331786 530404 331950 532754
rect 329108 530222 331950 530404
rect 329034 519950 331876 520116
rect 329034 517600 329180 519950
rect 331712 517600 331876 519950
rect 329034 517418 331876 517600
rect 352 511642 3128 511836
rect -800 511530 3128 511642
rect 352 511326 3128 511530
rect 380 510460 3156 510672
rect -800 510348 3156 510460
rect 380 510162 3156 510348
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 329208 498418 332050 498584
rect 329208 496068 329354 498418
rect 331886 496068 332050 498418
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 329208 495886 332050 496068
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 329170 484246 332012 484412
rect 329170 481896 329316 484246
rect 331848 481896 332012 484246
rect 329170 481714 332012 481896
rect 329096 471442 331938 471608
rect 329096 469092 329242 471442
rect 331774 469092 331938 471442
rect 329096 468910 331938 469092
rect 306 468420 3082 468584
rect -800 468308 3082 468420
rect 306 468074 3082 468308
rect 352 467238 3128 467468
rect -800 467126 3128 467238
rect 352 466958 3128 467126
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 329456 457886 332298 458052
rect 329456 455536 329602 457886
rect 332134 455536 332298 457886
rect 583520 455628 584800 455740
rect 329456 455354 332298 455536
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 329416 446162 332258 446328
rect 329416 443812 329562 446162
rect 332094 443812 332258 446162
rect 329416 443630 332258 443812
rect 342 425198 3118 425454
rect -800 425086 3118 425198
rect 342 424944 3118 425086
rect 350 424016 3126 424224
rect -800 423904 3126 424016
rect 350 423714 3126 423904
rect -800 422722 480 422834
rect 329496 422036 332338 422202
rect -800 421540 480 421652
rect -800 420358 480 420470
rect 329496 419686 329642 422036
rect 332174 419686 332338 422036
rect 329496 419504 332338 419686
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 329458 407864 332300 408030
rect 329458 405514 329604 407864
rect 332136 405514 332300 407864
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 329458 405332 332300 405514
rect 583520 405296 584800 405408
rect 329384 395060 332226 395226
rect 329384 392710 329530 395060
rect 332062 392710 332226 395060
rect 329384 392528 332226 392710
rect 329470 386250 332312 386416
rect 329470 383900 329616 386250
rect 332148 383900 332312 386250
rect 329470 383718 332312 383900
rect 370 381976 3146 382194
rect -800 381864 3146 381976
rect 370 381684 3146 381864
rect 408 380794 3184 381050
rect -800 380682 3184 380794
rect 408 380540 3184 380682
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 329432 372078 332274 372244
rect 329432 369728 329578 372078
rect 332110 369728 332274 372078
rect 329432 369546 332274 369728
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 329358 359274 332200 359440
rect 329358 356924 329504 359274
rect 332036 356924 332200 359274
rect 583520 358874 584800 358986
rect 329358 356742 332200 356924
rect 329078 347424 331920 347590
rect 329078 345074 329224 347424
rect 331756 345074 331920 347424
rect 329078 344892 331920 345074
rect 362 338754 3138 339018
rect -800 338642 3138 338754
rect 362 338508 3138 338642
rect 398 337572 3174 337772
rect -800 337460 3174 337572
rect 398 337262 3174 337460
rect -800 336278 480 336390
rect -800 335096 480 335208
rect 329004 334620 331846 334786
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 329004 332270 329150 334620
rect 331682 332270 331846 334620
rect 329004 332088 331846 332270
rect 329536 320098 332378 320264
rect 329536 317748 329682 320098
rect 332214 317748 332378 320098
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 329536 317566 332378 317748
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect 329498 310418 332340 310584
rect 329498 308068 329644 310418
rect 332176 308068 332340 310418
rect 329498 307886 332340 308068
rect 329460 299878 332302 300044
rect 329460 297528 329606 299878
rect 332138 297528 332302 299878
rect 329460 297346 332302 297528
rect 380 295532 3156 295794
rect -800 295420 3156 295532
rect 380 295284 3156 295420
rect 436 294350 3212 294640
rect -800 294238 3212 294350
rect 436 294130 3212 294238
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 329424 288774 332266 288940
rect 329424 286424 329570 288774
rect 332102 286424 332266 288774
rect 329424 286242 332266 286424
rect 329424 276394 332266 276560
rect 329424 274044 329570 276394
rect 332102 274044 332266 276394
rect 583520 275140 584800 275252
rect 329424 273862 332266 274044
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect 390 252510 3166 252784
rect -800 252398 3166 252510
rect 390 252274 3166 252398
rect 408 251328 3184 251648
rect -800 251216 3184 251328
rect 408 251138 3184 251216
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 329440 238186 332282 238352
rect 329440 235836 329586 238186
rect 332118 235836 332282 238186
rect 329440 235654 332282 235836
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 329658 222332 332500 222498
rect 329658 219982 329804 222332
rect 332336 219982 332500 222332
rect 329658 219800 332500 219982
rect -800 219064 1660 219688
rect -800 215278 9832 219064
rect -800 214888 1660 215278
rect -800 209150 1660 209688
rect -800 205364 9832 209150
rect 329860 205928 332702 206094
rect -800 204888 1660 205364
rect 329860 203578 330006 205928
rect 332538 203578 332702 205928
rect 329860 203396 332702 203578
rect 582340 191430 584800 196230
rect 329786 190930 332628 191096
rect 329786 188580 329932 190930
rect 332464 188580 332628 190930
rect 329786 188398 332628 188580
rect 582340 181430 584800 186230
rect -800 177066 1660 177688
rect -800 173280 9840 177066
rect 329748 176758 332590 176924
rect 329748 174408 329894 176758
rect 332426 174408 332590 176758
rect 329748 174226 332590 174408
rect -800 172888 1660 173280
rect -800 167178 1660 167688
rect -800 163392 9980 167178
rect 329674 163954 332516 164120
rect -800 162888 1660 163392
rect 329674 161604 329820 163954
rect 332352 161604 332516 163954
rect 329674 161422 332516 161604
rect 561626 151098 575864 151442
rect 582340 151098 584800 151630
rect 561626 150902 584800 151098
rect 561626 147496 562246 150902
rect 565960 147496 584800 150902
rect 561626 147312 584800 147496
rect 561626 147054 577510 147312
rect 561626 147032 573062 147054
rect 582340 146830 584800 147312
rect 329638 141454 332480 141620
rect 329638 139104 329784 141454
rect 332316 139104 332480 141454
rect 329638 138922 332480 139104
rect 574134 141070 577510 141090
rect 582340 141070 584800 141630
rect 574134 137968 584800 141070
rect 574190 137284 584800 137968
rect 582340 136830 584800 137284
rect 329490 129464 332332 129630
rect 329490 127114 329636 129464
rect 332168 127114 332332 129464
rect 329490 126932 332332 127114
rect 362 124888 3138 125174
rect -800 124776 3138 124888
rect 362 124664 3138 124776
rect 398 123706 3174 124002
rect -800 123594 3174 123706
rect 398 123492 3174 123594
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 329564 117808 332406 117974
rect 329564 115458 329710 117808
rect 332242 115458 332406 117808
rect 329564 115276 332406 115458
rect 329712 105634 332554 105800
rect 329712 103284 329858 105634
rect 332390 103284 332554 105634
rect 329712 103102 332554 103284
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect 329136 89918 331978 90084
rect 329136 87568 329282 89918
rect 331814 87568 331978 89918
rect 329136 87386 331978 87568
rect 390 81666 3166 82006
rect -800 81554 3166 81666
rect 390 81496 3166 81554
rect 408 80484 3184 80798
rect -800 80372 3184 80484
rect 408 80288 3184 80372
rect -800 79190 480 79302
rect -800 78008 480 78120
rect 329136 77330 331978 77496
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 329136 74980 329282 77330
rect 331814 74980 331978 77330
rect 329136 74798 331978 74980
rect 329136 64742 331978 64908
rect 329136 62392 329282 64742
rect 331814 62392 331978 64742
rect 329136 62210 331978 62392
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect 398 38444 3174 38718
rect -800 38332 3174 38444
rect 398 38208 3174 38332
rect 390 37262 3166 37492
rect -800 37150 3166 37262
rect 390 36982 3166 37150
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect 390 17022 3166 17302
rect -800 16910 3166 17022
rect 583520 16910 584800 17022
rect 390 16792 3166 16910
rect 426 15840 3202 16082
rect -800 15728 3202 15840
rect 583520 15728 584800 15840
rect 426 15572 3202 15728
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 329000 677548 331532 679898
rect 328962 663376 331494 665726
rect 329000 650632 331532 652982
rect 328962 636460 331494 638810
rect 329012 622110 331544 624460
rect 328974 607938 331506 610288
rect 329190 589392 331722 591742
rect 329152 575220 331684 577570
rect 329078 562416 331610 564766
rect 547626 551694 550246 553978
rect 329292 544576 331824 546926
rect 329254 530404 331786 532754
rect 329180 517600 331712 519950
rect 329354 496068 331886 498418
rect 329316 481896 331848 484246
rect 329242 469092 331774 471442
rect 329602 455536 332134 457886
rect 329562 443812 332094 446162
rect 329642 419686 332174 422036
rect 329604 405514 332136 407864
rect 329530 392710 332062 395060
rect 329616 383900 332148 386250
rect 329578 369728 332110 372078
rect 329504 356924 332036 359274
rect 329224 345074 331756 347424
rect 329150 332270 331682 334620
rect 329682 317748 332214 320098
rect 329644 308068 332176 310418
rect 329606 297528 332138 299878
rect 329570 286424 332102 288774
rect 329570 274044 332102 276394
rect 329586 235836 332118 238186
rect 329804 219982 332336 222332
rect 330006 203578 332538 205928
rect 329932 188580 332464 190930
rect 329894 174408 332426 176758
rect 329820 161604 332352 163954
rect 562246 147496 565960 150902
rect 329784 139104 332316 141454
rect 329636 127114 332168 129464
rect 329710 115458 332242 117808
rect 329858 103284 332390 105634
rect 329282 87568 331814 89918
rect 329282 74980 331814 77330
rect 329282 62392 331814 64742
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 165926 698488 169998 702300
rect 176336 698416 180408 702300
rect 217628 698310 221700 702300
rect 228108 698310 232180 702300
rect 319336 698382 323408 702300
rect 329748 698310 333820 702300
rect 328718 683614 333318 684348
rect 328540 682354 333318 683614
rect 327798 679898 333318 682354
rect 327798 677548 329000 679898
rect 331532 677548 333318 679898
rect 327798 674602 333318 677548
rect 327798 667938 333330 674602
rect 327582 665726 333330 667938
rect 327582 663376 328962 665726
rect 331494 663376 333330 665726
rect 327582 663094 333330 663376
rect 327578 661298 333330 663094
rect 328730 657432 333330 661298
rect 328718 656698 333330 657432
rect 328540 655438 333330 656698
rect 327798 652982 333330 655438
rect 327798 650632 329000 652982
rect 331532 650632 333330 652982
rect 327798 641022 333330 650632
rect 327582 638810 333330 641022
rect 21166 636852 22830 637056
rect 21166 602698 22844 636852
rect 327582 636460 328962 638810
rect 331494 636460 333330 638810
rect 327582 636178 333330 636460
rect 327578 634382 333330 636178
rect 328730 628176 333330 634382
rect 328552 626916 333330 628176
rect 327810 624460 333330 626916
rect 327810 622110 329012 624460
rect 331544 622110 333330 624460
rect 327810 612500 333330 622110
rect 327594 610288 333330 612500
rect 327594 607938 328974 610288
rect 331506 607938 333330 610288
rect 327594 607656 333330 607938
rect 327590 605842 333330 607656
rect 327810 605506 333330 605842
rect 18902 602608 37804 602698
rect 18902 602000 166796 602608
rect 328730 602000 333330 605506
rect 467664 602000 468934 612998
rect 482264 602000 482396 602122
rect 18902 598000 482396 602000
rect 18902 597946 166796 598000
rect 18902 597734 37804 597946
rect 328730 594198 333330 598000
rect 327988 591742 333330 594198
rect 327988 589392 329190 591742
rect 331722 589392 333330 591742
rect 327988 579782 333330 589392
rect 327772 577570 333330 579782
rect 327772 575220 329152 577570
rect 331684 575220 333330 577570
rect 327772 574938 333330 575220
rect 327768 573124 333330 574938
rect 327988 564766 333330 573124
rect 327988 562416 329078 564766
rect 331610 564032 333330 564766
rect 331610 562416 333518 564032
rect 327988 562112 333518 562416
rect 327984 560458 333518 562112
rect 328712 549382 333518 560458
rect 546990 553978 550846 554688
rect 546990 551694 547626 553978
rect 550246 551694 550846 553978
rect 546990 551096 550846 551694
rect 328090 546926 333518 549382
rect 328090 544576 329292 546926
rect 331824 545094 333518 546926
rect 331824 545048 333470 545094
rect 331824 544576 333432 545048
rect 328090 534966 333432 544576
rect 327874 532754 333432 534966
rect 327874 530404 329254 532754
rect 331786 530404 333432 532754
rect 327874 530122 333432 530404
rect 327870 528308 333432 530122
rect 24134 514000 24870 521360
rect 328090 519950 333432 528308
rect 328090 517600 329180 519950
rect 331712 519216 333432 519950
rect 331712 517600 333620 519216
rect 328090 517296 333620 517600
rect 328086 515642 333620 517296
rect 328730 514000 333620 515642
rect 533320 514000 535292 518462
rect 20000 513996 35040 514000
rect 58378 513996 125366 514000
rect 20000 513964 125366 513996
rect 141284 513964 550000 514000
rect 20000 510000 550000 513964
rect 328730 500898 333330 510000
rect 328730 500874 333580 500898
rect 328152 498418 333580 500874
rect 328152 496068 329354 498418
rect 331886 496586 333580 498418
rect 331886 496540 333532 496586
rect 331886 496068 333494 496540
rect 328152 486458 333494 496068
rect 327936 484246 333494 486458
rect 327936 481896 329316 484246
rect 331848 481896 333494 484246
rect 327936 481614 333494 481896
rect 327932 479800 333494 481614
rect 328152 471442 333494 479800
rect 328152 469092 329242 471442
rect 331774 470708 333494 471442
rect 331774 469092 333682 470708
rect 328152 468788 333682 469092
rect 328148 467134 333682 468788
rect 328730 466804 333682 467134
rect 328730 464000 333330 466804
rect 452096 464000 466120 464052
rect 139118 460000 466120 464000
rect 282314 459978 289018 460000
rect 328400 457886 333332 460000
rect 452096 459956 466120 460000
rect 328400 455536 329602 457886
rect 332134 455536 333332 457886
rect 328400 455342 333332 455536
rect 328400 453774 333434 455342
rect 328730 449552 333330 453774
rect 328360 446162 333330 449552
rect 328360 443812 329562 446162
rect 332094 443812 333330 446162
rect 328360 443618 333330 443812
rect 328360 442050 333394 443618
rect 328730 440000 333330 442050
rect 20000 439832 27174 440000
rect 84008 439832 452930 440000
rect 20000 436000 452930 439832
rect 328730 426590 333330 436000
rect 328440 424336 333330 426590
rect 328440 422036 333372 424336
rect 328440 419686 329642 422036
rect 332174 419686 333372 422036
rect 328440 419492 333372 419686
rect 328440 417678 333474 419492
rect 328440 410076 333330 417678
rect 328224 407864 333330 410076
rect 328224 405514 329604 407864
rect 332136 405514 333330 407864
rect 328224 405232 333330 405514
rect 328220 403418 333330 405232
rect 328440 395060 333330 403418
rect 328440 392710 329530 395060
rect 332062 392710 333330 395060
rect 328440 392406 333330 392710
rect 328436 389352 333330 392406
rect 328414 388550 333330 389352
rect 328414 386250 333346 388550
rect 328414 383900 329616 386250
rect 332148 383900 333346 386250
rect 328414 383706 333346 383900
rect 328414 381892 333448 383706
rect 328414 374290 333330 381892
rect 328198 372078 333330 374290
rect 328198 369728 329578 372078
rect 332110 369728 333330 372078
rect 328198 369446 333330 369728
rect 328194 367632 333330 369446
rect 328414 359274 333330 367632
rect 328414 356924 329504 359274
rect 332036 356924 333330 359274
rect 328414 356620 333330 356924
rect 328410 352716 333330 356620
rect 328730 350022 333330 352716
rect 328060 349636 333330 350022
rect 327844 347424 333330 349636
rect 327844 345074 329224 347424
rect 331756 345074 333330 347424
rect 327844 344792 333330 345074
rect 327840 342978 333330 344792
rect 21068 330134 21962 337076
rect 328060 334620 333330 342978
rect 328060 332270 329150 334620
rect 331682 332270 333330 334620
rect 328060 331966 333330 332270
rect 21068 330058 23302 330134
rect 19394 330000 24150 330058
rect 65158 330000 66540 330434
rect 125026 330000 128108 330466
rect 328056 330000 333330 331966
rect 19394 326000 552000 330000
rect 19394 325786 24150 326000
rect 328730 321652 333330 326000
rect 328296 320098 334194 321652
rect 328296 317748 329682 320098
rect 332214 317748 334194 320098
rect 328296 317288 334194 317748
rect 328296 316140 334296 317288
rect 328730 311986 333330 316140
rect 328730 310418 334764 311986
rect 328730 308068 329644 310418
rect 332176 308068 334764 310418
rect 328730 307622 334764 308068
rect 328730 306474 334866 307622
rect 328730 301466 333330 306474
rect 328730 299878 334906 301466
rect 328730 297528 329606 299878
rect 332138 297528 334906 299878
rect 328730 297102 334906 297528
rect 328730 295954 335008 297102
rect 328730 290518 333330 295954
rect 328730 288774 334764 290518
rect 328730 286424 329570 288774
rect 332102 286424 334764 288774
rect 328730 286154 334764 286424
rect 328730 285006 334866 286154
rect 328730 278294 333330 285006
rect 328730 276394 335048 278294
rect 328730 274044 329570 276394
rect 332102 274044 335048 276394
rect 328730 273930 335048 274044
rect 328730 272782 335150 273930
rect 328730 262902 333330 272782
rect 328730 258182 334628 262902
rect 328730 256376 334730 258182
rect 328730 254000 333330 256376
rect 398104 254000 427234 254030
rect 24000 253154 427234 254000
rect 24000 251940 428532 253154
rect 24000 250000 427234 251940
rect 328730 240394 333330 250000
rect 398104 249936 427234 250000
rect 328730 238186 333662 240394
rect 328730 235836 329586 238186
rect 332118 235836 333662 238186
rect 328730 235550 333662 235836
rect 328730 233736 333764 235550
rect 328730 224490 333330 233736
rect 328730 222332 334072 224490
rect 328730 219982 329804 222332
rect 332336 219982 334072 222332
rect 328730 219646 334072 219982
rect 328730 217832 334174 219646
rect 328730 208038 333330 217832
rect 328730 205928 334072 208038
rect 328730 203578 330006 205928
rect 332538 203578 334072 205928
rect 328730 203194 334072 203578
rect 328730 201380 334174 203194
rect 328730 193230 333330 201380
rect 328730 190930 333662 193230
rect 328730 188580 329932 190930
rect 332464 188580 333662 190930
rect 328730 188386 333662 188580
rect 328730 186572 333764 188386
rect 26884 151746 28684 181984
rect 328730 178970 333330 186572
rect 328514 176758 333330 178970
rect 328514 174408 329894 176758
rect 332426 174408 333330 176758
rect 328514 174126 333330 174408
rect 328510 172312 333330 174126
rect 328730 163954 333330 172312
rect 328730 161604 329820 163954
rect 332352 161604 333330 163954
rect 328730 161300 333330 161604
rect 34702 151746 36808 156612
rect 328726 151746 333432 161300
rect 14286 151604 379272 151746
rect 544358 151604 558746 151646
rect 14286 151578 558746 151604
rect 14286 150902 566372 151578
rect 14286 147496 562246 150902
rect 565960 147496 566372 150902
rect 14286 146826 566372 147496
rect 14286 146758 549092 146826
rect 557004 146816 566372 146826
rect 328726 143168 333432 146758
rect 375160 146620 549092 146758
rect 328462 141454 333432 143168
rect 328462 139104 329784 141454
rect 332316 139104 333432 141454
rect 328462 138940 333432 139104
rect 328458 138744 333432 138940
rect 328458 137816 333330 138744
rect 328730 130688 333330 137816
rect 328392 129464 333330 130688
rect 328392 127114 329636 129464
rect 332168 127114 333330 129464
rect 328392 126460 333330 127114
rect 328388 125336 333330 126460
rect 328730 119254 333330 125336
rect 328322 117808 333330 119254
rect 328322 115458 329710 117808
rect 332242 115458 333330 117808
rect 328322 115026 333330 115458
rect 328318 113902 333330 115026
rect 328730 106844 333330 113902
rect 328184 105634 333330 106844
rect 328184 103284 329858 105634
rect 332390 103284 333330 105634
rect 328184 102616 333330 103284
rect 328180 101492 333330 102616
rect 328730 91454 333330 101492
rect 328698 90952 333330 91454
rect 327608 89918 333954 90952
rect 327608 87568 329282 89918
rect 331814 87568 333954 89918
rect 327608 86900 333954 87568
rect 327604 86098 333954 86900
rect 328698 85802 333330 86098
rect 328730 78866 333330 85802
rect 328698 78364 333330 78866
rect 327608 77330 333954 78364
rect 327608 74980 329282 77330
rect 331814 74980 333954 77330
rect 327608 74312 333954 74980
rect 327604 73510 333954 74312
rect 328698 73214 333330 73510
rect 328730 66278 333330 73214
rect 328698 65776 333330 66278
rect 327608 64742 333954 65776
rect 327608 62392 329282 64742
rect 331814 62392 333954 64742
rect 327608 61724 333954 62392
rect 327604 60922 333954 61724
rect 328698 60626 333330 60922
rect 22000 55990 38348 56000
rect 52864 55990 54612 59938
rect 328730 56000 333330 60626
rect 103592 55990 199070 56000
rect 22000 55958 199070 55990
rect 208362 55958 352454 56000
rect 22000 52000 352454 55958
rect 191940 51646 215346 52000
rect 328730 48958 333330 52000
<< via4 >>
rect 547626 551694 550246 553978
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 165926 698488 169998 702300
rect 176336 698416 180408 702300
rect 217628 698310 221700 702300
rect 228108 698310 232180 702300
rect 319336 698382 323408 702300
rect 329748 698310 333820 702300
rect 20000 682000 558000 686000
rect 24260 662112 24882 682000
rect 56666 681854 58676 682000
rect 200674 681988 206622 682000
rect 281044 681932 288894 682000
rect 313172 681370 320000 682000
rect 378706 681892 386338 682000
rect 313114 674000 320000 681370
rect 313114 667938 318892 674000
rect 312956 664072 318892 667938
rect 312838 661298 318892 664072
rect 314104 657432 318786 661298
rect 314092 656698 318786 657432
rect 313914 655438 318786 656698
rect 313172 654454 318786 655438
rect 313114 647632 318786 654454
rect 473498 651952 474926 682000
rect 476044 681994 480744 682000
rect 313114 641022 318892 647632
rect 312956 637156 318892 641022
rect 312838 634382 318892 637156
rect 314104 628176 318786 634382
rect 313926 626916 318786 628176
rect 313184 625932 318786 626916
rect 313126 619110 318786 625932
rect 313126 612500 318904 619110
rect 312968 608634 318904 612500
rect 312850 605842 318904 608634
rect 313184 605506 318904 605842
rect 314104 594198 318786 605506
rect 313362 593214 318786 594198
rect 313304 586392 318786 593214
rect 313304 579782 319082 586392
rect 313146 575916 319082 579782
rect 313028 573124 319082 575916
rect 313362 572216 319082 573124
rect 313362 563090 318786 572216
rect 313244 562112 318786 563090
rect 313244 560458 318778 562112
rect 314020 555780 318778 560458
rect 511472 555824 520468 555836
rect 511472 555812 545988 555824
rect 511472 555780 550884 555812
rect 19816 553978 550884 555780
rect 19816 551694 547626 553978
rect 550246 551694 550884 553978
rect 19816 550272 550884 551694
rect 19816 550218 545988 550272
rect 19816 549956 520468 550218
rect 19816 549882 35040 549956
rect 58378 549952 520468 549956
rect 19816 549874 29458 549882
rect 58378 549874 512382 549952
rect 27312 536726 28130 549874
rect 314020 549382 318888 549874
rect 313464 548398 318888 549382
rect 313406 541576 318888 548398
rect 313406 534966 319184 541576
rect 458412 537880 462146 549874
rect 313248 531100 319184 534966
rect 313130 528308 319184 531100
rect 313464 527400 319184 528308
rect 313464 518274 318888 527400
rect 313346 517296 318888 518274
rect 313346 515642 318880 517296
rect 314104 512772 318880 515642
rect 314104 507240 318786 512772
rect 313774 500898 318848 507240
rect 313774 500874 318950 500898
rect 313526 499890 318950 500874
rect 313468 493068 318950 499890
rect 245920 490000 261942 490022
rect 313468 490000 319246 493068
rect 454318 490000 456470 490086
rect 18000 486144 456470 490000
rect 18000 486000 453686 486144
rect 33852 485518 34466 486000
rect 52314 485518 55228 486000
rect 245920 485980 261942 486000
rect 313310 482592 319246 486000
rect 313192 479800 319246 482592
rect 313526 478892 319246 479800
rect 454318 479534 456470 486144
rect 313526 469766 318950 478892
rect 454318 477172 469174 479534
rect 313408 468788 318950 469766
rect 313408 467134 318942 468788
rect 314104 466804 318942 467134
rect 314104 461276 318786 466804
rect 313774 460186 318786 461276
rect 313774 459358 318788 460186
rect 313716 454000 318890 459358
rect 139118 450000 453088 454000
rect 314104 449552 318786 450000
rect 313734 447634 318786 449552
rect 313676 442050 318850 447634
rect 314104 426590 318786 442050
rect 313814 424336 318786 426590
rect 313814 423508 318828 424336
rect 313756 410076 318930 423508
rect 313598 406210 318930 410076
rect 313480 405686 318930 406210
rect 313480 403418 318786 405686
rect 313814 393384 318786 403418
rect 313696 388550 318786 393384
rect 313696 387722 318802 388550
rect 313696 387062 318904 387722
rect 313730 374290 318904 387062
rect 313572 370424 318904 374290
rect 313454 369900 318904 370424
rect 313454 367632 318786 369900
rect 106616 363300 122898 363576
rect 19144 359160 122898 363300
rect 23398 356330 24108 359160
rect 118206 353918 122760 359160
rect 313788 357598 318786 367632
rect 313670 354000 318786 357598
rect 130354 353918 554000 354000
rect 118206 350000 554000 353918
rect 118206 349778 140834 350000
rect 313376 349636 318786 350000
rect 313218 345770 318786 349636
rect 313100 342978 318786 345770
rect 313434 332944 318786 342978
rect 313316 329970 318786 332944
rect 314104 321652 318786 329970
rect 313670 316140 319650 321652
rect 314104 311986 318786 316140
rect 314104 306474 320220 311986
rect 314104 301466 318786 306474
rect 314104 295954 320362 301466
rect 314104 290518 318786 295954
rect 314104 285006 320220 290518
rect 314104 278294 318786 285006
rect 314104 272782 320504 278294
rect 314104 270000 318786 272782
rect 396756 270000 431796 270076
rect 22000 266000 431796 270000
rect 42336 241032 44704 266000
rect 314104 262902 318786 266000
rect 396756 265968 431796 266000
rect 314104 256418 320084 262902
rect 430120 262496 430612 265968
rect 314104 256376 320080 256418
rect 42114 235962 44844 241032
rect 31480 233482 44844 235962
rect 31480 215264 32296 233482
rect 42114 233410 44844 233482
rect 314104 240394 318786 256376
rect 314104 233786 319118 240394
rect 314104 233736 319114 233786
rect 314104 224490 318786 233736
rect 314104 217882 319528 224490
rect 314104 217832 319524 217882
rect 314104 208038 318786 217832
rect 314104 201430 319528 208038
rect 314104 201380 319524 201430
rect 314104 193230 318786 201380
rect 314104 186622 319118 193230
rect 314104 186572 319114 186622
rect 314104 178970 318786 186572
rect 313888 175104 318786 178970
rect 313770 172312 318786 175104
rect 314104 162278 318786 172312
rect 313986 159536 318786 162278
rect 313986 143168 318782 159536
rect 313836 140422 318782 143168
rect 313836 139918 318786 140422
rect 313718 137816 318786 139918
rect 314104 130688 318786 137816
rect 313766 127438 318786 130688
rect 313648 125336 318786 127438
rect 314104 119254 318786 125336
rect 313696 116004 318786 119254
rect 313578 113902 318786 116004
rect 314104 106844 318786 113902
rect 313558 103594 318786 106844
rect 313440 101492 318786 103594
rect 314104 100000 318786 101492
rect 22000 96000 352454 100000
rect 45206 95926 51744 96000
rect 314104 91454 318786 96000
rect 314072 90952 318786 91454
rect 312982 87878 319410 90952
rect 312864 86098 319410 87878
rect 314072 85802 318786 86098
rect 314104 78866 318786 85802
rect 314072 78364 318786 78866
rect 312982 75290 319410 78364
rect 312864 73510 319410 75290
rect 314072 73214 318786 73510
rect 314104 66278 318786 73214
rect 314072 65776 318786 66278
rect 312982 62702 319410 65776
rect 312864 60922 319410 62702
rect 314072 60626 318786 60922
rect 314104 48958 318786 60626
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use pll_full_buffered2  pll_full_buffered2_0
timestamp 1647885998
transform 1 0 31278 0 1 174612
box -3258 0 88322 40874
use filter_buffered  filter_buffered_0
timestamp 1647885941
transform 1 0 46104 0 1 59356
box -2 0 89610 28900
use DIGITAL_BUFFER_v1  DIGITAL_BUFFER_v1_0
timestamp 1647886866
transform 1 0 409398 0 1 90248
box -940 -1820 87350 1165
use ashish  ashish_0
timestamp 1647888148
transform 1 0 406076 0 1 64768
box -2100 -2540 8350 2594
use div_pd_buffered  div_pd_buffered_0
timestamp 1647885998
transform 1 0 23112 0 1 341826
box -1894 -6452 88296 14680
use divider_buffered  divider_buffered_0
timestamp 1647885998
transform 1 0 429804 0 1 252392
box -1492 -3136 88296 10326
use cp_buffered  cp_buffered_0
timestamp 1647885941
transform 1 0 27122 0 1 525962
box -2796 -7196 88288 10904
use pd_buffered  pd_buffered_0
timestamp 1647885998
transform 1 0 27206 0 1 454596
box -1894 -6512 88296 8906
use ro_divider_buffered  ro_divider_buffered_0
timestamp 1647885998
transform 1 0 471678 0 1 468106
box -5944 -21716 87550 24552
use pll_full_buffered1  pll_full_buffered1_1
timestamp 1647885998
transform 1 0 23954 0 1 630304
box -2122 0 88318 31910
use ro_complete_buffered  ro_complete_buffered_0
timestamp 1647885998
transform 1 0 474094 0 1 631512
box -5924 -21716 87550 20544
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
