magic
tech sky130A
timestamp 1641017053
<< nwell >>
rect 150 303 280 310
rect 2210 303 2345 340
rect 4150 303 4285 340
rect 6400 303 6535 340
rect 9305 303 9440 340
rect 11250 303 11385 340
rect 12945 303 13080 340
rect 15130 303 15265 340
rect 17310 303 17445 340
rect 19495 303 19630 340
rect 20705 303 20840 340
rect 150 55 21181 303
rect -60 -905 30735 -545
<< nmos >>
rect 231 -120 246 -70
rect 356 -120 371 -70
rect 416 -120 431 -70
rect 476 -120 491 -70
rect 536 -120 551 -70
rect 661 -120 676 -70
rect 721 -120 736 -70
rect 781 -120 796 -70
rect 841 -120 856 -70
rect 906 -120 921 -70
rect 966 -120 981 -70
rect 1026 -120 1041 -70
rect 1086 -120 1101 -70
rect 1146 -120 1161 -70
rect 1206 -120 1221 -70
rect 1266 -120 1281 -70
rect 1326 -120 1341 -70
rect 1391 -120 1406 -70
rect 1451 -120 1466 -70
rect 1511 -120 1526 -70
rect 1571 -120 1586 -70
rect 1696 -120 1711 -70
rect 1756 -120 1771 -70
rect 1816 -120 1831 -70
rect 1876 -120 1891 -70
rect 1941 -120 1956 -70
rect 2001 -120 2016 -70
rect 2061 -120 2076 -70
rect 2121 -120 2136 -70
rect 2181 -120 2196 -70
rect 2241 -120 2256 -70
rect 2301 -120 2316 -70
rect 2361 -120 2376 -70
rect 2426 -120 2441 -70
rect 2486 -120 2501 -70
rect 2546 -120 2561 -70
rect 2606 -120 2621 -70
rect 2666 -120 2681 -70
rect 2726 -120 2741 -70
rect 2786 -120 2801 -70
rect 2846 -120 2861 -70
rect 2911 -120 2926 -70
rect 2971 -120 2986 -70
rect 3031 -120 3046 -70
rect 3091 -120 3106 -70
rect 3151 -120 3166 -70
rect 3211 -120 3226 -70
rect 3271 -120 3286 -70
rect 3331 -120 3346 -70
rect 3396 -120 3411 -70
rect 3456 -120 3471 -70
rect 3516 -120 3531 -70
rect 3576 -120 3591 -70
rect 3636 -120 3651 -70
rect 3696 -120 3711 -70
rect 3756 -120 3771 -70
rect 3816 -120 3831 -70
rect 3881 -120 3896 -70
rect 3941 -120 3956 -70
rect 4001 -120 4016 -70
rect 4061 -120 4076 -70
rect 4121 -120 4136 -70
rect 4181 -120 4196 -70
rect 4241 -120 4256 -70
rect 4301 -120 4316 -70
rect 4366 -120 4381 -70
rect 4426 -120 4441 -70
rect 4486 -120 4501 -70
rect 4546 -120 4561 -70
rect 4606 -120 4621 -70
rect 4666 -120 4681 -70
rect 4726 -120 4741 -70
rect 4786 -120 4801 -70
rect 4851 -120 4866 -70
rect 4911 -120 4926 -70
rect 4971 -120 4986 -70
rect 5031 -120 5046 -70
rect 5091 -120 5106 -70
rect 5151 -120 5166 -70
rect 5211 -120 5226 -70
rect 5271 -120 5286 -70
rect 5336 -120 5351 -70
rect 5396 -120 5411 -70
rect 5456 -120 5471 -70
rect 5516 -120 5531 -70
rect 5641 -120 5656 -70
rect 5701 -120 5716 -70
rect 5761 -120 5776 -70
rect 5821 -120 5836 -70
rect 5886 -120 5901 -70
rect 5946 -120 5961 -70
rect 6006 -120 6021 -70
rect 6066 -120 6081 -70
rect 6126 -120 6141 -70
rect 6186 -120 6201 -70
rect 6246 -120 6261 -70
rect 6306 -120 6321 -70
rect 6371 -120 6386 -70
rect 6431 -120 6446 -70
rect 6491 -120 6506 -70
rect 6551 -120 6566 -70
rect 6611 -120 6626 -70
rect 6671 -120 6686 -70
rect 6731 -120 6746 -70
rect 6791 -120 6806 -70
rect 6856 -120 6871 -70
rect 6916 -120 6931 -70
rect 6976 -120 6991 -70
rect 7036 -120 7051 -70
rect 7096 -120 7111 -70
rect 7156 -120 7171 -70
rect 7216 -120 7231 -70
rect 7276 -120 7291 -70
rect 7336 -120 7351 -70
rect 7396 -120 7411 -70
rect 7456 -120 7471 -70
rect 7516 -120 7531 -70
rect 7576 -120 7591 -70
rect 7636 -120 7651 -70
rect 7696 -120 7711 -70
rect 7756 -120 7771 -70
rect 7821 -120 7836 -70
rect 7881 -120 7896 -70
rect 7941 -120 7956 -70
rect 8001 -120 8016 -70
rect 8061 -120 8076 -70
rect 8121 -120 8136 -70
rect 8181 -120 8196 -70
rect 8241 -120 8256 -70
rect 8306 -120 8321 -70
rect 8366 -120 8381 -70
rect 8426 -120 8441 -70
rect 8486 -120 8501 -70
rect 8546 -120 8561 -70
rect 8606 -120 8621 -70
rect 8666 -120 8681 -70
rect 8726 -120 8741 -70
rect 8791 -120 8806 -70
rect 8851 -120 8866 -70
rect 8911 -120 8926 -70
rect 8971 -120 8986 -70
rect 9031 -120 9046 -70
rect 9091 -120 9106 -70
rect 9151 -120 9166 -70
rect 9211 -120 9226 -70
rect 9276 -120 9291 -70
rect 9336 -120 9351 -70
rect 9396 -120 9411 -70
rect 9456 -120 9471 -70
rect 9521 -120 9536 -70
rect 9581 -120 9596 -70
rect 9641 -120 9656 -70
rect 9701 -120 9716 -70
rect 9766 -120 9781 -70
rect 9826 -120 9841 -70
rect 9886 -120 9901 -70
rect 9946 -120 9961 -70
rect 10006 -120 10021 -70
rect 10066 -120 10081 -70
rect 10126 -120 10141 -70
rect 10186 -120 10201 -70
rect 10251 -120 10266 -70
rect 10311 -120 10326 -70
rect 10371 -120 10386 -70
rect 10431 -120 10446 -70
rect 10491 -120 10506 -70
rect 10551 -120 10566 -70
rect 10611 -120 10626 -70
rect 10671 -120 10686 -70
rect 10736 -120 10751 -70
rect 10796 -120 10811 -70
rect 10856 -120 10871 -70
rect 10916 -120 10931 -70
rect 10976 -120 10991 -70
rect 11036 -120 11051 -70
rect 11096 -120 11111 -70
rect 11156 -120 11171 -70
rect 11221 -120 11236 -70
rect 11281 -120 11296 -70
rect 11341 -120 11356 -70
rect 11401 -120 11416 -70
rect 11461 -120 11476 -70
rect 11521 -120 11536 -70
rect 11581 -120 11596 -70
rect 11641 -120 11656 -70
rect 11706 -120 11721 -70
rect 11766 -120 11781 -70
rect 11826 -120 11841 -70
rect 11886 -120 11901 -70
rect 11946 -120 11961 -70
rect 12006 -120 12021 -70
rect 12066 -120 12081 -70
rect 12126 -120 12141 -70
rect 12191 -120 12206 -70
rect 12251 -120 12266 -70
rect 12311 -120 12326 -70
rect 12371 -120 12386 -70
rect 12431 -120 12446 -70
rect 12491 -120 12506 -70
rect 12551 -120 12566 -70
rect 12611 -120 12626 -70
rect 12676 -120 12691 -70
rect 12736 -120 12751 -70
rect 12796 -120 12811 -70
rect 12856 -120 12871 -70
rect 12916 -120 12931 -70
rect 12976 -120 12991 -70
rect 13036 -120 13051 -70
rect 13096 -120 13111 -70
rect 13161 -120 13176 -70
rect 13221 -120 13236 -70
rect 13281 -120 13296 -70
rect 13341 -120 13356 -70
rect 13401 -120 13416 -70
rect 13461 -120 13476 -70
rect 13521 -120 13536 -70
rect 13581 -120 13596 -70
rect 13646 -120 13661 -70
rect 13706 -120 13721 -70
rect 13766 -120 13781 -70
rect 13826 -120 13841 -70
rect 13886 -120 13901 -70
rect 13946 -120 13961 -70
rect 14006 -120 14021 -70
rect 14066 -120 14081 -70
rect 14131 -120 14146 -70
rect 14191 -120 14206 -70
rect 14251 -120 14266 -70
rect 14311 -120 14326 -70
rect 14371 -120 14386 -70
rect 14431 -120 14446 -70
rect 14491 -120 14506 -70
rect 14551 -120 14566 -70
rect 14616 -120 14631 -70
rect 14676 -120 14691 -70
rect 14736 -120 14751 -70
rect 14796 -120 14811 -70
rect 14856 -120 14871 -70
rect 14916 -120 14931 -70
rect 14976 -120 14991 -70
rect 15036 -120 15051 -70
rect 15101 -120 15116 -70
rect 15161 -120 15176 -70
rect 15221 -120 15236 -70
rect 15281 -120 15296 -70
rect 15341 -120 15356 -70
rect 15401 -120 15416 -70
rect 15461 -120 15476 -70
rect 15521 -120 15536 -70
rect 15586 -120 15601 -70
rect 15646 -120 15661 -70
rect 15706 -120 15721 -70
rect 15766 -120 15781 -70
rect 15826 -120 15841 -70
rect 15886 -120 15901 -70
rect 15946 -120 15961 -70
rect 16006 -120 16021 -70
rect 16071 -120 16086 -70
rect 16131 -120 16146 -70
rect 16191 -120 16206 -70
rect 16251 -120 16266 -70
rect 16311 -120 16326 -70
rect 16371 -120 16386 -70
rect 16431 -120 16446 -70
rect 16491 -120 16506 -70
rect 16556 -120 16571 -70
rect 16616 -120 16631 -70
rect 16676 -120 16691 -70
rect 16736 -120 16751 -70
rect 16796 -120 16811 -70
rect 16856 -120 16871 -70
rect 16916 -120 16931 -70
rect 16976 -120 16991 -70
rect 17041 -120 17056 -70
rect 17101 -120 17116 -70
rect 17161 -120 17176 -70
rect 17221 -120 17236 -70
rect 17281 -120 17296 -70
rect 17341 -120 17356 -70
rect 17401 -120 17416 -70
rect 17461 -120 17476 -70
rect 17526 -120 17541 -70
rect 17586 -120 17601 -70
rect 17646 -120 17661 -70
rect 17706 -120 17721 -70
rect 17766 -120 17781 -70
rect 17826 -120 17841 -70
rect 17886 -120 17901 -70
rect 17946 -120 17961 -70
rect 18011 -120 18026 -70
rect 18071 -120 18086 -70
rect 18131 -120 18146 -70
rect 18191 -120 18206 -70
rect 18251 -120 18266 -70
rect 18311 -120 18326 -70
rect 18371 -120 18386 -70
rect 18431 -120 18446 -70
rect 18496 -120 18511 -70
rect 18556 -120 18571 -70
rect 18616 -120 18631 -70
rect 18676 -120 18691 -70
rect 18736 -120 18751 -70
rect 18796 -120 18811 -70
rect 18856 -120 18871 -70
rect 18916 -120 18931 -70
rect 18981 -120 18996 -70
rect 19041 -120 19056 -70
rect 19101 -120 19116 -70
rect 19161 -120 19176 -70
rect 19221 -120 19236 -70
rect 19281 -120 19296 -70
rect 19341 -120 19356 -70
rect 19401 -120 19416 -70
rect 19466 -120 19481 -70
rect 19526 -120 19541 -70
rect 19586 -120 19601 -70
rect 19646 -120 19661 -70
rect 19706 -120 19721 -70
rect 19766 -120 19781 -70
rect 19826 -120 19841 -70
rect 19886 -120 19901 -70
rect 19951 -120 19966 -70
rect 20011 -120 20026 -70
rect 20071 -120 20086 -70
rect 20131 -120 20146 -70
rect 20191 -120 20206 -70
rect 20251 -120 20266 -70
rect 20311 -120 20326 -70
rect 20371 -120 20386 -70
rect 20436 -120 20451 -70
rect 20496 -120 20511 -70
rect 20556 -120 20571 -70
rect 20616 -120 20631 -70
rect 20676 -120 20691 -70
rect 20736 -120 20751 -70
rect 20796 -120 20811 -70
rect 20856 -120 20871 -70
rect 20921 -120 20936 -70
rect 20981 -120 20996 -70
rect 21041 -120 21056 -70
rect 21101 -120 21116 -70
rect 0 -420 15 -320
rect 60 -420 75 -320
rect 120 -420 135 -320
rect 180 -420 195 -320
rect 240 -420 255 -320
rect 300 -420 315 -320
rect 360 -420 375 -320
rect 420 -420 435 -320
rect 480 -420 495 -320
rect 540 -420 555 -320
rect 600 -420 615 -320
rect 660 -420 675 -320
rect 720 -420 735 -320
rect 780 -420 795 -320
rect 840 -420 855 -320
rect 900 -420 915 -320
rect 960 -420 975 -320
rect 1020 -420 1035 -320
rect 1080 -420 1095 -320
rect 1140 -420 1155 -320
rect 1200 -420 1215 -320
rect 1260 -420 1275 -320
rect 1320 -420 1335 -320
rect 1380 -420 1395 -320
rect 1440 -420 1455 -320
rect 1500 -420 1515 -320
rect 1560 -420 1575 -320
rect 1620 -420 1635 -320
rect 1680 -420 1695 -320
rect 1740 -420 1755 -320
rect 1800 -420 1815 -320
rect 1860 -420 1875 -320
rect 1920 -420 1935 -320
rect 1980 -420 1995 -320
rect 2040 -420 2055 -320
rect 2100 -420 2115 -320
rect 2160 -420 2175 -320
rect 2220 -420 2235 -320
rect 2280 -420 2295 -320
rect 2340 -420 2355 -320
rect 2400 -420 2415 -320
rect 2460 -420 2475 -320
rect 2520 -420 2535 -320
rect 2580 -420 2595 -320
rect 2640 -420 2655 -320
rect 2700 -420 2715 -320
rect 2760 -420 2775 -320
rect 2820 -420 2835 -320
rect 2880 -420 2895 -320
rect 2940 -420 2955 -320
rect 3000 -420 3015 -320
rect 3060 -420 3075 -320
rect 3120 -420 3135 -320
rect 3180 -420 3195 -320
rect 3240 -420 3255 -320
rect 3300 -420 3315 -320
rect 3360 -420 3375 -320
rect 3420 -420 3435 -320
rect 3480 -420 3495 -320
rect 3540 -420 3555 -320
rect 3600 -420 3615 -320
rect 3660 -420 3675 -320
rect 3720 -420 3735 -320
rect 3780 -420 3795 -320
rect 3840 -420 3855 -320
rect 3900 -420 3915 -320
rect 3960 -420 3975 -320
rect 4020 -420 4035 -320
rect 4080 -420 4095 -320
rect 4140 -420 4155 -320
rect 4200 -420 4215 -320
rect 4260 -420 4275 -320
rect 4320 -420 4335 -320
rect 4380 -420 4395 -320
rect 4440 -420 4455 -320
rect 4500 -420 4515 -320
rect 4560 -420 4575 -320
rect 4620 -420 4635 -320
rect 4680 -420 4695 -320
rect 4740 -420 4755 -320
rect 4800 -420 4815 -320
rect 4860 -420 4875 -320
rect 4920 -420 4935 -320
rect 4980 -420 4995 -320
rect 5040 -420 5055 -320
rect 5100 -420 5115 -320
rect 5160 -420 5175 -320
rect 5220 -420 5235 -320
rect 5280 -420 5295 -320
rect 5340 -420 5355 -320
rect 5400 -420 5415 -320
rect 5460 -420 5475 -320
rect 5520 -420 5535 -320
rect 5580 -420 5595 -320
rect 5640 -420 5655 -320
rect 5700 -420 5715 -320
rect 5760 -420 5775 -320
rect 5820 -420 5835 -320
rect 5880 -420 5895 -320
rect 5940 -420 5955 -320
rect 6000 -420 6015 -320
rect 6060 -420 6075 -320
rect 6120 -420 6135 -320
rect 6180 -420 6195 -320
rect 6240 -420 6255 -320
rect 6300 -420 6315 -320
rect 6360 -420 6375 -320
rect 6420 -420 6435 -320
rect 6480 -420 6495 -320
rect 6540 -420 6555 -320
rect 6600 -420 6615 -320
rect 6660 -420 6675 -320
rect 6720 -420 6735 -320
rect 6780 -420 6795 -320
rect 6840 -420 6855 -320
rect 6900 -420 6915 -320
rect 6960 -420 6975 -320
rect 7020 -420 7035 -320
rect 7080 -420 7095 -320
rect 7140 -420 7155 -320
rect 7200 -420 7215 -320
rect 7260 -420 7275 -320
rect 7320 -420 7335 -320
rect 7380 -420 7395 -320
rect 7440 -420 7455 -320
rect 7500 -420 7515 -320
rect 7560 -420 7575 -320
rect 7620 -420 7635 -320
rect 7680 -420 7695 -320
rect 7740 -420 7755 -320
rect 7800 -420 7815 -320
rect 7860 -420 7875 -320
rect 7920 -420 7935 -320
rect 7980 -420 7995 -320
rect 8040 -420 8055 -320
rect 8100 -420 8115 -320
rect 8160 -420 8175 -320
rect 8220 -420 8235 -320
rect 8280 -420 8295 -320
rect 8340 -420 8355 -320
rect 8400 -420 8415 -320
rect 8460 -420 8475 -320
rect 8520 -420 8535 -320
rect 8580 -420 8595 -320
rect 8640 -420 8655 -320
rect 8700 -420 8715 -320
rect 8760 -420 8775 -320
rect 8820 -420 8835 -320
rect 8880 -420 8895 -320
rect 8940 -420 8955 -320
rect 9000 -420 9015 -320
rect 9060 -420 9075 -320
rect 9120 -420 9135 -320
rect 9180 -420 9195 -320
rect 9240 -420 9255 -320
rect 9300 -420 9315 -320
rect 9360 -420 9375 -320
rect 9420 -420 9435 -320
rect 9480 -420 9495 -320
rect 9540 -420 9555 -320
rect 9600 -420 9615 -320
rect 9660 -420 9675 -320
rect 9720 -420 9735 -320
rect 9780 -420 9795 -320
rect 9840 -420 9855 -320
rect 9900 -420 9915 -320
rect 9960 -420 9975 -320
rect 10020 -420 10035 -320
rect 10080 -420 10095 -320
rect 10140 -420 10155 -320
rect 10200 -420 10215 -320
rect 10260 -420 10275 -320
rect 10320 -420 10335 -320
rect 10380 -420 10395 -320
rect 10440 -420 10455 -320
rect 10500 -420 10515 -320
rect 10560 -420 10575 -320
rect 10620 -420 10635 -320
rect 10680 -420 10695 -320
rect 10740 -420 10755 -320
rect 10800 -420 10815 -320
rect 10860 -420 10875 -320
rect 10920 -420 10935 -320
rect 10980 -420 10995 -320
rect 11040 -420 11055 -320
rect 11100 -420 11115 -320
rect 11160 -420 11175 -320
rect 11220 -420 11235 -320
rect 11280 -420 11295 -320
rect 11340 -420 11355 -320
rect 11400 -420 11415 -320
rect 11460 -420 11475 -320
rect 11520 -420 11535 -320
rect 11580 -420 11595 -320
rect 11640 -420 11655 -320
rect 11700 -420 11715 -320
rect 11760 -420 11775 -320
rect 11820 -420 11835 -320
rect 11880 -420 11895 -320
rect 11940 -420 11955 -320
rect 12000 -420 12015 -320
rect 12060 -420 12075 -320
rect 12120 -420 12135 -320
rect 12180 -420 12195 -320
rect 12240 -420 12255 -320
rect 12300 -420 12315 -320
rect 12360 -420 12375 -320
rect 12420 -420 12435 -320
rect 12480 -420 12495 -320
rect 12540 -420 12555 -320
rect 12600 -420 12615 -320
rect 12660 -420 12675 -320
rect 12720 -420 12735 -320
rect 12780 -420 12795 -320
rect 12840 -420 12855 -320
rect 12900 -420 12915 -320
rect 12960 -420 12975 -320
rect 13020 -420 13035 -320
rect 13080 -420 13095 -320
rect 13140 -420 13155 -320
rect 13200 -420 13215 -320
rect 13260 -420 13275 -320
rect 13320 -420 13335 -320
rect 13380 -420 13395 -320
rect 13440 -420 13455 -320
rect 13500 -420 13515 -320
rect 13560 -420 13575 -320
rect 13620 -420 13635 -320
rect 13680 -420 13695 -320
rect 13740 -420 13755 -320
rect 13800 -420 13815 -320
rect 13860 -420 13875 -320
rect 13920 -420 13935 -320
rect 13980 -420 13995 -320
rect 14040 -420 14055 -320
rect 14100 -420 14115 -320
rect 14160 -420 14175 -320
rect 14220 -420 14235 -320
rect 14280 -420 14295 -320
rect 14340 -420 14355 -320
rect 14400 -420 14415 -320
rect 14460 -420 14475 -320
rect 14520 -420 14535 -320
rect 14580 -420 14595 -320
rect 14640 -420 14655 -320
rect 14700 -420 14715 -320
rect 14760 -420 14775 -320
rect 14820 -420 14835 -320
rect 14880 -420 14895 -320
rect 14940 -420 14955 -320
rect 15000 -420 15015 -320
rect 15060 -420 15075 -320
rect 15120 -420 15135 -320
rect 15180 -420 15195 -320
rect 15240 -420 15255 -320
rect 15300 -420 15315 -320
rect 15360 -420 15375 -320
rect 15420 -420 15435 -320
rect 15480 -420 15495 -320
rect 15540 -420 15555 -320
rect 15600 -420 15615 -320
rect 15660 -420 15675 -320
rect 15720 -420 15735 -320
rect 15780 -420 15795 -320
rect 15840 -420 15855 -320
rect 15900 -420 15915 -320
rect 15960 -420 15975 -320
rect 16020 -420 16035 -320
rect 16080 -420 16095 -320
rect 16140 -420 16155 -320
rect 16200 -420 16215 -320
rect 16260 -420 16275 -320
rect 16320 -420 16335 -320
rect 16380 -420 16395 -320
rect 16440 -420 16455 -320
rect 16500 -420 16515 -320
rect 16560 -420 16575 -320
rect 16620 -420 16635 -320
rect 16680 -420 16695 -320
rect 16740 -420 16755 -320
rect 16800 -420 16815 -320
rect 16860 -420 16875 -320
rect 16920 -420 16935 -320
rect 16980 -420 16995 -320
rect 17040 -420 17055 -320
rect 17100 -420 17115 -320
rect 17160 -420 17175 -320
rect 17220 -420 17235 -320
rect 17280 -420 17295 -320
rect 17340 -420 17355 -320
rect 17400 -420 17415 -320
rect 17460 -420 17475 -320
rect 17520 -420 17535 -320
rect 17580 -420 17595 -320
rect 17640 -420 17655 -320
rect 17700 -420 17715 -320
rect 17760 -420 17775 -320
rect 17820 -420 17835 -320
rect 17880 -420 17895 -320
rect 17940 -420 17955 -320
rect 18000 -420 18015 -320
rect 18060 -420 18075 -320
rect 18120 -420 18135 -320
rect 18180 -420 18195 -320
rect 18240 -420 18255 -320
rect 18300 -420 18315 -320
rect 18360 -420 18375 -320
rect 18420 -420 18435 -320
rect 18480 -420 18495 -320
rect 18540 -420 18555 -320
rect 18600 -420 18615 -320
rect 18660 -420 18675 -320
rect 18720 -420 18735 -320
rect 18780 -420 18795 -320
rect 18840 -420 18855 -320
rect 18900 -420 18915 -320
rect 18960 -420 18975 -320
rect 19020 -420 19035 -320
rect 19080 -420 19095 -320
rect 19140 -420 19155 -320
rect 19200 -420 19215 -320
rect 19260 -420 19275 -320
rect 19320 -420 19335 -320
rect 19380 -420 19395 -320
rect 19440 -420 19455 -320
rect 19500 -420 19515 -320
rect 19560 -420 19575 -320
rect 19620 -420 19635 -320
rect 19680 -420 19695 -320
rect 19740 -420 19755 -320
rect 19800 -420 19815 -320
rect 19860 -420 19875 -320
rect 19920 -420 19935 -320
rect 19980 -420 19995 -320
rect 20040 -420 20055 -320
rect 20100 -420 20115 -320
rect 20160 -420 20175 -320
rect 20220 -420 20235 -320
rect 20280 -420 20295 -320
rect 20340 -420 20355 -320
rect 20400 -420 20415 -320
rect 20460 -420 20475 -320
rect 20520 -420 20535 -320
rect 20580 -420 20595 -320
rect 20640 -420 20655 -320
rect 20700 -420 20715 -320
rect 20760 -420 20775 -320
rect 20820 -420 20835 -320
rect 20880 -420 20895 -320
rect 20940 -420 20955 -320
rect 21000 -420 21015 -320
rect 21060 -420 21075 -320
rect 21120 -420 21135 -320
rect 21180 -420 21195 -320
rect 21240 -420 21255 -320
rect 21300 -420 21315 -320
rect 21360 -420 21375 -320
rect 21420 -420 21435 -320
rect 21480 -420 21495 -320
rect 21540 -420 21555 -320
rect 21600 -420 21615 -320
rect 21660 -420 21675 -320
rect 21720 -420 21735 -320
rect 21780 -420 21795 -320
rect 21840 -420 21855 -320
rect 21900 -420 21915 -320
rect 21960 -420 21975 -320
rect 22020 -420 22035 -320
rect 22080 -420 22095 -320
rect 22140 -420 22155 -320
rect 22200 -420 22215 -320
rect 22260 -420 22275 -320
rect 22320 -420 22335 -320
rect 22380 -420 22395 -320
rect 22440 -420 22455 -320
rect 22500 -420 22515 -320
rect 22560 -420 22575 -320
rect 22620 -420 22635 -320
rect 22680 -420 22695 -320
rect 22740 -420 22755 -320
rect 22800 -420 22815 -320
rect 22860 -420 22875 -320
rect 22920 -420 22935 -320
rect 22980 -420 22995 -320
rect 23040 -420 23055 -320
rect 23100 -420 23115 -320
rect 23160 -420 23175 -320
rect 23220 -420 23235 -320
rect 23280 -420 23295 -320
rect 23340 -420 23355 -320
rect 23400 -420 23415 -320
rect 23460 -420 23475 -320
rect 23520 -420 23535 -320
rect 23580 -420 23595 -320
rect 23640 -420 23655 -320
rect 23700 -420 23715 -320
rect 23760 -420 23775 -320
rect 23820 -420 23835 -320
rect 23880 -420 23895 -320
rect 23940 -420 23955 -320
rect 24000 -420 24015 -320
rect 24060 -420 24075 -320
rect 24120 -420 24135 -320
rect 24180 -420 24195 -320
rect 24240 -420 24255 -320
rect 24300 -420 24315 -320
rect 24360 -420 24375 -320
rect 24420 -420 24435 -320
rect 24480 -420 24495 -320
rect 24540 -420 24555 -320
rect 24600 -420 24615 -320
rect 24660 -420 24675 -320
rect 24720 -420 24735 -320
rect 24780 -420 24795 -320
rect 24840 -420 24855 -320
rect 24900 -420 24915 -320
rect 24960 -420 24975 -320
rect 25020 -420 25035 -320
rect 25080 -420 25095 -320
rect 25140 -420 25155 -320
rect 25200 -420 25215 -320
rect 25260 -420 25275 -320
rect 25320 -420 25335 -320
rect 25380 -420 25395 -320
rect 25440 -420 25455 -320
rect 25500 -420 25515 -320
rect 25560 -420 25575 -320
rect 25620 -420 25635 -320
rect 25680 -420 25695 -320
rect 25740 -420 25755 -320
rect 25800 -420 25815 -320
rect 25860 -420 25875 -320
rect 25920 -420 25935 -320
rect 25980 -420 25995 -320
rect 26040 -420 26055 -320
rect 26100 -420 26115 -320
rect 26160 -420 26175 -320
rect 26220 -420 26235 -320
rect 26280 -420 26295 -320
rect 26340 -420 26355 -320
rect 26400 -420 26415 -320
rect 26460 -420 26475 -320
rect 26520 -420 26535 -320
rect 26580 -420 26595 -320
rect 26640 -420 26655 -320
rect 26700 -420 26715 -320
rect 26760 -420 26775 -320
rect 26820 -420 26835 -320
rect 26880 -420 26895 -320
rect 26940 -420 26955 -320
rect 27000 -420 27015 -320
rect 27060 -420 27075 -320
rect 27120 -420 27135 -320
rect 27180 -420 27195 -320
rect 27240 -420 27255 -320
rect 27300 -420 27315 -320
rect 27360 -420 27375 -320
rect 27420 -420 27435 -320
rect 27480 -420 27495 -320
rect 27540 -420 27555 -320
rect 27600 -420 27615 -320
rect 27660 -420 27675 -320
rect 27720 -420 27735 -320
rect 27780 -420 27795 -320
rect 27840 -420 27855 -320
rect 27900 -420 27915 -320
rect 27960 -420 27975 -320
rect 28020 -420 28035 -320
rect 28080 -420 28095 -320
rect 28140 -420 28155 -320
rect 28200 -420 28215 -320
rect 28260 -420 28275 -320
rect 28320 -420 28335 -320
rect 28380 -420 28395 -320
rect 28440 -420 28455 -320
rect 28500 -420 28515 -320
rect 28560 -420 28575 -320
rect 28620 -420 28635 -320
rect 28680 -420 28695 -320
rect 28740 -420 28755 -320
rect 28800 -420 28815 -320
rect 28860 -420 28875 -320
rect 28920 -420 28935 -320
rect 28980 -420 28995 -320
rect 29040 -420 29055 -320
rect 29100 -420 29115 -320
rect 29160 -420 29175 -320
rect 29220 -420 29235 -320
rect 29280 -420 29295 -320
rect 29340 -420 29355 -320
rect 29400 -420 29415 -320
rect 29460 -420 29475 -320
rect 29520 -420 29535 -320
rect 29580 -420 29595 -320
rect 29640 -420 29655 -320
rect 29700 -420 29715 -320
rect 29760 -420 29775 -320
rect 29820 -420 29835 -320
rect 29880 -420 29895 -320
rect 29940 -420 29955 -320
rect 30000 -420 30015 -320
rect 30060 -420 30075 -320
rect 30120 -420 30135 -320
rect 30180 -420 30195 -320
rect 30240 -420 30255 -320
rect 30300 -420 30315 -320
rect 30360 -420 30375 -320
rect 30420 -420 30435 -320
rect 30480 -420 30495 -320
rect 30540 -420 30555 -320
rect 30600 -420 30615 -320
rect 30660 -420 30675 -320
<< pmos >>
rect 231 85 246 185
rect 356 85 371 185
rect 416 85 431 185
rect 476 85 491 185
rect 536 85 551 185
rect 661 85 676 185
rect 721 85 736 185
rect 781 85 796 185
rect 841 85 856 185
rect 906 85 921 185
rect 966 85 981 185
rect 1026 85 1041 185
rect 1086 85 1101 185
rect 1146 85 1161 185
rect 1206 85 1221 185
rect 1266 85 1281 185
rect 1326 85 1341 185
rect 1391 85 1406 185
rect 1451 85 1466 185
rect 1511 85 1526 185
rect 1571 85 1586 185
rect 1696 85 1711 185
rect 1756 85 1771 185
rect 1816 85 1831 185
rect 1876 85 1891 185
rect 1941 85 1956 185
rect 2001 85 2016 185
rect 2061 85 2076 185
rect 2121 85 2136 185
rect 2181 85 2196 185
rect 2241 85 2256 185
rect 2301 85 2316 185
rect 2361 85 2376 185
rect 2426 85 2441 185
rect 2486 85 2501 185
rect 2546 85 2561 185
rect 2606 85 2621 185
rect 2666 85 2681 185
rect 2726 85 2741 185
rect 2786 85 2801 185
rect 2846 85 2861 185
rect 2911 85 2926 185
rect 2971 85 2986 185
rect 3031 85 3046 185
rect 3091 85 3106 185
rect 3151 85 3166 185
rect 3211 85 3226 185
rect 3271 85 3286 185
rect 3331 85 3346 185
rect 3396 85 3411 185
rect 3456 85 3471 185
rect 3516 85 3531 185
rect 3576 85 3591 185
rect 3636 85 3651 185
rect 3696 85 3711 185
rect 3756 85 3771 185
rect 3816 85 3831 185
rect 3881 85 3896 185
rect 3941 85 3956 185
rect 4001 85 4016 185
rect 4061 85 4076 185
rect 4121 85 4136 185
rect 4181 85 4196 185
rect 4241 85 4256 185
rect 4301 85 4316 185
rect 4366 85 4381 185
rect 4426 85 4441 185
rect 4486 85 4501 185
rect 4546 85 4561 185
rect 4606 85 4621 185
rect 4666 85 4681 185
rect 4726 85 4741 185
rect 4786 85 4801 185
rect 4851 85 4866 185
rect 4911 85 4926 185
rect 4971 85 4986 185
rect 5031 85 5046 185
rect 5091 85 5106 185
rect 5151 85 5166 185
rect 5211 85 5226 185
rect 5271 85 5286 185
rect 5336 85 5351 185
rect 5396 85 5411 185
rect 5456 85 5471 185
rect 5516 85 5531 185
rect 5641 85 5656 185
rect 5701 85 5716 185
rect 5761 85 5776 185
rect 5821 85 5836 185
rect 5886 85 5901 185
rect 5946 85 5961 185
rect 6006 85 6021 185
rect 6066 85 6081 185
rect 6126 85 6141 185
rect 6186 85 6201 185
rect 6246 85 6261 185
rect 6306 85 6321 185
rect 6371 85 6386 185
rect 6431 85 6446 185
rect 6491 85 6506 185
rect 6551 85 6566 185
rect 6611 85 6626 185
rect 6671 85 6686 185
rect 6731 85 6746 185
rect 6791 85 6806 185
rect 6856 85 6871 185
rect 6916 85 6931 185
rect 6976 85 6991 185
rect 7036 85 7051 185
rect 7096 85 7111 185
rect 7156 85 7171 185
rect 7216 85 7231 185
rect 7276 85 7291 185
rect 7336 85 7351 185
rect 7396 85 7411 185
rect 7456 85 7471 185
rect 7516 85 7531 185
rect 7576 85 7591 185
rect 7636 85 7651 185
rect 7696 85 7711 185
rect 7756 85 7771 185
rect 7821 85 7836 185
rect 7881 85 7896 185
rect 7941 85 7956 185
rect 8001 85 8016 185
rect 8061 85 8076 185
rect 8121 85 8136 185
rect 8181 85 8196 185
rect 8241 85 8256 185
rect 8306 85 8321 185
rect 8366 85 8381 185
rect 8426 85 8441 185
rect 8486 85 8501 185
rect 8546 85 8561 185
rect 8606 85 8621 185
rect 8666 85 8681 185
rect 8726 85 8741 185
rect 8791 85 8806 185
rect 8851 85 8866 185
rect 8911 85 8926 185
rect 8971 85 8986 185
rect 9031 85 9046 185
rect 9091 85 9106 185
rect 9151 85 9166 185
rect 9211 85 9226 185
rect 9276 85 9291 185
rect 9336 85 9351 185
rect 9396 85 9411 185
rect 9456 85 9471 185
rect 9521 85 9536 185
rect 9581 85 9596 185
rect 9641 85 9656 185
rect 9701 85 9716 185
rect 9766 85 9781 185
rect 9826 85 9841 185
rect 9886 85 9901 185
rect 9946 85 9961 185
rect 10006 85 10021 185
rect 10066 85 10081 185
rect 10126 85 10141 185
rect 10186 85 10201 185
rect 10251 85 10266 185
rect 10311 85 10326 185
rect 10371 85 10386 185
rect 10431 85 10446 185
rect 10491 85 10506 185
rect 10551 85 10566 185
rect 10611 85 10626 185
rect 10671 85 10686 185
rect 10736 85 10751 185
rect 10796 85 10811 185
rect 10856 85 10871 185
rect 10916 85 10931 185
rect 10976 85 10991 185
rect 11036 85 11051 185
rect 11096 85 11111 185
rect 11156 85 11171 185
rect 11221 85 11236 185
rect 11281 85 11296 185
rect 11341 85 11356 185
rect 11401 85 11416 185
rect 11461 85 11476 185
rect 11521 85 11536 185
rect 11581 85 11596 185
rect 11641 85 11656 185
rect 11706 85 11721 185
rect 11766 85 11781 185
rect 11826 85 11841 185
rect 11886 85 11901 185
rect 11946 85 11961 185
rect 12006 85 12021 185
rect 12066 85 12081 185
rect 12126 85 12141 185
rect 12191 85 12206 185
rect 12251 85 12266 185
rect 12311 85 12326 185
rect 12371 85 12386 185
rect 12431 85 12446 185
rect 12491 85 12506 185
rect 12551 85 12566 185
rect 12611 85 12626 185
rect 12676 85 12691 185
rect 12736 85 12751 185
rect 12796 85 12811 185
rect 12856 85 12871 185
rect 12916 85 12931 185
rect 12976 85 12991 185
rect 13036 85 13051 185
rect 13096 85 13111 185
rect 13161 85 13176 185
rect 13221 85 13236 185
rect 13281 85 13296 185
rect 13341 85 13356 185
rect 13401 85 13416 185
rect 13461 85 13476 185
rect 13521 85 13536 185
rect 13581 85 13596 185
rect 13646 85 13661 185
rect 13706 85 13721 185
rect 13766 85 13781 185
rect 13826 85 13841 185
rect 13886 85 13901 185
rect 13946 85 13961 185
rect 14006 85 14021 185
rect 14066 85 14081 185
rect 14131 85 14146 185
rect 14191 85 14206 185
rect 14251 85 14266 185
rect 14311 85 14326 185
rect 14371 85 14386 185
rect 14431 85 14446 185
rect 14491 85 14506 185
rect 14551 85 14566 185
rect 14616 85 14631 185
rect 14676 85 14691 185
rect 14736 85 14751 185
rect 14796 85 14811 185
rect 14856 85 14871 185
rect 14916 85 14931 185
rect 14976 85 14991 185
rect 15036 85 15051 185
rect 15101 85 15116 185
rect 15161 85 15176 185
rect 15221 85 15236 185
rect 15281 85 15296 185
rect 15341 85 15356 185
rect 15401 85 15416 185
rect 15461 85 15476 185
rect 15521 85 15536 185
rect 15586 85 15601 185
rect 15646 85 15661 185
rect 15706 85 15721 185
rect 15766 85 15781 185
rect 15826 85 15841 185
rect 15886 85 15901 185
rect 15946 85 15961 185
rect 16006 85 16021 185
rect 16071 85 16086 185
rect 16131 85 16146 185
rect 16191 85 16206 185
rect 16251 85 16266 185
rect 16311 85 16326 185
rect 16371 85 16386 185
rect 16431 85 16446 185
rect 16491 85 16506 185
rect 16556 85 16571 185
rect 16616 85 16631 185
rect 16676 85 16691 185
rect 16736 85 16751 185
rect 16796 85 16811 185
rect 16856 85 16871 185
rect 16916 85 16931 185
rect 16976 85 16991 185
rect 17041 85 17056 185
rect 17101 85 17116 185
rect 17161 85 17176 185
rect 17221 85 17236 185
rect 17281 85 17296 185
rect 17341 85 17356 185
rect 17401 85 17416 185
rect 17461 85 17476 185
rect 17526 85 17541 185
rect 17586 85 17601 185
rect 17646 85 17661 185
rect 17706 85 17721 185
rect 17766 85 17781 185
rect 17826 85 17841 185
rect 17886 85 17901 185
rect 17946 85 17961 185
rect 18011 85 18026 185
rect 18071 85 18086 185
rect 18131 85 18146 185
rect 18191 85 18206 185
rect 18251 85 18266 185
rect 18311 85 18326 185
rect 18371 85 18386 185
rect 18431 85 18446 185
rect 18496 85 18511 185
rect 18556 85 18571 185
rect 18616 85 18631 185
rect 18676 85 18691 185
rect 18736 85 18751 185
rect 18796 85 18811 185
rect 18856 85 18871 185
rect 18916 85 18931 185
rect 18981 85 18996 185
rect 19041 85 19056 185
rect 19101 85 19116 185
rect 19161 85 19176 185
rect 19221 85 19236 185
rect 19281 85 19296 185
rect 19341 85 19356 185
rect 19401 85 19416 185
rect 19466 85 19481 185
rect 19526 85 19541 185
rect 19586 85 19601 185
rect 19646 85 19661 185
rect 19706 85 19721 185
rect 19766 85 19781 185
rect 19826 85 19841 185
rect 19886 85 19901 185
rect 19951 85 19966 185
rect 20011 85 20026 185
rect 20071 85 20086 185
rect 20131 85 20146 185
rect 20191 85 20206 185
rect 20251 85 20266 185
rect 20311 85 20326 185
rect 20371 85 20386 185
rect 20436 85 20451 185
rect 20496 85 20511 185
rect 20556 85 20571 185
rect 20616 85 20631 185
rect 20676 85 20691 185
rect 20736 85 20751 185
rect 20796 85 20811 185
rect 20856 85 20871 185
rect 20921 85 20936 185
rect 20981 85 20996 185
rect 21041 85 21056 185
rect 21101 85 21116 185
rect 0 -770 15 -575
rect 60 -770 75 -575
rect 120 -770 135 -575
rect 180 -770 195 -575
rect 240 -770 255 -575
rect 300 -770 315 -575
rect 360 -770 375 -575
rect 420 -770 435 -575
rect 480 -770 495 -575
rect 540 -770 555 -575
rect 600 -770 615 -575
rect 660 -770 675 -575
rect 720 -770 735 -575
rect 780 -770 795 -575
rect 840 -770 855 -575
rect 900 -770 915 -575
rect 960 -770 975 -575
rect 1020 -770 1035 -575
rect 1080 -770 1095 -575
rect 1140 -770 1155 -575
rect 1200 -770 1215 -575
rect 1260 -770 1275 -575
rect 1320 -770 1335 -575
rect 1380 -770 1395 -575
rect 1440 -770 1455 -575
rect 1500 -770 1515 -575
rect 1560 -770 1575 -575
rect 1620 -770 1635 -575
rect 1680 -770 1695 -575
rect 1740 -770 1755 -575
rect 1800 -770 1815 -575
rect 1860 -770 1875 -575
rect 1920 -770 1935 -575
rect 1980 -770 1995 -575
rect 2040 -770 2055 -575
rect 2100 -770 2115 -575
rect 2160 -770 2175 -575
rect 2220 -770 2235 -575
rect 2280 -770 2295 -575
rect 2340 -770 2355 -575
rect 2400 -770 2415 -575
rect 2460 -770 2475 -575
rect 2520 -770 2535 -575
rect 2580 -770 2595 -575
rect 2640 -770 2655 -575
rect 2700 -770 2715 -575
rect 2760 -770 2775 -575
rect 2820 -770 2835 -575
rect 2880 -770 2895 -575
rect 2940 -770 2955 -575
rect 3000 -770 3015 -575
rect 3060 -770 3075 -575
rect 3120 -770 3135 -575
rect 3180 -770 3195 -575
rect 3240 -770 3255 -575
rect 3300 -770 3315 -575
rect 3360 -770 3375 -575
rect 3420 -770 3435 -575
rect 3480 -770 3495 -575
rect 3540 -770 3555 -575
rect 3600 -770 3615 -575
rect 3660 -770 3675 -575
rect 3720 -770 3735 -575
rect 3780 -770 3795 -575
rect 3840 -770 3855 -575
rect 3900 -770 3915 -575
rect 3960 -770 3975 -575
rect 4020 -770 4035 -575
rect 4080 -770 4095 -575
rect 4140 -770 4155 -575
rect 4200 -770 4215 -575
rect 4260 -770 4275 -575
rect 4320 -770 4335 -575
rect 4380 -770 4395 -575
rect 4440 -770 4455 -575
rect 4500 -770 4515 -575
rect 4560 -770 4575 -575
rect 4620 -770 4635 -575
rect 4680 -770 4695 -575
rect 4740 -770 4755 -575
rect 4800 -770 4815 -575
rect 4860 -770 4875 -575
rect 4920 -770 4935 -575
rect 4980 -770 4995 -575
rect 5040 -770 5055 -575
rect 5100 -770 5115 -575
rect 5160 -770 5175 -575
rect 5220 -770 5235 -575
rect 5280 -770 5295 -575
rect 5340 -770 5355 -575
rect 5400 -770 5415 -575
rect 5460 -770 5475 -575
rect 5520 -770 5535 -575
rect 5580 -770 5595 -575
rect 5640 -770 5655 -575
rect 5700 -770 5715 -575
rect 5760 -770 5775 -575
rect 5820 -770 5835 -575
rect 5880 -770 5895 -575
rect 5940 -770 5955 -575
rect 6000 -770 6015 -575
rect 6060 -770 6075 -575
rect 6120 -770 6135 -575
rect 6180 -770 6195 -575
rect 6240 -770 6255 -575
rect 6300 -770 6315 -575
rect 6360 -770 6375 -575
rect 6420 -770 6435 -575
rect 6480 -770 6495 -575
rect 6540 -770 6555 -575
rect 6600 -770 6615 -575
rect 6660 -770 6675 -575
rect 6720 -770 6735 -575
rect 6780 -770 6795 -575
rect 6840 -770 6855 -575
rect 6900 -770 6915 -575
rect 6960 -770 6975 -575
rect 7020 -770 7035 -575
rect 7080 -770 7095 -575
rect 7140 -770 7155 -575
rect 7200 -770 7215 -575
rect 7260 -770 7275 -575
rect 7320 -770 7335 -575
rect 7380 -770 7395 -575
rect 7440 -770 7455 -575
rect 7500 -770 7515 -575
rect 7560 -770 7575 -575
rect 7620 -770 7635 -575
rect 7680 -770 7695 -575
rect 7740 -770 7755 -575
rect 7800 -770 7815 -575
rect 7860 -770 7875 -575
rect 7920 -770 7935 -575
rect 7980 -770 7995 -575
rect 8040 -770 8055 -575
rect 8100 -770 8115 -575
rect 8160 -770 8175 -575
rect 8220 -770 8235 -575
rect 8280 -770 8295 -575
rect 8340 -770 8355 -575
rect 8400 -770 8415 -575
rect 8460 -770 8475 -575
rect 8520 -770 8535 -575
rect 8580 -770 8595 -575
rect 8640 -770 8655 -575
rect 8700 -770 8715 -575
rect 8760 -770 8775 -575
rect 8820 -770 8835 -575
rect 8880 -770 8895 -575
rect 8940 -770 8955 -575
rect 9000 -770 9015 -575
rect 9060 -770 9075 -575
rect 9120 -770 9135 -575
rect 9180 -770 9195 -575
rect 9240 -770 9255 -575
rect 9300 -770 9315 -575
rect 9360 -770 9375 -575
rect 9420 -770 9435 -575
rect 9480 -770 9495 -575
rect 9540 -770 9555 -575
rect 9600 -770 9615 -575
rect 9660 -770 9675 -575
rect 9720 -770 9735 -575
rect 9780 -770 9795 -575
rect 9840 -770 9855 -575
rect 9900 -770 9915 -575
rect 9960 -770 9975 -575
rect 10020 -770 10035 -575
rect 10080 -770 10095 -575
rect 10140 -770 10155 -575
rect 10200 -770 10215 -575
rect 10260 -770 10275 -575
rect 10320 -770 10335 -575
rect 10380 -770 10395 -575
rect 10440 -770 10455 -575
rect 10500 -770 10515 -575
rect 10560 -770 10575 -575
rect 10620 -770 10635 -575
rect 10680 -770 10695 -575
rect 10740 -770 10755 -575
rect 10800 -770 10815 -575
rect 10860 -770 10875 -575
rect 10920 -770 10935 -575
rect 10980 -770 10995 -575
rect 11040 -770 11055 -575
rect 11100 -770 11115 -575
rect 11160 -770 11175 -575
rect 11220 -770 11235 -575
rect 11280 -770 11295 -575
rect 11340 -770 11355 -575
rect 11400 -770 11415 -575
rect 11460 -770 11475 -575
rect 11520 -770 11535 -575
rect 11580 -770 11595 -575
rect 11640 -770 11655 -575
rect 11700 -770 11715 -575
rect 11760 -770 11775 -575
rect 11820 -770 11835 -575
rect 11880 -770 11895 -575
rect 11940 -770 11955 -575
rect 12000 -770 12015 -575
rect 12060 -770 12075 -575
rect 12120 -770 12135 -575
rect 12180 -770 12195 -575
rect 12240 -770 12255 -575
rect 12300 -770 12315 -575
rect 12360 -770 12375 -575
rect 12420 -770 12435 -575
rect 12480 -770 12495 -575
rect 12540 -770 12555 -575
rect 12600 -770 12615 -575
rect 12660 -770 12675 -575
rect 12720 -770 12735 -575
rect 12780 -770 12795 -575
rect 12840 -770 12855 -575
rect 12900 -770 12915 -575
rect 12960 -770 12975 -575
rect 13020 -770 13035 -575
rect 13080 -770 13095 -575
rect 13140 -770 13155 -575
rect 13200 -770 13215 -575
rect 13260 -770 13275 -575
rect 13320 -770 13335 -575
rect 13380 -770 13395 -575
rect 13440 -770 13455 -575
rect 13500 -770 13515 -575
rect 13560 -770 13575 -575
rect 13620 -770 13635 -575
rect 13680 -770 13695 -575
rect 13740 -770 13755 -575
rect 13800 -770 13815 -575
rect 13860 -770 13875 -575
rect 13920 -770 13935 -575
rect 13980 -770 13995 -575
rect 14040 -770 14055 -575
rect 14100 -770 14115 -575
rect 14160 -770 14175 -575
rect 14220 -770 14235 -575
rect 14280 -770 14295 -575
rect 14340 -770 14355 -575
rect 14400 -770 14415 -575
rect 14460 -770 14475 -575
rect 14520 -770 14535 -575
rect 14580 -770 14595 -575
rect 14640 -770 14655 -575
rect 14700 -770 14715 -575
rect 14760 -770 14775 -575
rect 14820 -770 14835 -575
rect 14880 -770 14895 -575
rect 14940 -770 14955 -575
rect 15000 -770 15015 -575
rect 15060 -770 15075 -575
rect 15120 -770 15135 -575
rect 15180 -770 15195 -575
rect 15240 -770 15255 -575
rect 15300 -770 15315 -575
rect 15360 -770 15375 -575
rect 15420 -770 15435 -575
rect 15480 -770 15495 -575
rect 15540 -770 15555 -575
rect 15600 -770 15615 -575
rect 15660 -770 15675 -575
rect 15720 -770 15735 -575
rect 15780 -770 15795 -575
rect 15840 -770 15855 -575
rect 15900 -770 15915 -575
rect 15960 -770 15975 -575
rect 16020 -770 16035 -575
rect 16080 -770 16095 -575
rect 16140 -770 16155 -575
rect 16200 -770 16215 -575
rect 16260 -770 16275 -575
rect 16320 -770 16335 -575
rect 16380 -770 16395 -575
rect 16440 -770 16455 -575
rect 16500 -770 16515 -575
rect 16560 -770 16575 -575
rect 16620 -770 16635 -575
rect 16680 -770 16695 -575
rect 16740 -770 16755 -575
rect 16800 -770 16815 -575
rect 16860 -770 16875 -575
rect 16920 -770 16935 -575
rect 16980 -770 16995 -575
rect 17040 -770 17055 -575
rect 17100 -770 17115 -575
rect 17160 -770 17175 -575
rect 17220 -770 17235 -575
rect 17280 -770 17295 -575
rect 17340 -770 17355 -575
rect 17400 -770 17415 -575
rect 17460 -770 17475 -575
rect 17520 -770 17535 -575
rect 17580 -770 17595 -575
rect 17640 -770 17655 -575
rect 17700 -770 17715 -575
rect 17760 -770 17775 -575
rect 17820 -770 17835 -575
rect 17880 -770 17895 -575
rect 17940 -770 17955 -575
rect 18000 -770 18015 -575
rect 18060 -770 18075 -575
rect 18120 -770 18135 -575
rect 18180 -770 18195 -575
rect 18240 -770 18255 -575
rect 18300 -770 18315 -575
rect 18360 -770 18375 -575
rect 18420 -770 18435 -575
rect 18480 -770 18495 -575
rect 18540 -770 18555 -575
rect 18600 -770 18615 -575
rect 18660 -770 18675 -575
rect 18720 -770 18735 -575
rect 18780 -770 18795 -575
rect 18840 -770 18855 -575
rect 18900 -770 18915 -575
rect 18960 -770 18975 -575
rect 19020 -770 19035 -575
rect 19080 -770 19095 -575
rect 19140 -770 19155 -575
rect 19200 -770 19215 -575
rect 19260 -770 19275 -575
rect 19320 -770 19335 -575
rect 19380 -770 19395 -575
rect 19440 -770 19455 -575
rect 19500 -770 19515 -575
rect 19560 -770 19575 -575
rect 19620 -770 19635 -575
rect 19680 -770 19695 -575
rect 19740 -770 19755 -575
rect 19800 -770 19815 -575
rect 19860 -770 19875 -575
rect 19920 -770 19935 -575
rect 19980 -770 19995 -575
rect 20040 -770 20055 -575
rect 20100 -770 20115 -575
rect 20160 -770 20175 -575
rect 20220 -770 20235 -575
rect 20280 -770 20295 -575
rect 20340 -770 20355 -575
rect 20400 -770 20415 -575
rect 20460 -770 20475 -575
rect 20520 -770 20535 -575
rect 20580 -770 20595 -575
rect 20640 -770 20655 -575
rect 20700 -770 20715 -575
rect 20760 -770 20775 -575
rect 20820 -770 20835 -575
rect 20880 -770 20895 -575
rect 20940 -770 20955 -575
rect 21000 -770 21015 -575
rect 21060 -770 21075 -575
rect 21120 -770 21135 -575
rect 21180 -770 21195 -575
rect 21240 -770 21255 -575
rect 21300 -770 21315 -575
rect 21360 -770 21375 -575
rect 21420 -770 21435 -575
rect 21480 -770 21495 -575
rect 21540 -770 21555 -575
rect 21600 -770 21615 -575
rect 21660 -770 21675 -575
rect 21720 -770 21735 -575
rect 21780 -770 21795 -575
rect 21840 -770 21855 -575
rect 21900 -770 21915 -575
rect 21960 -770 21975 -575
rect 22020 -770 22035 -575
rect 22080 -770 22095 -575
rect 22140 -770 22155 -575
rect 22200 -770 22215 -575
rect 22260 -770 22275 -575
rect 22320 -770 22335 -575
rect 22380 -770 22395 -575
rect 22440 -770 22455 -575
rect 22500 -770 22515 -575
rect 22560 -770 22575 -575
rect 22620 -770 22635 -575
rect 22680 -770 22695 -575
rect 22740 -770 22755 -575
rect 22800 -770 22815 -575
rect 22860 -770 22875 -575
rect 22920 -770 22935 -575
rect 22980 -770 22995 -575
rect 23040 -770 23055 -575
rect 23100 -770 23115 -575
rect 23160 -770 23175 -575
rect 23220 -770 23235 -575
rect 23280 -770 23295 -575
rect 23340 -770 23355 -575
rect 23400 -770 23415 -575
rect 23460 -770 23475 -575
rect 23520 -770 23535 -575
rect 23580 -770 23595 -575
rect 23640 -770 23655 -575
rect 23700 -770 23715 -575
rect 23760 -770 23775 -575
rect 23820 -770 23835 -575
rect 23880 -770 23895 -575
rect 23940 -770 23955 -575
rect 24000 -770 24015 -575
rect 24060 -770 24075 -575
rect 24120 -770 24135 -575
rect 24180 -770 24195 -575
rect 24240 -770 24255 -575
rect 24300 -770 24315 -575
rect 24360 -770 24375 -575
rect 24420 -770 24435 -575
rect 24480 -770 24495 -575
rect 24540 -770 24555 -575
rect 24600 -770 24615 -575
rect 24660 -770 24675 -575
rect 24720 -770 24735 -575
rect 24780 -770 24795 -575
rect 24840 -770 24855 -575
rect 24900 -770 24915 -575
rect 24960 -770 24975 -575
rect 25020 -770 25035 -575
rect 25080 -770 25095 -575
rect 25140 -770 25155 -575
rect 25200 -770 25215 -575
rect 25260 -770 25275 -575
rect 25320 -770 25335 -575
rect 25380 -770 25395 -575
rect 25440 -770 25455 -575
rect 25500 -770 25515 -575
rect 25560 -770 25575 -575
rect 25620 -770 25635 -575
rect 25680 -770 25695 -575
rect 25740 -770 25755 -575
rect 25800 -770 25815 -575
rect 25860 -770 25875 -575
rect 25920 -770 25935 -575
rect 25980 -770 25995 -575
rect 26040 -770 26055 -575
rect 26100 -770 26115 -575
rect 26160 -770 26175 -575
rect 26220 -770 26235 -575
rect 26280 -770 26295 -575
rect 26340 -770 26355 -575
rect 26400 -770 26415 -575
rect 26460 -770 26475 -575
rect 26520 -770 26535 -575
rect 26580 -770 26595 -575
rect 26640 -770 26655 -575
rect 26700 -770 26715 -575
rect 26760 -770 26775 -575
rect 26820 -770 26835 -575
rect 26880 -770 26895 -575
rect 26940 -770 26955 -575
rect 27000 -770 27015 -575
rect 27060 -770 27075 -575
rect 27120 -770 27135 -575
rect 27180 -770 27195 -575
rect 27240 -770 27255 -575
rect 27300 -770 27315 -575
rect 27360 -770 27375 -575
rect 27420 -770 27435 -575
rect 27480 -770 27495 -575
rect 27540 -770 27555 -575
rect 27600 -770 27615 -575
rect 27660 -770 27675 -575
rect 27720 -770 27735 -575
rect 27780 -770 27795 -575
rect 27840 -770 27855 -575
rect 27900 -770 27915 -575
rect 27960 -770 27975 -575
rect 28020 -770 28035 -575
rect 28080 -770 28095 -575
rect 28140 -770 28155 -575
rect 28200 -770 28215 -575
rect 28260 -770 28275 -575
rect 28320 -770 28335 -575
rect 28380 -770 28395 -575
rect 28440 -770 28455 -575
rect 28500 -770 28515 -575
rect 28560 -770 28575 -575
rect 28620 -770 28635 -575
rect 28680 -770 28695 -575
rect 28740 -770 28755 -575
rect 28800 -770 28815 -575
rect 28860 -770 28875 -575
rect 28920 -770 28935 -575
rect 28980 -770 28995 -575
rect 29040 -770 29055 -575
rect 29100 -770 29115 -575
rect 29160 -770 29175 -575
rect 29220 -770 29235 -575
rect 29280 -770 29295 -575
rect 29340 -770 29355 -575
rect 29400 -770 29415 -575
rect 29460 -770 29475 -575
rect 29520 -770 29535 -575
rect 29580 -770 29595 -575
rect 29640 -770 29655 -575
rect 29700 -770 29715 -575
rect 29760 -770 29775 -575
rect 29820 -770 29835 -575
rect 29880 -770 29895 -575
rect 29940 -770 29955 -575
rect 30000 -770 30015 -575
rect 30060 -770 30075 -575
rect 30120 -770 30135 -575
rect 30180 -770 30195 -575
rect 30240 -770 30255 -575
rect 30300 -770 30315 -575
rect 30360 -770 30375 -575
rect 30420 -770 30435 -575
rect 30480 -770 30495 -575
rect 30540 -770 30555 -575
rect 30600 -770 30615 -575
rect 30660 -770 30675 -575
<< ndiff >>
rect 191 -85 231 -70
rect 191 -110 196 -85
rect 221 -110 231 -85
rect 191 -120 231 -110
rect 246 -85 286 -70
rect 246 -110 256 -85
rect 281 -110 286 -85
rect 246 -120 286 -110
rect 316 -85 356 -70
rect 316 -110 321 -85
rect 346 -110 356 -85
rect 316 -120 356 -110
rect 371 -85 416 -70
rect 371 -110 381 -85
rect 406 -110 416 -85
rect 371 -120 416 -110
rect 431 -85 476 -70
rect 431 -110 441 -85
rect 466 -110 476 -85
rect 431 -120 476 -110
rect 491 -85 536 -70
rect 491 -110 501 -85
rect 526 -110 536 -85
rect 491 -120 536 -110
rect 551 -85 591 -70
rect 551 -110 561 -85
rect 586 -110 591 -85
rect 551 -120 591 -110
rect 621 -85 661 -70
rect 621 -110 626 -85
rect 651 -110 661 -85
rect 621 -120 661 -110
rect 676 -85 721 -70
rect 676 -110 686 -85
rect 711 -110 721 -85
rect 676 -120 721 -110
rect 736 -85 781 -70
rect 736 -110 746 -85
rect 771 -110 781 -85
rect 736 -120 781 -110
rect 796 -85 841 -70
rect 796 -110 806 -85
rect 831 -110 841 -85
rect 796 -120 841 -110
rect 856 -85 906 -70
rect 856 -110 871 -85
rect 896 -110 906 -85
rect 856 -120 906 -110
rect 921 -85 966 -70
rect 921 -110 931 -85
rect 956 -110 966 -85
rect 921 -120 966 -110
rect 981 -85 1026 -70
rect 981 -110 991 -85
rect 1016 -110 1026 -85
rect 981 -120 1026 -110
rect 1041 -85 1086 -70
rect 1041 -110 1051 -85
rect 1076 -110 1086 -85
rect 1041 -120 1086 -110
rect 1101 -85 1146 -70
rect 1101 -110 1111 -85
rect 1136 -110 1146 -85
rect 1101 -120 1146 -110
rect 1161 -85 1206 -70
rect 1161 -110 1171 -85
rect 1196 -110 1206 -85
rect 1161 -120 1206 -110
rect 1221 -85 1266 -70
rect 1221 -110 1231 -85
rect 1256 -110 1266 -85
rect 1221 -120 1266 -110
rect 1281 -85 1326 -70
rect 1281 -110 1291 -85
rect 1316 -110 1326 -85
rect 1281 -120 1326 -110
rect 1341 -85 1391 -70
rect 1341 -110 1356 -85
rect 1381 -110 1391 -85
rect 1341 -120 1391 -110
rect 1406 -85 1451 -70
rect 1406 -110 1416 -85
rect 1441 -110 1451 -85
rect 1406 -120 1451 -110
rect 1466 -85 1511 -70
rect 1466 -110 1476 -85
rect 1501 -110 1511 -85
rect 1466 -120 1511 -110
rect 1526 -85 1571 -70
rect 1526 -110 1536 -85
rect 1561 -110 1571 -85
rect 1526 -120 1571 -110
rect 1586 -85 1626 -70
rect 1586 -110 1596 -85
rect 1621 -110 1626 -85
rect 1586 -120 1626 -110
rect 1656 -85 1696 -70
rect 1656 -110 1661 -85
rect 1686 -110 1696 -85
rect 1656 -120 1696 -110
rect 1711 -85 1756 -70
rect 1711 -110 1721 -85
rect 1746 -110 1756 -85
rect 1711 -120 1756 -110
rect 1771 -85 1816 -70
rect 1771 -110 1781 -85
rect 1806 -110 1816 -85
rect 1771 -120 1816 -110
rect 1831 -85 1876 -70
rect 1831 -110 1841 -85
rect 1866 -110 1876 -85
rect 1831 -120 1876 -110
rect 1891 -85 1941 -70
rect 1891 -110 1906 -85
rect 1931 -110 1941 -85
rect 1891 -120 1941 -110
rect 1956 -85 2001 -70
rect 1956 -110 1966 -85
rect 1991 -110 2001 -85
rect 1956 -120 2001 -110
rect 2016 -85 2061 -70
rect 2016 -110 2026 -85
rect 2051 -110 2061 -85
rect 2016 -120 2061 -110
rect 2076 -85 2121 -70
rect 2076 -110 2086 -85
rect 2111 -110 2121 -85
rect 2076 -120 2121 -110
rect 2136 -85 2181 -70
rect 2136 -110 2146 -85
rect 2171 -110 2181 -85
rect 2136 -120 2181 -110
rect 2196 -85 2241 -70
rect 2196 -110 2206 -85
rect 2231 -110 2241 -85
rect 2196 -120 2241 -110
rect 2256 -85 2301 -70
rect 2256 -110 2266 -85
rect 2291 -110 2301 -85
rect 2256 -120 2301 -110
rect 2316 -85 2361 -70
rect 2316 -110 2326 -85
rect 2351 -110 2361 -85
rect 2316 -120 2361 -110
rect 2376 -85 2426 -70
rect 2376 -110 2391 -85
rect 2416 -110 2426 -85
rect 2376 -120 2426 -110
rect 2441 -85 2486 -70
rect 2441 -110 2451 -85
rect 2476 -110 2486 -85
rect 2441 -120 2486 -110
rect 2501 -85 2546 -70
rect 2501 -110 2511 -85
rect 2536 -110 2546 -85
rect 2501 -120 2546 -110
rect 2561 -85 2606 -70
rect 2561 -110 2571 -85
rect 2596 -110 2606 -85
rect 2561 -120 2606 -110
rect 2621 -85 2666 -70
rect 2621 -110 2631 -85
rect 2656 -110 2666 -85
rect 2621 -120 2666 -110
rect 2681 -85 2726 -70
rect 2681 -110 2691 -85
rect 2716 -110 2726 -85
rect 2681 -120 2726 -110
rect 2741 -85 2786 -70
rect 2741 -110 2751 -85
rect 2776 -110 2786 -85
rect 2741 -120 2786 -110
rect 2801 -85 2846 -70
rect 2801 -110 2811 -85
rect 2836 -110 2846 -85
rect 2801 -120 2846 -110
rect 2861 -85 2911 -70
rect 2861 -110 2876 -85
rect 2901 -110 2911 -85
rect 2861 -120 2911 -110
rect 2926 -85 2971 -70
rect 2926 -110 2936 -85
rect 2961 -110 2971 -85
rect 2926 -120 2971 -110
rect 2986 -85 3031 -70
rect 2986 -110 2996 -85
rect 3021 -110 3031 -85
rect 2986 -120 3031 -110
rect 3046 -85 3091 -70
rect 3046 -110 3056 -85
rect 3081 -110 3091 -85
rect 3046 -120 3091 -110
rect 3106 -85 3151 -70
rect 3106 -110 3116 -85
rect 3141 -110 3151 -85
rect 3106 -120 3151 -110
rect 3166 -85 3211 -70
rect 3166 -110 3176 -85
rect 3201 -110 3211 -85
rect 3166 -120 3211 -110
rect 3226 -85 3271 -70
rect 3226 -110 3236 -85
rect 3261 -110 3271 -85
rect 3226 -120 3271 -110
rect 3286 -85 3331 -70
rect 3286 -110 3296 -85
rect 3321 -110 3331 -85
rect 3286 -120 3331 -110
rect 3346 -85 3396 -70
rect 3346 -110 3361 -85
rect 3386 -110 3396 -85
rect 3346 -120 3396 -110
rect 3411 -85 3456 -70
rect 3411 -110 3421 -85
rect 3446 -110 3456 -85
rect 3411 -120 3456 -110
rect 3471 -85 3516 -70
rect 3471 -110 3481 -85
rect 3506 -110 3516 -85
rect 3471 -120 3516 -110
rect 3531 -85 3576 -70
rect 3531 -110 3541 -85
rect 3566 -110 3576 -85
rect 3531 -120 3576 -110
rect 3591 -85 3636 -70
rect 3591 -110 3601 -85
rect 3626 -110 3636 -85
rect 3591 -120 3636 -110
rect 3651 -85 3696 -70
rect 3651 -110 3661 -85
rect 3686 -110 3696 -85
rect 3651 -120 3696 -110
rect 3711 -85 3756 -70
rect 3711 -110 3721 -85
rect 3746 -110 3756 -85
rect 3711 -120 3756 -110
rect 3771 -85 3816 -70
rect 3771 -110 3781 -85
rect 3806 -110 3816 -85
rect 3771 -120 3816 -110
rect 3831 -85 3881 -70
rect 3831 -110 3846 -85
rect 3871 -110 3881 -85
rect 3831 -120 3881 -110
rect 3896 -85 3941 -70
rect 3896 -110 3906 -85
rect 3931 -110 3941 -85
rect 3896 -120 3941 -110
rect 3956 -85 4001 -70
rect 3956 -110 3966 -85
rect 3991 -110 4001 -85
rect 3956 -120 4001 -110
rect 4016 -85 4061 -70
rect 4016 -110 4026 -85
rect 4051 -110 4061 -85
rect 4016 -120 4061 -110
rect 4076 -85 4121 -70
rect 4076 -110 4086 -85
rect 4111 -110 4121 -85
rect 4076 -120 4121 -110
rect 4136 -85 4181 -70
rect 4136 -110 4146 -85
rect 4171 -110 4181 -85
rect 4136 -120 4181 -110
rect 4196 -85 4241 -70
rect 4196 -110 4206 -85
rect 4231 -110 4241 -85
rect 4196 -120 4241 -110
rect 4256 -85 4301 -70
rect 4256 -110 4266 -85
rect 4291 -110 4301 -85
rect 4256 -120 4301 -110
rect 4316 -85 4366 -70
rect 4316 -110 4331 -85
rect 4356 -110 4366 -85
rect 4316 -120 4366 -110
rect 4381 -85 4426 -70
rect 4381 -110 4391 -85
rect 4416 -110 4426 -85
rect 4381 -120 4426 -110
rect 4441 -85 4486 -70
rect 4441 -110 4451 -85
rect 4476 -110 4486 -85
rect 4441 -120 4486 -110
rect 4501 -85 4546 -70
rect 4501 -110 4511 -85
rect 4536 -110 4546 -85
rect 4501 -120 4546 -110
rect 4561 -85 4606 -70
rect 4561 -110 4571 -85
rect 4596 -110 4606 -85
rect 4561 -120 4606 -110
rect 4621 -85 4666 -70
rect 4621 -110 4631 -85
rect 4656 -110 4666 -85
rect 4621 -120 4666 -110
rect 4681 -85 4726 -70
rect 4681 -110 4691 -85
rect 4716 -110 4726 -85
rect 4681 -120 4726 -110
rect 4741 -85 4786 -70
rect 4741 -110 4751 -85
rect 4776 -110 4786 -85
rect 4741 -120 4786 -110
rect 4801 -85 4851 -70
rect 4801 -110 4816 -85
rect 4841 -110 4851 -85
rect 4801 -120 4851 -110
rect 4866 -85 4911 -70
rect 4866 -110 4876 -85
rect 4901 -110 4911 -85
rect 4866 -120 4911 -110
rect 4926 -85 4971 -70
rect 4926 -110 4936 -85
rect 4961 -110 4971 -85
rect 4926 -120 4971 -110
rect 4986 -85 5031 -70
rect 4986 -110 4996 -85
rect 5021 -110 5031 -85
rect 4986 -120 5031 -110
rect 5046 -85 5091 -70
rect 5046 -110 5056 -85
rect 5081 -110 5091 -85
rect 5046 -120 5091 -110
rect 5106 -85 5151 -70
rect 5106 -110 5116 -85
rect 5141 -110 5151 -85
rect 5106 -120 5151 -110
rect 5166 -85 5211 -70
rect 5166 -110 5176 -85
rect 5201 -110 5211 -85
rect 5166 -120 5211 -110
rect 5226 -85 5271 -70
rect 5226 -110 5236 -85
rect 5261 -110 5271 -85
rect 5226 -120 5271 -110
rect 5286 -85 5336 -70
rect 5286 -110 5301 -85
rect 5326 -110 5336 -85
rect 5286 -120 5336 -110
rect 5351 -85 5396 -70
rect 5351 -110 5361 -85
rect 5386 -110 5396 -85
rect 5351 -120 5396 -110
rect 5411 -85 5456 -70
rect 5411 -110 5421 -85
rect 5446 -110 5456 -85
rect 5411 -120 5456 -110
rect 5471 -85 5516 -70
rect 5471 -110 5481 -85
rect 5506 -110 5516 -85
rect 5471 -120 5516 -110
rect 5531 -85 5571 -70
rect 5531 -110 5541 -85
rect 5566 -110 5571 -85
rect 5531 -120 5571 -110
rect 5601 -85 5641 -70
rect 5601 -110 5606 -85
rect 5631 -110 5641 -85
rect 5601 -120 5641 -110
rect 5656 -85 5701 -70
rect 5656 -110 5666 -85
rect 5691 -110 5701 -85
rect 5656 -120 5701 -110
rect 5716 -85 5761 -70
rect 5716 -110 5726 -85
rect 5751 -110 5761 -85
rect 5716 -120 5761 -110
rect 5776 -85 5821 -70
rect 5776 -110 5786 -85
rect 5811 -110 5821 -85
rect 5776 -120 5821 -110
rect 5836 -85 5886 -70
rect 5836 -110 5851 -85
rect 5876 -110 5886 -85
rect 5836 -120 5886 -110
rect 5901 -85 5946 -70
rect 5901 -110 5911 -85
rect 5936 -110 5946 -85
rect 5901 -120 5946 -110
rect 5961 -85 6006 -70
rect 5961 -110 5971 -85
rect 5996 -110 6006 -85
rect 5961 -120 6006 -110
rect 6021 -85 6066 -70
rect 6021 -110 6031 -85
rect 6056 -110 6066 -85
rect 6021 -120 6066 -110
rect 6081 -85 6126 -70
rect 6081 -110 6091 -85
rect 6116 -110 6126 -85
rect 6081 -120 6126 -110
rect 6141 -85 6186 -70
rect 6141 -110 6151 -85
rect 6176 -110 6186 -85
rect 6141 -120 6186 -110
rect 6201 -85 6246 -70
rect 6201 -110 6211 -85
rect 6236 -110 6246 -85
rect 6201 -120 6246 -110
rect 6261 -85 6306 -70
rect 6261 -110 6271 -85
rect 6296 -110 6306 -85
rect 6261 -120 6306 -110
rect 6321 -85 6371 -70
rect 6321 -110 6336 -85
rect 6361 -110 6371 -85
rect 6321 -120 6371 -110
rect 6386 -85 6431 -70
rect 6386 -110 6396 -85
rect 6421 -110 6431 -85
rect 6386 -120 6431 -110
rect 6446 -85 6491 -70
rect 6446 -110 6456 -85
rect 6481 -110 6491 -85
rect 6446 -120 6491 -110
rect 6506 -85 6551 -70
rect 6506 -110 6516 -85
rect 6541 -110 6551 -85
rect 6506 -120 6551 -110
rect 6566 -85 6611 -70
rect 6566 -110 6576 -85
rect 6601 -110 6611 -85
rect 6566 -120 6611 -110
rect 6626 -85 6671 -70
rect 6626 -110 6636 -85
rect 6661 -110 6671 -85
rect 6626 -120 6671 -110
rect 6686 -85 6731 -70
rect 6686 -110 6696 -85
rect 6721 -110 6731 -85
rect 6686 -120 6731 -110
rect 6746 -85 6791 -70
rect 6746 -110 6756 -85
rect 6781 -110 6791 -85
rect 6746 -120 6791 -110
rect 6806 -85 6856 -70
rect 6806 -110 6821 -85
rect 6846 -110 6856 -85
rect 6806 -120 6856 -110
rect 6871 -85 6916 -70
rect 6871 -110 6881 -85
rect 6906 -110 6916 -85
rect 6871 -120 6916 -110
rect 6931 -85 6976 -70
rect 6931 -110 6941 -85
rect 6966 -110 6976 -85
rect 6931 -120 6976 -110
rect 6991 -85 7036 -70
rect 6991 -110 7001 -85
rect 7026 -110 7036 -85
rect 6991 -120 7036 -110
rect 7051 -85 7096 -70
rect 7051 -110 7061 -85
rect 7086 -110 7096 -85
rect 7051 -120 7096 -110
rect 7111 -85 7156 -70
rect 7111 -110 7121 -85
rect 7146 -110 7156 -85
rect 7111 -120 7156 -110
rect 7171 -85 7216 -70
rect 7171 -110 7181 -85
rect 7206 -110 7216 -85
rect 7171 -120 7216 -110
rect 7231 -85 7276 -70
rect 7231 -110 7241 -85
rect 7266 -110 7276 -85
rect 7231 -120 7276 -110
rect 7291 -85 7336 -70
rect 7291 -110 7301 -85
rect 7326 -110 7336 -85
rect 7291 -120 7336 -110
rect 7351 -85 7396 -70
rect 7351 -110 7361 -85
rect 7386 -110 7396 -85
rect 7351 -120 7396 -110
rect 7411 -85 7456 -70
rect 7411 -110 7421 -85
rect 7446 -110 7456 -85
rect 7411 -120 7456 -110
rect 7471 -85 7516 -70
rect 7471 -110 7481 -85
rect 7506 -110 7516 -85
rect 7471 -120 7516 -110
rect 7531 -85 7576 -70
rect 7531 -110 7541 -85
rect 7566 -110 7576 -85
rect 7531 -120 7576 -110
rect 7591 -85 7636 -70
rect 7591 -110 7601 -85
rect 7626 -110 7636 -85
rect 7591 -120 7636 -110
rect 7651 -85 7696 -70
rect 7651 -110 7661 -85
rect 7686 -110 7696 -85
rect 7651 -120 7696 -110
rect 7711 -85 7756 -70
rect 7711 -110 7721 -85
rect 7746 -110 7756 -85
rect 7711 -120 7756 -110
rect 7771 -85 7821 -70
rect 7771 -110 7786 -85
rect 7811 -110 7821 -85
rect 7771 -120 7821 -110
rect 7836 -85 7881 -70
rect 7836 -110 7846 -85
rect 7871 -110 7881 -85
rect 7836 -120 7881 -110
rect 7896 -85 7941 -70
rect 7896 -110 7906 -85
rect 7931 -110 7941 -85
rect 7896 -120 7941 -110
rect 7956 -85 8001 -70
rect 7956 -110 7966 -85
rect 7991 -110 8001 -85
rect 7956 -120 8001 -110
rect 8016 -85 8061 -70
rect 8016 -110 8026 -85
rect 8051 -110 8061 -85
rect 8016 -120 8061 -110
rect 8076 -85 8121 -70
rect 8076 -110 8086 -85
rect 8111 -110 8121 -85
rect 8076 -120 8121 -110
rect 8136 -85 8181 -70
rect 8136 -110 8146 -85
rect 8171 -110 8181 -85
rect 8136 -120 8181 -110
rect 8196 -85 8241 -70
rect 8196 -110 8206 -85
rect 8231 -110 8241 -85
rect 8196 -120 8241 -110
rect 8256 -85 8306 -70
rect 8256 -110 8271 -85
rect 8296 -110 8306 -85
rect 8256 -120 8306 -110
rect 8321 -85 8366 -70
rect 8321 -110 8331 -85
rect 8356 -110 8366 -85
rect 8321 -120 8366 -110
rect 8381 -85 8426 -70
rect 8381 -110 8391 -85
rect 8416 -110 8426 -85
rect 8381 -120 8426 -110
rect 8441 -85 8486 -70
rect 8441 -110 8451 -85
rect 8476 -110 8486 -85
rect 8441 -120 8486 -110
rect 8501 -85 8546 -70
rect 8501 -110 8511 -85
rect 8536 -110 8546 -85
rect 8501 -120 8546 -110
rect 8561 -85 8606 -70
rect 8561 -110 8571 -85
rect 8596 -110 8606 -85
rect 8561 -120 8606 -110
rect 8621 -85 8666 -70
rect 8621 -110 8631 -85
rect 8656 -110 8666 -85
rect 8621 -120 8666 -110
rect 8681 -85 8726 -70
rect 8681 -110 8691 -85
rect 8716 -110 8726 -85
rect 8681 -120 8726 -110
rect 8741 -85 8791 -70
rect 8741 -110 8756 -85
rect 8781 -110 8791 -85
rect 8741 -120 8791 -110
rect 8806 -85 8851 -70
rect 8806 -110 8816 -85
rect 8841 -110 8851 -85
rect 8806 -120 8851 -110
rect 8866 -85 8911 -70
rect 8866 -110 8876 -85
rect 8901 -110 8911 -85
rect 8866 -120 8911 -110
rect 8926 -85 8971 -70
rect 8926 -110 8936 -85
rect 8961 -110 8971 -85
rect 8926 -120 8971 -110
rect 8986 -85 9031 -70
rect 8986 -110 8996 -85
rect 9021 -110 9031 -85
rect 8986 -120 9031 -110
rect 9046 -85 9091 -70
rect 9046 -110 9056 -85
rect 9081 -110 9091 -85
rect 9046 -120 9091 -110
rect 9106 -85 9151 -70
rect 9106 -110 9116 -85
rect 9141 -110 9151 -85
rect 9106 -120 9151 -110
rect 9166 -85 9211 -70
rect 9166 -110 9176 -85
rect 9201 -110 9211 -85
rect 9166 -120 9211 -110
rect 9226 -85 9276 -70
rect 9226 -110 9241 -85
rect 9266 -110 9276 -85
rect 9226 -120 9276 -110
rect 9291 -85 9336 -70
rect 9291 -110 9301 -85
rect 9326 -110 9336 -85
rect 9291 -120 9336 -110
rect 9351 -85 9396 -70
rect 9351 -110 9361 -85
rect 9386 -110 9396 -85
rect 9351 -120 9396 -110
rect 9411 -85 9456 -70
rect 9411 -110 9421 -85
rect 9446 -110 9456 -85
rect 9411 -120 9456 -110
rect 9471 -85 9521 -70
rect 9471 -110 9486 -85
rect 9511 -110 9521 -85
rect 9471 -120 9521 -110
rect 9536 -85 9581 -70
rect 9536 -110 9546 -85
rect 9571 -110 9581 -85
rect 9536 -120 9581 -110
rect 9596 -85 9641 -70
rect 9596 -110 9606 -85
rect 9631 -110 9641 -85
rect 9596 -120 9641 -110
rect 9656 -85 9701 -70
rect 9656 -110 9666 -85
rect 9691 -110 9701 -85
rect 9656 -120 9701 -110
rect 9716 -85 9766 -70
rect 9716 -110 9731 -85
rect 9756 -110 9766 -85
rect 9716 -120 9766 -110
rect 9781 -85 9826 -70
rect 9781 -110 9791 -85
rect 9816 -110 9826 -85
rect 9781 -120 9826 -110
rect 9841 -85 9886 -70
rect 9841 -110 9851 -85
rect 9876 -110 9886 -85
rect 9841 -120 9886 -110
rect 9901 -85 9946 -70
rect 9901 -110 9911 -85
rect 9936 -110 9946 -85
rect 9901 -120 9946 -110
rect 9961 -85 10006 -70
rect 9961 -110 9971 -85
rect 9996 -110 10006 -85
rect 9961 -120 10006 -110
rect 10021 -85 10066 -70
rect 10021 -110 10031 -85
rect 10056 -110 10066 -85
rect 10021 -120 10066 -110
rect 10081 -85 10126 -70
rect 10081 -110 10091 -85
rect 10116 -110 10126 -85
rect 10081 -120 10126 -110
rect 10141 -85 10186 -70
rect 10141 -110 10151 -85
rect 10176 -110 10186 -85
rect 10141 -120 10186 -110
rect 10201 -85 10251 -70
rect 10201 -110 10216 -85
rect 10241 -110 10251 -85
rect 10201 -120 10251 -110
rect 10266 -85 10311 -70
rect 10266 -110 10276 -85
rect 10301 -110 10311 -85
rect 10266 -120 10311 -110
rect 10326 -85 10371 -70
rect 10326 -110 10336 -85
rect 10361 -110 10371 -85
rect 10326 -120 10371 -110
rect 10386 -85 10431 -70
rect 10386 -110 10396 -85
rect 10421 -110 10431 -85
rect 10386 -120 10431 -110
rect 10446 -85 10491 -70
rect 10446 -110 10456 -85
rect 10481 -110 10491 -85
rect 10446 -120 10491 -110
rect 10506 -85 10551 -70
rect 10506 -110 10516 -85
rect 10541 -110 10551 -85
rect 10506 -120 10551 -110
rect 10566 -85 10611 -70
rect 10566 -110 10576 -85
rect 10601 -110 10611 -85
rect 10566 -120 10611 -110
rect 10626 -85 10671 -70
rect 10626 -110 10636 -85
rect 10661 -110 10671 -85
rect 10626 -120 10671 -110
rect 10686 -85 10736 -70
rect 10686 -110 10701 -85
rect 10726 -110 10736 -85
rect 10686 -120 10736 -110
rect 10751 -85 10796 -70
rect 10751 -110 10761 -85
rect 10786 -110 10796 -85
rect 10751 -120 10796 -110
rect 10811 -85 10856 -70
rect 10811 -110 10821 -85
rect 10846 -110 10856 -85
rect 10811 -120 10856 -110
rect 10871 -85 10916 -70
rect 10871 -110 10881 -85
rect 10906 -110 10916 -85
rect 10871 -120 10916 -110
rect 10931 -85 10976 -70
rect 10931 -110 10941 -85
rect 10966 -110 10976 -85
rect 10931 -120 10976 -110
rect 10991 -85 11036 -70
rect 10991 -110 11001 -85
rect 11026 -110 11036 -85
rect 10991 -120 11036 -110
rect 11051 -85 11096 -70
rect 11051 -110 11061 -85
rect 11086 -110 11096 -85
rect 11051 -120 11096 -110
rect 11111 -85 11156 -70
rect 11111 -110 11121 -85
rect 11146 -110 11156 -85
rect 11111 -120 11156 -110
rect 11171 -85 11221 -70
rect 11171 -110 11186 -85
rect 11211 -110 11221 -85
rect 11171 -120 11221 -110
rect 11236 -85 11281 -70
rect 11236 -110 11246 -85
rect 11271 -110 11281 -85
rect 11236 -120 11281 -110
rect 11296 -85 11341 -70
rect 11296 -110 11306 -85
rect 11331 -110 11341 -85
rect 11296 -120 11341 -110
rect 11356 -85 11401 -70
rect 11356 -110 11366 -85
rect 11391 -110 11401 -85
rect 11356 -120 11401 -110
rect 11416 -85 11461 -70
rect 11416 -110 11426 -85
rect 11451 -110 11461 -85
rect 11416 -120 11461 -110
rect 11476 -85 11521 -70
rect 11476 -110 11486 -85
rect 11511 -110 11521 -85
rect 11476 -120 11521 -110
rect 11536 -85 11581 -70
rect 11536 -110 11546 -85
rect 11571 -110 11581 -85
rect 11536 -120 11581 -110
rect 11596 -85 11641 -70
rect 11596 -110 11606 -85
rect 11631 -110 11641 -85
rect 11596 -120 11641 -110
rect 11656 -85 11706 -70
rect 11656 -110 11671 -85
rect 11696 -110 11706 -85
rect 11656 -120 11706 -110
rect 11721 -85 11766 -70
rect 11721 -110 11731 -85
rect 11756 -110 11766 -85
rect 11721 -120 11766 -110
rect 11781 -85 11826 -70
rect 11781 -110 11791 -85
rect 11816 -110 11826 -85
rect 11781 -120 11826 -110
rect 11841 -85 11886 -70
rect 11841 -110 11851 -85
rect 11876 -110 11886 -85
rect 11841 -120 11886 -110
rect 11901 -85 11946 -70
rect 11901 -110 11911 -85
rect 11936 -110 11946 -85
rect 11901 -120 11946 -110
rect 11961 -85 12006 -70
rect 11961 -110 11971 -85
rect 11996 -110 12006 -85
rect 11961 -120 12006 -110
rect 12021 -85 12066 -70
rect 12021 -110 12031 -85
rect 12056 -110 12066 -85
rect 12021 -120 12066 -110
rect 12081 -85 12126 -70
rect 12081 -110 12091 -85
rect 12116 -110 12126 -85
rect 12081 -120 12126 -110
rect 12141 -85 12191 -70
rect 12141 -110 12156 -85
rect 12181 -110 12191 -85
rect 12141 -120 12191 -110
rect 12206 -85 12251 -70
rect 12206 -110 12216 -85
rect 12241 -110 12251 -85
rect 12206 -120 12251 -110
rect 12266 -85 12311 -70
rect 12266 -110 12276 -85
rect 12301 -110 12311 -85
rect 12266 -120 12311 -110
rect 12326 -85 12371 -70
rect 12326 -110 12336 -85
rect 12361 -110 12371 -85
rect 12326 -120 12371 -110
rect 12386 -85 12431 -70
rect 12386 -110 12396 -85
rect 12421 -110 12431 -85
rect 12386 -120 12431 -110
rect 12446 -85 12491 -70
rect 12446 -110 12456 -85
rect 12481 -110 12491 -85
rect 12446 -120 12491 -110
rect 12506 -85 12551 -70
rect 12506 -110 12516 -85
rect 12541 -110 12551 -85
rect 12506 -120 12551 -110
rect 12566 -85 12611 -70
rect 12566 -110 12576 -85
rect 12601 -110 12611 -85
rect 12566 -120 12611 -110
rect 12626 -85 12676 -70
rect 12626 -110 12641 -85
rect 12666 -110 12676 -85
rect 12626 -120 12676 -110
rect 12691 -85 12736 -70
rect 12691 -110 12701 -85
rect 12726 -110 12736 -85
rect 12691 -120 12736 -110
rect 12751 -85 12796 -70
rect 12751 -110 12761 -85
rect 12786 -110 12796 -85
rect 12751 -120 12796 -110
rect 12811 -85 12856 -70
rect 12811 -110 12821 -85
rect 12846 -110 12856 -85
rect 12811 -120 12856 -110
rect 12871 -85 12916 -70
rect 12871 -110 12881 -85
rect 12906 -110 12916 -85
rect 12871 -120 12916 -110
rect 12931 -85 12976 -70
rect 12931 -110 12941 -85
rect 12966 -110 12976 -85
rect 12931 -120 12976 -110
rect 12991 -85 13036 -70
rect 12991 -110 13001 -85
rect 13026 -110 13036 -85
rect 12991 -120 13036 -110
rect 13051 -85 13096 -70
rect 13051 -110 13061 -85
rect 13086 -110 13096 -85
rect 13051 -120 13096 -110
rect 13111 -85 13161 -70
rect 13111 -110 13126 -85
rect 13151 -110 13161 -85
rect 13111 -120 13161 -110
rect 13176 -85 13221 -70
rect 13176 -110 13186 -85
rect 13211 -110 13221 -85
rect 13176 -120 13221 -110
rect 13236 -85 13281 -70
rect 13236 -110 13246 -85
rect 13271 -110 13281 -85
rect 13236 -120 13281 -110
rect 13296 -85 13341 -70
rect 13296 -110 13306 -85
rect 13331 -110 13341 -85
rect 13296 -120 13341 -110
rect 13356 -85 13401 -70
rect 13356 -110 13366 -85
rect 13391 -110 13401 -85
rect 13356 -120 13401 -110
rect 13416 -85 13461 -70
rect 13416 -110 13426 -85
rect 13451 -110 13461 -85
rect 13416 -120 13461 -110
rect 13476 -85 13521 -70
rect 13476 -110 13486 -85
rect 13511 -110 13521 -85
rect 13476 -120 13521 -110
rect 13536 -85 13581 -70
rect 13536 -110 13546 -85
rect 13571 -110 13581 -85
rect 13536 -120 13581 -110
rect 13596 -85 13646 -70
rect 13596 -110 13611 -85
rect 13636 -110 13646 -85
rect 13596 -120 13646 -110
rect 13661 -85 13706 -70
rect 13661 -110 13671 -85
rect 13696 -110 13706 -85
rect 13661 -120 13706 -110
rect 13721 -85 13766 -70
rect 13721 -110 13731 -85
rect 13756 -110 13766 -85
rect 13721 -120 13766 -110
rect 13781 -85 13826 -70
rect 13781 -110 13791 -85
rect 13816 -110 13826 -85
rect 13781 -120 13826 -110
rect 13841 -85 13886 -70
rect 13841 -110 13851 -85
rect 13876 -110 13886 -85
rect 13841 -120 13886 -110
rect 13901 -85 13946 -70
rect 13901 -110 13911 -85
rect 13936 -110 13946 -85
rect 13901 -120 13946 -110
rect 13961 -85 14006 -70
rect 13961 -110 13971 -85
rect 13996 -110 14006 -85
rect 13961 -120 14006 -110
rect 14021 -85 14066 -70
rect 14021 -110 14031 -85
rect 14056 -110 14066 -85
rect 14021 -120 14066 -110
rect 14081 -85 14131 -70
rect 14081 -110 14096 -85
rect 14121 -110 14131 -85
rect 14081 -120 14131 -110
rect 14146 -85 14191 -70
rect 14146 -110 14156 -85
rect 14181 -110 14191 -85
rect 14146 -120 14191 -110
rect 14206 -85 14251 -70
rect 14206 -110 14216 -85
rect 14241 -110 14251 -85
rect 14206 -120 14251 -110
rect 14266 -85 14311 -70
rect 14266 -110 14276 -85
rect 14301 -110 14311 -85
rect 14266 -120 14311 -110
rect 14326 -85 14371 -70
rect 14326 -110 14336 -85
rect 14361 -110 14371 -85
rect 14326 -120 14371 -110
rect 14386 -85 14431 -70
rect 14386 -110 14396 -85
rect 14421 -110 14431 -85
rect 14386 -120 14431 -110
rect 14446 -85 14491 -70
rect 14446 -110 14456 -85
rect 14481 -110 14491 -85
rect 14446 -120 14491 -110
rect 14506 -85 14551 -70
rect 14506 -110 14516 -85
rect 14541 -110 14551 -85
rect 14506 -120 14551 -110
rect 14566 -85 14616 -70
rect 14566 -110 14581 -85
rect 14606 -110 14616 -85
rect 14566 -120 14616 -110
rect 14631 -85 14676 -70
rect 14631 -110 14641 -85
rect 14666 -110 14676 -85
rect 14631 -120 14676 -110
rect 14691 -85 14736 -70
rect 14691 -110 14701 -85
rect 14726 -110 14736 -85
rect 14691 -120 14736 -110
rect 14751 -85 14796 -70
rect 14751 -110 14761 -85
rect 14786 -110 14796 -85
rect 14751 -120 14796 -110
rect 14811 -85 14856 -70
rect 14811 -110 14821 -85
rect 14846 -110 14856 -85
rect 14811 -120 14856 -110
rect 14871 -85 14916 -70
rect 14871 -110 14881 -85
rect 14906 -110 14916 -85
rect 14871 -120 14916 -110
rect 14931 -85 14976 -70
rect 14931 -110 14941 -85
rect 14966 -110 14976 -85
rect 14931 -120 14976 -110
rect 14991 -85 15036 -70
rect 14991 -110 15001 -85
rect 15026 -110 15036 -85
rect 14991 -120 15036 -110
rect 15051 -85 15101 -70
rect 15051 -110 15066 -85
rect 15091 -110 15101 -85
rect 15051 -120 15101 -110
rect 15116 -85 15161 -70
rect 15116 -110 15126 -85
rect 15151 -110 15161 -85
rect 15116 -120 15161 -110
rect 15176 -85 15221 -70
rect 15176 -110 15186 -85
rect 15211 -110 15221 -85
rect 15176 -120 15221 -110
rect 15236 -85 15281 -70
rect 15236 -110 15246 -85
rect 15271 -110 15281 -85
rect 15236 -120 15281 -110
rect 15296 -85 15341 -70
rect 15296 -110 15306 -85
rect 15331 -110 15341 -85
rect 15296 -120 15341 -110
rect 15356 -85 15401 -70
rect 15356 -110 15366 -85
rect 15391 -110 15401 -85
rect 15356 -120 15401 -110
rect 15416 -85 15461 -70
rect 15416 -110 15426 -85
rect 15451 -110 15461 -85
rect 15416 -120 15461 -110
rect 15476 -85 15521 -70
rect 15476 -110 15486 -85
rect 15511 -110 15521 -85
rect 15476 -120 15521 -110
rect 15536 -85 15586 -70
rect 15536 -110 15551 -85
rect 15576 -110 15586 -85
rect 15536 -120 15586 -110
rect 15601 -85 15646 -70
rect 15601 -110 15611 -85
rect 15636 -110 15646 -85
rect 15601 -120 15646 -110
rect 15661 -85 15706 -70
rect 15661 -110 15671 -85
rect 15696 -110 15706 -85
rect 15661 -120 15706 -110
rect 15721 -85 15766 -70
rect 15721 -110 15731 -85
rect 15756 -110 15766 -85
rect 15721 -120 15766 -110
rect 15781 -85 15826 -70
rect 15781 -110 15791 -85
rect 15816 -110 15826 -85
rect 15781 -120 15826 -110
rect 15841 -85 15886 -70
rect 15841 -110 15851 -85
rect 15876 -110 15886 -85
rect 15841 -120 15886 -110
rect 15901 -85 15946 -70
rect 15901 -110 15911 -85
rect 15936 -110 15946 -85
rect 15901 -120 15946 -110
rect 15961 -85 16006 -70
rect 15961 -110 15971 -85
rect 15996 -110 16006 -85
rect 15961 -120 16006 -110
rect 16021 -85 16071 -70
rect 16021 -110 16036 -85
rect 16061 -110 16071 -85
rect 16021 -120 16071 -110
rect 16086 -85 16131 -70
rect 16086 -110 16096 -85
rect 16121 -110 16131 -85
rect 16086 -120 16131 -110
rect 16146 -85 16191 -70
rect 16146 -110 16156 -85
rect 16181 -110 16191 -85
rect 16146 -120 16191 -110
rect 16206 -85 16251 -70
rect 16206 -110 16216 -85
rect 16241 -110 16251 -85
rect 16206 -120 16251 -110
rect 16266 -85 16311 -70
rect 16266 -110 16276 -85
rect 16301 -110 16311 -85
rect 16266 -120 16311 -110
rect 16326 -85 16371 -70
rect 16326 -110 16336 -85
rect 16361 -110 16371 -85
rect 16326 -120 16371 -110
rect 16386 -85 16431 -70
rect 16386 -110 16396 -85
rect 16421 -110 16431 -85
rect 16386 -120 16431 -110
rect 16446 -85 16491 -70
rect 16446 -110 16456 -85
rect 16481 -110 16491 -85
rect 16446 -120 16491 -110
rect 16506 -85 16556 -70
rect 16506 -110 16521 -85
rect 16546 -110 16556 -85
rect 16506 -120 16556 -110
rect 16571 -85 16616 -70
rect 16571 -110 16581 -85
rect 16606 -110 16616 -85
rect 16571 -120 16616 -110
rect 16631 -85 16676 -70
rect 16631 -110 16641 -85
rect 16666 -110 16676 -85
rect 16631 -120 16676 -110
rect 16691 -85 16736 -70
rect 16691 -110 16701 -85
rect 16726 -110 16736 -85
rect 16691 -120 16736 -110
rect 16751 -85 16796 -70
rect 16751 -110 16761 -85
rect 16786 -110 16796 -85
rect 16751 -120 16796 -110
rect 16811 -85 16856 -70
rect 16811 -110 16821 -85
rect 16846 -110 16856 -85
rect 16811 -120 16856 -110
rect 16871 -85 16916 -70
rect 16871 -110 16881 -85
rect 16906 -110 16916 -85
rect 16871 -120 16916 -110
rect 16931 -85 16976 -70
rect 16931 -110 16941 -85
rect 16966 -110 16976 -85
rect 16931 -120 16976 -110
rect 16991 -85 17041 -70
rect 16991 -110 17006 -85
rect 17031 -110 17041 -85
rect 16991 -120 17041 -110
rect 17056 -85 17101 -70
rect 17056 -110 17066 -85
rect 17091 -110 17101 -85
rect 17056 -120 17101 -110
rect 17116 -85 17161 -70
rect 17116 -110 17126 -85
rect 17151 -110 17161 -85
rect 17116 -120 17161 -110
rect 17176 -85 17221 -70
rect 17176 -110 17186 -85
rect 17211 -110 17221 -85
rect 17176 -120 17221 -110
rect 17236 -85 17281 -70
rect 17236 -110 17246 -85
rect 17271 -110 17281 -85
rect 17236 -120 17281 -110
rect 17296 -85 17341 -70
rect 17296 -110 17306 -85
rect 17331 -110 17341 -85
rect 17296 -120 17341 -110
rect 17356 -85 17401 -70
rect 17356 -110 17366 -85
rect 17391 -110 17401 -85
rect 17356 -120 17401 -110
rect 17416 -85 17461 -70
rect 17416 -110 17426 -85
rect 17451 -110 17461 -85
rect 17416 -120 17461 -110
rect 17476 -85 17526 -70
rect 17476 -110 17491 -85
rect 17516 -110 17526 -85
rect 17476 -120 17526 -110
rect 17541 -85 17586 -70
rect 17541 -110 17551 -85
rect 17576 -110 17586 -85
rect 17541 -120 17586 -110
rect 17601 -85 17646 -70
rect 17601 -110 17611 -85
rect 17636 -110 17646 -85
rect 17601 -120 17646 -110
rect 17661 -85 17706 -70
rect 17661 -110 17671 -85
rect 17696 -110 17706 -85
rect 17661 -120 17706 -110
rect 17721 -85 17766 -70
rect 17721 -110 17731 -85
rect 17756 -110 17766 -85
rect 17721 -120 17766 -110
rect 17781 -85 17826 -70
rect 17781 -110 17791 -85
rect 17816 -110 17826 -85
rect 17781 -120 17826 -110
rect 17841 -85 17886 -70
rect 17841 -110 17851 -85
rect 17876 -110 17886 -85
rect 17841 -120 17886 -110
rect 17901 -85 17946 -70
rect 17901 -110 17911 -85
rect 17936 -110 17946 -85
rect 17901 -120 17946 -110
rect 17961 -85 18011 -70
rect 17961 -110 17976 -85
rect 18001 -110 18011 -85
rect 17961 -120 18011 -110
rect 18026 -85 18071 -70
rect 18026 -110 18036 -85
rect 18061 -110 18071 -85
rect 18026 -120 18071 -110
rect 18086 -85 18131 -70
rect 18086 -110 18096 -85
rect 18121 -110 18131 -85
rect 18086 -120 18131 -110
rect 18146 -85 18191 -70
rect 18146 -110 18156 -85
rect 18181 -110 18191 -85
rect 18146 -120 18191 -110
rect 18206 -85 18251 -70
rect 18206 -110 18216 -85
rect 18241 -110 18251 -85
rect 18206 -120 18251 -110
rect 18266 -85 18311 -70
rect 18266 -110 18276 -85
rect 18301 -110 18311 -85
rect 18266 -120 18311 -110
rect 18326 -85 18371 -70
rect 18326 -110 18336 -85
rect 18361 -110 18371 -85
rect 18326 -120 18371 -110
rect 18386 -85 18431 -70
rect 18386 -110 18396 -85
rect 18421 -110 18431 -85
rect 18386 -120 18431 -110
rect 18446 -85 18496 -70
rect 18446 -110 18461 -85
rect 18486 -110 18496 -85
rect 18446 -120 18496 -110
rect 18511 -85 18556 -70
rect 18511 -110 18521 -85
rect 18546 -110 18556 -85
rect 18511 -120 18556 -110
rect 18571 -85 18616 -70
rect 18571 -110 18581 -85
rect 18606 -110 18616 -85
rect 18571 -120 18616 -110
rect 18631 -85 18676 -70
rect 18631 -110 18641 -85
rect 18666 -110 18676 -85
rect 18631 -120 18676 -110
rect 18691 -85 18736 -70
rect 18691 -110 18701 -85
rect 18726 -110 18736 -85
rect 18691 -120 18736 -110
rect 18751 -85 18796 -70
rect 18751 -110 18761 -85
rect 18786 -110 18796 -85
rect 18751 -120 18796 -110
rect 18811 -85 18856 -70
rect 18811 -110 18821 -85
rect 18846 -110 18856 -85
rect 18811 -120 18856 -110
rect 18871 -85 18916 -70
rect 18871 -110 18881 -85
rect 18906 -110 18916 -85
rect 18871 -120 18916 -110
rect 18931 -85 18981 -70
rect 18931 -110 18946 -85
rect 18971 -110 18981 -85
rect 18931 -120 18981 -110
rect 18996 -85 19041 -70
rect 18996 -110 19006 -85
rect 19031 -110 19041 -85
rect 18996 -120 19041 -110
rect 19056 -85 19101 -70
rect 19056 -110 19066 -85
rect 19091 -110 19101 -85
rect 19056 -120 19101 -110
rect 19116 -85 19161 -70
rect 19116 -110 19126 -85
rect 19151 -110 19161 -85
rect 19116 -120 19161 -110
rect 19176 -85 19221 -70
rect 19176 -110 19186 -85
rect 19211 -110 19221 -85
rect 19176 -120 19221 -110
rect 19236 -85 19281 -70
rect 19236 -110 19246 -85
rect 19271 -110 19281 -85
rect 19236 -120 19281 -110
rect 19296 -85 19341 -70
rect 19296 -110 19306 -85
rect 19331 -110 19341 -85
rect 19296 -120 19341 -110
rect 19356 -85 19401 -70
rect 19356 -110 19366 -85
rect 19391 -110 19401 -85
rect 19356 -120 19401 -110
rect 19416 -85 19466 -70
rect 19416 -110 19431 -85
rect 19456 -110 19466 -85
rect 19416 -120 19466 -110
rect 19481 -85 19526 -70
rect 19481 -110 19491 -85
rect 19516 -110 19526 -85
rect 19481 -120 19526 -110
rect 19541 -85 19586 -70
rect 19541 -110 19551 -85
rect 19576 -110 19586 -85
rect 19541 -120 19586 -110
rect 19601 -85 19646 -70
rect 19601 -110 19611 -85
rect 19636 -110 19646 -85
rect 19601 -120 19646 -110
rect 19661 -85 19706 -70
rect 19661 -110 19671 -85
rect 19696 -110 19706 -85
rect 19661 -120 19706 -110
rect 19721 -85 19766 -70
rect 19721 -110 19731 -85
rect 19756 -110 19766 -85
rect 19721 -120 19766 -110
rect 19781 -85 19826 -70
rect 19781 -110 19791 -85
rect 19816 -110 19826 -85
rect 19781 -120 19826 -110
rect 19841 -85 19886 -70
rect 19841 -110 19851 -85
rect 19876 -110 19886 -85
rect 19841 -120 19886 -110
rect 19901 -85 19951 -70
rect 19901 -110 19916 -85
rect 19941 -110 19951 -85
rect 19901 -120 19951 -110
rect 19966 -85 20011 -70
rect 19966 -110 19976 -85
rect 20001 -110 20011 -85
rect 19966 -120 20011 -110
rect 20026 -85 20071 -70
rect 20026 -110 20036 -85
rect 20061 -110 20071 -85
rect 20026 -120 20071 -110
rect 20086 -85 20131 -70
rect 20086 -110 20096 -85
rect 20121 -110 20131 -85
rect 20086 -120 20131 -110
rect 20146 -85 20191 -70
rect 20146 -110 20156 -85
rect 20181 -110 20191 -85
rect 20146 -120 20191 -110
rect 20206 -85 20251 -70
rect 20206 -110 20216 -85
rect 20241 -110 20251 -85
rect 20206 -120 20251 -110
rect 20266 -85 20311 -70
rect 20266 -110 20276 -85
rect 20301 -110 20311 -85
rect 20266 -120 20311 -110
rect 20326 -85 20371 -70
rect 20326 -110 20336 -85
rect 20361 -110 20371 -85
rect 20326 -120 20371 -110
rect 20386 -85 20436 -70
rect 20386 -110 20401 -85
rect 20426 -110 20436 -85
rect 20386 -120 20436 -110
rect 20451 -85 20496 -70
rect 20451 -110 20461 -85
rect 20486 -110 20496 -85
rect 20451 -120 20496 -110
rect 20511 -85 20556 -70
rect 20511 -110 20521 -85
rect 20546 -110 20556 -85
rect 20511 -120 20556 -110
rect 20571 -85 20616 -70
rect 20571 -110 20581 -85
rect 20606 -110 20616 -85
rect 20571 -120 20616 -110
rect 20631 -85 20676 -70
rect 20631 -110 20641 -85
rect 20666 -110 20676 -85
rect 20631 -120 20676 -110
rect 20691 -85 20736 -70
rect 20691 -110 20701 -85
rect 20726 -110 20736 -85
rect 20691 -120 20736 -110
rect 20751 -85 20796 -70
rect 20751 -110 20761 -85
rect 20786 -110 20796 -85
rect 20751 -120 20796 -110
rect 20811 -85 20856 -70
rect 20811 -110 20821 -85
rect 20846 -110 20856 -85
rect 20811 -120 20856 -110
rect 20871 -85 20921 -70
rect 20871 -110 20886 -85
rect 20911 -110 20921 -85
rect 20871 -120 20921 -110
rect 20936 -85 20981 -70
rect 20936 -110 20946 -85
rect 20971 -110 20981 -85
rect 20936 -120 20981 -110
rect 20996 -85 21041 -70
rect 20996 -110 21006 -85
rect 21031 -110 21041 -85
rect 20996 -120 21041 -110
rect 21056 -85 21101 -70
rect 21056 -110 21066 -85
rect 21091 -110 21101 -85
rect 21056 -120 21101 -110
rect 21116 -85 21156 -70
rect 21116 -110 21126 -85
rect 21151 -110 21156 -85
rect 21116 -120 21156 -110
rect -40 -335 0 -320
rect -40 -360 -35 -335
rect -10 -360 0 -335
rect -40 -380 0 -360
rect -40 -405 -35 -380
rect -10 -405 0 -380
rect -40 -420 0 -405
rect 15 -335 60 -320
rect 15 -360 25 -335
rect 50 -360 60 -335
rect 15 -380 60 -360
rect 15 -405 25 -380
rect 50 -405 60 -380
rect 15 -420 60 -405
rect 75 -335 120 -320
rect 75 -360 85 -335
rect 110 -360 120 -335
rect 75 -380 120 -360
rect 75 -405 85 -380
rect 110 -405 120 -380
rect 75 -420 120 -405
rect 135 -335 180 -320
rect 135 -360 145 -335
rect 170 -360 180 -335
rect 135 -380 180 -360
rect 135 -405 145 -380
rect 170 -405 180 -380
rect 135 -420 180 -405
rect 195 -335 240 -320
rect 195 -360 205 -335
rect 230 -360 240 -335
rect 195 -380 240 -360
rect 195 -405 205 -380
rect 230 -405 240 -380
rect 195 -420 240 -405
rect 255 -335 300 -320
rect 255 -360 265 -335
rect 290 -360 300 -335
rect 255 -380 300 -360
rect 255 -405 265 -380
rect 290 -405 300 -380
rect 255 -420 300 -405
rect 315 -335 360 -320
rect 315 -360 325 -335
rect 350 -360 360 -335
rect 315 -380 360 -360
rect 315 -405 325 -380
rect 350 -405 360 -380
rect 315 -420 360 -405
rect 375 -335 420 -320
rect 375 -360 385 -335
rect 410 -360 420 -335
rect 375 -380 420 -360
rect 375 -405 385 -380
rect 410 -405 420 -380
rect 375 -420 420 -405
rect 435 -335 480 -320
rect 435 -360 445 -335
rect 470 -360 480 -335
rect 435 -380 480 -360
rect 435 -405 445 -380
rect 470 -405 480 -380
rect 435 -420 480 -405
rect 495 -335 540 -320
rect 495 -360 505 -335
rect 530 -360 540 -335
rect 495 -380 540 -360
rect 495 -405 505 -380
rect 530 -405 540 -380
rect 495 -420 540 -405
rect 555 -335 600 -320
rect 555 -360 565 -335
rect 590 -360 600 -335
rect 555 -380 600 -360
rect 555 -405 565 -380
rect 590 -405 600 -380
rect 555 -420 600 -405
rect 615 -335 660 -320
rect 615 -360 625 -335
rect 650 -360 660 -335
rect 615 -380 660 -360
rect 615 -405 625 -380
rect 650 -405 660 -380
rect 615 -420 660 -405
rect 675 -335 720 -320
rect 675 -360 685 -335
rect 710 -360 720 -335
rect 675 -380 720 -360
rect 675 -405 685 -380
rect 710 -405 720 -380
rect 675 -420 720 -405
rect 735 -335 780 -320
rect 735 -360 745 -335
rect 770 -360 780 -335
rect 735 -380 780 -360
rect 735 -405 745 -380
rect 770 -405 780 -380
rect 735 -420 780 -405
rect 795 -335 840 -320
rect 795 -360 805 -335
rect 830 -360 840 -335
rect 795 -380 840 -360
rect 795 -405 805 -380
rect 830 -405 840 -380
rect 795 -420 840 -405
rect 855 -335 900 -320
rect 855 -360 865 -335
rect 890 -360 900 -335
rect 855 -380 900 -360
rect 855 -405 865 -380
rect 890 -405 900 -380
rect 855 -420 900 -405
rect 915 -335 960 -320
rect 915 -360 925 -335
rect 950 -360 960 -335
rect 915 -380 960 -360
rect 915 -405 925 -380
rect 950 -405 960 -380
rect 915 -420 960 -405
rect 975 -335 1020 -320
rect 975 -360 985 -335
rect 1010 -360 1020 -335
rect 975 -380 1020 -360
rect 975 -405 985 -380
rect 1010 -405 1020 -380
rect 975 -420 1020 -405
rect 1035 -335 1080 -320
rect 1035 -360 1045 -335
rect 1070 -360 1080 -335
rect 1035 -380 1080 -360
rect 1035 -405 1045 -380
rect 1070 -405 1080 -380
rect 1035 -420 1080 -405
rect 1095 -335 1140 -320
rect 1095 -360 1105 -335
rect 1130 -360 1140 -335
rect 1095 -380 1140 -360
rect 1095 -405 1105 -380
rect 1130 -405 1140 -380
rect 1095 -420 1140 -405
rect 1155 -335 1200 -320
rect 1155 -360 1165 -335
rect 1190 -360 1200 -335
rect 1155 -380 1200 -360
rect 1155 -405 1165 -380
rect 1190 -405 1200 -380
rect 1155 -420 1200 -405
rect 1215 -335 1260 -320
rect 1215 -360 1225 -335
rect 1250 -360 1260 -335
rect 1215 -380 1260 -360
rect 1215 -405 1225 -380
rect 1250 -405 1260 -380
rect 1215 -420 1260 -405
rect 1275 -335 1320 -320
rect 1275 -360 1285 -335
rect 1310 -360 1320 -335
rect 1275 -380 1320 -360
rect 1275 -405 1285 -380
rect 1310 -405 1320 -380
rect 1275 -420 1320 -405
rect 1335 -335 1380 -320
rect 1335 -360 1345 -335
rect 1370 -360 1380 -335
rect 1335 -380 1380 -360
rect 1335 -405 1345 -380
rect 1370 -405 1380 -380
rect 1335 -420 1380 -405
rect 1395 -335 1440 -320
rect 1395 -360 1405 -335
rect 1430 -360 1440 -335
rect 1395 -380 1440 -360
rect 1395 -405 1405 -380
rect 1430 -405 1440 -380
rect 1395 -420 1440 -405
rect 1455 -335 1500 -320
rect 1455 -360 1465 -335
rect 1490 -360 1500 -335
rect 1455 -380 1500 -360
rect 1455 -405 1465 -380
rect 1490 -405 1500 -380
rect 1455 -420 1500 -405
rect 1515 -335 1560 -320
rect 1515 -360 1525 -335
rect 1550 -360 1560 -335
rect 1515 -380 1560 -360
rect 1515 -405 1525 -380
rect 1550 -405 1560 -380
rect 1515 -420 1560 -405
rect 1575 -335 1620 -320
rect 1575 -360 1585 -335
rect 1610 -360 1620 -335
rect 1575 -380 1620 -360
rect 1575 -405 1585 -380
rect 1610 -405 1620 -380
rect 1575 -420 1620 -405
rect 1635 -335 1680 -320
rect 1635 -360 1645 -335
rect 1670 -360 1680 -335
rect 1635 -380 1680 -360
rect 1635 -405 1645 -380
rect 1670 -405 1680 -380
rect 1635 -420 1680 -405
rect 1695 -335 1740 -320
rect 1695 -360 1705 -335
rect 1730 -360 1740 -335
rect 1695 -380 1740 -360
rect 1695 -405 1705 -380
rect 1730 -405 1740 -380
rect 1695 -420 1740 -405
rect 1755 -335 1800 -320
rect 1755 -360 1765 -335
rect 1790 -360 1800 -335
rect 1755 -380 1800 -360
rect 1755 -405 1765 -380
rect 1790 -405 1800 -380
rect 1755 -420 1800 -405
rect 1815 -335 1860 -320
rect 1815 -360 1825 -335
rect 1850 -360 1860 -335
rect 1815 -380 1860 -360
rect 1815 -405 1825 -380
rect 1850 -405 1860 -380
rect 1815 -420 1860 -405
rect 1875 -335 1920 -320
rect 1875 -360 1885 -335
rect 1910 -360 1920 -335
rect 1875 -380 1920 -360
rect 1875 -405 1885 -380
rect 1910 -405 1920 -380
rect 1875 -420 1920 -405
rect 1935 -335 1980 -320
rect 1935 -360 1945 -335
rect 1970 -360 1980 -335
rect 1935 -380 1980 -360
rect 1935 -405 1945 -380
rect 1970 -405 1980 -380
rect 1935 -420 1980 -405
rect 1995 -335 2040 -320
rect 1995 -360 2005 -335
rect 2030 -360 2040 -335
rect 1995 -380 2040 -360
rect 1995 -405 2005 -380
rect 2030 -405 2040 -380
rect 1995 -420 2040 -405
rect 2055 -335 2100 -320
rect 2055 -360 2065 -335
rect 2090 -360 2100 -335
rect 2055 -380 2100 -360
rect 2055 -405 2065 -380
rect 2090 -405 2100 -380
rect 2055 -420 2100 -405
rect 2115 -335 2160 -320
rect 2115 -360 2125 -335
rect 2150 -360 2160 -335
rect 2115 -380 2160 -360
rect 2115 -405 2125 -380
rect 2150 -405 2160 -380
rect 2115 -420 2160 -405
rect 2175 -335 2220 -320
rect 2175 -360 2185 -335
rect 2210 -360 2220 -335
rect 2175 -380 2220 -360
rect 2175 -405 2185 -380
rect 2210 -405 2220 -380
rect 2175 -420 2220 -405
rect 2235 -335 2280 -320
rect 2235 -360 2245 -335
rect 2270 -360 2280 -335
rect 2235 -380 2280 -360
rect 2235 -405 2245 -380
rect 2270 -405 2280 -380
rect 2235 -420 2280 -405
rect 2295 -335 2340 -320
rect 2295 -360 2305 -335
rect 2330 -360 2340 -335
rect 2295 -380 2340 -360
rect 2295 -405 2305 -380
rect 2330 -405 2340 -380
rect 2295 -420 2340 -405
rect 2355 -335 2400 -320
rect 2355 -360 2365 -335
rect 2390 -360 2400 -335
rect 2355 -380 2400 -360
rect 2355 -405 2365 -380
rect 2390 -405 2400 -380
rect 2355 -420 2400 -405
rect 2415 -335 2460 -320
rect 2415 -360 2425 -335
rect 2450 -360 2460 -335
rect 2415 -380 2460 -360
rect 2415 -405 2425 -380
rect 2450 -405 2460 -380
rect 2415 -420 2460 -405
rect 2475 -335 2520 -320
rect 2475 -360 2485 -335
rect 2510 -360 2520 -335
rect 2475 -380 2520 -360
rect 2475 -405 2485 -380
rect 2510 -405 2520 -380
rect 2475 -420 2520 -405
rect 2535 -335 2580 -320
rect 2535 -360 2545 -335
rect 2570 -360 2580 -335
rect 2535 -380 2580 -360
rect 2535 -405 2545 -380
rect 2570 -405 2580 -380
rect 2535 -420 2580 -405
rect 2595 -335 2640 -320
rect 2595 -360 2605 -335
rect 2630 -360 2640 -335
rect 2595 -380 2640 -360
rect 2595 -405 2605 -380
rect 2630 -405 2640 -380
rect 2595 -420 2640 -405
rect 2655 -335 2700 -320
rect 2655 -360 2665 -335
rect 2690 -360 2700 -335
rect 2655 -380 2700 -360
rect 2655 -405 2665 -380
rect 2690 -405 2700 -380
rect 2655 -420 2700 -405
rect 2715 -335 2760 -320
rect 2715 -360 2725 -335
rect 2750 -360 2760 -335
rect 2715 -380 2760 -360
rect 2715 -405 2725 -380
rect 2750 -405 2760 -380
rect 2715 -420 2760 -405
rect 2775 -335 2820 -320
rect 2775 -360 2785 -335
rect 2810 -360 2820 -335
rect 2775 -380 2820 -360
rect 2775 -405 2785 -380
rect 2810 -405 2820 -380
rect 2775 -420 2820 -405
rect 2835 -335 2880 -320
rect 2835 -360 2845 -335
rect 2870 -360 2880 -335
rect 2835 -380 2880 -360
rect 2835 -405 2845 -380
rect 2870 -405 2880 -380
rect 2835 -420 2880 -405
rect 2895 -335 2940 -320
rect 2895 -360 2905 -335
rect 2930 -360 2940 -335
rect 2895 -380 2940 -360
rect 2895 -405 2905 -380
rect 2930 -405 2940 -380
rect 2895 -420 2940 -405
rect 2955 -335 3000 -320
rect 2955 -360 2965 -335
rect 2990 -360 3000 -335
rect 2955 -380 3000 -360
rect 2955 -405 2965 -380
rect 2990 -405 3000 -380
rect 2955 -420 3000 -405
rect 3015 -335 3060 -320
rect 3015 -360 3025 -335
rect 3050 -360 3060 -335
rect 3015 -380 3060 -360
rect 3015 -405 3025 -380
rect 3050 -405 3060 -380
rect 3015 -420 3060 -405
rect 3075 -335 3120 -320
rect 3075 -360 3085 -335
rect 3110 -360 3120 -335
rect 3075 -380 3120 -360
rect 3075 -405 3085 -380
rect 3110 -405 3120 -380
rect 3075 -420 3120 -405
rect 3135 -335 3180 -320
rect 3135 -360 3145 -335
rect 3170 -360 3180 -335
rect 3135 -380 3180 -360
rect 3135 -405 3145 -380
rect 3170 -405 3180 -380
rect 3135 -420 3180 -405
rect 3195 -335 3240 -320
rect 3195 -360 3205 -335
rect 3230 -360 3240 -335
rect 3195 -380 3240 -360
rect 3195 -405 3205 -380
rect 3230 -405 3240 -380
rect 3195 -420 3240 -405
rect 3255 -335 3300 -320
rect 3255 -360 3265 -335
rect 3290 -360 3300 -335
rect 3255 -380 3300 -360
rect 3255 -405 3265 -380
rect 3290 -405 3300 -380
rect 3255 -420 3300 -405
rect 3315 -335 3360 -320
rect 3315 -360 3325 -335
rect 3350 -360 3360 -335
rect 3315 -380 3360 -360
rect 3315 -405 3325 -380
rect 3350 -405 3360 -380
rect 3315 -420 3360 -405
rect 3375 -335 3420 -320
rect 3375 -360 3385 -335
rect 3410 -360 3420 -335
rect 3375 -380 3420 -360
rect 3375 -405 3385 -380
rect 3410 -405 3420 -380
rect 3375 -420 3420 -405
rect 3435 -335 3480 -320
rect 3435 -360 3445 -335
rect 3470 -360 3480 -335
rect 3435 -380 3480 -360
rect 3435 -405 3445 -380
rect 3470 -405 3480 -380
rect 3435 -420 3480 -405
rect 3495 -335 3540 -320
rect 3495 -360 3505 -335
rect 3530 -360 3540 -335
rect 3495 -380 3540 -360
rect 3495 -405 3505 -380
rect 3530 -405 3540 -380
rect 3495 -420 3540 -405
rect 3555 -335 3600 -320
rect 3555 -360 3565 -335
rect 3590 -360 3600 -335
rect 3555 -380 3600 -360
rect 3555 -405 3565 -380
rect 3590 -405 3600 -380
rect 3555 -420 3600 -405
rect 3615 -335 3660 -320
rect 3615 -360 3625 -335
rect 3650 -360 3660 -335
rect 3615 -380 3660 -360
rect 3615 -405 3625 -380
rect 3650 -405 3660 -380
rect 3615 -420 3660 -405
rect 3675 -335 3720 -320
rect 3675 -360 3685 -335
rect 3710 -360 3720 -335
rect 3675 -380 3720 -360
rect 3675 -405 3685 -380
rect 3710 -405 3720 -380
rect 3675 -420 3720 -405
rect 3735 -335 3780 -320
rect 3735 -360 3745 -335
rect 3770 -360 3780 -335
rect 3735 -380 3780 -360
rect 3735 -405 3745 -380
rect 3770 -405 3780 -380
rect 3735 -420 3780 -405
rect 3795 -335 3840 -320
rect 3795 -360 3805 -335
rect 3830 -360 3840 -335
rect 3795 -380 3840 -360
rect 3795 -405 3805 -380
rect 3830 -405 3840 -380
rect 3795 -420 3840 -405
rect 3855 -335 3900 -320
rect 3855 -360 3865 -335
rect 3890 -360 3900 -335
rect 3855 -380 3900 -360
rect 3855 -405 3865 -380
rect 3890 -405 3900 -380
rect 3855 -420 3900 -405
rect 3915 -335 3960 -320
rect 3915 -360 3925 -335
rect 3950 -360 3960 -335
rect 3915 -380 3960 -360
rect 3915 -405 3925 -380
rect 3950 -405 3960 -380
rect 3915 -420 3960 -405
rect 3975 -335 4020 -320
rect 3975 -360 3985 -335
rect 4010 -360 4020 -335
rect 3975 -380 4020 -360
rect 3975 -405 3985 -380
rect 4010 -405 4020 -380
rect 3975 -420 4020 -405
rect 4035 -335 4080 -320
rect 4035 -360 4045 -335
rect 4070 -360 4080 -335
rect 4035 -380 4080 -360
rect 4035 -405 4045 -380
rect 4070 -405 4080 -380
rect 4035 -420 4080 -405
rect 4095 -335 4140 -320
rect 4095 -360 4105 -335
rect 4130 -360 4140 -335
rect 4095 -380 4140 -360
rect 4095 -405 4105 -380
rect 4130 -405 4140 -380
rect 4095 -420 4140 -405
rect 4155 -335 4200 -320
rect 4155 -360 4165 -335
rect 4190 -360 4200 -335
rect 4155 -380 4200 -360
rect 4155 -405 4165 -380
rect 4190 -405 4200 -380
rect 4155 -420 4200 -405
rect 4215 -335 4260 -320
rect 4215 -360 4225 -335
rect 4250 -360 4260 -335
rect 4215 -380 4260 -360
rect 4215 -405 4225 -380
rect 4250 -405 4260 -380
rect 4215 -420 4260 -405
rect 4275 -335 4320 -320
rect 4275 -360 4285 -335
rect 4310 -360 4320 -335
rect 4275 -380 4320 -360
rect 4275 -405 4285 -380
rect 4310 -405 4320 -380
rect 4275 -420 4320 -405
rect 4335 -335 4380 -320
rect 4335 -360 4345 -335
rect 4370 -360 4380 -335
rect 4335 -380 4380 -360
rect 4335 -405 4345 -380
rect 4370 -405 4380 -380
rect 4335 -420 4380 -405
rect 4395 -335 4440 -320
rect 4395 -360 4405 -335
rect 4430 -360 4440 -335
rect 4395 -380 4440 -360
rect 4395 -405 4405 -380
rect 4430 -405 4440 -380
rect 4395 -420 4440 -405
rect 4455 -335 4500 -320
rect 4455 -360 4465 -335
rect 4490 -360 4500 -335
rect 4455 -380 4500 -360
rect 4455 -405 4465 -380
rect 4490 -405 4500 -380
rect 4455 -420 4500 -405
rect 4515 -335 4560 -320
rect 4515 -360 4525 -335
rect 4550 -360 4560 -335
rect 4515 -380 4560 -360
rect 4515 -405 4525 -380
rect 4550 -405 4560 -380
rect 4515 -420 4560 -405
rect 4575 -335 4620 -320
rect 4575 -360 4585 -335
rect 4610 -360 4620 -335
rect 4575 -380 4620 -360
rect 4575 -405 4585 -380
rect 4610 -405 4620 -380
rect 4575 -420 4620 -405
rect 4635 -335 4680 -320
rect 4635 -360 4645 -335
rect 4670 -360 4680 -335
rect 4635 -380 4680 -360
rect 4635 -405 4645 -380
rect 4670 -405 4680 -380
rect 4635 -420 4680 -405
rect 4695 -335 4740 -320
rect 4695 -360 4705 -335
rect 4730 -360 4740 -335
rect 4695 -380 4740 -360
rect 4695 -405 4705 -380
rect 4730 -405 4740 -380
rect 4695 -420 4740 -405
rect 4755 -335 4800 -320
rect 4755 -360 4765 -335
rect 4790 -360 4800 -335
rect 4755 -380 4800 -360
rect 4755 -405 4765 -380
rect 4790 -405 4800 -380
rect 4755 -420 4800 -405
rect 4815 -335 4860 -320
rect 4815 -360 4825 -335
rect 4850 -360 4860 -335
rect 4815 -380 4860 -360
rect 4815 -405 4825 -380
rect 4850 -405 4860 -380
rect 4815 -420 4860 -405
rect 4875 -335 4920 -320
rect 4875 -360 4885 -335
rect 4910 -360 4920 -335
rect 4875 -380 4920 -360
rect 4875 -405 4885 -380
rect 4910 -405 4920 -380
rect 4875 -420 4920 -405
rect 4935 -335 4980 -320
rect 4935 -360 4945 -335
rect 4970 -360 4980 -335
rect 4935 -380 4980 -360
rect 4935 -405 4945 -380
rect 4970 -405 4980 -380
rect 4935 -420 4980 -405
rect 4995 -335 5040 -320
rect 4995 -360 5005 -335
rect 5030 -360 5040 -335
rect 4995 -380 5040 -360
rect 4995 -405 5005 -380
rect 5030 -405 5040 -380
rect 4995 -420 5040 -405
rect 5055 -335 5100 -320
rect 5055 -360 5065 -335
rect 5090 -360 5100 -335
rect 5055 -380 5100 -360
rect 5055 -405 5065 -380
rect 5090 -405 5100 -380
rect 5055 -420 5100 -405
rect 5115 -335 5160 -320
rect 5115 -360 5125 -335
rect 5150 -360 5160 -335
rect 5115 -380 5160 -360
rect 5115 -405 5125 -380
rect 5150 -405 5160 -380
rect 5115 -420 5160 -405
rect 5175 -335 5220 -320
rect 5175 -360 5185 -335
rect 5210 -360 5220 -335
rect 5175 -380 5220 -360
rect 5175 -405 5185 -380
rect 5210 -405 5220 -380
rect 5175 -420 5220 -405
rect 5235 -335 5280 -320
rect 5235 -360 5245 -335
rect 5270 -360 5280 -335
rect 5235 -380 5280 -360
rect 5235 -405 5245 -380
rect 5270 -405 5280 -380
rect 5235 -420 5280 -405
rect 5295 -335 5340 -320
rect 5295 -360 5305 -335
rect 5330 -360 5340 -335
rect 5295 -380 5340 -360
rect 5295 -405 5305 -380
rect 5330 -405 5340 -380
rect 5295 -420 5340 -405
rect 5355 -335 5400 -320
rect 5355 -360 5365 -335
rect 5390 -360 5400 -335
rect 5355 -380 5400 -360
rect 5355 -405 5365 -380
rect 5390 -405 5400 -380
rect 5355 -420 5400 -405
rect 5415 -335 5460 -320
rect 5415 -360 5425 -335
rect 5450 -360 5460 -335
rect 5415 -380 5460 -360
rect 5415 -405 5425 -380
rect 5450 -405 5460 -380
rect 5415 -420 5460 -405
rect 5475 -335 5520 -320
rect 5475 -360 5485 -335
rect 5510 -360 5520 -335
rect 5475 -380 5520 -360
rect 5475 -405 5485 -380
rect 5510 -405 5520 -380
rect 5475 -420 5520 -405
rect 5535 -335 5580 -320
rect 5535 -360 5545 -335
rect 5570 -360 5580 -335
rect 5535 -380 5580 -360
rect 5535 -405 5545 -380
rect 5570 -405 5580 -380
rect 5535 -420 5580 -405
rect 5595 -335 5640 -320
rect 5595 -360 5605 -335
rect 5630 -360 5640 -335
rect 5595 -380 5640 -360
rect 5595 -405 5605 -380
rect 5630 -405 5640 -380
rect 5595 -420 5640 -405
rect 5655 -335 5700 -320
rect 5655 -360 5665 -335
rect 5690 -360 5700 -335
rect 5655 -380 5700 -360
rect 5655 -405 5665 -380
rect 5690 -405 5700 -380
rect 5655 -420 5700 -405
rect 5715 -335 5760 -320
rect 5715 -360 5725 -335
rect 5750 -360 5760 -335
rect 5715 -380 5760 -360
rect 5715 -405 5725 -380
rect 5750 -405 5760 -380
rect 5715 -420 5760 -405
rect 5775 -335 5820 -320
rect 5775 -360 5785 -335
rect 5810 -360 5820 -335
rect 5775 -380 5820 -360
rect 5775 -405 5785 -380
rect 5810 -405 5820 -380
rect 5775 -420 5820 -405
rect 5835 -335 5880 -320
rect 5835 -360 5845 -335
rect 5870 -360 5880 -335
rect 5835 -380 5880 -360
rect 5835 -405 5845 -380
rect 5870 -405 5880 -380
rect 5835 -420 5880 -405
rect 5895 -335 5940 -320
rect 5895 -360 5905 -335
rect 5930 -360 5940 -335
rect 5895 -380 5940 -360
rect 5895 -405 5905 -380
rect 5930 -405 5940 -380
rect 5895 -420 5940 -405
rect 5955 -335 6000 -320
rect 5955 -360 5965 -335
rect 5990 -360 6000 -335
rect 5955 -380 6000 -360
rect 5955 -405 5965 -380
rect 5990 -405 6000 -380
rect 5955 -420 6000 -405
rect 6015 -335 6060 -320
rect 6015 -360 6025 -335
rect 6050 -360 6060 -335
rect 6015 -380 6060 -360
rect 6015 -405 6025 -380
rect 6050 -405 6060 -380
rect 6015 -420 6060 -405
rect 6075 -335 6120 -320
rect 6075 -360 6085 -335
rect 6110 -360 6120 -335
rect 6075 -380 6120 -360
rect 6075 -405 6085 -380
rect 6110 -405 6120 -380
rect 6075 -420 6120 -405
rect 6135 -335 6180 -320
rect 6135 -360 6145 -335
rect 6170 -360 6180 -335
rect 6135 -380 6180 -360
rect 6135 -405 6145 -380
rect 6170 -405 6180 -380
rect 6135 -420 6180 -405
rect 6195 -335 6240 -320
rect 6195 -360 6205 -335
rect 6230 -360 6240 -335
rect 6195 -380 6240 -360
rect 6195 -405 6205 -380
rect 6230 -405 6240 -380
rect 6195 -420 6240 -405
rect 6255 -335 6300 -320
rect 6255 -360 6265 -335
rect 6290 -360 6300 -335
rect 6255 -380 6300 -360
rect 6255 -405 6265 -380
rect 6290 -405 6300 -380
rect 6255 -420 6300 -405
rect 6315 -335 6360 -320
rect 6315 -360 6325 -335
rect 6350 -360 6360 -335
rect 6315 -380 6360 -360
rect 6315 -405 6325 -380
rect 6350 -405 6360 -380
rect 6315 -420 6360 -405
rect 6375 -335 6420 -320
rect 6375 -360 6385 -335
rect 6410 -360 6420 -335
rect 6375 -380 6420 -360
rect 6375 -405 6385 -380
rect 6410 -405 6420 -380
rect 6375 -420 6420 -405
rect 6435 -335 6480 -320
rect 6435 -360 6445 -335
rect 6470 -360 6480 -335
rect 6435 -380 6480 -360
rect 6435 -405 6445 -380
rect 6470 -405 6480 -380
rect 6435 -420 6480 -405
rect 6495 -335 6540 -320
rect 6495 -360 6505 -335
rect 6530 -360 6540 -335
rect 6495 -380 6540 -360
rect 6495 -405 6505 -380
rect 6530 -405 6540 -380
rect 6495 -420 6540 -405
rect 6555 -335 6600 -320
rect 6555 -360 6565 -335
rect 6590 -360 6600 -335
rect 6555 -380 6600 -360
rect 6555 -405 6565 -380
rect 6590 -405 6600 -380
rect 6555 -420 6600 -405
rect 6615 -335 6660 -320
rect 6615 -360 6625 -335
rect 6650 -360 6660 -335
rect 6615 -380 6660 -360
rect 6615 -405 6625 -380
rect 6650 -405 6660 -380
rect 6615 -420 6660 -405
rect 6675 -335 6720 -320
rect 6675 -360 6685 -335
rect 6710 -360 6720 -335
rect 6675 -380 6720 -360
rect 6675 -405 6685 -380
rect 6710 -405 6720 -380
rect 6675 -420 6720 -405
rect 6735 -335 6780 -320
rect 6735 -360 6745 -335
rect 6770 -360 6780 -335
rect 6735 -380 6780 -360
rect 6735 -405 6745 -380
rect 6770 -405 6780 -380
rect 6735 -420 6780 -405
rect 6795 -335 6840 -320
rect 6795 -360 6805 -335
rect 6830 -360 6840 -335
rect 6795 -380 6840 -360
rect 6795 -405 6805 -380
rect 6830 -405 6840 -380
rect 6795 -420 6840 -405
rect 6855 -335 6900 -320
rect 6855 -360 6865 -335
rect 6890 -360 6900 -335
rect 6855 -380 6900 -360
rect 6855 -405 6865 -380
rect 6890 -405 6900 -380
rect 6855 -420 6900 -405
rect 6915 -335 6960 -320
rect 6915 -360 6925 -335
rect 6950 -360 6960 -335
rect 6915 -380 6960 -360
rect 6915 -405 6925 -380
rect 6950 -405 6960 -380
rect 6915 -420 6960 -405
rect 6975 -335 7020 -320
rect 6975 -360 6985 -335
rect 7010 -360 7020 -335
rect 6975 -380 7020 -360
rect 6975 -405 6985 -380
rect 7010 -405 7020 -380
rect 6975 -420 7020 -405
rect 7035 -335 7080 -320
rect 7035 -360 7045 -335
rect 7070 -360 7080 -335
rect 7035 -380 7080 -360
rect 7035 -405 7045 -380
rect 7070 -405 7080 -380
rect 7035 -420 7080 -405
rect 7095 -335 7140 -320
rect 7095 -360 7105 -335
rect 7130 -360 7140 -335
rect 7095 -380 7140 -360
rect 7095 -405 7105 -380
rect 7130 -405 7140 -380
rect 7095 -420 7140 -405
rect 7155 -335 7200 -320
rect 7155 -360 7165 -335
rect 7190 -360 7200 -335
rect 7155 -380 7200 -360
rect 7155 -405 7165 -380
rect 7190 -405 7200 -380
rect 7155 -420 7200 -405
rect 7215 -335 7260 -320
rect 7215 -360 7225 -335
rect 7250 -360 7260 -335
rect 7215 -380 7260 -360
rect 7215 -405 7225 -380
rect 7250 -405 7260 -380
rect 7215 -420 7260 -405
rect 7275 -335 7320 -320
rect 7275 -360 7285 -335
rect 7310 -360 7320 -335
rect 7275 -380 7320 -360
rect 7275 -405 7285 -380
rect 7310 -405 7320 -380
rect 7275 -420 7320 -405
rect 7335 -335 7380 -320
rect 7335 -360 7345 -335
rect 7370 -360 7380 -335
rect 7335 -380 7380 -360
rect 7335 -405 7345 -380
rect 7370 -405 7380 -380
rect 7335 -420 7380 -405
rect 7395 -335 7440 -320
rect 7395 -360 7405 -335
rect 7430 -360 7440 -335
rect 7395 -380 7440 -360
rect 7395 -405 7405 -380
rect 7430 -405 7440 -380
rect 7395 -420 7440 -405
rect 7455 -335 7500 -320
rect 7455 -360 7465 -335
rect 7490 -360 7500 -335
rect 7455 -380 7500 -360
rect 7455 -405 7465 -380
rect 7490 -405 7500 -380
rect 7455 -420 7500 -405
rect 7515 -335 7560 -320
rect 7515 -360 7525 -335
rect 7550 -360 7560 -335
rect 7515 -380 7560 -360
rect 7515 -405 7525 -380
rect 7550 -405 7560 -380
rect 7515 -420 7560 -405
rect 7575 -335 7620 -320
rect 7575 -360 7585 -335
rect 7610 -360 7620 -335
rect 7575 -380 7620 -360
rect 7575 -405 7585 -380
rect 7610 -405 7620 -380
rect 7575 -420 7620 -405
rect 7635 -335 7680 -320
rect 7635 -360 7645 -335
rect 7670 -360 7680 -335
rect 7635 -380 7680 -360
rect 7635 -405 7645 -380
rect 7670 -405 7680 -380
rect 7635 -420 7680 -405
rect 7695 -335 7740 -320
rect 7695 -360 7705 -335
rect 7730 -360 7740 -335
rect 7695 -380 7740 -360
rect 7695 -405 7705 -380
rect 7730 -405 7740 -380
rect 7695 -420 7740 -405
rect 7755 -335 7800 -320
rect 7755 -360 7765 -335
rect 7790 -360 7800 -335
rect 7755 -380 7800 -360
rect 7755 -405 7765 -380
rect 7790 -405 7800 -380
rect 7755 -420 7800 -405
rect 7815 -335 7860 -320
rect 7815 -360 7825 -335
rect 7850 -360 7860 -335
rect 7815 -380 7860 -360
rect 7815 -405 7825 -380
rect 7850 -405 7860 -380
rect 7815 -420 7860 -405
rect 7875 -335 7920 -320
rect 7875 -360 7885 -335
rect 7910 -360 7920 -335
rect 7875 -380 7920 -360
rect 7875 -405 7885 -380
rect 7910 -405 7920 -380
rect 7875 -420 7920 -405
rect 7935 -335 7980 -320
rect 7935 -360 7945 -335
rect 7970 -360 7980 -335
rect 7935 -380 7980 -360
rect 7935 -405 7945 -380
rect 7970 -405 7980 -380
rect 7935 -420 7980 -405
rect 7995 -335 8040 -320
rect 7995 -360 8005 -335
rect 8030 -360 8040 -335
rect 7995 -380 8040 -360
rect 7995 -405 8005 -380
rect 8030 -405 8040 -380
rect 7995 -420 8040 -405
rect 8055 -335 8100 -320
rect 8055 -360 8065 -335
rect 8090 -360 8100 -335
rect 8055 -380 8100 -360
rect 8055 -405 8065 -380
rect 8090 -405 8100 -380
rect 8055 -420 8100 -405
rect 8115 -335 8160 -320
rect 8115 -360 8125 -335
rect 8150 -360 8160 -335
rect 8115 -380 8160 -360
rect 8115 -405 8125 -380
rect 8150 -405 8160 -380
rect 8115 -420 8160 -405
rect 8175 -335 8220 -320
rect 8175 -360 8185 -335
rect 8210 -360 8220 -335
rect 8175 -380 8220 -360
rect 8175 -405 8185 -380
rect 8210 -405 8220 -380
rect 8175 -420 8220 -405
rect 8235 -335 8280 -320
rect 8235 -360 8245 -335
rect 8270 -360 8280 -335
rect 8235 -380 8280 -360
rect 8235 -405 8245 -380
rect 8270 -405 8280 -380
rect 8235 -420 8280 -405
rect 8295 -335 8340 -320
rect 8295 -360 8305 -335
rect 8330 -360 8340 -335
rect 8295 -380 8340 -360
rect 8295 -405 8305 -380
rect 8330 -405 8340 -380
rect 8295 -420 8340 -405
rect 8355 -335 8400 -320
rect 8355 -360 8365 -335
rect 8390 -360 8400 -335
rect 8355 -380 8400 -360
rect 8355 -405 8365 -380
rect 8390 -405 8400 -380
rect 8355 -420 8400 -405
rect 8415 -335 8460 -320
rect 8415 -360 8425 -335
rect 8450 -360 8460 -335
rect 8415 -380 8460 -360
rect 8415 -405 8425 -380
rect 8450 -405 8460 -380
rect 8415 -420 8460 -405
rect 8475 -335 8520 -320
rect 8475 -360 8485 -335
rect 8510 -360 8520 -335
rect 8475 -380 8520 -360
rect 8475 -405 8485 -380
rect 8510 -405 8520 -380
rect 8475 -420 8520 -405
rect 8535 -335 8580 -320
rect 8535 -360 8545 -335
rect 8570 -360 8580 -335
rect 8535 -380 8580 -360
rect 8535 -405 8545 -380
rect 8570 -405 8580 -380
rect 8535 -420 8580 -405
rect 8595 -335 8640 -320
rect 8595 -360 8605 -335
rect 8630 -360 8640 -335
rect 8595 -380 8640 -360
rect 8595 -405 8605 -380
rect 8630 -405 8640 -380
rect 8595 -420 8640 -405
rect 8655 -335 8700 -320
rect 8655 -360 8665 -335
rect 8690 -360 8700 -335
rect 8655 -380 8700 -360
rect 8655 -405 8665 -380
rect 8690 -405 8700 -380
rect 8655 -420 8700 -405
rect 8715 -335 8760 -320
rect 8715 -360 8725 -335
rect 8750 -360 8760 -335
rect 8715 -380 8760 -360
rect 8715 -405 8725 -380
rect 8750 -405 8760 -380
rect 8715 -420 8760 -405
rect 8775 -335 8820 -320
rect 8775 -360 8785 -335
rect 8810 -360 8820 -335
rect 8775 -380 8820 -360
rect 8775 -405 8785 -380
rect 8810 -405 8820 -380
rect 8775 -420 8820 -405
rect 8835 -335 8880 -320
rect 8835 -360 8845 -335
rect 8870 -360 8880 -335
rect 8835 -380 8880 -360
rect 8835 -405 8845 -380
rect 8870 -405 8880 -380
rect 8835 -420 8880 -405
rect 8895 -335 8940 -320
rect 8895 -360 8905 -335
rect 8930 -360 8940 -335
rect 8895 -380 8940 -360
rect 8895 -405 8905 -380
rect 8930 -405 8940 -380
rect 8895 -420 8940 -405
rect 8955 -335 9000 -320
rect 8955 -360 8965 -335
rect 8990 -360 9000 -335
rect 8955 -380 9000 -360
rect 8955 -405 8965 -380
rect 8990 -405 9000 -380
rect 8955 -420 9000 -405
rect 9015 -335 9060 -320
rect 9015 -360 9025 -335
rect 9050 -360 9060 -335
rect 9015 -380 9060 -360
rect 9015 -405 9025 -380
rect 9050 -405 9060 -380
rect 9015 -420 9060 -405
rect 9075 -335 9120 -320
rect 9075 -360 9085 -335
rect 9110 -360 9120 -335
rect 9075 -380 9120 -360
rect 9075 -405 9085 -380
rect 9110 -405 9120 -380
rect 9075 -420 9120 -405
rect 9135 -335 9180 -320
rect 9135 -360 9145 -335
rect 9170 -360 9180 -335
rect 9135 -380 9180 -360
rect 9135 -405 9145 -380
rect 9170 -405 9180 -380
rect 9135 -420 9180 -405
rect 9195 -335 9240 -320
rect 9195 -360 9205 -335
rect 9230 -360 9240 -335
rect 9195 -380 9240 -360
rect 9195 -405 9205 -380
rect 9230 -405 9240 -380
rect 9195 -420 9240 -405
rect 9255 -335 9300 -320
rect 9255 -360 9265 -335
rect 9290 -360 9300 -335
rect 9255 -380 9300 -360
rect 9255 -405 9265 -380
rect 9290 -405 9300 -380
rect 9255 -420 9300 -405
rect 9315 -335 9360 -320
rect 9315 -360 9325 -335
rect 9350 -360 9360 -335
rect 9315 -380 9360 -360
rect 9315 -405 9325 -380
rect 9350 -405 9360 -380
rect 9315 -420 9360 -405
rect 9375 -335 9420 -320
rect 9375 -360 9385 -335
rect 9410 -360 9420 -335
rect 9375 -380 9420 -360
rect 9375 -405 9385 -380
rect 9410 -405 9420 -380
rect 9375 -420 9420 -405
rect 9435 -335 9480 -320
rect 9435 -360 9445 -335
rect 9470 -360 9480 -335
rect 9435 -380 9480 -360
rect 9435 -405 9445 -380
rect 9470 -405 9480 -380
rect 9435 -420 9480 -405
rect 9495 -335 9540 -320
rect 9495 -360 9505 -335
rect 9530 -360 9540 -335
rect 9495 -380 9540 -360
rect 9495 -405 9505 -380
rect 9530 -405 9540 -380
rect 9495 -420 9540 -405
rect 9555 -335 9600 -320
rect 9555 -360 9565 -335
rect 9590 -360 9600 -335
rect 9555 -380 9600 -360
rect 9555 -405 9565 -380
rect 9590 -405 9600 -380
rect 9555 -420 9600 -405
rect 9615 -335 9660 -320
rect 9615 -360 9625 -335
rect 9650 -360 9660 -335
rect 9615 -380 9660 -360
rect 9615 -405 9625 -380
rect 9650 -405 9660 -380
rect 9615 -420 9660 -405
rect 9675 -335 9720 -320
rect 9675 -360 9685 -335
rect 9710 -360 9720 -335
rect 9675 -380 9720 -360
rect 9675 -405 9685 -380
rect 9710 -405 9720 -380
rect 9675 -420 9720 -405
rect 9735 -335 9780 -320
rect 9735 -360 9745 -335
rect 9770 -360 9780 -335
rect 9735 -380 9780 -360
rect 9735 -405 9745 -380
rect 9770 -405 9780 -380
rect 9735 -420 9780 -405
rect 9795 -335 9840 -320
rect 9795 -360 9805 -335
rect 9830 -360 9840 -335
rect 9795 -380 9840 -360
rect 9795 -405 9805 -380
rect 9830 -405 9840 -380
rect 9795 -420 9840 -405
rect 9855 -335 9900 -320
rect 9855 -360 9865 -335
rect 9890 -360 9900 -335
rect 9855 -380 9900 -360
rect 9855 -405 9865 -380
rect 9890 -405 9900 -380
rect 9855 -420 9900 -405
rect 9915 -335 9960 -320
rect 9915 -360 9925 -335
rect 9950 -360 9960 -335
rect 9915 -380 9960 -360
rect 9915 -405 9925 -380
rect 9950 -405 9960 -380
rect 9915 -420 9960 -405
rect 9975 -335 10020 -320
rect 9975 -360 9985 -335
rect 10010 -360 10020 -335
rect 9975 -380 10020 -360
rect 9975 -405 9985 -380
rect 10010 -405 10020 -380
rect 9975 -420 10020 -405
rect 10035 -335 10080 -320
rect 10035 -360 10045 -335
rect 10070 -360 10080 -335
rect 10035 -380 10080 -360
rect 10035 -405 10045 -380
rect 10070 -405 10080 -380
rect 10035 -420 10080 -405
rect 10095 -335 10140 -320
rect 10095 -360 10105 -335
rect 10130 -360 10140 -335
rect 10095 -380 10140 -360
rect 10095 -405 10105 -380
rect 10130 -405 10140 -380
rect 10095 -420 10140 -405
rect 10155 -335 10200 -320
rect 10155 -360 10165 -335
rect 10190 -360 10200 -335
rect 10155 -380 10200 -360
rect 10155 -405 10165 -380
rect 10190 -405 10200 -380
rect 10155 -420 10200 -405
rect 10215 -335 10260 -320
rect 10215 -360 10225 -335
rect 10250 -360 10260 -335
rect 10215 -380 10260 -360
rect 10215 -405 10225 -380
rect 10250 -405 10260 -380
rect 10215 -420 10260 -405
rect 10275 -335 10320 -320
rect 10275 -360 10285 -335
rect 10310 -360 10320 -335
rect 10275 -380 10320 -360
rect 10275 -405 10285 -380
rect 10310 -405 10320 -380
rect 10275 -420 10320 -405
rect 10335 -335 10380 -320
rect 10335 -360 10345 -335
rect 10370 -360 10380 -335
rect 10335 -380 10380 -360
rect 10335 -405 10345 -380
rect 10370 -405 10380 -380
rect 10335 -420 10380 -405
rect 10395 -335 10440 -320
rect 10395 -360 10405 -335
rect 10430 -360 10440 -335
rect 10395 -380 10440 -360
rect 10395 -405 10405 -380
rect 10430 -405 10440 -380
rect 10395 -420 10440 -405
rect 10455 -335 10500 -320
rect 10455 -360 10465 -335
rect 10490 -360 10500 -335
rect 10455 -380 10500 -360
rect 10455 -405 10465 -380
rect 10490 -405 10500 -380
rect 10455 -420 10500 -405
rect 10515 -335 10560 -320
rect 10515 -360 10525 -335
rect 10550 -360 10560 -335
rect 10515 -380 10560 -360
rect 10515 -405 10525 -380
rect 10550 -405 10560 -380
rect 10515 -420 10560 -405
rect 10575 -335 10620 -320
rect 10575 -360 10585 -335
rect 10610 -360 10620 -335
rect 10575 -380 10620 -360
rect 10575 -405 10585 -380
rect 10610 -405 10620 -380
rect 10575 -420 10620 -405
rect 10635 -335 10680 -320
rect 10635 -360 10645 -335
rect 10670 -360 10680 -335
rect 10635 -380 10680 -360
rect 10635 -405 10645 -380
rect 10670 -405 10680 -380
rect 10635 -420 10680 -405
rect 10695 -335 10740 -320
rect 10695 -360 10705 -335
rect 10730 -360 10740 -335
rect 10695 -380 10740 -360
rect 10695 -405 10705 -380
rect 10730 -405 10740 -380
rect 10695 -420 10740 -405
rect 10755 -335 10800 -320
rect 10755 -360 10765 -335
rect 10790 -360 10800 -335
rect 10755 -380 10800 -360
rect 10755 -405 10765 -380
rect 10790 -405 10800 -380
rect 10755 -420 10800 -405
rect 10815 -335 10860 -320
rect 10815 -360 10825 -335
rect 10850 -360 10860 -335
rect 10815 -380 10860 -360
rect 10815 -405 10825 -380
rect 10850 -405 10860 -380
rect 10815 -420 10860 -405
rect 10875 -335 10920 -320
rect 10875 -360 10885 -335
rect 10910 -360 10920 -335
rect 10875 -380 10920 -360
rect 10875 -405 10885 -380
rect 10910 -405 10920 -380
rect 10875 -420 10920 -405
rect 10935 -335 10980 -320
rect 10935 -360 10945 -335
rect 10970 -360 10980 -335
rect 10935 -380 10980 -360
rect 10935 -405 10945 -380
rect 10970 -405 10980 -380
rect 10935 -420 10980 -405
rect 10995 -335 11040 -320
rect 10995 -360 11005 -335
rect 11030 -360 11040 -335
rect 10995 -380 11040 -360
rect 10995 -405 11005 -380
rect 11030 -405 11040 -380
rect 10995 -420 11040 -405
rect 11055 -335 11100 -320
rect 11055 -360 11065 -335
rect 11090 -360 11100 -335
rect 11055 -380 11100 -360
rect 11055 -405 11065 -380
rect 11090 -405 11100 -380
rect 11055 -420 11100 -405
rect 11115 -335 11160 -320
rect 11115 -360 11125 -335
rect 11150 -360 11160 -335
rect 11115 -380 11160 -360
rect 11115 -405 11125 -380
rect 11150 -405 11160 -380
rect 11115 -420 11160 -405
rect 11175 -335 11220 -320
rect 11175 -360 11185 -335
rect 11210 -360 11220 -335
rect 11175 -380 11220 -360
rect 11175 -405 11185 -380
rect 11210 -405 11220 -380
rect 11175 -420 11220 -405
rect 11235 -335 11280 -320
rect 11235 -360 11245 -335
rect 11270 -360 11280 -335
rect 11235 -380 11280 -360
rect 11235 -405 11245 -380
rect 11270 -405 11280 -380
rect 11235 -420 11280 -405
rect 11295 -335 11340 -320
rect 11295 -360 11305 -335
rect 11330 -360 11340 -335
rect 11295 -380 11340 -360
rect 11295 -405 11305 -380
rect 11330 -405 11340 -380
rect 11295 -420 11340 -405
rect 11355 -335 11400 -320
rect 11355 -360 11365 -335
rect 11390 -360 11400 -335
rect 11355 -380 11400 -360
rect 11355 -405 11365 -380
rect 11390 -405 11400 -380
rect 11355 -420 11400 -405
rect 11415 -335 11460 -320
rect 11415 -360 11425 -335
rect 11450 -360 11460 -335
rect 11415 -380 11460 -360
rect 11415 -405 11425 -380
rect 11450 -405 11460 -380
rect 11415 -420 11460 -405
rect 11475 -335 11520 -320
rect 11475 -360 11485 -335
rect 11510 -360 11520 -335
rect 11475 -380 11520 -360
rect 11475 -405 11485 -380
rect 11510 -405 11520 -380
rect 11475 -420 11520 -405
rect 11535 -335 11580 -320
rect 11535 -360 11545 -335
rect 11570 -360 11580 -335
rect 11535 -380 11580 -360
rect 11535 -405 11545 -380
rect 11570 -405 11580 -380
rect 11535 -420 11580 -405
rect 11595 -335 11640 -320
rect 11595 -360 11605 -335
rect 11630 -360 11640 -335
rect 11595 -380 11640 -360
rect 11595 -405 11605 -380
rect 11630 -405 11640 -380
rect 11595 -420 11640 -405
rect 11655 -335 11700 -320
rect 11655 -360 11665 -335
rect 11690 -360 11700 -335
rect 11655 -380 11700 -360
rect 11655 -405 11665 -380
rect 11690 -405 11700 -380
rect 11655 -420 11700 -405
rect 11715 -335 11760 -320
rect 11715 -360 11725 -335
rect 11750 -360 11760 -335
rect 11715 -380 11760 -360
rect 11715 -405 11725 -380
rect 11750 -405 11760 -380
rect 11715 -420 11760 -405
rect 11775 -335 11820 -320
rect 11775 -360 11785 -335
rect 11810 -360 11820 -335
rect 11775 -380 11820 -360
rect 11775 -405 11785 -380
rect 11810 -405 11820 -380
rect 11775 -420 11820 -405
rect 11835 -335 11880 -320
rect 11835 -360 11845 -335
rect 11870 -360 11880 -335
rect 11835 -380 11880 -360
rect 11835 -405 11845 -380
rect 11870 -405 11880 -380
rect 11835 -420 11880 -405
rect 11895 -335 11940 -320
rect 11895 -360 11905 -335
rect 11930 -360 11940 -335
rect 11895 -380 11940 -360
rect 11895 -405 11905 -380
rect 11930 -405 11940 -380
rect 11895 -420 11940 -405
rect 11955 -335 12000 -320
rect 11955 -360 11965 -335
rect 11990 -360 12000 -335
rect 11955 -380 12000 -360
rect 11955 -405 11965 -380
rect 11990 -405 12000 -380
rect 11955 -420 12000 -405
rect 12015 -335 12060 -320
rect 12015 -360 12025 -335
rect 12050 -360 12060 -335
rect 12015 -380 12060 -360
rect 12015 -405 12025 -380
rect 12050 -405 12060 -380
rect 12015 -420 12060 -405
rect 12075 -335 12120 -320
rect 12075 -360 12085 -335
rect 12110 -360 12120 -335
rect 12075 -380 12120 -360
rect 12075 -405 12085 -380
rect 12110 -405 12120 -380
rect 12075 -420 12120 -405
rect 12135 -335 12180 -320
rect 12135 -360 12145 -335
rect 12170 -360 12180 -335
rect 12135 -380 12180 -360
rect 12135 -405 12145 -380
rect 12170 -405 12180 -380
rect 12135 -420 12180 -405
rect 12195 -335 12240 -320
rect 12195 -360 12205 -335
rect 12230 -360 12240 -335
rect 12195 -380 12240 -360
rect 12195 -405 12205 -380
rect 12230 -405 12240 -380
rect 12195 -420 12240 -405
rect 12255 -335 12300 -320
rect 12255 -360 12265 -335
rect 12290 -360 12300 -335
rect 12255 -380 12300 -360
rect 12255 -405 12265 -380
rect 12290 -405 12300 -380
rect 12255 -420 12300 -405
rect 12315 -335 12360 -320
rect 12315 -360 12325 -335
rect 12350 -360 12360 -335
rect 12315 -380 12360 -360
rect 12315 -405 12325 -380
rect 12350 -405 12360 -380
rect 12315 -420 12360 -405
rect 12375 -335 12420 -320
rect 12375 -360 12385 -335
rect 12410 -360 12420 -335
rect 12375 -380 12420 -360
rect 12375 -405 12385 -380
rect 12410 -405 12420 -380
rect 12375 -420 12420 -405
rect 12435 -335 12480 -320
rect 12435 -360 12445 -335
rect 12470 -360 12480 -335
rect 12435 -380 12480 -360
rect 12435 -405 12445 -380
rect 12470 -405 12480 -380
rect 12435 -420 12480 -405
rect 12495 -335 12540 -320
rect 12495 -360 12505 -335
rect 12530 -360 12540 -335
rect 12495 -380 12540 -360
rect 12495 -405 12505 -380
rect 12530 -405 12540 -380
rect 12495 -420 12540 -405
rect 12555 -335 12600 -320
rect 12555 -360 12565 -335
rect 12590 -360 12600 -335
rect 12555 -380 12600 -360
rect 12555 -405 12565 -380
rect 12590 -405 12600 -380
rect 12555 -420 12600 -405
rect 12615 -335 12660 -320
rect 12615 -360 12625 -335
rect 12650 -360 12660 -335
rect 12615 -380 12660 -360
rect 12615 -405 12625 -380
rect 12650 -405 12660 -380
rect 12615 -420 12660 -405
rect 12675 -335 12720 -320
rect 12675 -360 12685 -335
rect 12710 -360 12720 -335
rect 12675 -380 12720 -360
rect 12675 -405 12685 -380
rect 12710 -405 12720 -380
rect 12675 -420 12720 -405
rect 12735 -335 12780 -320
rect 12735 -360 12745 -335
rect 12770 -360 12780 -335
rect 12735 -380 12780 -360
rect 12735 -405 12745 -380
rect 12770 -405 12780 -380
rect 12735 -420 12780 -405
rect 12795 -335 12840 -320
rect 12795 -360 12805 -335
rect 12830 -360 12840 -335
rect 12795 -380 12840 -360
rect 12795 -405 12805 -380
rect 12830 -405 12840 -380
rect 12795 -420 12840 -405
rect 12855 -335 12900 -320
rect 12855 -360 12865 -335
rect 12890 -360 12900 -335
rect 12855 -380 12900 -360
rect 12855 -405 12865 -380
rect 12890 -405 12900 -380
rect 12855 -420 12900 -405
rect 12915 -335 12960 -320
rect 12915 -360 12925 -335
rect 12950 -360 12960 -335
rect 12915 -380 12960 -360
rect 12915 -405 12925 -380
rect 12950 -405 12960 -380
rect 12915 -420 12960 -405
rect 12975 -335 13020 -320
rect 12975 -360 12985 -335
rect 13010 -360 13020 -335
rect 12975 -380 13020 -360
rect 12975 -405 12985 -380
rect 13010 -405 13020 -380
rect 12975 -420 13020 -405
rect 13035 -335 13080 -320
rect 13035 -360 13045 -335
rect 13070 -360 13080 -335
rect 13035 -380 13080 -360
rect 13035 -405 13045 -380
rect 13070 -405 13080 -380
rect 13035 -420 13080 -405
rect 13095 -335 13140 -320
rect 13095 -360 13105 -335
rect 13130 -360 13140 -335
rect 13095 -380 13140 -360
rect 13095 -405 13105 -380
rect 13130 -405 13140 -380
rect 13095 -420 13140 -405
rect 13155 -335 13200 -320
rect 13155 -360 13165 -335
rect 13190 -360 13200 -335
rect 13155 -380 13200 -360
rect 13155 -405 13165 -380
rect 13190 -405 13200 -380
rect 13155 -420 13200 -405
rect 13215 -335 13260 -320
rect 13215 -360 13225 -335
rect 13250 -360 13260 -335
rect 13215 -380 13260 -360
rect 13215 -405 13225 -380
rect 13250 -405 13260 -380
rect 13215 -420 13260 -405
rect 13275 -335 13320 -320
rect 13275 -360 13285 -335
rect 13310 -360 13320 -335
rect 13275 -380 13320 -360
rect 13275 -405 13285 -380
rect 13310 -405 13320 -380
rect 13275 -420 13320 -405
rect 13335 -335 13380 -320
rect 13335 -360 13345 -335
rect 13370 -360 13380 -335
rect 13335 -380 13380 -360
rect 13335 -405 13345 -380
rect 13370 -405 13380 -380
rect 13335 -420 13380 -405
rect 13395 -335 13440 -320
rect 13395 -360 13405 -335
rect 13430 -360 13440 -335
rect 13395 -380 13440 -360
rect 13395 -405 13405 -380
rect 13430 -405 13440 -380
rect 13395 -420 13440 -405
rect 13455 -335 13500 -320
rect 13455 -360 13465 -335
rect 13490 -360 13500 -335
rect 13455 -380 13500 -360
rect 13455 -405 13465 -380
rect 13490 -405 13500 -380
rect 13455 -420 13500 -405
rect 13515 -335 13560 -320
rect 13515 -360 13525 -335
rect 13550 -360 13560 -335
rect 13515 -380 13560 -360
rect 13515 -405 13525 -380
rect 13550 -405 13560 -380
rect 13515 -420 13560 -405
rect 13575 -335 13620 -320
rect 13575 -360 13585 -335
rect 13610 -360 13620 -335
rect 13575 -380 13620 -360
rect 13575 -405 13585 -380
rect 13610 -405 13620 -380
rect 13575 -420 13620 -405
rect 13635 -335 13680 -320
rect 13635 -360 13645 -335
rect 13670 -360 13680 -335
rect 13635 -380 13680 -360
rect 13635 -405 13645 -380
rect 13670 -405 13680 -380
rect 13635 -420 13680 -405
rect 13695 -335 13740 -320
rect 13695 -360 13705 -335
rect 13730 -360 13740 -335
rect 13695 -380 13740 -360
rect 13695 -405 13705 -380
rect 13730 -405 13740 -380
rect 13695 -420 13740 -405
rect 13755 -335 13800 -320
rect 13755 -360 13765 -335
rect 13790 -360 13800 -335
rect 13755 -380 13800 -360
rect 13755 -405 13765 -380
rect 13790 -405 13800 -380
rect 13755 -420 13800 -405
rect 13815 -335 13860 -320
rect 13815 -360 13825 -335
rect 13850 -360 13860 -335
rect 13815 -380 13860 -360
rect 13815 -405 13825 -380
rect 13850 -405 13860 -380
rect 13815 -420 13860 -405
rect 13875 -335 13920 -320
rect 13875 -360 13885 -335
rect 13910 -360 13920 -335
rect 13875 -380 13920 -360
rect 13875 -405 13885 -380
rect 13910 -405 13920 -380
rect 13875 -420 13920 -405
rect 13935 -335 13980 -320
rect 13935 -360 13945 -335
rect 13970 -360 13980 -335
rect 13935 -380 13980 -360
rect 13935 -405 13945 -380
rect 13970 -405 13980 -380
rect 13935 -420 13980 -405
rect 13995 -335 14040 -320
rect 13995 -360 14005 -335
rect 14030 -360 14040 -335
rect 13995 -380 14040 -360
rect 13995 -405 14005 -380
rect 14030 -405 14040 -380
rect 13995 -420 14040 -405
rect 14055 -335 14100 -320
rect 14055 -360 14065 -335
rect 14090 -360 14100 -335
rect 14055 -380 14100 -360
rect 14055 -405 14065 -380
rect 14090 -405 14100 -380
rect 14055 -420 14100 -405
rect 14115 -335 14160 -320
rect 14115 -360 14125 -335
rect 14150 -360 14160 -335
rect 14115 -380 14160 -360
rect 14115 -405 14125 -380
rect 14150 -405 14160 -380
rect 14115 -420 14160 -405
rect 14175 -335 14220 -320
rect 14175 -360 14185 -335
rect 14210 -360 14220 -335
rect 14175 -380 14220 -360
rect 14175 -405 14185 -380
rect 14210 -405 14220 -380
rect 14175 -420 14220 -405
rect 14235 -335 14280 -320
rect 14235 -360 14245 -335
rect 14270 -360 14280 -335
rect 14235 -380 14280 -360
rect 14235 -405 14245 -380
rect 14270 -405 14280 -380
rect 14235 -420 14280 -405
rect 14295 -335 14340 -320
rect 14295 -360 14305 -335
rect 14330 -360 14340 -335
rect 14295 -380 14340 -360
rect 14295 -405 14305 -380
rect 14330 -405 14340 -380
rect 14295 -420 14340 -405
rect 14355 -335 14400 -320
rect 14355 -360 14365 -335
rect 14390 -360 14400 -335
rect 14355 -380 14400 -360
rect 14355 -405 14365 -380
rect 14390 -405 14400 -380
rect 14355 -420 14400 -405
rect 14415 -335 14460 -320
rect 14415 -360 14425 -335
rect 14450 -360 14460 -335
rect 14415 -380 14460 -360
rect 14415 -405 14425 -380
rect 14450 -405 14460 -380
rect 14415 -420 14460 -405
rect 14475 -335 14520 -320
rect 14475 -360 14485 -335
rect 14510 -360 14520 -335
rect 14475 -380 14520 -360
rect 14475 -405 14485 -380
rect 14510 -405 14520 -380
rect 14475 -420 14520 -405
rect 14535 -335 14580 -320
rect 14535 -360 14545 -335
rect 14570 -360 14580 -335
rect 14535 -380 14580 -360
rect 14535 -405 14545 -380
rect 14570 -405 14580 -380
rect 14535 -420 14580 -405
rect 14595 -335 14640 -320
rect 14595 -360 14605 -335
rect 14630 -360 14640 -335
rect 14595 -380 14640 -360
rect 14595 -405 14605 -380
rect 14630 -405 14640 -380
rect 14595 -420 14640 -405
rect 14655 -335 14700 -320
rect 14655 -360 14665 -335
rect 14690 -360 14700 -335
rect 14655 -380 14700 -360
rect 14655 -405 14665 -380
rect 14690 -405 14700 -380
rect 14655 -420 14700 -405
rect 14715 -335 14760 -320
rect 14715 -360 14725 -335
rect 14750 -360 14760 -335
rect 14715 -380 14760 -360
rect 14715 -405 14725 -380
rect 14750 -405 14760 -380
rect 14715 -420 14760 -405
rect 14775 -335 14820 -320
rect 14775 -360 14785 -335
rect 14810 -360 14820 -335
rect 14775 -380 14820 -360
rect 14775 -405 14785 -380
rect 14810 -405 14820 -380
rect 14775 -420 14820 -405
rect 14835 -335 14880 -320
rect 14835 -360 14845 -335
rect 14870 -360 14880 -335
rect 14835 -380 14880 -360
rect 14835 -405 14845 -380
rect 14870 -405 14880 -380
rect 14835 -420 14880 -405
rect 14895 -335 14940 -320
rect 14895 -360 14905 -335
rect 14930 -360 14940 -335
rect 14895 -380 14940 -360
rect 14895 -405 14905 -380
rect 14930 -405 14940 -380
rect 14895 -420 14940 -405
rect 14955 -335 15000 -320
rect 14955 -360 14965 -335
rect 14990 -360 15000 -335
rect 14955 -380 15000 -360
rect 14955 -405 14965 -380
rect 14990 -405 15000 -380
rect 14955 -420 15000 -405
rect 15015 -335 15060 -320
rect 15015 -360 15025 -335
rect 15050 -360 15060 -335
rect 15015 -380 15060 -360
rect 15015 -405 15025 -380
rect 15050 -405 15060 -380
rect 15015 -420 15060 -405
rect 15075 -335 15120 -320
rect 15075 -360 15085 -335
rect 15110 -360 15120 -335
rect 15075 -380 15120 -360
rect 15075 -405 15085 -380
rect 15110 -405 15120 -380
rect 15075 -420 15120 -405
rect 15135 -335 15180 -320
rect 15135 -360 15145 -335
rect 15170 -360 15180 -335
rect 15135 -380 15180 -360
rect 15135 -405 15145 -380
rect 15170 -405 15180 -380
rect 15135 -420 15180 -405
rect 15195 -335 15240 -320
rect 15195 -360 15205 -335
rect 15230 -360 15240 -335
rect 15195 -380 15240 -360
rect 15195 -405 15205 -380
rect 15230 -405 15240 -380
rect 15195 -420 15240 -405
rect 15255 -335 15300 -320
rect 15255 -360 15265 -335
rect 15290 -360 15300 -335
rect 15255 -380 15300 -360
rect 15255 -405 15265 -380
rect 15290 -405 15300 -380
rect 15255 -420 15300 -405
rect 15315 -335 15360 -320
rect 15315 -360 15325 -335
rect 15350 -360 15360 -335
rect 15315 -380 15360 -360
rect 15315 -405 15325 -380
rect 15350 -405 15360 -380
rect 15315 -420 15360 -405
rect 15375 -335 15420 -320
rect 15375 -360 15385 -335
rect 15410 -360 15420 -335
rect 15375 -380 15420 -360
rect 15375 -405 15385 -380
rect 15410 -405 15420 -380
rect 15375 -420 15420 -405
rect 15435 -335 15480 -320
rect 15435 -360 15445 -335
rect 15470 -360 15480 -335
rect 15435 -380 15480 -360
rect 15435 -405 15445 -380
rect 15470 -405 15480 -380
rect 15435 -420 15480 -405
rect 15495 -335 15540 -320
rect 15495 -360 15505 -335
rect 15530 -360 15540 -335
rect 15495 -380 15540 -360
rect 15495 -405 15505 -380
rect 15530 -405 15540 -380
rect 15495 -420 15540 -405
rect 15555 -335 15600 -320
rect 15555 -360 15565 -335
rect 15590 -360 15600 -335
rect 15555 -380 15600 -360
rect 15555 -405 15565 -380
rect 15590 -405 15600 -380
rect 15555 -420 15600 -405
rect 15615 -335 15660 -320
rect 15615 -360 15625 -335
rect 15650 -360 15660 -335
rect 15615 -380 15660 -360
rect 15615 -405 15625 -380
rect 15650 -405 15660 -380
rect 15615 -420 15660 -405
rect 15675 -335 15720 -320
rect 15675 -360 15685 -335
rect 15710 -360 15720 -335
rect 15675 -380 15720 -360
rect 15675 -405 15685 -380
rect 15710 -405 15720 -380
rect 15675 -420 15720 -405
rect 15735 -335 15780 -320
rect 15735 -360 15745 -335
rect 15770 -360 15780 -335
rect 15735 -380 15780 -360
rect 15735 -405 15745 -380
rect 15770 -405 15780 -380
rect 15735 -420 15780 -405
rect 15795 -335 15840 -320
rect 15795 -360 15805 -335
rect 15830 -360 15840 -335
rect 15795 -380 15840 -360
rect 15795 -405 15805 -380
rect 15830 -405 15840 -380
rect 15795 -420 15840 -405
rect 15855 -335 15900 -320
rect 15855 -360 15865 -335
rect 15890 -360 15900 -335
rect 15855 -380 15900 -360
rect 15855 -405 15865 -380
rect 15890 -405 15900 -380
rect 15855 -420 15900 -405
rect 15915 -335 15960 -320
rect 15915 -360 15925 -335
rect 15950 -360 15960 -335
rect 15915 -380 15960 -360
rect 15915 -405 15925 -380
rect 15950 -405 15960 -380
rect 15915 -420 15960 -405
rect 15975 -335 16020 -320
rect 15975 -360 15985 -335
rect 16010 -360 16020 -335
rect 15975 -380 16020 -360
rect 15975 -405 15985 -380
rect 16010 -405 16020 -380
rect 15975 -420 16020 -405
rect 16035 -335 16080 -320
rect 16035 -360 16045 -335
rect 16070 -360 16080 -335
rect 16035 -380 16080 -360
rect 16035 -405 16045 -380
rect 16070 -405 16080 -380
rect 16035 -420 16080 -405
rect 16095 -335 16140 -320
rect 16095 -360 16105 -335
rect 16130 -360 16140 -335
rect 16095 -380 16140 -360
rect 16095 -405 16105 -380
rect 16130 -405 16140 -380
rect 16095 -420 16140 -405
rect 16155 -335 16200 -320
rect 16155 -360 16165 -335
rect 16190 -360 16200 -335
rect 16155 -380 16200 -360
rect 16155 -405 16165 -380
rect 16190 -405 16200 -380
rect 16155 -420 16200 -405
rect 16215 -335 16260 -320
rect 16215 -360 16225 -335
rect 16250 -360 16260 -335
rect 16215 -380 16260 -360
rect 16215 -405 16225 -380
rect 16250 -405 16260 -380
rect 16215 -420 16260 -405
rect 16275 -335 16320 -320
rect 16275 -360 16285 -335
rect 16310 -360 16320 -335
rect 16275 -380 16320 -360
rect 16275 -405 16285 -380
rect 16310 -405 16320 -380
rect 16275 -420 16320 -405
rect 16335 -335 16380 -320
rect 16335 -360 16345 -335
rect 16370 -360 16380 -335
rect 16335 -380 16380 -360
rect 16335 -405 16345 -380
rect 16370 -405 16380 -380
rect 16335 -420 16380 -405
rect 16395 -335 16440 -320
rect 16395 -360 16405 -335
rect 16430 -360 16440 -335
rect 16395 -380 16440 -360
rect 16395 -405 16405 -380
rect 16430 -405 16440 -380
rect 16395 -420 16440 -405
rect 16455 -335 16500 -320
rect 16455 -360 16465 -335
rect 16490 -360 16500 -335
rect 16455 -380 16500 -360
rect 16455 -405 16465 -380
rect 16490 -405 16500 -380
rect 16455 -420 16500 -405
rect 16515 -335 16560 -320
rect 16515 -360 16525 -335
rect 16550 -360 16560 -335
rect 16515 -380 16560 -360
rect 16515 -405 16525 -380
rect 16550 -405 16560 -380
rect 16515 -420 16560 -405
rect 16575 -335 16620 -320
rect 16575 -360 16585 -335
rect 16610 -360 16620 -335
rect 16575 -380 16620 -360
rect 16575 -405 16585 -380
rect 16610 -405 16620 -380
rect 16575 -420 16620 -405
rect 16635 -335 16680 -320
rect 16635 -360 16645 -335
rect 16670 -360 16680 -335
rect 16635 -380 16680 -360
rect 16635 -405 16645 -380
rect 16670 -405 16680 -380
rect 16635 -420 16680 -405
rect 16695 -335 16740 -320
rect 16695 -360 16705 -335
rect 16730 -360 16740 -335
rect 16695 -380 16740 -360
rect 16695 -405 16705 -380
rect 16730 -405 16740 -380
rect 16695 -420 16740 -405
rect 16755 -335 16800 -320
rect 16755 -360 16765 -335
rect 16790 -360 16800 -335
rect 16755 -380 16800 -360
rect 16755 -405 16765 -380
rect 16790 -405 16800 -380
rect 16755 -420 16800 -405
rect 16815 -335 16860 -320
rect 16815 -360 16825 -335
rect 16850 -360 16860 -335
rect 16815 -380 16860 -360
rect 16815 -405 16825 -380
rect 16850 -405 16860 -380
rect 16815 -420 16860 -405
rect 16875 -335 16920 -320
rect 16875 -360 16885 -335
rect 16910 -360 16920 -335
rect 16875 -380 16920 -360
rect 16875 -405 16885 -380
rect 16910 -405 16920 -380
rect 16875 -420 16920 -405
rect 16935 -335 16980 -320
rect 16935 -360 16945 -335
rect 16970 -360 16980 -335
rect 16935 -380 16980 -360
rect 16935 -405 16945 -380
rect 16970 -405 16980 -380
rect 16935 -420 16980 -405
rect 16995 -335 17040 -320
rect 16995 -360 17005 -335
rect 17030 -360 17040 -335
rect 16995 -380 17040 -360
rect 16995 -405 17005 -380
rect 17030 -405 17040 -380
rect 16995 -420 17040 -405
rect 17055 -335 17100 -320
rect 17055 -360 17065 -335
rect 17090 -360 17100 -335
rect 17055 -380 17100 -360
rect 17055 -405 17065 -380
rect 17090 -405 17100 -380
rect 17055 -420 17100 -405
rect 17115 -335 17160 -320
rect 17115 -360 17125 -335
rect 17150 -360 17160 -335
rect 17115 -380 17160 -360
rect 17115 -405 17125 -380
rect 17150 -405 17160 -380
rect 17115 -420 17160 -405
rect 17175 -335 17220 -320
rect 17175 -360 17185 -335
rect 17210 -360 17220 -335
rect 17175 -380 17220 -360
rect 17175 -405 17185 -380
rect 17210 -405 17220 -380
rect 17175 -420 17220 -405
rect 17235 -335 17280 -320
rect 17235 -360 17245 -335
rect 17270 -360 17280 -335
rect 17235 -380 17280 -360
rect 17235 -405 17245 -380
rect 17270 -405 17280 -380
rect 17235 -420 17280 -405
rect 17295 -335 17340 -320
rect 17295 -360 17305 -335
rect 17330 -360 17340 -335
rect 17295 -380 17340 -360
rect 17295 -405 17305 -380
rect 17330 -405 17340 -380
rect 17295 -420 17340 -405
rect 17355 -335 17400 -320
rect 17355 -360 17365 -335
rect 17390 -360 17400 -335
rect 17355 -380 17400 -360
rect 17355 -405 17365 -380
rect 17390 -405 17400 -380
rect 17355 -420 17400 -405
rect 17415 -335 17460 -320
rect 17415 -360 17425 -335
rect 17450 -360 17460 -335
rect 17415 -380 17460 -360
rect 17415 -405 17425 -380
rect 17450 -405 17460 -380
rect 17415 -420 17460 -405
rect 17475 -335 17520 -320
rect 17475 -360 17485 -335
rect 17510 -360 17520 -335
rect 17475 -380 17520 -360
rect 17475 -405 17485 -380
rect 17510 -405 17520 -380
rect 17475 -420 17520 -405
rect 17535 -335 17580 -320
rect 17535 -360 17545 -335
rect 17570 -360 17580 -335
rect 17535 -380 17580 -360
rect 17535 -405 17545 -380
rect 17570 -405 17580 -380
rect 17535 -420 17580 -405
rect 17595 -335 17640 -320
rect 17595 -360 17605 -335
rect 17630 -360 17640 -335
rect 17595 -380 17640 -360
rect 17595 -405 17605 -380
rect 17630 -405 17640 -380
rect 17595 -420 17640 -405
rect 17655 -335 17700 -320
rect 17655 -360 17665 -335
rect 17690 -360 17700 -335
rect 17655 -380 17700 -360
rect 17655 -405 17665 -380
rect 17690 -405 17700 -380
rect 17655 -420 17700 -405
rect 17715 -335 17760 -320
rect 17715 -360 17725 -335
rect 17750 -360 17760 -335
rect 17715 -380 17760 -360
rect 17715 -405 17725 -380
rect 17750 -405 17760 -380
rect 17715 -420 17760 -405
rect 17775 -335 17820 -320
rect 17775 -360 17785 -335
rect 17810 -360 17820 -335
rect 17775 -380 17820 -360
rect 17775 -405 17785 -380
rect 17810 -405 17820 -380
rect 17775 -420 17820 -405
rect 17835 -335 17880 -320
rect 17835 -360 17845 -335
rect 17870 -360 17880 -335
rect 17835 -380 17880 -360
rect 17835 -405 17845 -380
rect 17870 -405 17880 -380
rect 17835 -420 17880 -405
rect 17895 -335 17940 -320
rect 17895 -360 17905 -335
rect 17930 -360 17940 -335
rect 17895 -380 17940 -360
rect 17895 -405 17905 -380
rect 17930 -405 17940 -380
rect 17895 -420 17940 -405
rect 17955 -335 18000 -320
rect 17955 -360 17965 -335
rect 17990 -360 18000 -335
rect 17955 -380 18000 -360
rect 17955 -405 17965 -380
rect 17990 -405 18000 -380
rect 17955 -420 18000 -405
rect 18015 -335 18060 -320
rect 18015 -360 18025 -335
rect 18050 -360 18060 -335
rect 18015 -380 18060 -360
rect 18015 -405 18025 -380
rect 18050 -405 18060 -380
rect 18015 -420 18060 -405
rect 18075 -335 18120 -320
rect 18075 -360 18085 -335
rect 18110 -360 18120 -335
rect 18075 -380 18120 -360
rect 18075 -405 18085 -380
rect 18110 -405 18120 -380
rect 18075 -420 18120 -405
rect 18135 -335 18180 -320
rect 18135 -360 18145 -335
rect 18170 -360 18180 -335
rect 18135 -380 18180 -360
rect 18135 -405 18145 -380
rect 18170 -405 18180 -380
rect 18135 -420 18180 -405
rect 18195 -335 18240 -320
rect 18195 -360 18205 -335
rect 18230 -360 18240 -335
rect 18195 -380 18240 -360
rect 18195 -405 18205 -380
rect 18230 -405 18240 -380
rect 18195 -420 18240 -405
rect 18255 -335 18300 -320
rect 18255 -360 18265 -335
rect 18290 -360 18300 -335
rect 18255 -380 18300 -360
rect 18255 -405 18265 -380
rect 18290 -405 18300 -380
rect 18255 -420 18300 -405
rect 18315 -335 18360 -320
rect 18315 -360 18325 -335
rect 18350 -360 18360 -335
rect 18315 -380 18360 -360
rect 18315 -405 18325 -380
rect 18350 -405 18360 -380
rect 18315 -420 18360 -405
rect 18375 -335 18420 -320
rect 18375 -360 18385 -335
rect 18410 -360 18420 -335
rect 18375 -380 18420 -360
rect 18375 -405 18385 -380
rect 18410 -405 18420 -380
rect 18375 -420 18420 -405
rect 18435 -335 18480 -320
rect 18435 -360 18445 -335
rect 18470 -360 18480 -335
rect 18435 -380 18480 -360
rect 18435 -405 18445 -380
rect 18470 -405 18480 -380
rect 18435 -420 18480 -405
rect 18495 -335 18540 -320
rect 18495 -360 18505 -335
rect 18530 -360 18540 -335
rect 18495 -380 18540 -360
rect 18495 -405 18505 -380
rect 18530 -405 18540 -380
rect 18495 -420 18540 -405
rect 18555 -335 18600 -320
rect 18555 -360 18565 -335
rect 18590 -360 18600 -335
rect 18555 -380 18600 -360
rect 18555 -405 18565 -380
rect 18590 -405 18600 -380
rect 18555 -420 18600 -405
rect 18615 -335 18660 -320
rect 18615 -360 18625 -335
rect 18650 -360 18660 -335
rect 18615 -380 18660 -360
rect 18615 -405 18625 -380
rect 18650 -405 18660 -380
rect 18615 -420 18660 -405
rect 18675 -335 18720 -320
rect 18675 -360 18685 -335
rect 18710 -360 18720 -335
rect 18675 -380 18720 -360
rect 18675 -405 18685 -380
rect 18710 -405 18720 -380
rect 18675 -420 18720 -405
rect 18735 -335 18780 -320
rect 18735 -360 18745 -335
rect 18770 -360 18780 -335
rect 18735 -380 18780 -360
rect 18735 -405 18745 -380
rect 18770 -405 18780 -380
rect 18735 -420 18780 -405
rect 18795 -335 18840 -320
rect 18795 -360 18805 -335
rect 18830 -360 18840 -335
rect 18795 -380 18840 -360
rect 18795 -405 18805 -380
rect 18830 -405 18840 -380
rect 18795 -420 18840 -405
rect 18855 -335 18900 -320
rect 18855 -360 18865 -335
rect 18890 -360 18900 -335
rect 18855 -380 18900 -360
rect 18855 -405 18865 -380
rect 18890 -405 18900 -380
rect 18855 -420 18900 -405
rect 18915 -335 18960 -320
rect 18915 -360 18925 -335
rect 18950 -360 18960 -335
rect 18915 -380 18960 -360
rect 18915 -405 18925 -380
rect 18950 -405 18960 -380
rect 18915 -420 18960 -405
rect 18975 -335 19020 -320
rect 18975 -360 18985 -335
rect 19010 -360 19020 -335
rect 18975 -380 19020 -360
rect 18975 -405 18985 -380
rect 19010 -405 19020 -380
rect 18975 -420 19020 -405
rect 19035 -335 19080 -320
rect 19035 -360 19045 -335
rect 19070 -360 19080 -335
rect 19035 -380 19080 -360
rect 19035 -405 19045 -380
rect 19070 -405 19080 -380
rect 19035 -420 19080 -405
rect 19095 -335 19140 -320
rect 19095 -360 19105 -335
rect 19130 -360 19140 -335
rect 19095 -380 19140 -360
rect 19095 -405 19105 -380
rect 19130 -405 19140 -380
rect 19095 -420 19140 -405
rect 19155 -335 19200 -320
rect 19155 -360 19165 -335
rect 19190 -360 19200 -335
rect 19155 -380 19200 -360
rect 19155 -405 19165 -380
rect 19190 -405 19200 -380
rect 19155 -420 19200 -405
rect 19215 -335 19260 -320
rect 19215 -360 19225 -335
rect 19250 -360 19260 -335
rect 19215 -380 19260 -360
rect 19215 -405 19225 -380
rect 19250 -405 19260 -380
rect 19215 -420 19260 -405
rect 19275 -335 19320 -320
rect 19275 -360 19285 -335
rect 19310 -360 19320 -335
rect 19275 -380 19320 -360
rect 19275 -405 19285 -380
rect 19310 -405 19320 -380
rect 19275 -420 19320 -405
rect 19335 -335 19380 -320
rect 19335 -360 19345 -335
rect 19370 -360 19380 -335
rect 19335 -380 19380 -360
rect 19335 -405 19345 -380
rect 19370 -405 19380 -380
rect 19335 -420 19380 -405
rect 19395 -335 19440 -320
rect 19395 -360 19405 -335
rect 19430 -360 19440 -335
rect 19395 -380 19440 -360
rect 19395 -405 19405 -380
rect 19430 -405 19440 -380
rect 19395 -420 19440 -405
rect 19455 -335 19500 -320
rect 19455 -360 19465 -335
rect 19490 -360 19500 -335
rect 19455 -380 19500 -360
rect 19455 -405 19465 -380
rect 19490 -405 19500 -380
rect 19455 -420 19500 -405
rect 19515 -335 19560 -320
rect 19515 -360 19525 -335
rect 19550 -360 19560 -335
rect 19515 -380 19560 -360
rect 19515 -405 19525 -380
rect 19550 -405 19560 -380
rect 19515 -420 19560 -405
rect 19575 -335 19620 -320
rect 19575 -360 19585 -335
rect 19610 -360 19620 -335
rect 19575 -380 19620 -360
rect 19575 -405 19585 -380
rect 19610 -405 19620 -380
rect 19575 -420 19620 -405
rect 19635 -335 19680 -320
rect 19635 -360 19645 -335
rect 19670 -360 19680 -335
rect 19635 -380 19680 -360
rect 19635 -405 19645 -380
rect 19670 -405 19680 -380
rect 19635 -420 19680 -405
rect 19695 -335 19740 -320
rect 19695 -360 19705 -335
rect 19730 -360 19740 -335
rect 19695 -380 19740 -360
rect 19695 -405 19705 -380
rect 19730 -405 19740 -380
rect 19695 -420 19740 -405
rect 19755 -335 19800 -320
rect 19755 -360 19765 -335
rect 19790 -360 19800 -335
rect 19755 -380 19800 -360
rect 19755 -405 19765 -380
rect 19790 -405 19800 -380
rect 19755 -420 19800 -405
rect 19815 -335 19860 -320
rect 19815 -360 19825 -335
rect 19850 -360 19860 -335
rect 19815 -380 19860 -360
rect 19815 -405 19825 -380
rect 19850 -405 19860 -380
rect 19815 -420 19860 -405
rect 19875 -335 19920 -320
rect 19875 -360 19885 -335
rect 19910 -360 19920 -335
rect 19875 -380 19920 -360
rect 19875 -405 19885 -380
rect 19910 -405 19920 -380
rect 19875 -420 19920 -405
rect 19935 -335 19980 -320
rect 19935 -360 19945 -335
rect 19970 -360 19980 -335
rect 19935 -380 19980 -360
rect 19935 -405 19945 -380
rect 19970 -405 19980 -380
rect 19935 -420 19980 -405
rect 19995 -335 20040 -320
rect 19995 -360 20005 -335
rect 20030 -360 20040 -335
rect 19995 -380 20040 -360
rect 19995 -405 20005 -380
rect 20030 -405 20040 -380
rect 19995 -420 20040 -405
rect 20055 -335 20100 -320
rect 20055 -360 20065 -335
rect 20090 -360 20100 -335
rect 20055 -380 20100 -360
rect 20055 -405 20065 -380
rect 20090 -405 20100 -380
rect 20055 -420 20100 -405
rect 20115 -335 20160 -320
rect 20115 -360 20125 -335
rect 20150 -360 20160 -335
rect 20115 -380 20160 -360
rect 20115 -405 20125 -380
rect 20150 -405 20160 -380
rect 20115 -420 20160 -405
rect 20175 -335 20220 -320
rect 20175 -360 20185 -335
rect 20210 -360 20220 -335
rect 20175 -380 20220 -360
rect 20175 -405 20185 -380
rect 20210 -405 20220 -380
rect 20175 -420 20220 -405
rect 20235 -335 20280 -320
rect 20235 -360 20245 -335
rect 20270 -360 20280 -335
rect 20235 -380 20280 -360
rect 20235 -405 20245 -380
rect 20270 -405 20280 -380
rect 20235 -420 20280 -405
rect 20295 -335 20340 -320
rect 20295 -360 20305 -335
rect 20330 -360 20340 -335
rect 20295 -380 20340 -360
rect 20295 -405 20305 -380
rect 20330 -405 20340 -380
rect 20295 -420 20340 -405
rect 20355 -335 20400 -320
rect 20355 -360 20365 -335
rect 20390 -360 20400 -335
rect 20355 -380 20400 -360
rect 20355 -405 20365 -380
rect 20390 -405 20400 -380
rect 20355 -420 20400 -405
rect 20415 -335 20460 -320
rect 20415 -360 20425 -335
rect 20450 -360 20460 -335
rect 20415 -380 20460 -360
rect 20415 -405 20425 -380
rect 20450 -405 20460 -380
rect 20415 -420 20460 -405
rect 20475 -335 20520 -320
rect 20475 -360 20485 -335
rect 20510 -360 20520 -335
rect 20475 -380 20520 -360
rect 20475 -405 20485 -380
rect 20510 -405 20520 -380
rect 20475 -420 20520 -405
rect 20535 -335 20580 -320
rect 20535 -360 20545 -335
rect 20570 -360 20580 -335
rect 20535 -380 20580 -360
rect 20535 -405 20545 -380
rect 20570 -405 20580 -380
rect 20535 -420 20580 -405
rect 20595 -335 20640 -320
rect 20595 -360 20605 -335
rect 20630 -360 20640 -335
rect 20595 -380 20640 -360
rect 20595 -405 20605 -380
rect 20630 -405 20640 -380
rect 20595 -420 20640 -405
rect 20655 -335 20700 -320
rect 20655 -360 20665 -335
rect 20690 -360 20700 -335
rect 20655 -380 20700 -360
rect 20655 -405 20665 -380
rect 20690 -405 20700 -380
rect 20655 -420 20700 -405
rect 20715 -335 20760 -320
rect 20715 -360 20725 -335
rect 20750 -360 20760 -335
rect 20715 -380 20760 -360
rect 20715 -405 20725 -380
rect 20750 -405 20760 -380
rect 20715 -420 20760 -405
rect 20775 -335 20820 -320
rect 20775 -360 20785 -335
rect 20810 -360 20820 -335
rect 20775 -380 20820 -360
rect 20775 -405 20785 -380
rect 20810 -405 20820 -380
rect 20775 -420 20820 -405
rect 20835 -335 20880 -320
rect 20835 -360 20845 -335
rect 20870 -360 20880 -335
rect 20835 -380 20880 -360
rect 20835 -405 20845 -380
rect 20870 -405 20880 -380
rect 20835 -420 20880 -405
rect 20895 -335 20940 -320
rect 20895 -360 20905 -335
rect 20930 -360 20940 -335
rect 20895 -380 20940 -360
rect 20895 -405 20905 -380
rect 20930 -405 20940 -380
rect 20895 -420 20940 -405
rect 20955 -335 21000 -320
rect 20955 -360 20965 -335
rect 20990 -360 21000 -335
rect 20955 -380 21000 -360
rect 20955 -405 20965 -380
rect 20990 -405 21000 -380
rect 20955 -420 21000 -405
rect 21015 -335 21060 -320
rect 21015 -360 21025 -335
rect 21050 -360 21060 -335
rect 21015 -380 21060 -360
rect 21015 -405 21025 -380
rect 21050 -405 21060 -380
rect 21015 -420 21060 -405
rect 21075 -335 21120 -320
rect 21075 -360 21085 -335
rect 21110 -360 21120 -335
rect 21075 -380 21120 -360
rect 21075 -405 21085 -380
rect 21110 -405 21120 -380
rect 21075 -420 21120 -405
rect 21135 -335 21180 -320
rect 21135 -360 21145 -335
rect 21170 -360 21180 -335
rect 21135 -380 21180 -360
rect 21135 -405 21145 -380
rect 21170 -405 21180 -380
rect 21135 -420 21180 -405
rect 21195 -335 21240 -320
rect 21195 -360 21205 -335
rect 21230 -360 21240 -335
rect 21195 -380 21240 -360
rect 21195 -405 21205 -380
rect 21230 -405 21240 -380
rect 21195 -420 21240 -405
rect 21255 -335 21300 -320
rect 21255 -360 21265 -335
rect 21290 -360 21300 -335
rect 21255 -380 21300 -360
rect 21255 -405 21265 -380
rect 21290 -405 21300 -380
rect 21255 -420 21300 -405
rect 21315 -335 21360 -320
rect 21315 -360 21325 -335
rect 21350 -360 21360 -335
rect 21315 -380 21360 -360
rect 21315 -405 21325 -380
rect 21350 -405 21360 -380
rect 21315 -420 21360 -405
rect 21375 -335 21420 -320
rect 21375 -360 21385 -335
rect 21410 -360 21420 -335
rect 21375 -380 21420 -360
rect 21375 -405 21385 -380
rect 21410 -405 21420 -380
rect 21375 -420 21420 -405
rect 21435 -335 21480 -320
rect 21435 -360 21445 -335
rect 21470 -360 21480 -335
rect 21435 -380 21480 -360
rect 21435 -405 21445 -380
rect 21470 -405 21480 -380
rect 21435 -420 21480 -405
rect 21495 -335 21540 -320
rect 21495 -360 21505 -335
rect 21530 -360 21540 -335
rect 21495 -380 21540 -360
rect 21495 -405 21505 -380
rect 21530 -405 21540 -380
rect 21495 -420 21540 -405
rect 21555 -335 21600 -320
rect 21555 -360 21565 -335
rect 21590 -360 21600 -335
rect 21555 -380 21600 -360
rect 21555 -405 21565 -380
rect 21590 -405 21600 -380
rect 21555 -420 21600 -405
rect 21615 -335 21660 -320
rect 21615 -360 21625 -335
rect 21650 -360 21660 -335
rect 21615 -380 21660 -360
rect 21615 -405 21625 -380
rect 21650 -405 21660 -380
rect 21615 -420 21660 -405
rect 21675 -335 21720 -320
rect 21675 -360 21685 -335
rect 21710 -360 21720 -335
rect 21675 -380 21720 -360
rect 21675 -405 21685 -380
rect 21710 -405 21720 -380
rect 21675 -420 21720 -405
rect 21735 -335 21780 -320
rect 21735 -360 21745 -335
rect 21770 -360 21780 -335
rect 21735 -380 21780 -360
rect 21735 -405 21745 -380
rect 21770 -405 21780 -380
rect 21735 -420 21780 -405
rect 21795 -335 21840 -320
rect 21795 -360 21805 -335
rect 21830 -360 21840 -335
rect 21795 -380 21840 -360
rect 21795 -405 21805 -380
rect 21830 -405 21840 -380
rect 21795 -420 21840 -405
rect 21855 -335 21900 -320
rect 21855 -360 21865 -335
rect 21890 -360 21900 -335
rect 21855 -380 21900 -360
rect 21855 -405 21865 -380
rect 21890 -405 21900 -380
rect 21855 -420 21900 -405
rect 21915 -335 21960 -320
rect 21915 -360 21925 -335
rect 21950 -360 21960 -335
rect 21915 -380 21960 -360
rect 21915 -405 21925 -380
rect 21950 -405 21960 -380
rect 21915 -420 21960 -405
rect 21975 -335 22020 -320
rect 21975 -360 21985 -335
rect 22010 -360 22020 -335
rect 21975 -380 22020 -360
rect 21975 -405 21985 -380
rect 22010 -405 22020 -380
rect 21975 -420 22020 -405
rect 22035 -335 22080 -320
rect 22035 -360 22045 -335
rect 22070 -360 22080 -335
rect 22035 -380 22080 -360
rect 22035 -405 22045 -380
rect 22070 -405 22080 -380
rect 22035 -420 22080 -405
rect 22095 -335 22140 -320
rect 22095 -360 22105 -335
rect 22130 -360 22140 -335
rect 22095 -380 22140 -360
rect 22095 -405 22105 -380
rect 22130 -405 22140 -380
rect 22095 -420 22140 -405
rect 22155 -335 22200 -320
rect 22155 -360 22165 -335
rect 22190 -360 22200 -335
rect 22155 -380 22200 -360
rect 22155 -405 22165 -380
rect 22190 -405 22200 -380
rect 22155 -420 22200 -405
rect 22215 -335 22260 -320
rect 22215 -360 22225 -335
rect 22250 -360 22260 -335
rect 22215 -380 22260 -360
rect 22215 -405 22225 -380
rect 22250 -405 22260 -380
rect 22215 -420 22260 -405
rect 22275 -335 22320 -320
rect 22275 -360 22285 -335
rect 22310 -360 22320 -335
rect 22275 -380 22320 -360
rect 22275 -405 22285 -380
rect 22310 -405 22320 -380
rect 22275 -420 22320 -405
rect 22335 -335 22380 -320
rect 22335 -360 22345 -335
rect 22370 -360 22380 -335
rect 22335 -380 22380 -360
rect 22335 -405 22345 -380
rect 22370 -405 22380 -380
rect 22335 -420 22380 -405
rect 22395 -335 22440 -320
rect 22395 -360 22405 -335
rect 22430 -360 22440 -335
rect 22395 -380 22440 -360
rect 22395 -405 22405 -380
rect 22430 -405 22440 -380
rect 22395 -420 22440 -405
rect 22455 -335 22500 -320
rect 22455 -360 22465 -335
rect 22490 -360 22500 -335
rect 22455 -380 22500 -360
rect 22455 -405 22465 -380
rect 22490 -405 22500 -380
rect 22455 -420 22500 -405
rect 22515 -335 22560 -320
rect 22515 -360 22525 -335
rect 22550 -360 22560 -335
rect 22515 -380 22560 -360
rect 22515 -405 22525 -380
rect 22550 -405 22560 -380
rect 22515 -420 22560 -405
rect 22575 -335 22620 -320
rect 22575 -360 22585 -335
rect 22610 -360 22620 -335
rect 22575 -380 22620 -360
rect 22575 -405 22585 -380
rect 22610 -405 22620 -380
rect 22575 -420 22620 -405
rect 22635 -335 22680 -320
rect 22635 -360 22645 -335
rect 22670 -360 22680 -335
rect 22635 -380 22680 -360
rect 22635 -405 22645 -380
rect 22670 -405 22680 -380
rect 22635 -420 22680 -405
rect 22695 -335 22740 -320
rect 22695 -360 22705 -335
rect 22730 -360 22740 -335
rect 22695 -380 22740 -360
rect 22695 -405 22705 -380
rect 22730 -405 22740 -380
rect 22695 -420 22740 -405
rect 22755 -335 22800 -320
rect 22755 -360 22765 -335
rect 22790 -360 22800 -335
rect 22755 -380 22800 -360
rect 22755 -405 22765 -380
rect 22790 -405 22800 -380
rect 22755 -420 22800 -405
rect 22815 -335 22860 -320
rect 22815 -360 22825 -335
rect 22850 -360 22860 -335
rect 22815 -380 22860 -360
rect 22815 -405 22825 -380
rect 22850 -405 22860 -380
rect 22815 -420 22860 -405
rect 22875 -335 22920 -320
rect 22875 -360 22885 -335
rect 22910 -360 22920 -335
rect 22875 -380 22920 -360
rect 22875 -405 22885 -380
rect 22910 -405 22920 -380
rect 22875 -420 22920 -405
rect 22935 -335 22980 -320
rect 22935 -360 22945 -335
rect 22970 -360 22980 -335
rect 22935 -380 22980 -360
rect 22935 -405 22945 -380
rect 22970 -405 22980 -380
rect 22935 -420 22980 -405
rect 22995 -335 23040 -320
rect 22995 -360 23005 -335
rect 23030 -360 23040 -335
rect 22995 -380 23040 -360
rect 22995 -405 23005 -380
rect 23030 -405 23040 -380
rect 22995 -420 23040 -405
rect 23055 -335 23100 -320
rect 23055 -360 23065 -335
rect 23090 -360 23100 -335
rect 23055 -380 23100 -360
rect 23055 -405 23065 -380
rect 23090 -405 23100 -380
rect 23055 -420 23100 -405
rect 23115 -335 23160 -320
rect 23115 -360 23125 -335
rect 23150 -360 23160 -335
rect 23115 -380 23160 -360
rect 23115 -405 23125 -380
rect 23150 -405 23160 -380
rect 23115 -420 23160 -405
rect 23175 -335 23220 -320
rect 23175 -360 23185 -335
rect 23210 -360 23220 -335
rect 23175 -380 23220 -360
rect 23175 -405 23185 -380
rect 23210 -405 23220 -380
rect 23175 -420 23220 -405
rect 23235 -335 23280 -320
rect 23235 -360 23245 -335
rect 23270 -360 23280 -335
rect 23235 -380 23280 -360
rect 23235 -405 23245 -380
rect 23270 -405 23280 -380
rect 23235 -420 23280 -405
rect 23295 -335 23340 -320
rect 23295 -360 23305 -335
rect 23330 -360 23340 -335
rect 23295 -380 23340 -360
rect 23295 -405 23305 -380
rect 23330 -405 23340 -380
rect 23295 -420 23340 -405
rect 23355 -335 23400 -320
rect 23355 -360 23365 -335
rect 23390 -360 23400 -335
rect 23355 -380 23400 -360
rect 23355 -405 23365 -380
rect 23390 -405 23400 -380
rect 23355 -420 23400 -405
rect 23415 -335 23460 -320
rect 23415 -360 23425 -335
rect 23450 -360 23460 -335
rect 23415 -380 23460 -360
rect 23415 -405 23425 -380
rect 23450 -405 23460 -380
rect 23415 -420 23460 -405
rect 23475 -335 23520 -320
rect 23475 -360 23485 -335
rect 23510 -360 23520 -335
rect 23475 -380 23520 -360
rect 23475 -405 23485 -380
rect 23510 -405 23520 -380
rect 23475 -420 23520 -405
rect 23535 -335 23580 -320
rect 23535 -360 23545 -335
rect 23570 -360 23580 -335
rect 23535 -380 23580 -360
rect 23535 -405 23545 -380
rect 23570 -405 23580 -380
rect 23535 -420 23580 -405
rect 23595 -335 23640 -320
rect 23595 -360 23605 -335
rect 23630 -360 23640 -335
rect 23595 -380 23640 -360
rect 23595 -405 23605 -380
rect 23630 -405 23640 -380
rect 23595 -420 23640 -405
rect 23655 -335 23700 -320
rect 23655 -360 23665 -335
rect 23690 -360 23700 -335
rect 23655 -380 23700 -360
rect 23655 -405 23665 -380
rect 23690 -405 23700 -380
rect 23655 -420 23700 -405
rect 23715 -335 23760 -320
rect 23715 -360 23725 -335
rect 23750 -360 23760 -335
rect 23715 -380 23760 -360
rect 23715 -405 23725 -380
rect 23750 -405 23760 -380
rect 23715 -420 23760 -405
rect 23775 -335 23820 -320
rect 23775 -360 23785 -335
rect 23810 -360 23820 -335
rect 23775 -380 23820 -360
rect 23775 -405 23785 -380
rect 23810 -405 23820 -380
rect 23775 -420 23820 -405
rect 23835 -335 23880 -320
rect 23835 -360 23845 -335
rect 23870 -360 23880 -335
rect 23835 -380 23880 -360
rect 23835 -405 23845 -380
rect 23870 -405 23880 -380
rect 23835 -420 23880 -405
rect 23895 -335 23940 -320
rect 23895 -360 23905 -335
rect 23930 -360 23940 -335
rect 23895 -380 23940 -360
rect 23895 -405 23905 -380
rect 23930 -405 23940 -380
rect 23895 -420 23940 -405
rect 23955 -335 24000 -320
rect 23955 -360 23965 -335
rect 23990 -360 24000 -335
rect 23955 -380 24000 -360
rect 23955 -405 23965 -380
rect 23990 -405 24000 -380
rect 23955 -420 24000 -405
rect 24015 -335 24060 -320
rect 24015 -360 24025 -335
rect 24050 -360 24060 -335
rect 24015 -380 24060 -360
rect 24015 -405 24025 -380
rect 24050 -405 24060 -380
rect 24015 -420 24060 -405
rect 24075 -335 24120 -320
rect 24075 -360 24085 -335
rect 24110 -360 24120 -335
rect 24075 -380 24120 -360
rect 24075 -405 24085 -380
rect 24110 -405 24120 -380
rect 24075 -420 24120 -405
rect 24135 -335 24180 -320
rect 24135 -360 24145 -335
rect 24170 -360 24180 -335
rect 24135 -380 24180 -360
rect 24135 -405 24145 -380
rect 24170 -405 24180 -380
rect 24135 -420 24180 -405
rect 24195 -335 24240 -320
rect 24195 -360 24205 -335
rect 24230 -360 24240 -335
rect 24195 -380 24240 -360
rect 24195 -405 24205 -380
rect 24230 -405 24240 -380
rect 24195 -420 24240 -405
rect 24255 -335 24300 -320
rect 24255 -360 24265 -335
rect 24290 -360 24300 -335
rect 24255 -380 24300 -360
rect 24255 -405 24265 -380
rect 24290 -405 24300 -380
rect 24255 -420 24300 -405
rect 24315 -335 24360 -320
rect 24315 -360 24325 -335
rect 24350 -360 24360 -335
rect 24315 -380 24360 -360
rect 24315 -405 24325 -380
rect 24350 -405 24360 -380
rect 24315 -420 24360 -405
rect 24375 -335 24420 -320
rect 24375 -360 24385 -335
rect 24410 -360 24420 -335
rect 24375 -380 24420 -360
rect 24375 -405 24385 -380
rect 24410 -405 24420 -380
rect 24375 -420 24420 -405
rect 24435 -335 24480 -320
rect 24435 -360 24445 -335
rect 24470 -360 24480 -335
rect 24435 -380 24480 -360
rect 24435 -405 24445 -380
rect 24470 -405 24480 -380
rect 24435 -420 24480 -405
rect 24495 -335 24540 -320
rect 24495 -360 24505 -335
rect 24530 -360 24540 -335
rect 24495 -380 24540 -360
rect 24495 -405 24505 -380
rect 24530 -405 24540 -380
rect 24495 -420 24540 -405
rect 24555 -335 24600 -320
rect 24555 -360 24565 -335
rect 24590 -360 24600 -335
rect 24555 -380 24600 -360
rect 24555 -405 24565 -380
rect 24590 -405 24600 -380
rect 24555 -420 24600 -405
rect 24615 -335 24660 -320
rect 24615 -360 24625 -335
rect 24650 -360 24660 -335
rect 24615 -380 24660 -360
rect 24615 -405 24625 -380
rect 24650 -405 24660 -380
rect 24615 -420 24660 -405
rect 24675 -335 24720 -320
rect 24675 -360 24685 -335
rect 24710 -360 24720 -335
rect 24675 -380 24720 -360
rect 24675 -405 24685 -380
rect 24710 -405 24720 -380
rect 24675 -420 24720 -405
rect 24735 -335 24780 -320
rect 24735 -360 24745 -335
rect 24770 -360 24780 -335
rect 24735 -380 24780 -360
rect 24735 -405 24745 -380
rect 24770 -405 24780 -380
rect 24735 -420 24780 -405
rect 24795 -335 24840 -320
rect 24795 -360 24805 -335
rect 24830 -360 24840 -335
rect 24795 -380 24840 -360
rect 24795 -405 24805 -380
rect 24830 -405 24840 -380
rect 24795 -420 24840 -405
rect 24855 -335 24900 -320
rect 24855 -360 24865 -335
rect 24890 -360 24900 -335
rect 24855 -380 24900 -360
rect 24855 -405 24865 -380
rect 24890 -405 24900 -380
rect 24855 -420 24900 -405
rect 24915 -335 24960 -320
rect 24915 -360 24925 -335
rect 24950 -360 24960 -335
rect 24915 -380 24960 -360
rect 24915 -405 24925 -380
rect 24950 -405 24960 -380
rect 24915 -420 24960 -405
rect 24975 -335 25020 -320
rect 24975 -360 24985 -335
rect 25010 -360 25020 -335
rect 24975 -380 25020 -360
rect 24975 -405 24985 -380
rect 25010 -405 25020 -380
rect 24975 -420 25020 -405
rect 25035 -335 25080 -320
rect 25035 -360 25045 -335
rect 25070 -360 25080 -335
rect 25035 -380 25080 -360
rect 25035 -405 25045 -380
rect 25070 -405 25080 -380
rect 25035 -420 25080 -405
rect 25095 -335 25140 -320
rect 25095 -360 25105 -335
rect 25130 -360 25140 -335
rect 25095 -380 25140 -360
rect 25095 -405 25105 -380
rect 25130 -405 25140 -380
rect 25095 -420 25140 -405
rect 25155 -335 25200 -320
rect 25155 -360 25165 -335
rect 25190 -360 25200 -335
rect 25155 -380 25200 -360
rect 25155 -405 25165 -380
rect 25190 -405 25200 -380
rect 25155 -420 25200 -405
rect 25215 -335 25260 -320
rect 25215 -360 25225 -335
rect 25250 -360 25260 -335
rect 25215 -380 25260 -360
rect 25215 -405 25225 -380
rect 25250 -405 25260 -380
rect 25215 -420 25260 -405
rect 25275 -335 25320 -320
rect 25275 -360 25285 -335
rect 25310 -360 25320 -335
rect 25275 -380 25320 -360
rect 25275 -405 25285 -380
rect 25310 -405 25320 -380
rect 25275 -420 25320 -405
rect 25335 -335 25380 -320
rect 25335 -360 25345 -335
rect 25370 -360 25380 -335
rect 25335 -380 25380 -360
rect 25335 -405 25345 -380
rect 25370 -405 25380 -380
rect 25335 -420 25380 -405
rect 25395 -335 25440 -320
rect 25395 -360 25405 -335
rect 25430 -360 25440 -335
rect 25395 -380 25440 -360
rect 25395 -405 25405 -380
rect 25430 -405 25440 -380
rect 25395 -420 25440 -405
rect 25455 -335 25500 -320
rect 25455 -360 25465 -335
rect 25490 -360 25500 -335
rect 25455 -380 25500 -360
rect 25455 -405 25465 -380
rect 25490 -405 25500 -380
rect 25455 -420 25500 -405
rect 25515 -335 25560 -320
rect 25515 -360 25525 -335
rect 25550 -360 25560 -335
rect 25515 -380 25560 -360
rect 25515 -405 25525 -380
rect 25550 -405 25560 -380
rect 25515 -420 25560 -405
rect 25575 -335 25620 -320
rect 25575 -360 25585 -335
rect 25610 -360 25620 -335
rect 25575 -380 25620 -360
rect 25575 -405 25585 -380
rect 25610 -405 25620 -380
rect 25575 -420 25620 -405
rect 25635 -335 25680 -320
rect 25635 -360 25645 -335
rect 25670 -360 25680 -335
rect 25635 -380 25680 -360
rect 25635 -405 25645 -380
rect 25670 -405 25680 -380
rect 25635 -420 25680 -405
rect 25695 -335 25740 -320
rect 25695 -360 25705 -335
rect 25730 -360 25740 -335
rect 25695 -380 25740 -360
rect 25695 -405 25705 -380
rect 25730 -405 25740 -380
rect 25695 -420 25740 -405
rect 25755 -335 25800 -320
rect 25755 -360 25765 -335
rect 25790 -360 25800 -335
rect 25755 -380 25800 -360
rect 25755 -405 25765 -380
rect 25790 -405 25800 -380
rect 25755 -420 25800 -405
rect 25815 -335 25860 -320
rect 25815 -360 25825 -335
rect 25850 -360 25860 -335
rect 25815 -380 25860 -360
rect 25815 -405 25825 -380
rect 25850 -405 25860 -380
rect 25815 -420 25860 -405
rect 25875 -335 25920 -320
rect 25875 -360 25885 -335
rect 25910 -360 25920 -335
rect 25875 -380 25920 -360
rect 25875 -405 25885 -380
rect 25910 -405 25920 -380
rect 25875 -420 25920 -405
rect 25935 -335 25980 -320
rect 25935 -360 25945 -335
rect 25970 -360 25980 -335
rect 25935 -380 25980 -360
rect 25935 -405 25945 -380
rect 25970 -405 25980 -380
rect 25935 -420 25980 -405
rect 25995 -335 26040 -320
rect 25995 -360 26005 -335
rect 26030 -360 26040 -335
rect 25995 -380 26040 -360
rect 25995 -405 26005 -380
rect 26030 -405 26040 -380
rect 25995 -420 26040 -405
rect 26055 -335 26100 -320
rect 26055 -360 26065 -335
rect 26090 -360 26100 -335
rect 26055 -380 26100 -360
rect 26055 -405 26065 -380
rect 26090 -405 26100 -380
rect 26055 -420 26100 -405
rect 26115 -335 26160 -320
rect 26115 -360 26125 -335
rect 26150 -360 26160 -335
rect 26115 -380 26160 -360
rect 26115 -405 26125 -380
rect 26150 -405 26160 -380
rect 26115 -420 26160 -405
rect 26175 -335 26220 -320
rect 26175 -360 26185 -335
rect 26210 -360 26220 -335
rect 26175 -380 26220 -360
rect 26175 -405 26185 -380
rect 26210 -405 26220 -380
rect 26175 -420 26220 -405
rect 26235 -335 26280 -320
rect 26235 -360 26245 -335
rect 26270 -360 26280 -335
rect 26235 -380 26280 -360
rect 26235 -405 26245 -380
rect 26270 -405 26280 -380
rect 26235 -420 26280 -405
rect 26295 -335 26340 -320
rect 26295 -360 26305 -335
rect 26330 -360 26340 -335
rect 26295 -380 26340 -360
rect 26295 -405 26305 -380
rect 26330 -405 26340 -380
rect 26295 -420 26340 -405
rect 26355 -335 26400 -320
rect 26355 -360 26365 -335
rect 26390 -360 26400 -335
rect 26355 -380 26400 -360
rect 26355 -405 26365 -380
rect 26390 -405 26400 -380
rect 26355 -420 26400 -405
rect 26415 -335 26460 -320
rect 26415 -360 26425 -335
rect 26450 -360 26460 -335
rect 26415 -380 26460 -360
rect 26415 -405 26425 -380
rect 26450 -405 26460 -380
rect 26415 -420 26460 -405
rect 26475 -335 26520 -320
rect 26475 -360 26485 -335
rect 26510 -360 26520 -335
rect 26475 -380 26520 -360
rect 26475 -405 26485 -380
rect 26510 -405 26520 -380
rect 26475 -420 26520 -405
rect 26535 -335 26580 -320
rect 26535 -360 26545 -335
rect 26570 -360 26580 -335
rect 26535 -380 26580 -360
rect 26535 -405 26545 -380
rect 26570 -405 26580 -380
rect 26535 -420 26580 -405
rect 26595 -335 26640 -320
rect 26595 -360 26605 -335
rect 26630 -360 26640 -335
rect 26595 -380 26640 -360
rect 26595 -405 26605 -380
rect 26630 -405 26640 -380
rect 26595 -420 26640 -405
rect 26655 -335 26700 -320
rect 26655 -360 26665 -335
rect 26690 -360 26700 -335
rect 26655 -380 26700 -360
rect 26655 -405 26665 -380
rect 26690 -405 26700 -380
rect 26655 -420 26700 -405
rect 26715 -335 26760 -320
rect 26715 -360 26725 -335
rect 26750 -360 26760 -335
rect 26715 -380 26760 -360
rect 26715 -405 26725 -380
rect 26750 -405 26760 -380
rect 26715 -420 26760 -405
rect 26775 -335 26820 -320
rect 26775 -360 26785 -335
rect 26810 -360 26820 -335
rect 26775 -380 26820 -360
rect 26775 -405 26785 -380
rect 26810 -405 26820 -380
rect 26775 -420 26820 -405
rect 26835 -335 26880 -320
rect 26835 -360 26845 -335
rect 26870 -360 26880 -335
rect 26835 -380 26880 -360
rect 26835 -405 26845 -380
rect 26870 -405 26880 -380
rect 26835 -420 26880 -405
rect 26895 -335 26940 -320
rect 26895 -360 26905 -335
rect 26930 -360 26940 -335
rect 26895 -380 26940 -360
rect 26895 -405 26905 -380
rect 26930 -405 26940 -380
rect 26895 -420 26940 -405
rect 26955 -335 27000 -320
rect 26955 -360 26965 -335
rect 26990 -360 27000 -335
rect 26955 -380 27000 -360
rect 26955 -405 26965 -380
rect 26990 -405 27000 -380
rect 26955 -420 27000 -405
rect 27015 -335 27060 -320
rect 27015 -360 27025 -335
rect 27050 -360 27060 -335
rect 27015 -380 27060 -360
rect 27015 -405 27025 -380
rect 27050 -405 27060 -380
rect 27015 -420 27060 -405
rect 27075 -335 27120 -320
rect 27075 -360 27085 -335
rect 27110 -360 27120 -335
rect 27075 -380 27120 -360
rect 27075 -405 27085 -380
rect 27110 -405 27120 -380
rect 27075 -420 27120 -405
rect 27135 -335 27180 -320
rect 27135 -360 27145 -335
rect 27170 -360 27180 -335
rect 27135 -380 27180 -360
rect 27135 -405 27145 -380
rect 27170 -405 27180 -380
rect 27135 -420 27180 -405
rect 27195 -335 27240 -320
rect 27195 -360 27205 -335
rect 27230 -360 27240 -335
rect 27195 -380 27240 -360
rect 27195 -405 27205 -380
rect 27230 -405 27240 -380
rect 27195 -420 27240 -405
rect 27255 -335 27300 -320
rect 27255 -360 27265 -335
rect 27290 -360 27300 -335
rect 27255 -380 27300 -360
rect 27255 -405 27265 -380
rect 27290 -405 27300 -380
rect 27255 -420 27300 -405
rect 27315 -335 27360 -320
rect 27315 -360 27325 -335
rect 27350 -360 27360 -335
rect 27315 -380 27360 -360
rect 27315 -405 27325 -380
rect 27350 -405 27360 -380
rect 27315 -420 27360 -405
rect 27375 -335 27420 -320
rect 27375 -360 27385 -335
rect 27410 -360 27420 -335
rect 27375 -380 27420 -360
rect 27375 -405 27385 -380
rect 27410 -405 27420 -380
rect 27375 -420 27420 -405
rect 27435 -335 27480 -320
rect 27435 -360 27445 -335
rect 27470 -360 27480 -335
rect 27435 -380 27480 -360
rect 27435 -405 27445 -380
rect 27470 -405 27480 -380
rect 27435 -420 27480 -405
rect 27495 -335 27540 -320
rect 27495 -360 27505 -335
rect 27530 -360 27540 -335
rect 27495 -380 27540 -360
rect 27495 -405 27505 -380
rect 27530 -405 27540 -380
rect 27495 -420 27540 -405
rect 27555 -335 27600 -320
rect 27555 -360 27565 -335
rect 27590 -360 27600 -335
rect 27555 -380 27600 -360
rect 27555 -405 27565 -380
rect 27590 -405 27600 -380
rect 27555 -420 27600 -405
rect 27615 -335 27660 -320
rect 27615 -360 27625 -335
rect 27650 -360 27660 -335
rect 27615 -380 27660 -360
rect 27615 -405 27625 -380
rect 27650 -405 27660 -380
rect 27615 -420 27660 -405
rect 27675 -335 27720 -320
rect 27675 -360 27685 -335
rect 27710 -360 27720 -335
rect 27675 -380 27720 -360
rect 27675 -405 27685 -380
rect 27710 -405 27720 -380
rect 27675 -420 27720 -405
rect 27735 -335 27780 -320
rect 27735 -360 27745 -335
rect 27770 -360 27780 -335
rect 27735 -380 27780 -360
rect 27735 -405 27745 -380
rect 27770 -405 27780 -380
rect 27735 -420 27780 -405
rect 27795 -335 27840 -320
rect 27795 -360 27805 -335
rect 27830 -360 27840 -335
rect 27795 -380 27840 -360
rect 27795 -405 27805 -380
rect 27830 -405 27840 -380
rect 27795 -420 27840 -405
rect 27855 -335 27900 -320
rect 27855 -360 27865 -335
rect 27890 -360 27900 -335
rect 27855 -380 27900 -360
rect 27855 -405 27865 -380
rect 27890 -405 27900 -380
rect 27855 -420 27900 -405
rect 27915 -335 27960 -320
rect 27915 -360 27925 -335
rect 27950 -360 27960 -335
rect 27915 -380 27960 -360
rect 27915 -405 27925 -380
rect 27950 -405 27960 -380
rect 27915 -420 27960 -405
rect 27975 -335 28020 -320
rect 27975 -360 27985 -335
rect 28010 -360 28020 -335
rect 27975 -380 28020 -360
rect 27975 -405 27985 -380
rect 28010 -405 28020 -380
rect 27975 -420 28020 -405
rect 28035 -335 28080 -320
rect 28035 -360 28045 -335
rect 28070 -360 28080 -335
rect 28035 -380 28080 -360
rect 28035 -405 28045 -380
rect 28070 -405 28080 -380
rect 28035 -420 28080 -405
rect 28095 -335 28140 -320
rect 28095 -360 28105 -335
rect 28130 -360 28140 -335
rect 28095 -380 28140 -360
rect 28095 -405 28105 -380
rect 28130 -405 28140 -380
rect 28095 -420 28140 -405
rect 28155 -335 28200 -320
rect 28155 -360 28165 -335
rect 28190 -360 28200 -335
rect 28155 -380 28200 -360
rect 28155 -405 28165 -380
rect 28190 -405 28200 -380
rect 28155 -420 28200 -405
rect 28215 -335 28260 -320
rect 28215 -360 28225 -335
rect 28250 -360 28260 -335
rect 28215 -380 28260 -360
rect 28215 -405 28225 -380
rect 28250 -405 28260 -380
rect 28215 -420 28260 -405
rect 28275 -335 28320 -320
rect 28275 -360 28285 -335
rect 28310 -360 28320 -335
rect 28275 -380 28320 -360
rect 28275 -405 28285 -380
rect 28310 -405 28320 -380
rect 28275 -420 28320 -405
rect 28335 -335 28380 -320
rect 28335 -360 28345 -335
rect 28370 -360 28380 -335
rect 28335 -380 28380 -360
rect 28335 -405 28345 -380
rect 28370 -405 28380 -380
rect 28335 -420 28380 -405
rect 28395 -335 28440 -320
rect 28395 -360 28405 -335
rect 28430 -360 28440 -335
rect 28395 -380 28440 -360
rect 28395 -405 28405 -380
rect 28430 -405 28440 -380
rect 28395 -420 28440 -405
rect 28455 -335 28500 -320
rect 28455 -360 28465 -335
rect 28490 -360 28500 -335
rect 28455 -380 28500 -360
rect 28455 -405 28465 -380
rect 28490 -405 28500 -380
rect 28455 -420 28500 -405
rect 28515 -335 28560 -320
rect 28515 -360 28525 -335
rect 28550 -360 28560 -335
rect 28515 -380 28560 -360
rect 28515 -405 28525 -380
rect 28550 -405 28560 -380
rect 28515 -420 28560 -405
rect 28575 -335 28620 -320
rect 28575 -360 28585 -335
rect 28610 -360 28620 -335
rect 28575 -380 28620 -360
rect 28575 -405 28585 -380
rect 28610 -405 28620 -380
rect 28575 -420 28620 -405
rect 28635 -335 28680 -320
rect 28635 -360 28645 -335
rect 28670 -360 28680 -335
rect 28635 -380 28680 -360
rect 28635 -405 28645 -380
rect 28670 -405 28680 -380
rect 28635 -420 28680 -405
rect 28695 -335 28740 -320
rect 28695 -360 28705 -335
rect 28730 -360 28740 -335
rect 28695 -380 28740 -360
rect 28695 -405 28705 -380
rect 28730 -405 28740 -380
rect 28695 -420 28740 -405
rect 28755 -335 28800 -320
rect 28755 -360 28765 -335
rect 28790 -360 28800 -335
rect 28755 -380 28800 -360
rect 28755 -405 28765 -380
rect 28790 -405 28800 -380
rect 28755 -420 28800 -405
rect 28815 -335 28860 -320
rect 28815 -360 28825 -335
rect 28850 -360 28860 -335
rect 28815 -380 28860 -360
rect 28815 -405 28825 -380
rect 28850 -405 28860 -380
rect 28815 -420 28860 -405
rect 28875 -335 28920 -320
rect 28875 -360 28885 -335
rect 28910 -360 28920 -335
rect 28875 -380 28920 -360
rect 28875 -405 28885 -380
rect 28910 -405 28920 -380
rect 28875 -420 28920 -405
rect 28935 -335 28980 -320
rect 28935 -360 28945 -335
rect 28970 -360 28980 -335
rect 28935 -380 28980 -360
rect 28935 -405 28945 -380
rect 28970 -405 28980 -380
rect 28935 -420 28980 -405
rect 28995 -335 29040 -320
rect 28995 -360 29005 -335
rect 29030 -360 29040 -335
rect 28995 -380 29040 -360
rect 28995 -405 29005 -380
rect 29030 -405 29040 -380
rect 28995 -420 29040 -405
rect 29055 -335 29100 -320
rect 29055 -360 29065 -335
rect 29090 -360 29100 -335
rect 29055 -380 29100 -360
rect 29055 -405 29065 -380
rect 29090 -405 29100 -380
rect 29055 -420 29100 -405
rect 29115 -335 29160 -320
rect 29115 -360 29125 -335
rect 29150 -360 29160 -335
rect 29115 -380 29160 -360
rect 29115 -405 29125 -380
rect 29150 -405 29160 -380
rect 29115 -420 29160 -405
rect 29175 -335 29220 -320
rect 29175 -360 29185 -335
rect 29210 -360 29220 -335
rect 29175 -380 29220 -360
rect 29175 -405 29185 -380
rect 29210 -405 29220 -380
rect 29175 -420 29220 -405
rect 29235 -335 29280 -320
rect 29235 -360 29245 -335
rect 29270 -360 29280 -335
rect 29235 -380 29280 -360
rect 29235 -405 29245 -380
rect 29270 -405 29280 -380
rect 29235 -420 29280 -405
rect 29295 -335 29340 -320
rect 29295 -360 29305 -335
rect 29330 -360 29340 -335
rect 29295 -380 29340 -360
rect 29295 -405 29305 -380
rect 29330 -405 29340 -380
rect 29295 -420 29340 -405
rect 29355 -335 29400 -320
rect 29355 -360 29365 -335
rect 29390 -360 29400 -335
rect 29355 -380 29400 -360
rect 29355 -405 29365 -380
rect 29390 -405 29400 -380
rect 29355 -420 29400 -405
rect 29415 -335 29460 -320
rect 29415 -360 29425 -335
rect 29450 -360 29460 -335
rect 29415 -380 29460 -360
rect 29415 -405 29425 -380
rect 29450 -405 29460 -380
rect 29415 -420 29460 -405
rect 29475 -335 29520 -320
rect 29475 -360 29485 -335
rect 29510 -360 29520 -335
rect 29475 -380 29520 -360
rect 29475 -405 29485 -380
rect 29510 -405 29520 -380
rect 29475 -420 29520 -405
rect 29535 -335 29580 -320
rect 29535 -360 29545 -335
rect 29570 -360 29580 -335
rect 29535 -380 29580 -360
rect 29535 -405 29545 -380
rect 29570 -405 29580 -380
rect 29535 -420 29580 -405
rect 29595 -335 29640 -320
rect 29595 -360 29605 -335
rect 29630 -360 29640 -335
rect 29595 -380 29640 -360
rect 29595 -405 29605 -380
rect 29630 -405 29640 -380
rect 29595 -420 29640 -405
rect 29655 -335 29700 -320
rect 29655 -360 29665 -335
rect 29690 -360 29700 -335
rect 29655 -380 29700 -360
rect 29655 -405 29665 -380
rect 29690 -405 29700 -380
rect 29655 -420 29700 -405
rect 29715 -335 29760 -320
rect 29715 -360 29725 -335
rect 29750 -360 29760 -335
rect 29715 -380 29760 -360
rect 29715 -405 29725 -380
rect 29750 -405 29760 -380
rect 29715 -420 29760 -405
rect 29775 -335 29820 -320
rect 29775 -360 29785 -335
rect 29810 -360 29820 -335
rect 29775 -380 29820 -360
rect 29775 -405 29785 -380
rect 29810 -405 29820 -380
rect 29775 -420 29820 -405
rect 29835 -335 29880 -320
rect 29835 -360 29845 -335
rect 29870 -360 29880 -335
rect 29835 -380 29880 -360
rect 29835 -405 29845 -380
rect 29870 -405 29880 -380
rect 29835 -420 29880 -405
rect 29895 -335 29940 -320
rect 29895 -360 29905 -335
rect 29930 -360 29940 -335
rect 29895 -380 29940 -360
rect 29895 -405 29905 -380
rect 29930 -405 29940 -380
rect 29895 -420 29940 -405
rect 29955 -335 30000 -320
rect 29955 -360 29965 -335
rect 29990 -360 30000 -335
rect 29955 -380 30000 -360
rect 29955 -405 29965 -380
rect 29990 -405 30000 -380
rect 29955 -420 30000 -405
rect 30015 -335 30060 -320
rect 30015 -360 30025 -335
rect 30050 -360 30060 -335
rect 30015 -380 30060 -360
rect 30015 -405 30025 -380
rect 30050 -405 30060 -380
rect 30015 -420 30060 -405
rect 30075 -335 30120 -320
rect 30075 -360 30085 -335
rect 30110 -360 30120 -335
rect 30075 -380 30120 -360
rect 30075 -405 30085 -380
rect 30110 -405 30120 -380
rect 30075 -420 30120 -405
rect 30135 -335 30180 -320
rect 30135 -360 30145 -335
rect 30170 -360 30180 -335
rect 30135 -380 30180 -360
rect 30135 -405 30145 -380
rect 30170 -405 30180 -380
rect 30135 -420 30180 -405
rect 30195 -335 30240 -320
rect 30195 -360 30205 -335
rect 30230 -360 30240 -335
rect 30195 -380 30240 -360
rect 30195 -405 30205 -380
rect 30230 -405 30240 -380
rect 30195 -420 30240 -405
rect 30255 -335 30300 -320
rect 30255 -360 30265 -335
rect 30290 -360 30300 -335
rect 30255 -380 30300 -360
rect 30255 -405 30265 -380
rect 30290 -405 30300 -380
rect 30255 -420 30300 -405
rect 30315 -335 30360 -320
rect 30315 -360 30325 -335
rect 30350 -360 30360 -335
rect 30315 -380 30360 -360
rect 30315 -405 30325 -380
rect 30350 -405 30360 -380
rect 30315 -420 30360 -405
rect 30375 -335 30420 -320
rect 30375 -360 30385 -335
rect 30410 -360 30420 -335
rect 30375 -380 30420 -360
rect 30375 -405 30385 -380
rect 30410 -405 30420 -380
rect 30375 -420 30420 -405
rect 30435 -335 30480 -320
rect 30435 -360 30445 -335
rect 30470 -360 30480 -335
rect 30435 -380 30480 -360
rect 30435 -405 30445 -380
rect 30470 -405 30480 -380
rect 30435 -420 30480 -405
rect 30495 -335 30540 -320
rect 30495 -360 30505 -335
rect 30530 -360 30540 -335
rect 30495 -380 30540 -360
rect 30495 -405 30505 -380
rect 30530 -405 30540 -380
rect 30495 -420 30540 -405
rect 30555 -335 30600 -320
rect 30555 -360 30565 -335
rect 30590 -360 30600 -335
rect 30555 -380 30600 -360
rect 30555 -405 30565 -380
rect 30590 -405 30600 -380
rect 30555 -420 30600 -405
rect 30615 -335 30660 -320
rect 30615 -360 30625 -335
rect 30650 -360 30660 -335
rect 30615 -380 30660 -360
rect 30615 -405 30625 -380
rect 30650 -405 30660 -380
rect 30615 -420 30660 -405
rect 30675 -335 30715 -320
rect 30675 -360 30685 -335
rect 30710 -360 30715 -335
rect 30675 -380 30715 -360
rect 30675 -405 30685 -380
rect 30710 -405 30715 -380
rect 30675 -420 30715 -405
<< pdiff >>
rect 436 265 476 275
rect 436 240 441 265
rect 466 240 476 265
rect 436 225 476 240
rect 741 265 781 275
rect 741 240 746 265
rect 771 240 781 265
rect 741 225 781 240
rect 986 265 1026 275
rect 986 240 991 265
rect 1016 240 1026 265
rect 986 225 1026 240
rect 1226 265 1266 275
rect 1226 240 1231 265
rect 1256 240 1266 265
rect 1226 225 1266 240
rect 1471 265 1511 275
rect 1471 240 1476 265
rect 1501 240 1511 265
rect 1471 225 1511 240
rect 1776 265 1816 275
rect 1776 240 1781 265
rect 1806 240 1816 265
rect 1776 225 1816 240
rect 2021 265 2061 275
rect 2021 240 2026 265
rect 2051 240 2061 265
rect 2506 265 2546 275
rect 2021 225 2061 240
rect 2506 240 2511 265
rect 2536 240 2546 265
rect 2506 225 2546 240
rect 2746 265 2786 275
rect 2746 240 2751 265
rect 2776 240 2786 265
rect 2746 225 2786 240
rect 2991 265 3031 275
rect 2991 240 2996 265
rect 3021 240 3031 265
rect 2991 225 3031 240
rect 3231 265 3271 275
rect 3231 240 3236 265
rect 3261 240 3271 265
rect 3231 225 3271 240
rect 3476 265 3516 275
rect 3476 240 3481 265
rect 3506 240 3516 265
rect 3476 225 3516 240
rect 3716 265 3756 275
rect 3716 240 3721 265
rect 3746 240 3756 265
rect 3716 225 3756 240
rect 3961 265 4001 275
rect 3961 240 3966 265
rect 3991 240 4001 265
rect 4446 265 4486 275
rect 3961 225 4001 240
rect 4446 240 4451 265
rect 4476 240 4486 265
rect 4446 225 4486 240
rect 4686 265 4726 275
rect 4686 240 4691 265
rect 4716 240 4726 265
rect 4686 225 4726 240
rect 4931 265 4971 275
rect 4931 240 4936 265
rect 4961 240 4971 265
rect 4931 225 4971 240
rect 5171 265 5211 275
rect 5171 240 5176 265
rect 5201 240 5211 265
rect 5171 225 5211 240
rect 5416 265 5456 275
rect 5416 240 5421 265
rect 5446 240 5456 265
rect 5416 225 5456 240
rect 5721 265 5761 275
rect 5721 240 5726 265
rect 5751 240 5761 265
rect 5721 225 5761 240
rect 5966 265 6006 275
rect 5966 240 5971 265
rect 5996 240 6006 265
rect 5966 225 6006 240
rect 6206 265 6246 275
rect 6206 240 6211 265
rect 6236 240 6246 265
rect 6691 265 6731 275
rect 6206 225 6246 240
rect 6691 240 6696 265
rect 6721 240 6731 265
rect 6691 225 6731 240
rect 6936 265 6976 275
rect 6936 240 6941 265
rect 6966 240 6976 265
rect 6936 225 6976 240
rect 7176 265 7216 275
rect 7176 240 7181 265
rect 7206 240 7216 265
rect 7176 225 7216 240
rect 7416 265 7456 275
rect 7416 240 7421 265
rect 7446 240 7456 265
rect 7416 225 7456 240
rect 7656 265 7696 275
rect 7656 240 7661 265
rect 7686 240 7696 265
rect 7656 225 7696 240
rect 7901 265 7941 275
rect 7901 240 7906 265
rect 7931 240 7941 265
rect 7901 225 7941 240
rect 8141 265 8181 275
rect 8141 240 8146 265
rect 8171 240 8181 265
rect 8141 225 8181 240
rect 8386 265 8426 275
rect 8386 240 8391 265
rect 8416 240 8426 265
rect 8386 225 8426 240
rect 8626 265 8666 275
rect 8626 240 8631 265
rect 8656 240 8666 265
rect 8626 225 8666 240
rect 8871 265 8911 275
rect 8871 240 8876 265
rect 8901 240 8911 265
rect 8871 225 8911 240
rect 9111 265 9151 275
rect 9111 240 9116 265
rect 9141 240 9151 265
rect 9601 265 9641 275
rect 9111 225 9151 240
rect 9601 240 9606 265
rect 9631 240 9641 265
rect 9601 225 9641 240
rect 9846 265 9886 275
rect 9846 240 9851 265
rect 9876 240 9886 265
rect 9846 225 9886 240
rect 10086 265 10126 275
rect 10086 240 10091 265
rect 10116 240 10126 265
rect 10086 225 10126 240
rect 10331 265 10371 275
rect 10331 240 10336 265
rect 10361 240 10371 265
rect 10331 225 10371 240
rect 10571 265 10611 275
rect 10571 240 10576 265
rect 10601 240 10611 265
rect 10571 225 10611 240
rect 10816 265 10856 275
rect 10816 240 10821 265
rect 10846 240 10856 265
rect 10816 225 10856 240
rect 11056 265 11096 275
rect 11056 240 11061 265
rect 11086 240 11096 265
rect 11541 265 11581 275
rect 11056 225 11096 240
rect 11541 240 11546 265
rect 11571 240 11581 265
rect 11541 225 11581 240
rect 11786 265 11826 275
rect 11786 240 11791 265
rect 11816 240 11826 265
rect 11786 225 11826 240
rect 12026 265 12066 275
rect 12026 240 12031 265
rect 12056 240 12066 265
rect 12026 225 12066 240
rect 12271 265 12311 275
rect 12271 240 12276 265
rect 12301 240 12311 265
rect 12271 225 12311 240
rect 12511 265 12551 275
rect 12511 240 12516 265
rect 12541 240 12551 265
rect 12511 225 12551 240
rect 12756 265 12796 275
rect 12756 240 12761 265
rect 12786 240 12796 265
rect 13241 265 13281 275
rect 12756 225 12796 240
rect 13241 240 13246 265
rect 13271 240 13281 265
rect 13241 225 13281 240
rect 13481 265 13521 275
rect 13481 240 13486 265
rect 13511 240 13521 265
rect 13481 225 13521 240
rect 13726 265 13766 275
rect 13726 240 13731 265
rect 13756 240 13766 265
rect 13726 225 13766 240
rect 13966 265 14006 275
rect 13966 240 13971 265
rect 13996 240 14006 265
rect 13966 225 14006 240
rect 14211 265 14251 275
rect 14211 240 14216 265
rect 14241 240 14251 265
rect 14211 225 14251 240
rect 14451 265 14491 275
rect 14451 240 14456 265
rect 14481 240 14491 265
rect 14451 225 14491 240
rect 14696 265 14736 275
rect 14696 240 14701 265
rect 14726 240 14736 265
rect 14696 225 14736 240
rect 14936 265 14976 275
rect 14936 240 14941 265
rect 14966 240 14976 265
rect 15421 265 15461 275
rect 14936 225 14976 240
rect 15421 240 15426 265
rect 15451 240 15461 265
rect 15421 225 15461 240
rect 15666 265 15706 275
rect 15666 240 15671 265
rect 15696 240 15706 265
rect 15666 225 15706 240
rect 15906 265 15946 275
rect 15906 240 15911 265
rect 15936 240 15946 265
rect 15906 225 15946 240
rect 16151 265 16191 275
rect 16151 240 16156 265
rect 16181 240 16191 265
rect 16151 225 16191 240
rect 16391 265 16431 275
rect 16391 240 16396 265
rect 16421 240 16431 265
rect 16391 225 16431 240
rect 16636 265 16676 275
rect 16636 240 16641 265
rect 16666 240 16676 265
rect 16636 225 16676 240
rect 16876 265 16916 275
rect 16876 240 16881 265
rect 16906 240 16916 265
rect 16876 225 16916 240
rect 17121 265 17161 275
rect 17121 240 17126 265
rect 17151 240 17161 265
rect 17606 265 17646 275
rect 17121 225 17161 240
rect 17606 240 17611 265
rect 17636 240 17646 265
rect 17606 225 17646 240
rect 17846 265 17886 275
rect 17846 240 17851 265
rect 17876 240 17886 265
rect 17846 225 17886 240
rect 18091 265 18131 275
rect 18091 240 18096 265
rect 18121 240 18131 265
rect 18091 225 18131 240
rect 18331 265 18371 275
rect 18331 240 18336 265
rect 18361 240 18371 265
rect 18331 225 18371 240
rect 18576 265 18616 275
rect 18576 240 18581 265
rect 18606 240 18616 265
rect 18576 225 18616 240
rect 18816 265 18856 275
rect 18816 240 18821 265
rect 18846 240 18856 265
rect 18816 225 18856 240
rect 19061 265 19101 275
rect 19061 240 19066 265
rect 19091 240 19101 265
rect 19061 225 19101 240
rect 19301 265 19341 275
rect 19301 240 19306 265
rect 19331 240 19341 265
rect 19786 265 19826 275
rect 19301 225 19341 240
rect 19786 240 19791 265
rect 19816 240 19826 265
rect 19786 225 19826 240
rect 20031 265 20071 275
rect 20031 240 20036 265
rect 20061 240 20071 265
rect 20031 225 20071 240
rect 20271 265 20311 275
rect 20271 240 20276 265
rect 20301 240 20311 265
rect 20271 225 20311 240
rect 20516 265 20556 275
rect 20516 240 20521 265
rect 20546 240 20556 265
rect 21001 265 21041 275
rect 20516 225 20556 240
rect 21001 240 21006 265
rect 21031 240 21041 265
rect 21001 225 21041 240
rect 191 165 231 185
rect 191 140 196 165
rect 221 140 231 165
rect 191 120 231 140
rect 191 95 196 120
rect 221 95 231 120
rect 191 85 231 95
rect 246 165 286 185
rect 246 140 256 165
rect 281 140 286 165
rect 246 120 286 140
rect 246 95 256 120
rect 281 95 286 120
rect 246 85 286 95
rect 316 165 356 185
rect 316 140 321 165
rect 346 140 356 165
rect 316 120 356 140
rect 316 95 321 120
rect 346 95 356 120
rect 316 85 356 95
rect 371 165 416 185
rect 371 140 381 165
rect 406 140 416 165
rect 371 120 416 140
rect 371 95 381 120
rect 406 95 416 120
rect 371 85 416 95
rect 431 165 476 185
rect 431 140 441 165
rect 466 140 476 165
rect 431 120 476 140
rect 431 95 441 120
rect 466 95 476 120
rect 431 85 476 95
rect 491 165 536 185
rect 491 140 501 165
rect 526 140 536 165
rect 491 120 536 140
rect 491 95 501 120
rect 526 95 536 120
rect 491 85 536 95
rect 551 165 591 185
rect 551 140 561 165
rect 586 140 591 165
rect 551 120 591 140
rect 551 95 561 120
rect 586 95 591 120
rect 551 85 591 95
rect 621 165 661 185
rect 621 140 626 165
rect 651 140 661 165
rect 621 120 661 140
rect 621 95 626 120
rect 651 95 661 120
rect 621 85 661 95
rect 676 165 721 185
rect 676 140 686 165
rect 711 140 721 165
rect 676 120 721 140
rect 676 95 686 120
rect 711 95 721 120
rect 676 85 721 95
rect 736 165 781 185
rect 736 140 746 165
rect 771 140 781 165
rect 736 120 781 140
rect 736 95 746 120
rect 771 95 781 120
rect 736 85 781 95
rect 796 165 841 185
rect 796 140 806 165
rect 831 140 841 165
rect 796 120 841 140
rect 796 95 806 120
rect 831 95 841 120
rect 796 85 841 95
rect 856 165 906 185
rect 856 140 871 165
rect 896 140 906 165
rect 856 120 906 140
rect 856 95 871 120
rect 896 95 906 120
rect 856 85 906 95
rect 921 165 966 185
rect 921 140 931 165
rect 956 140 966 165
rect 921 120 966 140
rect 921 95 931 120
rect 956 95 966 120
rect 921 85 966 95
rect 981 165 1026 185
rect 981 140 991 165
rect 1016 140 1026 165
rect 981 120 1026 140
rect 981 95 991 120
rect 1016 95 1026 120
rect 981 85 1026 95
rect 1041 165 1086 185
rect 1041 140 1051 165
rect 1076 140 1086 165
rect 1041 120 1086 140
rect 1041 95 1051 120
rect 1076 95 1086 120
rect 1041 85 1086 95
rect 1101 165 1146 185
rect 1101 140 1111 165
rect 1136 140 1146 165
rect 1101 120 1146 140
rect 1101 95 1111 120
rect 1136 95 1146 120
rect 1101 85 1146 95
rect 1161 165 1206 185
rect 1161 140 1171 165
rect 1196 140 1206 165
rect 1161 120 1206 140
rect 1161 95 1171 120
rect 1196 95 1206 120
rect 1161 85 1206 95
rect 1221 165 1266 185
rect 1221 140 1231 165
rect 1256 140 1266 165
rect 1221 120 1266 140
rect 1221 95 1231 120
rect 1256 95 1266 120
rect 1221 85 1266 95
rect 1281 165 1326 185
rect 1281 140 1291 165
rect 1316 140 1326 165
rect 1281 120 1326 140
rect 1281 95 1291 120
rect 1316 95 1326 120
rect 1281 85 1326 95
rect 1341 165 1391 185
rect 1341 140 1356 165
rect 1381 140 1391 165
rect 1341 120 1391 140
rect 1341 95 1356 120
rect 1381 95 1391 120
rect 1341 85 1391 95
rect 1406 165 1451 185
rect 1406 140 1416 165
rect 1441 140 1451 165
rect 1406 120 1451 140
rect 1406 95 1416 120
rect 1441 95 1451 120
rect 1406 85 1451 95
rect 1466 165 1511 185
rect 1466 140 1476 165
rect 1501 140 1511 165
rect 1466 120 1511 140
rect 1466 95 1476 120
rect 1501 95 1511 120
rect 1466 85 1511 95
rect 1526 165 1571 185
rect 1526 140 1536 165
rect 1561 140 1571 165
rect 1526 120 1571 140
rect 1526 95 1536 120
rect 1561 95 1571 120
rect 1526 85 1571 95
rect 1586 165 1626 185
rect 1586 140 1596 165
rect 1621 140 1626 165
rect 1586 120 1626 140
rect 1586 95 1596 120
rect 1621 95 1626 120
rect 1586 85 1626 95
rect 1656 165 1696 185
rect 1656 140 1661 165
rect 1686 140 1696 165
rect 1656 120 1696 140
rect 1656 95 1661 120
rect 1686 95 1696 120
rect 1656 85 1696 95
rect 1711 165 1756 185
rect 1711 140 1721 165
rect 1746 140 1756 165
rect 1711 120 1756 140
rect 1711 95 1721 120
rect 1746 95 1756 120
rect 1711 85 1756 95
rect 1771 165 1816 185
rect 1771 140 1781 165
rect 1806 140 1816 165
rect 1771 120 1816 140
rect 1771 95 1781 120
rect 1806 95 1816 120
rect 1771 85 1816 95
rect 1831 165 1876 185
rect 1831 140 1841 165
rect 1866 140 1876 165
rect 1831 120 1876 140
rect 1831 95 1841 120
rect 1866 95 1876 120
rect 1831 85 1876 95
rect 1891 165 1941 185
rect 1891 140 1906 165
rect 1931 140 1941 165
rect 1891 120 1941 140
rect 1891 95 1906 120
rect 1931 95 1941 120
rect 1891 85 1941 95
rect 1956 165 2001 185
rect 1956 140 1966 165
rect 1991 140 2001 165
rect 1956 120 2001 140
rect 1956 95 1966 120
rect 1991 95 2001 120
rect 1956 85 2001 95
rect 2016 165 2061 185
rect 2016 140 2026 165
rect 2051 140 2061 165
rect 2016 120 2061 140
rect 2016 95 2026 120
rect 2051 95 2061 120
rect 2016 85 2061 95
rect 2076 165 2121 185
rect 2076 140 2086 165
rect 2111 140 2121 165
rect 2076 120 2121 140
rect 2076 95 2086 120
rect 2111 95 2121 120
rect 2076 85 2121 95
rect 2136 165 2181 185
rect 2136 140 2146 165
rect 2171 140 2181 165
rect 2136 120 2181 140
rect 2136 95 2146 120
rect 2171 95 2181 120
rect 2136 85 2181 95
rect 2196 165 2241 185
rect 2196 140 2206 165
rect 2231 140 2241 165
rect 2196 120 2241 140
rect 2196 95 2206 120
rect 2231 95 2241 120
rect 2196 85 2241 95
rect 2256 165 2301 185
rect 2256 140 2266 165
rect 2291 140 2301 165
rect 2256 120 2301 140
rect 2256 95 2266 120
rect 2291 95 2301 120
rect 2256 85 2301 95
rect 2316 165 2361 185
rect 2316 140 2326 165
rect 2351 140 2361 165
rect 2316 120 2361 140
rect 2316 95 2326 120
rect 2351 95 2361 120
rect 2316 85 2361 95
rect 2376 165 2426 185
rect 2376 140 2391 165
rect 2416 140 2426 165
rect 2376 120 2426 140
rect 2376 95 2391 120
rect 2416 95 2426 120
rect 2376 85 2426 95
rect 2441 165 2486 185
rect 2441 140 2451 165
rect 2476 140 2486 165
rect 2441 120 2486 140
rect 2441 95 2451 120
rect 2476 95 2486 120
rect 2441 85 2486 95
rect 2501 165 2546 185
rect 2501 140 2511 165
rect 2536 140 2546 165
rect 2501 120 2546 140
rect 2501 95 2511 120
rect 2536 95 2546 120
rect 2501 85 2546 95
rect 2561 165 2606 185
rect 2561 140 2571 165
rect 2596 140 2606 165
rect 2561 120 2606 140
rect 2561 95 2571 120
rect 2596 95 2606 120
rect 2561 85 2606 95
rect 2621 165 2666 185
rect 2621 140 2631 165
rect 2656 140 2666 165
rect 2621 120 2666 140
rect 2621 95 2631 120
rect 2656 95 2666 120
rect 2621 85 2666 95
rect 2681 165 2726 185
rect 2681 140 2691 165
rect 2716 140 2726 165
rect 2681 120 2726 140
rect 2681 95 2691 120
rect 2716 95 2726 120
rect 2681 85 2726 95
rect 2741 165 2786 185
rect 2741 140 2751 165
rect 2776 140 2786 165
rect 2741 120 2786 140
rect 2741 95 2751 120
rect 2776 95 2786 120
rect 2741 85 2786 95
rect 2801 165 2846 185
rect 2801 140 2811 165
rect 2836 140 2846 165
rect 2801 120 2846 140
rect 2801 95 2811 120
rect 2836 95 2846 120
rect 2801 85 2846 95
rect 2861 165 2911 185
rect 2861 140 2876 165
rect 2901 140 2911 165
rect 2861 120 2911 140
rect 2861 95 2876 120
rect 2901 95 2911 120
rect 2861 85 2911 95
rect 2926 165 2971 185
rect 2926 140 2936 165
rect 2961 140 2971 165
rect 2926 120 2971 140
rect 2926 95 2936 120
rect 2961 95 2971 120
rect 2926 85 2971 95
rect 2986 165 3031 185
rect 2986 140 2996 165
rect 3021 140 3031 165
rect 2986 120 3031 140
rect 2986 95 2996 120
rect 3021 95 3031 120
rect 2986 85 3031 95
rect 3046 165 3091 185
rect 3046 140 3056 165
rect 3081 140 3091 165
rect 3046 120 3091 140
rect 3046 95 3056 120
rect 3081 95 3091 120
rect 3046 85 3091 95
rect 3106 165 3151 185
rect 3106 140 3116 165
rect 3141 140 3151 165
rect 3106 120 3151 140
rect 3106 95 3116 120
rect 3141 95 3151 120
rect 3106 85 3151 95
rect 3166 165 3211 185
rect 3166 140 3176 165
rect 3201 140 3211 165
rect 3166 120 3211 140
rect 3166 95 3176 120
rect 3201 95 3211 120
rect 3166 85 3211 95
rect 3226 165 3271 185
rect 3226 140 3236 165
rect 3261 140 3271 165
rect 3226 120 3271 140
rect 3226 95 3236 120
rect 3261 95 3271 120
rect 3226 85 3271 95
rect 3286 165 3331 185
rect 3286 140 3296 165
rect 3321 140 3331 165
rect 3286 120 3331 140
rect 3286 95 3296 120
rect 3321 95 3331 120
rect 3286 85 3331 95
rect 3346 165 3396 185
rect 3346 140 3361 165
rect 3386 140 3396 165
rect 3346 120 3396 140
rect 3346 95 3361 120
rect 3386 95 3396 120
rect 3346 85 3396 95
rect 3411 165 3456 185
rect 3411 140 3421 165
rect 3446 140 3456 165
rect 3411 120 3456 140
rect 3411 95 3421 120
rect 3446 95 3456 120
rect 3411 85 3456 95
rect 3471 165 3516 185
rect 3471 140 3481 165
rect 3506 140 3516 165
rect 3471 120 3516 140
rect 3471 95 3481 120
rect 3506 95 3516 120
rect 3471 85 3516 95
rect 3531 165 3576 185
rect 3531 140 3541 165
rect 3566 140 3576 165
rect 3531 120 3576 140
rect 3531 95 3541 120
rect 3566 95 3576 120
rect 3531 85 3576 95
rect 3591 165 3636 185
rect 3591 140 3601 165
rect 3626 140 3636 165
rect 3591 120 3636 140
rect 3591 95 3601 120
rect 3626 95 3636 120
rect 3591 85 3636 95
rect 3651 165 3696 185
rect 3651 140 3661 165
rect 3686 140 3696 165
rect 3651 120 3696 140
rect 3651 95 3661 120
rect 3686 95 3696 120
rect 3651 85 3696 95
rect 3711 165 3756 185
rect 3711 140 3721 165
rect 3746 140 3756 165
rect 3711 120 3756 140
rect 3711 95 3721 120
rect 3746 95 3756 120
rect 3711 85 3756 95
rect 3771 165 3816 185
rect 3771 140 3781 165
rect 3806 140 3816 165
rect 3771 120 3816 140
rect 3771 95 3781 120
rect 3806 95 3816 120
rect 3771 85 3816 95
rect 3831 165 3881 185
rect 3831 140 3846 165
rect 3871 140 3881 165
rect 3831 120 3881 140
rect 3831 95 3846 120
rect 3871 95 3881 120
rect 3831 85 3881 95
rect 3896 165 3941 185
rect 3896 140 3906 165
rect 3931 140 3941 165
rect 3896 120 3941 140
rect 3896 95 3906 120
rect 3931 95 3941 120
rect 3896 85 3941 95
rect 3956 165 4001 185
rect 3956 140 3966 165
rect 3991 140 4001 165
rect 3956 120 4001 140
rect 3956 95 3966 120
rect 3991 95 4001 120
rect 3956 85 4001 95
rect 4016 165 4061 185
rect 4016 140 4026 165
rect 4051 140 4061 165
rect 4016 120 4061 140
rect 4016 95 4026 120
rect 4051 95 4061 120
rect 4016 85 4061 95
rect 4076 165 4121 185
rect 4076 140 4086 165
rect 4111 140 4121 165
rect 4076 120 4121 140
rect 4076 95 4086 120
rect 4111 95 4121 120
rect 4076 85 4121 95
rect 4136 165 4181 185
rect 4136 140 4146 165
rect 4171 140 4181 165
rect 4136 120 4181 140
rect 4136 95 4146 120
rect 4171 95 4181 120
rect 4136 85 4181 95
rect 4196 165 4241 185
rect 4196 140 4206 165
rect 4231 140 4241 165
rect 4196 120 4241 140
rect 4196 95 4206 120
rect 4231 95 4241 120
rect 4196 85 4241 95
rect 4256 165 4301 185
rect 4256 140 4266 165
rect 4291 140 4301 165
rect 4256 120 4301 140
rect 4256 95 4266 120
rect 4291 95 4301 120
rect 4256 85 4301 95
rect 4316 165 4366 185
rect 4316 140 4331 165
rect 4356 140 4366 165
rect 4316 120 4366 140
rect 4316 95 4331 120
rect 4356 95 4366 120
rect 4316 85 4366 95
rect 4381 165 4426 185
rect 4381 140 4391 165
rect 4416 140 4426 165
rect 4381 120 4426 140
rect 4381 95 4391 120
rect 4416 95 4426 120
rect 4381 85 4426 95
rect 4441 165 4486 185
rect 4441 140 4451 165
rect 4476 140 4486 165
rect 4441 120 4486 140
rect 4441 95 4451 120
rect 4476 95 4486 120
rect 4441 85 4486 95
rect 4501 165 4546 185
rect 4501 140 4511 165
rect 4536 140 4546 165
rect 4501 120 4546 140
rect 4501 95 4511 120
rect 4536 95 4546 120
rect 4501 85 4546 95
rect 4561 165 4606 185
rect 4561 140 4571 165
rect 4596 140 4606 165
rect 4561 120 4606 140
rect 4561 95 4571 120
rect 4596 95 4606 120
rect 4561 85 4606 95
rect 4621 165 4666 185
rect 4621 140 4631 165
rect 4656 140 4666 165
rect 4621 120 4666 140
rect 4621 95 4631 120
rect 4656 95 4666 120
rect 4621 85 4666 95
rect 4681 165 4726 185
rect 4681 140 4691 165
rect 4716 140 4726 165
rect 4681 120 4726 140
rect 4681 95 4691 120
rect 4716 95 4726 120
rect 4681 85 4726 95
rect 4741 165 4786 185
rect 4741 140 4751 165
rect 4776 140 4786 165
rect 4741 120 4786 140
rect 4741 95 4751 120
rect 4776 95 4786 120
rect 4741 85 4786 95
rect 4801 165 4851 185
rect 4801 140 4816 165
rect 4841 140 4851 165
rect 4801 120 4851 140
rect 4801 95 4816 120
rect 4841 95 4851 120
rect 4801 85 4851 95
rect 4866 165 4911 185
rect 4866 140 4876 165
rect 4901 140 4911 165
rect 4866 120 4911 140
rect 4866 95 4876 120
rect 4901 95 4911 120
rect 4866 85 4911 95
rect 4926 165 4971 185
rect 4926 140 4936 165
rect 4961 140 4971 165
rect 4926 120 4971 140
rect 4926 95 4936 120
rect 4961 95 4971 120
rect 4926 85 4971 95
rect 4986 165 5031 185
rect 4986 140 4996 165
rect 5021 140 5031 165
rect 4986 120 5031 140
rect 4986 95 4996 120
rect 5021 95 5031 120
rect 4986 85 5031 95
rect 5046 165 5091 185
rect 5046 140 5056 165
rect 5081 140 5091 165
rect 5046 120 5091 140
rect 5046 95 5056 120
rect 5081 95 5091 120
rect 5046 85 5091 95
rect 5106 165 5151 185
rect 5106 140 5116 165
rect 5141 140 5151 165
rect 5106 120 5151 140
rect 5106 95 5116 120
rect 5141 95 5151 120
rect 5106 85 5151 95
rect 5166 165 5211 185
rect 5166 140 5176 165
rect 5201 140 5211 165
rect 5166 120 5211 140
rect 5166 95 5176 120
rect 5201 95 5211 120
rect 5166 85 5211 95
rect 5226 165 5271 185
rect 5226 140 5236 165
rect 5261 140 5271 165
rect 5226 120 5271 140
rect 5226 95 5236 120
rect 5261 95 5271 120
rect 5226 85 5271 95
rect 5286 165 5336 185
rect 5286 140 5301 165
rect 5326 140 5336 165
rect 5286 120 5336 140
rect 5286 95 5301 120
rect 5326 95 5336 120
rect 5286 85 5336 95
rect 5351 165 5396 185
rect 5351 140 5361 165
rect 5386 140 5396 165
rect 5351 120 5396 140
rect 5351 95 5361 120
rect 5386 95 5396 120
rect 5351 85 5396 95
rect 5411 165 5456 185
rect 5411 140 5421 165
rect 5446 140 5456 165
rect 5411 120 5456 140
rect 5411 95 5421 120
rect 5446 95 5456 120
rect 5411 85 5456 95
rect 5471 165 5516 185
rect 5471 140 5481 165
rect 5506 140 5516 165
rect 5471 120 5516 140
rect 5471 95 5481 120
rect 5506 95 5516 120
rect 5471 85 5516 95
rect 5531 165 5571 185
rect 5531 140 5541 165
rect 5566 140 5571 165
rect 5531 120 5571 140
rect 5531 95 5541 120
rect 5566 95 5571 120
rect 5531 85 5571 95
rect 5601 165 5641 185
rect 5601 140 5606 165
rect 5631 140 5641 165
rect 5601 120 5641 140
rect 5601 95 5606 120
rect 5631 95 5641 120
rect 5601 85 5641 95
rect 5656 165 5701 185
rect 5656 140 5666 165
rect 5691 140 5701 165
rect 5656 120 5701 140
rect 5656 95 5666 120
rect 5691 95 5701 120
rect 5656 85 5701 95
rect 5716 165 5761 185
rect 5716 140 5726 165
rect 5751 140 5761 165
rect 5716 120 5761 140
rect 5716 95 5726 120
rect 5751 95 5761 120
rect 5716 85 5761 95
rect 5776 165 5821 185
rect 5776 140 5786 165
rect 5811 140 5821 165
rect 5776 120 5821 140
rect 5776 95 5786 120
rect 5811 95 5821 120
rect 5776 85 5821 95
rect 5836 165 5886 185
rect 5836 140 5851 165
rect 5876 140 5886 165
rect 5836 120 5886 140
rect 5836 95 5851 120
rect 5876 95 5886 120
rect 5836 85 5886 95
rect 5901 165 5946 185
rect 5901 140 5911 165
rect 5936 140 5946 165
rect 5901 120 5946 140
rect 5901 95 5911 120
rect 5936 95 5946 120
rect 5901 85 5946 95
rect 5961 165 6006 185
rect 5961 140 5971 165
rect 5996 140 6006 165
rect 5961 120 6006 140
rect 5961 95 5971 120
rect 5996 95 6006 120
rect 5961 85 6006 95
rect 6021 165 6066 185
rect 6021 140 6031 165
rect 6056 140 6066 165
rect 6021 120 6066 140
rect 6021 95 6031 120
rect 6056 95 6066 120
rect 6021 85 6066 95
rect 6081 165 6126 185
rect 6081 140 6091 165
rect 6116 140 6126 165
rect 6081 120 6126 140
rect 6081 95 6091 120
rect 6116 95 6126 120
rect 6081 85 6126 95
rect 6141 165 6186 185
rect 6141 140 6151 165
rect 6176 140 6186 165
rect 6141 120 6186 140
rect 6141 95 6151 120
rect 6176 95 6186 120
rect 6141 85 6186 95
rect 6201 165 6246 185
rect 6201 140 6211 165
rect 6236 140 6246 165
rect 6201 120 6246 140
rect 6201 95 6211 120
rect 6236 95 6246 120
rect 6201 85 6246 95
rect 6261 165 6306 185
rect 6261 140 6271 165
rect 6296 140 6306 165
rect 6261 120 6306 140
rect 6261 95 6271 120
rect 6296 95 6306 120
rect 6261 85 6306 95
rect 6321 165 6371 185
rect 6321 140 6336 165
rect 6361 140 6371 165
rect 6321 120 6371 140
rect 6321 95 6336 120
rect 6361 95 6371 120
rect 6321 85 6371 95
rect 6386 165 6431 185
rect 6386 140 6396 165
rect 6421 140 6431 165
rect 6386 120 6431 140
rect 6386 95 6396 120
rect 6421 95 6431 120
rect 6386 85 6431 95
rect 6446 165 6491 185
rect 6446 140 6456 165
rect 6481 140 6491 165
rect 6446 120 6491 140
rect 6446 95 6456 120
rect 6481 95 6491 120
rect 6446 85 6491 95
rect 6506 165 6551 185
rect 6506 140 6516 165
rect 6541 140 6551 165
rect 6506 120 6551 140
rect 6506 95 6516 120
rect 6541 95 6551 120
rect 6506 85 6551 95
rect 6566 165 6611 185
rect 6566 140 6576 165
rect 6601 140 6611 165
rect 6566 120 6611 140
rect 6566 95 6576 120
rect 6601 95 6611 120
rect 6566 85 6611 95
rect 6626 165 6671 185
rect 6626 140 6636 165
rect 6661 140 6671 165
rect 6626 120 6671 140
rect 6626 95 6636 120
rect 6661 95 6671 120
rect 6626 85 6671 95
rect 6686 165 6731 185
rect 6686 140 6696 165
rect 6721 140 6731 165
rect 6686 120 6731 140
rect 6686 95 6696 120
rect 6721 95 6731 120
rect 6686 85 6731 95
rect 6746 165 6791 185
rect 6746 140 6756 165
rect 6781 140 6791 165
rect 6746 120 6791 140
rect 6746 95 6756 120
rect 6781 95 6791 120
rect 6746 85 6791 95
rect 6806 165 6856 185
rect 6806 140 6821 165
rect 6846 140 6856 165
rect 6806 120 6856 140
rect 6806 95 6821 120
rect 6846 95 6856 120
rect 6806 85 6856 95
rect 6871 165 6916 185
rect 6871 140 6881 165
rect 6906 140 6916 165
rect 6871 120 6916 140
rect 6871 95 6881 120
rect 6906 95 6916 120
rect 6871 85 6916 95
rect 6931 165 6976 185
rect 6931 140 6941 165
rect 6966 140 6976 165
rect 6931 120 6976 140
rect 6931 95 6941 120
rect 6966 95 6976 120
rect 6931 85 6976 95
rect 6991 165 7036 185
rect 6991 140 7001 165
rect 7026 140 7036 165
rect 6991 120 7036 140
rect 6991 95 7001 120
rect 7026 95 7036 120
rect 6991 85 7036 95
rect 7051 165 7096 185
rect 7051 140 7061 165
rect 7086 140 7096 165
rect 7051 120 7096 140
rect 7051 95 7061 120
rect 7086 95 7096 120
rect 7051 85 7096 95
rect 7111 165 7156 185
rect 7111 140 7121 165
rect 7146 140 7156 165
rect 7111 120 7156 140
rect 7111 95 7121 120
rect 7146 95 7156 120
rect 7111 85 7156 95
rect 7171 165 7216 185
rect 7171 140 7181 165
rect 7206 140 7216 165
rect 7171 120 7216 140
rect 7171 95 7181 120
rect 7206 95 7216 120
rect 7171 85 7216 95
rect 7231 165 7276 185
rect 7231 140 7241 165
rect 7266 140 7276 165
rect 7231 120 7276 140
rect 7231 95 7241 120
rect 7266 95 7276 120
rect 7231 85 7276 95
rect 7291 165 7336 185
rect 7291 140 7301 165
rect 7326 140 7336 165
rect 7291 120 7336 140
rect 7291 95 7301 120
rect 7326 95 7336 120
rect 7291 85 7336 95
rect 7351 165 7396 185
rect 7351 140 7361 165
rect 7386 140 7396 165
rect 7351 120 7396 140
rect 7351 95 7361 120
rect 7386 95 7396 120
rect 7351 85 7396 95
rect 7411 165 7456 185
rect 7411 140 7421 165
rect 7446 140 7456 165
rect 7411 120 7456 140
rect 7411 95 7421 120
rect 7446 95 7456 120
rect 7411 85 7456 95
rect 7471 165 7516 185
rect 7471 140 7481 165
rect 7506 140 7516 165
rect 7471 120 7516 140
rect 7471 95 7481 120
rect 7506 95 7516 120
rect 7471 85 7516 95
rect 7531 165 7576 185
rect 7531 140 7541 165
rect 7566 140 7576 165
rect 7531 120 7576 140
rect 7531 95 7541 120
rect 7566 95 7576 120
rect 7531 85 7576 95
rect 7591 165 7636 185
rect 7591 140 7601 165
rect 7626 140 7636 165
rect 7591 120 7636 140
rect 7591 95 7601 120
rect 7626 95 7636 120
rect 7591 85 7636 95
rect 7651 165 7696 185
rect 7651 140 7661 165
rect 7686 140 7696 165
rect 7651 120 7696 140
rect 7651 95 7661 120
rect 7686 95 7696 120
rect 7651 85 7696 95
rect 7711 165 7756 185
rect 7711 140 7721 165
rect 7746 140 7756 165
rect 7711 120 7756 140
rect 7711 95 7721 120
rect 7746 95 7756 120
rect 7711 85 7756 95
rect 7771 165 7821 185
rect 7771 140 7786 165
rect 7811 140 7821 165
rect 7771 120 7821 140
rect 7771 95 7786 120
rect 7811 95 7821 120
rect 7771 85 7821 95
rect 7836 165 7881 185
rect 7836 140 7846 165
rect 7871 140 7881 165
rect 7836 120 7881 140
rect 7836 95 7846 120
rect 7871 95 7881 120
rect 7836 85 7881 95
rect 7896 165 7941 185
rect 7896 140 7906 165
rect 7931 140 7941 165
rect 7896 120 7941 140
rect 7896 95 7906 120
rect 7931 95 7941 120
rect 7896 85 7941 95
rect 7956 165 8001 185
rect 7956 140 7966 165
rect 7991 140 8001 165
rect 7956 120 8001 140
rect 7956 95 7966 120
rect 7991 95 8001 120
rect 7956 85 8001 95
rect 8016 165 8061 185
rect 8016 140 8026 165
rect 8051 140 8061 165
rect 8016 120 8061 140
rect 8016 95 8026 120
rect 8051 95 8061 120
rect 8016 85 8061 95
rect 8076 165 8121 185
rect 8076 140 8086 165
rect 8111 140 8121 165
rect 8076 120 8121 140
rect 8076 95 8086 120
rect 8111 95 8121 120
rect 8076 85 8121 95
rect 8136 165 8181 185
rect 8136 140 8146 165
rect 8171 140 8181 165
rect 8136 120 8181 140
rect 8136 95 8146 120
rect 8171 95 8181 120
rect 8136 85 8181 95
rect 8196 165 8241 185
rect 8196 140 8206 165
rect 8231 140 8241 165
rect 8196 120 8241 140
rect 8196 95 8206 120
rect 8231 95 8241 120
rect 8196 85 8241 95
rect 8256 165 8306 185
rect 8256 140 8271 165
rect 8296 140 8306 165
rect 8256 120 8306 140
rect 8256 95 8271 120
rect 8296 95 8306 120
rect 8256 85 8306 95
rect 8321 165 8366 185
rect 8321 140 8331 165
rect 8356 140 8366 165
rect 8321 120 8366 140
rect 8321 95 8331 120
rect 8356 95 8366 120
rect 8321 85 8366 95
rect 8381 165 8426 185
rect 8381 140 8391 165
rect 8416 140 8426 165
rect 8381 120 8426 140
rect 8381 95 8391 120
rect 8416 95 8426 120
rect 8381 85 8426 95
rect 8441 165 8486 185
rect 8441 140 8451 165
rect 8476 140 8486 165
rect 8441 120 8486 140
rect 8441 95 8451 120
rect 8476 95 8486 120
rect 8441 85 8486 95
rect 8501 165 8546 185
rect 8501 140 8511 165
rect 8536 140 8546 165
rect 8501 120 8546 140
rect 8501 95 8511 120
rect 8536 95 8546 120
rect 8501 85 8546 95
rect 8561 165 8606 185
rect 8561 140 8571 165
rect 8596 140 8606 165
rect 8561 120 8606 140
rect 8561 95 8571 120
rect 8596 95 8606 120
rect 8561 85 8606 95
rect 8621 165 8666 185
rect 8621 140 8631 165
rect 8656 140 8666 165
rect 8621 120 8666 140
rect 8621 95 8631 120
rect 8656 95 8666 120
rect 8621 85 8666 95
rect 8681 165 8726 185
rect 8681 140 8691 165
rect 8716 140 8726 165
rect 8681 120 8726 140
rect 8681 95 8691 120
rect 8716 95 8726 120
rect 8681 85 8726 95
rect 8741 165 8791 185
rect 8741 140 8756 165
rect 8781 140 8791 165
rect 8741 120 8791 140
rect 8741 95 8756 120
rect 8781 95 8791 120
rect 8741 85 8791 95
rect 8806 165 8851 185
rect 8806 140 8816 165
rect 8841 140 8851 165
rect 8806 120 8851 140
rect 8806 95 8816 120
rect 8841 95 8851 120
rect 8806 85 8851 95
rect 8866 165 8911 185
rect 8866 140 8876 165
rect 8901 140 8911 165
rect 8866 120 8911 140
rect 8866 95 8876 120
rect 8901 95 8911 120
rect 8866 85 8911 95
rect 8926 165 8971 185
rect 8926 140 8936 165
rect 8961 140 8971 165
rect 8926 120 8971 140
rect 8926 95 8936 120
rect 8961 95 8971 120
rect 8926 85 8971 95
rect 8986 165 9031 185
rect 8986 140 8996 165
rect 9021 140 9031 165
rect 8986 120 9031 140
rect 8986 95 8996 120
rect 9021 95 9031 120
rect 8986 85 9031 95
rect 9046 165 9091 185
rect 9046 140 9056 165
rect 9081 140 9091 165
rect 9046 120 9091 140
rect 9046 95 9056 120
rect 9081 95 9091 120
rect 9046 85 9091 95
rect 9106 165 9151 185
rect 9106 140 9116 165
rect 9141 140 9151 165
rect 9106 120 9151 140
rect 9106 95 9116 120
rect 9141 95 9151 120
rect 9106 85 9151 95
rect 9166 165 9211 185
rect 9166 140 9176 165
rect 9201 140 9211 165
rect 9166 120 9211 140
rect 9166 95 9176 120
rect 9201 95 9211 120
rect 9166 85 9211 95
rect 9226 165 9276 185
rect 9226 140 9241 165
rect 9266 140 9276 165
rect 9226 120 9276 140
rect 9226 95 9241 120
rect 9266 95 9276 120
rect 9226 85 9276 95
rect 9291 165 9336 185
rect 9291 140 9301 165
rect 9326 140 9336 165
rect 9291 120 9336 140
rect 9291 95 9301 120
rect 9326 95 9336 120
rect 9291 85 9336 95
rect 9351 165 9396 185
rect 9351 140 9361 165
rect 9386 140 9396 165
rect 9351 120 9396 140
rect 9351 95 9361 120
rect 9386 95 9396 120
rect 9351 85 9396 95
rect 9411 165 9456 185
rect 9411 140 9421 165
rect 9446 140 9456 165
rect 9411 120 9456 140
rect 9411 95 9421 120
rect 9446 95 9456 120
rect 9411 85 9456 95
rect 9471 165 9521 185
rect 9471 140 9486 165
rect 9511 140 9521 165
rect 9471 120 9521 140
rect 9471 95 9486 120
rect 9511 95 9521 120
rect 9471 85 9521 95
rect 9536 165 9581 185
rect 9536 140 9546 165
rect 9571 140 9581 165
rect 9536 120 9581 140
rect 9536 95 9546 120
rect 9571 95 9581 120
rect 9536 85 9581 95
rect 9596 165 9641 185
rect 9596 140 9606 165
rect 9631 140 9641 165
rect 9596 120 9641 140
rect 9596 95 9606 120
rect 9631 95 9641 120
rect 9596 85 9641 95
rect 9656 165 9701 185
rect 9656 140 9666 165
rect 9691 140 9701 165
rect 9656 120 9701 140
rect 9656 95 9666 120
rect 9691 95 9701 120
rect 9656 85 9701 95
rect 9716 165 9766 185
rect 9716 140 9731 165
rect 9756 140 9766 165
rect 9716 120 9766 140
rect 9716 95 9731 120
rect 9756 95 9766 120
rect 9716 85 9766 95
rect 9781 165 9826 185
rect 9781 140 9791 165
rect 9816 140 9826 165
rect 9781 120 9826 140
rect 9781 95 9791 120
rect 9816 95 9826 120
rect 9781 85 9826 95
rect 9841 165 9886 185
rect 9841 140 9851 165
rect 9876 140 9886 165
rect 9841 120 9886 140
rect 9841 95 9851 120
rect 9876 95 9886 120
rect 9841 85 9886 95
rect 9901 165 9946 185
rect 9901 140 9911 165
rect 9936 140 9946 165
rect 9901 120 9946 140
rect 9901 95 9911 120
rect 9936 95 9946 120
rect 9901 85 9946 95
rect 9961 165 10006 185
rect 9961 140 9971 165
rect 9996 140 10006 165
rect 9961 120 10006 140
rect 9961 95 9971 120
rect 9996 95 10006 120
rect 9961 85 10006 95
rect 10021 165 10066 185
rect 10021 140 10031 165
rect 10056 140 10066 165
rect 10021 120 10066 140
rect 10021 95 10031 120
rect 10056 95 10066 120
rect 10021 85 10066 95
rect 10081 165 10126 185
rect 10081 140 10091 165
rect 10116 140 10126 165
rect 10081 120 10126 140
rect 10081 95 10091 120
rect 10116 95 10126 120
rect 10081 85 10126 95
rect 10141 165 10186 185
rect 10141 140 10151 165
rect 10176 140 10186 165
rect 10141 120 10186 140
rect 10141 95 10151 120
rect 10176 95 10186 120
rect 10141 85 10186 95
rect 10201 165 10251 185
rect 10201 140 10216 165
rect 10241 140 10251 165
rect 10201 120 10251 140
rect 10201 95 10216 120
rect 10241 95 10251 120
rect 10201 85 10251 95
rect 10266 165 10311 185
rect 10266 140 10276 165
rect 10301 140 10311 165
rect 10266 120 10311 140
rect 10266 95 10276 120
rect 10301 95 10311 120
rect 10266 85 10311 95
rect 10326 165 10371 185
rect 10326 140 10336 165
rect 10361 140 10371 165
rect 10326 120 10371 140
rect 10326 95 10336 120
rect 10361 95 10371 120
rect 10326 85 10371 95
rect 10386 165 10431 185
rect 10386 140 10396 165
rect 10421 140 10431 165
rect 10386 120 10431 140
rect 10386 95 10396 120
rect 10421 95 10431 120
rect 10386 85 10431 95
rect 10446 165 10491 185
rect 10446 140 10456 165
rect 10481 140 10491 165
rect 10446 120 10491 140
rect 10446 95 10456 120
rect 10481 95 10491 120
rect 10446 85 10491 95
rect 10506 165 10551 185
rect 10506 140 10516 165
rect 10541 140 10551 165
rect 10506 120 10551 140
rect 10506 95 10516 120
rect 10541 95 10551 120
rect 10506 85 10551 95
rect 10566 165 10611 185
rect 10566 140 10576 165
rect 10601 140 10611 165
rect 10566 120 10611 140
rect 10566 95 10576 120
rect 10601 95 10611 120
rect 10566 85 10611 95
rect 10626 165 10671 185
rect 10626 140 10636 165
rect 10661 140 10671 165
rect 10626 120 10671 140
rect 10626 95 10636 120
rect 10661 95 10671 120
rect 10626 85 10671 95
rect 10686 165 10736 185
rect 10686 140 10701 165
rect 10726 140 10736 165
rect 10686 120 10736 140
rect 10686 95 10701 120
rect 10726 95 10736 120
rect 10686 85 10736 95
rect 10751 165 10796 185
rect 10751 140 10761 165
rect 10786 140 10796 165
rect 10751 120 10796 140
rect 10751 95 10761 120
rect 10786 95 10796 120
rect 10751 85 10796 95
rect 10811 165 10856 185
rect 10811 140 10821 165
rect 10846 140 10856 165
rect 10811 120 10856 140
rect 10811 95 10821 120
rect 10846 95 10856 120
rect 10811 85 10856 95
rect 10871 165 10916 185
rect 10871 140 10881 165
rect 10906 140 10916 165
rect 10871 120 10916 140
rect 10871 95 10881 120
rect 10906 95 10916 120
rect 10871 85 10916 95
rect 10931 165 10976 185
rect 10931 140 10941 165
rect 10966 140 10976 165
rect 10931 120 10976 140
rect 10931 95 10941 120
rect 10966 95 10976 120
rect 10931 85 10976 95
rect 10991 165 11036 185
rect 10991 140 11001 165
rect 11026 140 11036 165
rect 10991 120 11036 140
rect 10991 95 11001 120
rect 11026 95 11036 120
rect 10991 85 11036 95
rect 11051 165 11096 185
rect 11051 140 11061 165
rect 11086 140 11096 165
rect 11051 120 11096 140
rect 11051 95 11061 120
rect 11086 95 11096 120
rect 11051 85 11096 95
rect 11111 165 11156 185
rect 11111 140 11121 165
rect 11146 140 11156 165
rect 11111 120 11156 140
rect 11111 95 11121 120
rect 11146 95 11156 120
rect 11111 85 11156 95
rect 11171 165 11221 185
rect 11171 140 11186 165
rect 11211 140 11221 165
rect 11171 120 11221 140
rect 11171 95 11186 120
rect 11211 95 11221 120
rect 11171 85 11221 95
rect 11236 165 11281 185
rect 11236 140 11246 165
rect 11271 140 11281 165
rect 11236 120 11281 140
rect 11236 95 11246 120
rect 11271 95 11281 120
rect 11236 85 11281 95
rect 11296 165 11341 185
rect 11296 140 11306 165
rect 11331 140 11341 165
rect 11296 120 11341 140
rect 11296 95 11306 120
rect 11331 95 11341 120
rect 11296 85 11341 95
rect 11356 165 11401 185
rect 11356 140 11366 165
rect 11391 140 11401 165
rect 11356 120 11401 140
rect 11356 95 11366 120
rect 11391 95 11401 120
rect 11356 85 11401 95
rect 11416 165 11461 185
rect 11416 140 11426 165
rect 11451 140 11461 165
rect 11416 120 11461 140
rect 11416 95 11426 120
rect 11451 95 11461 120
rect 11416 85 11461 95
rect 11476 165 11521 185
rect 11476 140 11486 165
rect 11511 140 11521 165
rect 11476 120 11521 140
rect 11476 95 11486 120
rect 11511 95 11521 120
rect 11476 85 11521 95
rect 11536 165 11581 185
rect 11536 140 11546 165
rect 11571 140 11581 165
rect 11536 120 11581 140
rect 11536 95 11546 120
rect 11571 95 11581 120
rect 11536 85 11581 95
rect 11596 165 11641 185
rect 11596 140 11606 165
rect 11631 140 11641 165
rect 11596 120 11641 140
rect 11596 95 11606 120
rect 11631 95 11641 120
rect 11596 85 11641 95
rect 11656 165 11706 185
rect 11656 140 11671 165
rect 11696 140 11706 165
rect 11656 120 11706 140
rect 11656 95 11671 120
rect 11696 95 11706 120
rect 11656 85 11706 95
rect 11721 165 11766 185
rect 11721 140 11731 165
rect 11756 140 11766 165
rect 11721 120 11766 140
rect 11721 95 11731 120
rect 11756 95 11766 120
rect 11721 85 11766 95
rect 11781 165 11826 185
rect 11781 140 11791 165
rect 11816 140 11826 165
rect 11781 120 11826 140
rect 11781 95 11791 120
rect 11816 95 11826 120
rect 11781 85 11826 95
rect 11841 165 11886 185
rect 11841 140 11851 165
rect 11876 140 11886 165
rect 11841 120 11886 140
rect 11841 95 11851 120
rect 11876 95 11886 120
rect 11841 85 11886 95
rect 11901 165 11946 185
rect 11901 140 11911 165
rect 11936 140 11946 165
rect 11901 120 11946 140
rect 11901 95 11911 120
rect 11936 95 11946 120
rect 11901 85 11946 95
rect 11961 165 12006 185
rect 11961 140 11971 165
rect 11996 140 12006 165
rect 11961 120 12006 140
rect 11961 95 11971 120
rect 11996 95 12006 120
rect 11961 85 12006 95
rect 12021 165 12066 185
rect 12021 140 12031 165
rect 12056 140 12066 165
rect 12021 120 12066 140
rect 12021 95 12031 120
rect 12056 95 12066 120
rect 12021 85 12066 95
rect 12081 165 12126 185
rect 12081 140 12091 165
rect 12116 140 12126 165
rect 12081 120 12126 140
rect 12081 95 12091 120
rect 12116 95 12126 120
rect 12081 85 12126 95
rect 12141 165 12191 185
rect 12141 140 12156 165
rect 12181 140 12191 165
rect 12141 120 12191 140
rect 12141 95 12156 120
rect 12181 95 12191 120
rect 12141 85 12191 95
rect 12206 165 12251 185
rect 12206 140 12216 165
rect 12241 140 12251 165
rect 12206 120 12251 140
rect 12206 95 12216 120
rect 12241 95 12251 120
rect 12206 85 12251 95
rect 12266 165 12311 185
rect 12266 140 12276 165
rect 12301 140 12311 165
rect 12266 120 12311 140
rect 12266 95 12276 120
rect 12301 95 12311 120
rect 12266 85 12311 95
rect 12326 165 12371 185
rect 12326 140 12336 165
rect 12361 140 12371 165
rect 12326 120 12371 140
rect 12326 95 12336 120
rect 12361 95 12371 120
rect 12326 85 12371 95
rect 12386 165 12431 185
rect 12386 140 12396 165
rect 12421 140 12431 165
rect 12386 120 12431 140
rect 12386 95 12396 120
rect 12421 95 12431 120
rect 12386 85 12431 95
rect 12446 165 12491 185
rect 12446 140 12456 165
rect 12481 140 12491 165
rect 12446 120 12491 140
rect 12446 95 12456 120
rect 12481 95 12491 120
rect 12446 85 12491 95
rect 12506 165 12551 185
rect 12506 140 12516 165
rect 12541 140 12551 165
rect 12506 120 12551 140
rect 12506 95 12516 120
rect 12541 95 12551 120
rect 12506 85 12551 95
rect 12566 165 12611 185
rect 12566 140 12576 165
rect 12601 140 12611 165
rect 12566 120 12611 140
rect 12566 95 12576 120
rect 12601 95 12611 120
rect 12566 85 12611 95
rect 12626 165 12676 185
rect 12626 140 12641 165
rect 12666 140 12676 165
rect 12626 120 12676 140
rect 12626 95 12641 120
rect 12666 95 12676 120
rect 12626 85 12676 95
rect 12691 165 12736 185
rect 12691 140 12701 165
rect 12726 140 12736 165
rect 12691 120 12736 140
rect 12691 95 12701 120
rect 12726 95 12736 120
rect 12691 85 12736 95
rect 12751 165 12796 185
rect 12751 140 12761 165
rect 12786 140 12796 165
rect 12751 120 12796 140
rect 12751 95 12761 120
rect 12786 95 12796 120
rect 12751 85 12796 95
rect 12811 165 12856 185
rect 12811 140 12821 165
rect 12846 140 12856 165
rect 12811 120 12856 140
rect 12811 95 12821 120
rect 12846 95 12856 120
rect 12811 85 12856 95
rect 12871 165 12916 185
rect 12871 140 12881 165
rect 12906 140 12916 165
rect 12871 120 12916 140
rect 12871 95 12881 120
rect 12906 95 12916 120
rect 12871 85 12916 95
rect 12931 165 12976 185
rect 12931 140 12941 165
rect 12966 140 12976 165
rect 12931 120 12976 140
rect 12931 95 12941 120
rect 12966 95 12976 120
rect 12931 85 12976 95
rect 12991 165 13036 185
rect 12991 140 13001 165
rect 13026 140 13036 165
rect 12991 120 13036 140
rect 12991 95 13001 120
rect 13026 95 13036 120
rect 12991 85 13036 95
rect 13051 165 13096 185
rect 13051 140 13061 165
rect 13086 140 13096 165
rect 13051 120 13096 140
rect 13051 95 13061 120
rect 13086 95 13096 120
rect 13051 85 13096 95
rect 13111 165 13161 185
rect 13111 140 13126 165
rect 13151 140 13161 165
rect 13111 120 13161 140
rect 13111 95 13126 120
rect 13151 95 13161 120
rect 13111 85 13161 95
rect 13176 165 13221 185
rect 13176 140 13186 165
rect 13211 140 13221 165
rect 13176 120 13221 140
rect 13176 95 13186 120
rect 13211 95 13221 120
rect 13176 85 13221 95
rect 13236 165 13281 185
rect 13236 140 13246 165
rect 13271 140 13281 165
rect 13236 120 13281 140
rect 13236 95 13246 120
rect 13271 95 13281 120
rect 13236 85 13281 95
rect 13296 165 13341 185
rect 13296 140 13306 165
rect 13331 140 13341 165
rect 13296 120 13341 140
rect 13296 95 13306 120
rect 13331 95 13341 120
rect 13296 85 13341 95
rect 13356 165 13401 185
rect 13356 140 13366 165
rect 13391 140 13401 165
rect 13356 120 13401 140
rect 13356 95 13366 120
rect 13391 95 13401 120
rect 13356 85 13401 95
rect 13416 165 13461 185
rect 13416 140 13426 165
rect 13451 140 13461 165
rect 13416 120 13461 140
rect 13416 95 13426 120
rect 13451 95 13461 120
rect 13416 85 13461 95
rect 13476 165 13521 185
rect 13476 140 13486 165
rect 13511 140 13521 165
rect 13476 120 13521 140
rect 13476 95 13486 120
rect 13511 95 13521 120
rect 13476 85 13521 95
rect 13536 165 13581 185
rect 13536 140 13546 165
rect 13571 140 13581 165
rect 13536 120 13581 140
rect 13536 95 13546 120
rect 13571 95 13581 120
rect 13536 85 13581 95
rect 13596 165 13646 185
rect 13596 140 13611 165
rect 13636 140 13646 165
rect 13596 120 13646 140
rect 13596 95 13611 120
rect 13636 95 13646 120
rect 13596 85 13646 95
rect 13661 165 13706 185
rect 13661 140 13671 165
rect 13696 140 13706 165
rect 13661 120 13706 140
rect 13661 95 13671 120
rect 13696 95 13706 120
rect 13661 85 13706 95
rect 13721 165 13766 185
rect 13721 140 13731 165
rect 13756 140 13766 165
rect 13721 120 13766 140
rect 13721 95 13731 120
rect 13756 95 13766 120
rect 13721 85 13766 95
rect 13781 165 13826 185
rect 13781 140 13791 165
rect 13816 140 13826 165
rect 13781 120 13826 140
rect 13781 95 13791 120
rect 13816 95 13826 120
rect 13781 85 13826 95
rect 13841 165 13886 185
rect 13841 140 13851 165
rect 13876 140 13886 165
rect 13841 120 13886 140
rect 13841 95 13851 120
rect 13876 95 13886 120
rect 13841 85 13886 95
rect 13901 165 13946 185
rect 13901 140 13911 165
rect 13936 140 13946 165
rect 13901 120 13946 140
rect 13901 95 13911 120
rect 13936 95 13946 120
rect 13901 85 13946 95
rect 13961 165 14006 185
rect 13961 140 13971 165
rect 13996 140 14006 165
rect 13961 120 14006 140
rect 13961 95 13971 120
rect 13996 95 14006 120
rect 13961 85 14006 95
rect 14021 165 14066 185
rect 14021 140 14031 165
rect 14056 140 14066 165
rect 14021 120 14066 140
rect 14021 95 14031 120
rect 14056 95 14066 120
rect 14021 85 14066 95
rect 14081 165 14131 185
rect 14081 140 14096 165
rect 14121 140 14131 165
rect 14081 120 14131 140
rect 14081 95 14096 120
rect 14121 95 14131 120
rect 14081 85 14131 95
rect 14146 165 14191 185
rect 14146 140 14156 165
rect 14181 140 14191 165
rect 14146 120 14191 140
rect 14146 95 14156 120
rect 14181 95 14191 120
rect 14146 85 14191 95
rect 14206 165 14251 185
rect 14206 140 14216 165
rect 14241 140 14251 165
rect 14206 120 14251 140
rect 14206 95 14216 120
rect 14241 95 14251 120
rect 14206 85 14251 95
rect 14266 165 14311 185
rect 14266 140 14276 165
rect 14301 140 14311 165
rect 14266 120 14311 140
rect 14266 95 14276 120
rect 14301 95 14311 120
rect 14266 85 14311 95
rect 14326 165 14371 185
rect 14326 140 14336 165
rect 14361 140 14371 165
rect 14326 120 14371 140
rect 14326 95 14336 120
rect 14361 95 14371 120
rect 14326 85 14371 95
rect 14386 165 14431 185
rect 14386 140 14396 165
rect 14421 140 14431 165
rect 14386 120 14431 140
rect 14386 95 14396 120
rect 14421 95 14431 120
rect 14386 85 14431 95
rect 14446 165 14491 185
rect 14446 140 14456 165
rect 14481 140 14491 165
rect 14446 120 14491 140
rect 14446 95 14456 120
rect 14481 95 14491 120
rect 14446 85 14491 95
rect 14506 165 14551 185
rect 14506 140 14516 165
rect 14541 140 14551 165
rect 14506 120 14551 140
rect 14506 95 14516 120
rect 14541 95 14551 120
rect 14506 85 14551 95
rect 14566 165 14616 185
rect 14566 140 14581 165
rect 14606 140 14616 165
rect 14566 120 14616 140
rect 14566 95 14581 120
rect 14606 95 14616 120
rect 14566 85 14616 95
rect 14631 165 14676 185
rect 14631 140 14641 165
rect 14666 140 14676 165
rect 14631 120 14676 140
rect 14631 95 14641 120
rect 14666 95 14676 120
rect 14631 85 14676 95
rect 14691 165 14736 185
rect 14691 140 14701 165
rect 14726 140 14736 165
rect 14691 120 14736 140
rect 14691 95 14701 120
rect 14726 95 14736 120
rect 14691 85 14736 95
rect 14751 165 14796 185
rect 14751 140 14761 165
rect 14786 140 14796 165
rect 14751 120 14796 140
rect 14751 95 14761 120
rect 14786 95 14796 120
rect 14751 85 14796 95
rect 14811 165 14856 185
rect 14811 140 14821 165
rect 14846 140 14856 165
rect 14811 120 14856 140
rect 14811 95 14821 120
rect 14846 95 14856 120
rect 14811 85 14856 95
rect 14871 165 14916 185
rect 14871 140 14881 165
rect 14906 140 14916 165
rect 14871 120 14916 140
rect 14871 95 14881 120
rect 14906 95 14916 120
rect 14871 85 14916 95
rect 14931 165 14976 185
rect 14931 140 14941 165
rect 14966 140 14976 165
rect 14931 120 14976 140
rect 14931 95 14941 120
rect 14966 95 14976 120
rect 14931 85 14976 95
rect 14991 165 15036 185
rect 14991 140 15001 165
rect 15026 140 15036 165
rect 14991 120 15036 140
rect 14991 95 15001 120
rect 15026 95 15036 120
rect 14991 85 15036 95
rect 15051 165 15101 185
rect 15051 140 15066 165
rect 15091 140 15101 165
rect 15051 120 15101 140
rect 15051 95 15066 120
rect 15091 95 15101 120
rect 15051 85 15101 95
rect 15116 165 15161 185
rect 15116 140 15126 165
rect 15151 140 15161 165
rect 15116 120 15161 140
rect 15116 95 15126 120
rect 15151 95 15161 120
rect 15116 85 15161 95
rect 15176 165 15221 185
rect 15176 140 15186 165
rect 15211 140 15221 165
rect 15176 120 15221 140
rect 15176 95 15186 120
rect 15211 95 15221 120
rect 15176 85 15221 95
rect 15236 165 15281 185
rect 15236 140 15246 165
rect 15271 140 15281 165
rect 15236 120 15281 140
rect 15236 95 15246 120
rect 15271 95 15281 120
rect 15236 85 15281 95
rect 15296 165 15341 185
rect 15296 140 15306 165
rect 15331 140 15341 165
rect 15296 120 15341 140
rect 15296 95 15306 120
rect 15331 95 15341 120
rect 15296 85 15341 95
rect 15356 165 15401 185
rect 15356 140 15366 165
rect 15391 140 15401 165
rect 15356 120 15401 140
rect 15356 95 15366 120
rect 15391 95 15401 120
rect 15356 85 15401 95
rect 15416 165 15461 185
rect 15416 140 15426 165
rect 15451 140 15461 165
rect 15416 120 15461 140
rect 15416 95 15426 120
rect 15451 95 15461 120
rect 15416 85 15461 95
rect 15476 165 15521 185
rect 15476 140 15486 165
rect 15511 140 15521 165
rect 15476 120 15521 140
rect 15476 95 15486 120
rect 15511 95 15521 120
rect 15476 85 15521 95
rect 15536 165 15586 185
rect 15536 140 15551 165
rect 15576 140 15586 165
rect 15536 120 15586 140
rect 15536 95 15551 120
rect 15576 95 15586 120
rect 15536 85 15586 95
rect 15601 165 15646 185
rect 15601 140 15611 165
rect 15636 140 15646 165
rect 15601 120 15646 140
rect 15601 95 15611 120
rect 15636 95 15646 120
rect 15601 85 15646 95
rect 15661 165 15706 185
rect 15661 140 15671 165
rect 15696 140 15706 165
rect 15661 120 15706 140
rect 15661 95 15671 120
rect 15696 95 15706 120
rect 15661 85 15706 95
rect 15721 165 15766 185
rect 15721 140 15731 165
rect 15756 140 15766 165
rect 15721 120 15766 140
rect 15721 95 15731 120
rect 15756 95 15766 120
rect 15721 85 15766 95
rect 15781 165 15826 185
rect 15781 140 15791 165
rect 15816 140 15826 165
rect 15781 120 15826 140
rect 15781 95 15791 120
rect 15816 95 15826 120
rect 15781 85 15826 95
rect 15841 165 15886 185
rect 15841 140 15851 165
rect 15876 140 15886 165
rect 15841 120 15886 140
rect 15841 95 15851 120
rect 15876 95 15886 120
rect 15841 85 15886 95
rect 15901 165 15946 185
rect 15901 140 15911 165
rect 15936 140 15946 165
rect 15901 120 15946 140
rect 15901 95 15911 120
rect 15936 95 15946 120
rect 15901 85 15946 95
rect 15961 165 16006 185
rect 15961 140 15971 165
rect 15996 140 16006 165
rect 15961 120 16006 140
rect 15961 95 15971 120
rect 15996 95 16006 120
rect 15961 85 16006 95
rect 16021 165 16071 185
rect 16021 140 16036 165
rect 16061 140 16071 165
rect 16021 120 16071 140
rect 16021 95 16036 120
rect 16061 95 16071 120
rect 16021 85 16071 95
rect 16086 165 16131 185
rect 16086 140 16096 165
rect 16121 140 16131 165
rect 16086 120 16131 140
rect 16086 95 16096 120
rect 16121 95 16131 120
rect 16086 85 16131 95
rect 16146 165 16191 185
rect 16146 140 16156 165
rect 16181 140 16191 165
rect 16146 120 16191 140
rect 16146 95 16156 120
rect 16181 95 16191 120
rect 16146 85 16191 95
rect 16206 165 16251 185
rect 16206 140 16216 165
rect 16241 140 16251 165
rect 16206 120 16251 140
rect 16206 95 16216 120
rect 16241 95 16251 120
rect 16206 85 16251 95
rect 16266 165 16311 185
rect 16266 140 16276 165
rect 16301 140 16311 165
rect 16266 120 16311 140
rect 16266 95 16276 120
rect 16301 95 16311 120
rect 16266 85 16311 95
rect 16326 165 16371 185
rect 16326 140 16336 165
rect 16361 140 16371 165
rect 16326 120 16371 140
rect 16326 95 16336 120
rect 16361 95 16371 120
rect 16326 85 16371 95
rect 16386 165 16431 185
rect 16386 140 16396 165
rect 16421 140 16431 165
rect 16386 120 16431 140
rect 16386 95 16396 120
rect 16421 95 16431 120
rect 16386 85 16431 95
rect 16446 165 16491 185
rect 16446 140 16456 165
rect 16481 140 16491 165
rect 16446 120 16491 140
rect 16446 95 16456 120
rect 16481 95 16491 120
rect 16446 85 16491 95
rect 16506 165 16556 185
rect 16506 140 16521 165
rect 16546 140 16556 165
rect 16506 120 16556 140
rect 16506 95 16521 120
rect 16546 95 16556 120
rect 16506 85 16556 95
rect 16571 165 16616 185
rect 16571 140 16581 165
rect 16606 140 16616 165
rect 16571 120 16616 140
rect 16571 95 16581 120
rect 16606 95 16616 120
rect 16571 85 16616 95
rect 16631 165 16676 185
rect 16631 140 16641 165
rect 16666 140 16676 165
rect 16631 120 16676 140
rect 16631 95 16641 120
rect 16666 95 16676 120
rect 16631 85 16676 95
rect 16691 165 16736 185
rect 16691 140 16701 165
rect 16726 140 16736 165
rect 16691 120 16736 140
rect 16691 95 16701 120
rect 16726 95 16736 120
rect 16691 85 16736 95
rect 16751 165 16796 185
rect 16751 140 16761 165
rect 16786 140 16796 165
rect 16751 120 16796 140
rect 16751 95 16761 120
rect 16786 95 16796 120
rect 16751 85 16796 95
rect 16811 165 16856 185
rect 16811 140 16821 165
rect 16846 140 16856 165
rect 16811 120 16856 140
rect 16811 95 16821 120
rect 16846 95 16856 120
rect 16811 85 16856 95
rect 16871 165 16916 185
rect 16871 140 16881 165
rect 16906 140 16916 165
rect 16871 120 16916 140
rect 16871 95 16881 120
rect 16906 95 16916 120
rect 16871 85 16916 95
rect 16931 165 16976 185
rect 16931 140 16941 165
rect 16966 140 16976 165
rect 16931 120 16976 140
rect 16931 95 16941 120
rect 16966 95 16976 120
rect 16931 85 16976 95
rect 16991 165 17041 185
rect 16991 140 17006 165
rect 17031 140 17041 165
rect 16991 120 17041 140
rect 16991 95 17006 120
rect 17031 95 17041 120
rect 16991 85 17041 95
rect 17056 165 17101 185
rect 17056 140 17066 165
rect 17091 140 17101 165
rect 17056 120 17101 140
rect 17056 95 17066 120
rect 17091 95 17101 120
rect 17056 85 17101 95
rect 17116 165 17161 185
rect 17116 140 17126 165
rect 17151 140 17161 165
rect 17116 120 17161 140
rect 17116 95 17126 120
rect 17151 95 17161 120
rect 17116 85 17161 95
rect 17176 165 17221 185
rect 17176 140 17186 165
rect 17211 140 17221 165
rect 17176 120 17221 140
rect 17176 95 17186 120
rect 17211 95 17221 120
rect 17176 85 17221 95
rect 17236 165 17281 185
rect 17236 140 17246 165
rect 17271 140 17281 165
rect 17236 120 17281 140
rect 17236 95 17246 120
rect 17271 95 17281 120
rect 17236 85 17281 95
rect 17296 165 17341 185
rect 17296 140 17306 165
rect 17331 140 17341 165
rect 17296 120 17341 140
rect 17296 95 17306 120
rect 17331 95 17341 120
rect 17296 85 17341 95
rect 17356 165 17401 185
rect 17356 140 17366 165
rect 17391 140 17401 165
rect 17356 120 17401 140
rect 17356 95 17366 120
rect 17391 95 17401 120
rect 17356 85 17401 95
rect 17416 165 17461 185
rect 17416 140 17426 165
rect 17451 140 17461 165
rect 17416 120 17461 140
rect 17416 95 17426 120
rect 17451 95 17461 120
rect 17416 85 17461 95
rect 17476 165 17526 185
rect 17476 140 17491 165
rect 17516 140 17526 165
rect 17476 120 17526 140
rect 17476 95 17491 120
rect 17516 95 17526 120
rect 17476 85 17526 95
rect 17541 165 17586 185
rect 17541 140 17551 165
rect 17576 140 17586 165
rect 17541 120 17586 140
rect 17541 95 17551 120
rect 17576 95 17586 120
rect 17541 85 17586 95
rect 17601 165 17646 185
rect 17601 140 17611 165
rect 17636 140 17646 165
rect 17601 120 17646 140
rect 17601 95 17611 120
rect 17636 95 17646 120
rect 17601 85 17646 95
rect 17661 165 17706 185
rect 17661 140 17671 165
rect 17696 140 17706 165
rect 17661 120 17706 140
rect 17661 95 17671 120
rect 17696 95 17706 120
rect 17661 85 17706 95
rect 17721 165 17766 185
rect 17721 140 17731 165
rect 17756 140 17766 165
rect 17721 120 17766 140
rect 17721 95 17731 120
rect 17756 95 17766 120
rect 17721 85 17766 95
rect 17781 165 17826 185
rect 17781 140 17791 165
rect 17816 140 17826 165
rect 17781 120 17826 140
rect 17781 95 17791 120
rect 17816 95 17826 120
rect 17781 85 17826 95
rect 17841 165 17886 185
rect 17841 140 17851 165
rect 17876 140 17886 165
rect 17841 120 17886 140
rect 17841 95 17851 120
rect 17876 95 17886 120
rect 17841 85 17886 95
rect 17901 165 17946 185
rect 17901 140 17911 165
rect 17936 140 17946 165
rect 17901 120 17946 140
rect 17901 95 17911 120
rect 17936 95 17946 120
rect 17901 85 17946 95
rect 17961 165 18011 185
rect 17961 140 17976 165
rect 18001 140 18011 165
rect 17961 120 18011 140
rect 17961 95 17976 120
rect 18001 95 18011 120
rect 17961 85 18011 95
rect 18026 165 18071 185
rect 18026 140 18036 165
rect 18061 140 18071 165
rect 18026 120 18071 140
rect 18026 95 18036 120
rect 18061 95 18071 120
rect 18026 85 18071 95
rect 18086 165 18131 185
rect 18086 140 18096 165
rect 18121 140 18131 165
rect 18086 120 18131 140
rect 18086 95 18096 120
rect 18121 95 18131 120
rect 18086 85 18131 95
rect 18146 165 18191 185
rect 18146 140 18156 165
rect 18181 140 18191 165
rect 18146 120 18191 140
rect 18146 95 18156 120
rect 18181 95 18191 120
rect 18146 85 18191 95
rect 18206 165 18251 185
rect 18206 140 18216 165
rect 18241 140 18251 165
rect 18206 120 18251 140
rect 18206 95 18216 120
rect 18241 95 18251 120
rect 18206 85 18251 95
rect 18266 165 18311 185
rect 18266 140 18276 165
rect 18301 140 18311 165
rect 18266 120 18311 140
rect 18266 95 18276 120
rect 18301 95 18311 120
rect 18266 85 18311 95
rect 18326 165 18371 185
rect 18326 140 18336 165
rect 18361 140 18371 165
rect 18326 120 18371 140
rect 18326 95 18336 120
rect 18361 95 18371 120
rect 18326 85 18371 95
rect 18386 165 18431 185
rect 18386 140 18396 165
rect 18421 140 18431 165
rect 18386 120 18431 140
rect 18386 95 18396 120
rect 18421 95 18431 120
rect 18386 85 18431 95
rect 18446 165 18496 185
rect 18446 140 18461 165
rect 18486 140 18496 165
rect 18446 120 18496 140
rect 18446 95 18461 120
rect 18486 95 18496 120
rect 18446 85 18496 95
rect 18511 165 18556 185
rect 18511 140 18521 165
rect 18546 140 18556 165
rect 18511 120 18556 140
rect 18511 95 18521 120
rect 18546 95 18556 120
rect 18511 85 18556 95
rect 18571 165 18616 185
rect 18571 140 18581 165
rect 18606 140 18616 165
rect 18571 120 18616 140
rect 18571 95 18581 120
rect 18606 95 18616 120
rect 18571 85 18616 95
rect 18631 165 18676 185
rect 18631 140 18641 165
rect 18666 140 18676 165
rect 18631 120 18676 140
rect 18631 95 18641 120
rect 18666 95 18676 120
rect 18631 85 18676 95
rect 18691 165 18736 185
rect 18691 140 18701 165
rect 18726 140 18736 165
rect 18691 120 18736 140
rect 18691 95 18701 120
rect 18726 95 18736 120
rect 18691 85 18736 95
rect 18751 165 18796 185
rect 18751 140 18761 165
rect 18786 140 18796 165
rect 18751 120 18796 140
rect 18751 95 18761 120
rect 18786 95 18796 120
rect 18751 85 18796 95
rect 18811 165 18856 185
rect 18811 140 18821 165
rect 18846 140 18856 165
rect 18811 120 18856 140
rect 18811 95 18821 120
rect 18846 95 18856 120
rect 18811 85 18856 95
rect 18871 165 18916 185
rect 18871 140 18881 165
rect 18906 140 18916 165
rect 18871 120 18916 140
rect 18871 95 18881 120
rect 18906 95 18916 120
rect 18871 85 18916 95
rect 18931 165 18981 185
rect 18931 140 18946 165
rect 18971 140 18981 165
rect 18931 120 18981 140
rect 18931 95 18946 120
rect 18971 95 18981 120
rect 18931 85 18981 95
rect 18996 165 19041 185
rect 18996 140 19006 165
rect 19031 140 19041 165
rect 18996 120 19041 140
rect 18996 95 19006 120
rect 19031 95 19041 120
rect 18996 85 19041 95
rect 19056 165 19101 185
rect 19056 140 19066 165
rect 19091 140 19101 165
rect 19056 120 19101 140
rect 19056 95 19066 120
rect 19091 95 19101 120
rect 19056 85 19101 95
rect 19116 165 19161 185
rect 19116 140 19126 165
rect 19151 140 19161 165
rect 19116 120 19161 140
rect 19116 95 19126 120
rect 19151 95 19161 120
rect 19116 85 19161 95
rect 19176 165 19221 185
rect 19176 140 19186 165
rect 19211 140 19221 165
rect 19176 120 19221 140
rect 19176 95 19186 120
rect 19211 95 19221 120
rect 19176 85 19221 95
rect 19236 165 19281 185
rect 19236 140 19246 165
rect 19271 140 19281 165
rect 19236 120 19281 140
rect 19236 95 19246 120
rect 19271 95 19281 120
rect 19236 85 19281 95
rect 19296 165 19341 185
rect 19296 140 19306 165
rect 19331 140 19341 165
rect 19296 120 19341 140
rect 19296 95 19306 120
rect 19331 95 19341 120
rect 19296 85 19341 95
rect 19356 165 19401 185
rect 19356 140 19366 165
rect 19391 140 19401 165
rect 19356 120 19401 140
rect 19356 95 19366 120
rect 19391 95 19401 120
rect 19356 85 19401 95
rect 19416 165 19466 185
rect 19416 140 19431 165
rect 19456 140 19466 165
rect 19416 120 19466 140
rect 19416 95 19431 120
rect 19456 95 19466 120
rect 19416 85 19466 95
rect 19481 165 19526 185
rect 19481 140 19491 165
rect 19516 140 19526 165
rect 19481 120 19526 140
rect 19481 95 19491 120
rect 19516 95 19526 120
rect 19481 85 19526 95
rect 19541 165 19586 185
rect 19541 140 19551 165
rect 19576 140 19586 165
rect 19541 120 19586 140
rect 19541 95 19551 120
rect 19576 95 19586 120
rect 19541 85 19586 95
rect 19601 165 19646 185
rect 19601 140 19611 165
rect 19636 140 19646 165
rect 19601 120 19646 140
rect 19601 95 19611 120
rect 19636 95 19646 120
rect 19601 85 19646 95
rect 19661 165 19706 185
rect 19661 140 19671 165
rect 19696 140 19706 165
rect 19661 120 19706 140
rect 19661 95 19671 120
rect 19696 95 19706 120
rect 19661 85 19706 95
rect 19721 165 19766 185
rect 19721 140 19731 165
rect 19756 140 19766 165
rect 19721 120 19766 140
rect 19721 95 19731 120
rect 19756 95 19766 120
rect 19721 85 19766 95
rect 19781 165 19826 185
rect 19781 140 19791 165
rect 19816 140 19826 165
rect 19781 120 19826 140
rect 19781 95 19791 120
rect 19816 95 19826 120
rect 19781 85 19826 95
rect 19841 165 19886 185
rect 19841 140 19851 165
rect 19876 140 19886 165
rect 19841 120 19886 140
rect 19841 95 19851 120
rect 19876 95 19886 120
rect 19841 85 19886 95
rect 19901 165 19951 185
rect 19901 140 19916 165
rect 19941 140 19951 165
rect 19901 120 19951 140
rect 19901 95 19916 120
rect 19941 95 19951 120
rect 19901 85 19951 95
rect 19966 165 20011 185
rect 19966 140 19976 165
rect 20001 140 20011 165
rect 19966 120 20011 140
rect 19966 95 19976 120
rect 20001 95 20011 120
rect 19966 85 20011 95
rect 20026 165 20071 185
rect 20026 140 20036 165
rect 20061 140 20071 165
rect 20026 120 20071 140
rect 20026 95 20036 120
rect 20061 95 20071 120
rect 20026 85 20071 95
rect 20086 165 20131 185
rect 20086 140 20096 165
rect 20121 140 20131 165
rect 20086 120 20131 140
rect 20086 95 20096 120
rect 20121 95 20131 120
rect 20086 85 20131 95
rect 20146 165 20191 185
rect 20146 140 20156 165
rect 20181 140 20191 165
rect 20146 120 20191 140
rect 20146 95 20156 120
rect 20181 95 20191 120
rect 20146 85 20191 95
rect 20206 165 20251 185
rect 20206 140 20216 165
rect 20241 140 20251 165
rect 20206 120 20251 140
rect 20206 95 20216 120
rect 20241 95 20251 120
rect 20206 85 20251 95
rect 20266 165 20311 185
rect 20266 140 20276 165
rect 20301 140 20311 165
rect 20266 120 20311 140
rect 20266 95 20276 120
rect 20301 95 20311 120
rect 20266 85 20311 95
rect 20326 165 20371 185
rect 20326 140 20336 165
rect 20361 140 20371 165
rect 20326 120 20371 140
rect 20326 95 20336 120
rect 20361 95 20371 120
rect 20326 85 20371 95
rect 20386 165 20436 185
rect 20386 140 20401 165
rect 20426 140 20436 165
rect 20386 120 20436 140
rect 20386 95 20401 120
rect 20426 95 20436 120
rect 20386 85 20436 95
rect 20451 165 20496 185
rect 20451 140 20461 165
rect 20486 140 20496 165
rect 20451 120 20496 140
rect 20451 95 20461 120
rect 20486 95 20496 120
rect 20451 85 20496 95
rect 20511 165 20556 185
rect 20511 140 20521 165
rect 20546 140 20556 165
rect 20511 120 20556 140
rect 20511 95 20521 120
rect 20546 95 20556 120
rect 20511 85 20556 95
rect 20571 165 20616 185
rect 20571 140 20581 165
rect 20606 140 20616 165
rect 20571 120 20616 140
rect 20571 95 20581 120
rect 20606 95 20616 120
rect 20571 85 20616 95
rect 20631 165 20676 185
rect 20631 140 20641 165
rect 20666 140 20676 165
rect 20631 120 20676 140
rect 20631 95 20641 120
rect 20666 95 20676 120
rect 20631 85 20676 95
rect 20691 165 20736 185
rect 20691 140 20701 165
rect 20726 140 20736 165
rect 20691 120 20736 140
rect 20691 95 20701 120
rect 20726 95 20736 120
rect 20691 85 20736 95
rect 20751 165 20796 185
rect 20751 140 20761 165
rect 20786 140 20796 165
rect 20751 120 20796 140
rect 20751 95 20761 120
rect 20786 95 20796 120
rect 20751 85 20796 95
rect 20811 165 20856 185
rect 20811 140 20821 165
rect 20846 140 20856 165
rect 20811 120 20856 140
rect 20811 95 20821 120
rect 20846 95 20856 120
rect 20811 85 20856 95
rect 20871 165 20921 185
rect 20871 140 20886 165
rect 20911 140 20921 165
rect 20871 120 20921 140
rect 20871 95 20886 120
rect 20911 95 20921 120
rect 20871 85 20921 95
rect 20936 165 20981 185
rect 20936 140 20946 165
rect 20971 140 20981 165
rect 20936 120 20981 140
rect 20936 95 20946 120
rect 20971 95 20981 120
rect 20936 85 20981 95
rect 20996 165 21041 185
rect 20996 140 21006 165
rect 21031 140 21041 165
rect 20996 120 21041 140
rect 20996 95 21006 120
rect 21031 95 21041 120
rect 20996 85 21041 95
rect 21056 165 21101 185
rect 21056 140 21066 165
rect 21091 140 21101 165
rect 21056 120 21101 140
rect 21056 95 21066 120
rect 21091 95 21101 120
rect 21056 85 21101 95
rect 21116 165 21156 185
rect 21116 140 21126 165
rect 21151 140 21156 165
rect 21116 120 21156 140
rect 21116 95 21126 120
rect 21151 95 21156 120
rect 21116 85 21156 95
rect -40 -585 0 -575
rect -40 -610 -35 -585
rect -10 -610 0 -585
rect -40 -630 0 -610
rect -40 -655 -35 -630
rect -10 -655 0 -630
rect -40 -675 0 -655
rect -40 -700 -35 -675
rect -10 -700 0 -675
rect -40 -725 0 -700
rect -40 -750 -35 -725
rect -10 -750 0 -725
rect -40 -770 0 -750
rect 15 -585 60 -575
rect 15 -610 25 -585
rect 50 -610 60 -585
rect 15 -630 60 -610
rect 15 -655 25 -630
rect 50 -655 60 -630
rect 15 -675 60 -655
rect 15 -700 25 -675
rect 50 -700 60 -675
rect 15 -725 60 -700
rect 15 -750 25 -725
rect 50 -750 60 -725
rect 15 -770 60 -750
rect 75 -585 120 -575
rect 75 -610 85 -585
rect 110 -610 120 -585
rect 75 -630 120 -610
rect 75 -655 85 -630
rect 110 -655 120 -630
rect 75 -675 120 -655
rect 75 -700 85 -675
rect 110 -700 120 -675
rect 75 -725 120 -700
rect 75 -750 85 -725
rect 110 -750 120 -725
rect 75 -770 120 -750
rect 135 -585 180 -575
rect 135 -610 145 -585
rect 170 -610 180 -585
rect 135 -630 180 -610
rect 135 -655 145 -630
rect 170 -655 180 -630
rect 135 -675 180 -655
rect 135 -700 145 -675
rect 170 -700 180 -675
rect 135 -725 180 -700
rect 135 -750 145 -725
rect 170 -750 180 -725
rect 135 -770 180 -750
rect 195 -585 240 -575
rect 195 -610 205 -585
rect 230 -610 240 -585
rect 195 -630 240 -610
rect 195 -655 205 -630
rect 230 -655 240 -630
rect 195 -675 240 -655
rect 195 -700 205 -675
rect 230 -700 240 -675
rect 195 -725 240 -700
rect 195 -750 205 -725
rect 230 -750 240 -725
rect 195 -770 240 -750
rect 255 -585 300 -575
rect 255 -610 265 -585
rect 290 -610 300 -585
rect 255 -630 300 -610
rect 255 -655 265 -630
rect 290 -655 300 -630
rect 255 -675 300 -655
rect 255 -700 265 -675
rect 290 -700 300 -675
rect 255 -725 300 -700
rect 255 -750 265 -725
rect 290 -750 300 -725
rect 255 -770 300 -750
rect 315 -585 360 -575
rect 315 -610 325 -585
rect 350 -610 360 -585
rect 315 -630 360 -610
rect 315 -655 325 -630
rect 350 -655 360 -630
rect 315 -675 360 -655
rect 315 -700 325 -675
rect 350 -700 360 -675
rect 315 -725 360 -700
rect 315 -750 325 -725
rect 350 -750 360 -725
rect 315 -770 360 -750
rect 375 -585 420 -575
rect 375 -610 385 -585
rect 410 -610 420 -585
rect 375 -630 420 -610
rect 375 -655 385 -630
rect 410 -655 420 -630
rect 375 -675 420 -655
rect 375 -700 385 -675
rect 410 -700 420 -675
rect 375 -725 420 -700
rect 375 -750 385 -725
rect 410 -750 420 -725
rect 375 -770 420 -750
rect 435 -585 480 -575
rect 435 -610 445 -585
rect 470 -610 480 -585
rect 435 -630 480 -610
rect 435 -655 445 -630
rect 470 -655 480 -630
rect 435 -675 480 -655
rect 435 -700 445 -675
rect 470 -700 480 -675
rect 435 -725 480 -700
rect 435 -750 445 -725
rect 470 -750 480 -725
rect 435 -770 480 -750
rect 495 -585 540 -575
rect 495 -610 505 -585
rect 530 -610 540 -585
rect 495 -630 540 -610
rect 495 -655 505 -630
rect 530 -655 540 -630
rect 495 -675 540 -655
rect 495 -700 505 -675
rect 530 -700 540 -675
rect 495 -725 540 -700
rect 495 -750 505 -725
rect 530 -750 540 -725
rect 495 -770 540 -750
rect 555 -585 600 -575
rect 555 -610 565 -585
rect 590 -610 600 -585
rect 555 -630 600 -610
rect 555 -655 565 -630
rect 590 -655 600 -630
rect 555 -675 600 -655
rect 555 -700 565 -675
rect 590 -700 600 -675
rect 555 -725 600 -700
rect 555 -750 565 -725
rect 590 -750 600 -725
rect 555 -770 600 -750
rect 615 -585 660 -575
rect 615 -610 625 -585
rect 650 -610 660 -585
rect 615 -630 660 -610
rect 615 -655 625 -630
rect 650 -655 660 -630
rect 615 -675 660 -655
rect 615 -700 625 -675
rect 650 -700 660 -675
rect 615 -725 660 -700
rect 615 -750 625 -725
rect 650 -750 660 -725
rect 615 -770 660 -750
rect 675 -585 720 -575
rect 675 -610 685 -585
rect 710 -610 720 -585
rect 675 -630 720 -610
rect 675 -655 685 -630
rect 710 -655 720 -630
rect 675 -675 720 -655
rect 675 -700 685 -675
rect 710 -700 720 -675
rect 675 -725 720 -700
rect 675 -750 685 -725
rect 710 -750 720 -725
rect 675 -770 720 -750
rect 735 -585 780 -575
rect 735 -610 745 -585
rect 770 -610 780 -585
rect 735 -630 780 -610
rect 735 -655 745 -630
rect 770 -655 780 -630
rect 735 -675 780 -655
rect 735 -700 745 -675
rect 770 -700 780 -675
rect 735 -725 780 -700
rect 735 -750 745 -725
rect 770 -750 780 -725
rect 735 -770 780 -750
rect 795 -585 840 -575
rect 795 -610 805 -585
rect 830 -610 840 -585
rect 795 -630 840 -610
rect 795 -655 805 -630
rect 830 -655 840 -630
rect 795 -675 840 -655
rect 795 -700 805 -675
rect 830 -700 840 -675
rect 795 -725 840 -700
rect 795 -750 805 -725
rect 830 -750 840 -725
rect 795 -770 840 -750
rect 855 -585 900 -575
rect 855 -610 865 -585
rect 890 -610 900 -585
rect 855 -630 900 -610
rect 855 -655 865 -630
rect 890 -655 900 -630
rect 855 -675 900 -655
rect 855 -700 865 -675
rect 890 -700 900 -675
rect 855 -725 900 -700
rect 855 -750 865 -725
rect 890 -750 900 -725
rect 855 -770 900 -750
rect 915 -585 960 -575
rect 915 -610 925 -585
rect 950 -610 960 -585
rect 915 -630 960 -610
rect 915 -655 925 -630
rect 950 -655 960 -630
rect 915 -675 960 -655
rect 915 -700 925 -675
rect 950 -700 960 -675
rect 915 -725 960 -700
rect 915 -750 925 -725
rect 950 -750 960 -725
rect 915 -770 960 -750
rect 975 -585 1020 -575
rect 975 -610 985 -585
rect 1010 -610 1020 -585
rect 975 -630 1020 -610
rect 975 -655 985 -630
rect 1010 -655 1020 -630
rect 975 -675 1020 -655
rect 975 -700 985 -675
rect 1010 -700 1020 -675
rect 975 -725 1020 -700
rect 975 -750 985 -725
rect 1010 -750 1020 -725
rect 975 -770 1020 -750
rect 1035 -585 1080 -575
rect 1035 -610 1045 -585
rect 1070 -610 1080 -585
rect 1035 -630 1080 -610
rect 1035 -655 1045 -630
rect 1070 -655 1080 -630
rect 1035 -675 1080 -655
rect 1035 -700 1045 -675
rect 1070 -700 1080 -675
rect 1035 -725 1080 -700
rect 1035 -750 1045 -725
rect 1070 -750 1080 -725
rect 1035 -770 1080 -750
rect 1095 -585 1140 -575
rect 1095 -610 1105 -585
rect 1130 -610 1140 -585
rect 1095 -630 1140 -610
rect 1095 -655 1105 -630
rect 1130 -655 1140 -630
rect 1095 -675 1140 -655
rect 1095 -700 1105 -675
rect 1130 -700 1140 -675
rect 1095 -725 1140 -700
rect 1095 -750 1105 -725
rect 1130 -750 1140 -725
rect 1095 -770 1140 -750
rect 1155 -585 1200 -575
rect 1155 -610 1165 -585
rect 1190 -610 1200 -585
rect 1155 -630 1200 -610
rect 1155 -655 1165 -630
rect 1190 -655 1200 -630
rect 1155 -675 1200 -655
rect 1155 -700 1165 -675
rect 1190 -700 1200 -675
rect 1155 -725 1200 -700
rect 1155 -750 1165 -725
rect 1190 -750 1200 -725
rect 1155 -770 1200 -750
rect 1215 -585 1260 -575
rect 1215 -610 1225 -585
rect 1250 -610 1260 -585
rect 1215 -630 1260 -610
rect 1215 -655 1225 -630
rect 1250 -655 1260 -630
rect 1215 -675 1260 -655
rect 1215 -700 1225 -675
rect 1250 -700 1260 -675
rect 1215 -725 1260 -700
rect 1215 -750 1225 -725
rect 1250 -750 1260 -725
rect 1215 -770 1260 -750
rect 1275 -585 1320 -575
rect 1275 -610 1285 -585
rect 1310 -610 1320 -585
rect 1275 -630 1320 -610
rect 1275 -655 1285 -630
rect 1310 -655 1320 -630
rect 1275 -675 1320 -655
rect 1275 -700 1285 -675
rect 1310 -700 1320 -675
rect 1275 -725 1320 -700
rect 1275 -750 1285 -725
rect 1310 -750 1320 -725
rect 1275 -770 1320 -750
rect 1335 -585 1380 -575
rect 1335 -610 1345 -585
rect 1370 -610 1380 -585
rect 1335 -630 1380 -610
rect 1335 -655 1345 -630
rect 1370 -655 1380 -630
rect 1335 -675 1380 -655
rect 1335 -700 1345 -675
rect 1370 -700 1380 -675
rect 1335 -725 1380 -700
rect 1335 -750 1345 -725
rect 1370 -750 1380 -725
rect 1335 -770 1380 -750
rect 1395 -585 1440 -575
rect 1395 -610 1405 -585
rect 1430 -610 1440 -585
rect 1395 -630 1440 -610
rect 1395 -655 1405 -630
rect 1430 -655 1440 -630
rect 1395 -675 1440 -655
rect 1395 -700 1405 -675
rect 1430 -700 1440 -675
rect 1395 -725 1440 -700
rect 1395 -750 1405 -725
rect 1430 -750 1440 -725
rect 1395 -770 1440 -750
rect 1455 -585 1500 -575
rect 1455 -610 1465 -585
rect 1490 -610 1500 -585
rect 1455 -630 1500 -610
rect 1455 -655 1465 -630
rect 1490 -655 1500 -630
rect 1455 -675 1500 -655
rect 1455 -700 1465 -675
rect 1490 -700 1500 -675
rect 1455 -725 1500 -700
rect 1455 -750 1465 -725
rect 1490 -750 1500 -725
rect 1455 -770 1500 -750
rect 1515 -585 1560 -575
rect 1515 -610 1525 -585
rect 1550 -610 1560 -585
rect 1515 -630 1560 -610
rect 1515 -655 1525 -630
rect 1550 -655 1560 -630
rect 1515 -675 1560 -655
rect 1515 -700 1525 -675
rect 1550 -700 1560 -675
rect 1515 -725 1560 -700
rect 1515 -750 1525 -725
rect 1550 -750 1560 -725
rect 1515 -770 1560 -750
rect 1575 -585 1620 -575
rect 1575 -610 1585 -585
rect 1610 -610 1620 -585
rect 1575 -630 1620 -610
rect 1575 -655 1585 -630
rect 1610 -655 1620 -630
rect 1575 -675 1620 -655
rect 1575 -700 1585 -675
rect 1610 -700 1620 -675
rect 1575 -725 1620 -700
rect 1575 -750 1585 -725
rect 1610 -750 1620 -725
rect 1575 -770 1620 -750
rect 1635 -585 1680 -575
rect 1635 -610 1645 -585
rect 1670 -610 1680 -585
rect 1635 -630 1680 -610
rect 1635 -655 1645 -630
rect 1670 -655 1680 -630
rect 1635 -675 1680 -655
rect 1635 -700 1645 -675
rect 1670 -700 1680 -675
rect 1635 -725 1680 -700
rect 1635 -750 1645 -725
rect 1670 -750 1680 -725
rect 1635 -770 1680 -750
rect 1695 -585 1740 -575
rect 1695 -610 1705 -585
rect 1730 -610 1740 -585
rect 1695 -630 1740 -610
rect 1695 -655 1705 -630
rect 1730 -655 1740 -630
rect 1695 -675 1740 -655
rect 1695 -700 1705 -675
rect 1730 -700 1740 -675
rect 1695 -725 1740 -700
rect 1695 -750 1705 -725
rect 1730 -750 1740 -725
rect 1695 -770 1740 -750
rect 1755 -585 1800 -575
rect 1755 -610 1765 -585
rect 1790 -610 1800 -585
rect 1755 -630 1800 -610
rect 1755 -655 1765 -630
rect 1790 -655 1800 -630
rect 1755 -675 1800 -655
rect 1755 -700 1765 -675
rect 1790 -700 1800 -675
rect 1755 -725 1800 -700
rect 1755 -750 1765 -725
rect 1790 -750 1800 -725
rect 1755 -770 1800 -750
rect 1815 -585 1860 -575
rect 1815 -610 1825 -585
rect 1850 -610 1860 -585
rect 1815 -630 1860 -610
rect 1815 -655 1825 -630
rect 1850 -655 1860 -630
rect 1815 -675 1860 -655
rect 1815 -700 1825 -675
rect 1850 -700 1860 -675
rect 1815 -725 1860 -700
rect 1815 -750 1825 -725
rect 1850 -750 1860 -725
rect 1815 -770 1860 -750
rect 1875 -585 1920 -575
rect 1875 -610 1885 -585
rect 1910 -610 1920 -585
rect 1875 -630 1920 -610
rect 1875 -655 1885 -630
rect 1910 -655 1920 -630
rect 1875 -675 1920 -655
rect 1875 -700 1885 -675
rect 1910 -700 1920 -675
rect 1875 -725 1920 -700
rect 1875 -750 1885 -725
rect 1910 -750 1920 -725
rect 1875 -770 1920 -750
rect 1935 -585 1980 -575
rect 1935 -610 1945 -585
rect 1970 -610 1980 -585
rect 1935 -630 1980 -610
rect 1935 -655 1945 -630
rect 1970 -655 1980 -630
rect 1935 -675 1980 -655
rect 1935 -700 1945 -675
rect 1970 -700 1980 -675
rect 1935 -725 1980 -700
rect 1935 -750 1945 -725
rect 1970 -750 1980 -725
rect 1935 -770 1980 -750
rect 1995 -585 2040 -575
rect 1995 -610 2005 -585
rect 2030 -610 2040 -585
rect 1995 -630 2040 -610
rect 1995 -655 2005 -630
rect 2030 -655 2040 -630
rect 1995 -675 2040 -655
rect 1995 -700 2005 -675
rect 2030 -700 2040 -675
rect 1995 -725 2040 -700
rect 1995 -750 2005 -725
rect 2030 -750 2040 -725
rect 1995 -770 2040 -750
rect 2055 -585 2100 -575
rect 2055 -610 2065 -585
rect 2090 -610 2100 -585
rect 2055 -630 2100 -610
rect 2055 -655 2065 -630
rect 2090 -655 2100 -630
rect 2055 -675 2100 -655
rect 2055 -700 2065 -675
rect 2090 -700 2100 -675
rect 2055 -725 2100 -700
rect 2055 -750 2065 -725
rect 2090 -750 2100 -725
rect 2055 -770 2100 -750
rect 2115 -585 2160 -575
rect 2115 -610 2125 -585
rect 2150 -610 2160 -585
rect 2115 -630 2160 -610
rect 2115 -655 2125 -630
rect 2150 -655 2160 -630
rect 2115 -675 2160 -655
rect 2115 -700 2125 -675
rect 2150 -700 2160 -675
rect 2115 -725 2160 -700
rect 2115 -750 2125 -725
rect 2150 -750 2160 -725
rect 2115 -770 2160 -750
rect 2175 -585 2220 -575
rect 2175 -610 2185 -585
rect 2210 -610 2220 -585
rect 2175 -630 2220 -610
rect 2175 -655 2185 -630
rect 2210 -655 2220 -630
rect 2175 -675 2220 -655
rect 2175 -700 2185 -675
rect 2210 -700 2220 -675
rect 2175 -725 2220 -700
rect 2175 -750 2185 -725
rect 2210 -750 2220 -725
rect 2175 -770 2220 -750
rect 2235 -585 2280 -575
rect 2235 -610 2245 -585
rect 2270 -610 2280 -585
rect 2235 -630 2280 -610
rect 2235 -655 2245 -630
rect 2270 -655 2280 -630
rect 2235 -675 2280 -655
rect 2235 -700 2245 -675
rect 2270 -700 2280 -675
rect 2235 -725 2280 -700
rect 2235 -750 2245 -725
rect 2270 -750 2280 -725
rect 2235 -770 2280 -750
rect 2295 -585 2340 -575
rect 2295 -610 2305 -585
rect 2330 -610 2340 -585
rect 2295 -630 2340 -610
rect 2295 -655 2305 -630
rect 2330 -655 2340 -630
rect 2295 -675 2340 -655
rect 2295 -700 2305 -675
rect 2330 -700 2340 -675
rect 2295 -725 2340 -700
rect 2295 -750 2305 -725
rect 2330 -750 2340 -725
rect 2295 -770 2340 -750
rect 2355 -585 2400 -575
rect 2355 -610 2365 -585
rect 2390 -610 2400 -585
rect 2355 -630 2400 -610
rect 2355 -655 2365 -630
rect 2390 -655 2400 -630
rect 2355 -675 2400 -655
rect 2355 -700 2365 -675
rect 2390 -700 2400 -675
rect 2355 -725 2400 -700
rect 2355 -750 2365 -725
rect 2390 -750 2400 -725
rect 2355 -770 2400 -750
rect 2415 -585 2460 -575
rect 2415 -610 2425 -585
rect 2450 -610 2460 -585
rect 2415 -630 2460 -610
rect 2415 -655 2425 -630
rect 2450 -655 2460 -630
rect 2415 -675 2460 -655
rect 2415 -700 2425 -675
rect 2450 -700 2460 -675
rect 2415 -725 2460 -700
rect 2415 -750 2425 -725
rect 2450 -750 2460 -725
rect 2415 -770 2460 -750
rect 2475 -585 2520 -575
rect 2475 -610 2485 -585
rect 2510 -610 2520 -585
rect 2475 -630 2520 -610
rect 2475 -655 2485 -630
rect 2510 -655 2520 -630
rect 2475 -675 2520 -655
rect 2475 -700 2485 -675
rect 2510 -700 2520 -675
rect 2475 -725 2520 -700
rect 2475 -750 2485 -725
rect 2510 -750 2520 -725
rect 2475 -770 2520 -750
rect 2535 -585 2580 -575
rect 2535 -610 2545 -585
rect 2570 -610 2580 -585
rect 2535 -630 2580 -610
rect 2535 -655 2545 -630
rect 2570 -655 2580 -630
rect 2535 -675 2580 -655
rect 2535 -700 2545 -675
rect 2570 -700 2580 -675
rect 2535 -725 2580 -700
rect 2535 -750 2545 -725
rect 2570 -750 2580 -725
rect 2535 -770 2580 -750
rect 2595 -585 2640 -575
rect 2595 -610 2605 -585
rect 2630 -610 2640 -585
rect 2595 -630 2640 -610
rect 2595 -655 2605 -630
rect 2630 -655 2640 -630
rect 2595 -675 2640 -655
rect 2595 -700 2605 -675
rect 2630 -700 2640 -675
rect 2595 -725 2640 -700
rect 2595 -750 2605 -725
rect 2630 -750 2640 -725
rect 2595 -770 2640 -750
rect 2655 -585 2700 -575
rect 2655 -610 2665 -585
rect 2690 -610 2700 -585
rect 2655 -630 2700 -610
rect 2655 -655 2665 -630
rect 2690 -655 2700 -630
rect 2655 -675 2700 -655
rect 2655 -700 2665 -675
rect 2690 -700 2700 -675
rect 2655 -725 2700 -700
rect 2655 -750 2665 -725
rect 2690 -750 2700 -725
rect 2655 -770 2700 -750
rect 2715 -585 2760 -575
rect 2715 -610 2725 -585
rect 2750 -610 2760 -585
rect 2715 -630 2760 -610
rect 2715 -655 2725 -630
rect 2750 -655 2760 -630
rect 2715 -675 2760 -655
rect 2715 -700 2725 -675
rect 2750 -700 2760 -675
rect 2715 -725 2760 -700
rect 2715 -750 2725 -725
rect 2750 -750 2760 -725
rect 2715 -770 2760 -750
rect 2775 -585 2820 -575
rect 2775 -610 2785 -585
rect 2810 -610 2820 -585
rect 2775 -630 2820 -610
rect 2775 -655 2785 -630
rect 2810 -655 2820 -630
rect 2775 -675 2820 -655
rect 2775 -700 2785 -675
rect 2810 -700 2820 -675
rect 2775 -725 2820 -700
rect 2775 -750 2785 -725
rect 2810 -750 2820 -725
rect 2775 -770 2820 -750
rect 2835 -585 2880 -575
rect 2835 -610 2845 -585
rect 2870 -610 2880 -585
rect 2835 -630 2880 -610
rect 2835 -655 2845 -630
rect 2870 -655 2880 -630
rect 2835 -675 2880 -655
rect 2835 -700 2845 -675
rect 2870 -700 2880 -675
rect 2835 -725 2880 -700
rect 2835 -750 2845 -725
rect 2870 -750 2880 -725
rect 2835 -770 2880 -750
rect 2895 -585 2940 -575
rect 2895 -610 2905 -585
rect 2930 -610 2940 -585
rect 2895 -630 2940 -610
rect 2895 -655 2905 -630
rect 2930 -655 2940 -630
rect 2895 -675 2940 -655
rect 2895 -700 2905 -675
rect 2930 -700 2940 -675
rect 2895 -725 2940 -700
rect 2895 -750 2905 -725
rect 2930 -750 2940 -725
rect 2895 -770 2940 -750
rect 2955 -585 3000 -575
rect 2955 -610 2965 -585
rect 2990 -610 3000 -585
rect 2955 -630 3000 -610
rect 2955 -655 2965 -630
rect 2990 -655 3000 -630
rect 2955 -675 3000 -655
rect 2955 -700 2965 -675
rect 2990 -700 3000 -675
rect 2955 -725 3000 -700
rect 2955 -750 2965 -725
rect 2990 -750 3000 -725
rect 2955 -770 3000 -750
rect 3015 -585 3060 -575
rect 3015 -610 3025 -585
rect 3050 -610 3060 -585
rect 3015 -630 3060 -610
rect 3015 -655 3025 -630
rect 3050 -655 3060 -630
rect 3015 -675 3060 -655
rect 3015 -700 3025 -675
rect 3050 -700 3060 -675
rect 3015 -725 3060 -700
rect 3015 -750 3025 -725
rect 3050 -750 3060 -725
rect 3015 -770 3060 -750
rect 3075 -585 3120 -575
rect 3075 -610 3085 -585
rect 3110 -610 3120 -585
rect 3075 -630 3120 -610
rect 3075 -655 3085 -630
rect 3110 -655 3120 -630
rect 3075 -675 3120 -655
rect 3075 -700 3085 -675
rect 3110 -700 3120 -675
rect 3075 -725 3120 -700
rect 3075 -750 3085 -725
rect 3110 -750 3120 -725
rect 3075 -770 3120 -750
rect 3135 -585 3180 -575
rect 3135 -610 3145 -585
rect 3170 -610 3180 -585
rect 3135 -630 3180 -610
rect 3135 -655 3145 -630
rect 3170 -655 3180 -630
rect 3135 -675 3180 -655
rect 3135 -700 3145 -675
rect 3170 -700 3180 -675
rect 3135 -725 3180 -700
rect 3135 -750 3145 -725
rect 3170 -750 3180 -725
rect 3135 -770 3180 -750
rect 3195 -585 3240 -575
rect 3195 -610 3205 -585
rect 3230 -610 3240 -585
rect 3195 -630 3240 -610
rect 3195 -655 3205 -630
rect 3230 -655 3240 -630
rect 3195 -675 3240 -655
rect 3195 -700 3205 -675
rect 3230 -700 3240 -675
rect 3195 -725 3240 -700
rect 3195 -750 3205 -725
rect 3230 -750 3240 -725
rect 3195 -770 3240 -750
rect 3255 -585 3300 -575
rect 3255 -610 3265 -585
rect 3290 -610 3300 -585
rect 3255 -630 3300 -610
rect 3255 -655 3265 -630
rect 3290 -655 3300 -630
rect 3255 -675 3300 -655
rect 3255 -700 3265 -675
rect 3290 -700 3300 -675
rect 3255 -725 3300 -700
rect 3255 -750 3265 -725
rect 3290 -750 3300 -725
rect 3255 -770 3300 -750
rect 3315 -585 3360 -575
rect 3315 -610 3325 -585
rect 3350 -610 3360 -585
rect 3315 -630 3360 -610
rect 3315 -655 3325 -630
rect 3350 -655 3360 -630
rect 3315 -675 3360 -655
rect 3315 -700 3325 -675
rect 3350 -700 3360 -675
rect 3315 -725 3360 -700
rect 3315 -750 3325 -725
rect 3350 -750 3360 -725
rect 3315 -770 3360 -750
rect 3375 -585 3420 -575
rect 3375 -610 3385 -585
rect 3410 -610 3420 -585
rect 3375 -630 3420 -610
rect 3375 -655 3385 -630
rect 3410 -655 3420 -630
rect 3375 -675 3420 -655
rect 3375 -700 3385 -675
rect 3410 -700 3420 -675
rect 3375 -725 3420 -700
rect 3375 -750 3385 -725
rect 3410 -750 3420 -725
rect 3375 -770 3420 -750
rect 3435 -585 3480 -575
rect 3435 -610 3445 -585
rect 3470 -610 3480 -585
rect 3435 -630 3480 -610
rect 3435 -655 3445 -630
rect 3470 -655 3480 -630
rect 3435 -675 3480 -655
rect 3435 -700 3445 -675
rect 3470 -700 3480 -675
rect 3435 -725 3480 -700
rect 3435 -750 3445 -725
rect 3470 -750 3480 -725
rect 3435 -770 3480 -750
rect 3495 -585 3540 -575
rect 3495 -610 3505 -585
rect 3530 -610 3540 -585
rect 3495 -630 3540 -610
rect 3495 -655 3505 -630
rect 3530 -655 3540 -630
rect 3495 -675 3540 -655
rect 3495 -700 3505 -675
rect 3530 -700 3540 -675
rect 3495 -725 3540 -700
rect 3495 -750 3505 -725
rect 3530 -750 3540 -725
rect 3495 -770 3540 -750
rect 3555 -585 3600 -575
rect 3555 -610 3565 -585
rect 3590 -610 3600 -585
rect 3555 -630 3600 -610
rect 3555 -655 3565 -630
rect 3590 -655 3600 -630
rect 3555 -675 3600 -655
rect 3555 -700 3565 -675
rect 3590 -700 3600 -675
rect 3555 -725 3600 -700
rect 3555 -750 3565 -725
rect 3590 -750 3600 -725
rect 3555 -770 3600 -750
rect 3615 -585 3660 -575
rect 3615 -610 3625 -585
rect 3650 -610 3660 -585
rect 3615 -630 3660 -610
rect 3615 -655 3625 -630
rect 3650 -655 3660 -630
rect 3615 -675 3660 -655
rect 3615 -700 3625 -675
rect 3650 -700 3660 -675
rect 3615 -725 3660 -700
rect 3615 -750 3625 -725
rect 3650 -750 3660 -725
rect 3615 -770 3660 -750
rect 3675 -585 3720 -575
rect 3675 -610 3685 -585
rect 3710 -610 3720 -585
rect 3675 -630 3720 -610
rect 3675 -655 3685 -630
rect 3710 -655 3720 -630
rect 3675 -675 3720 -655
rect 3675 -700 3685 -675
rect 3710 -700 3720 -675
rect 3675 -725 3720 -700
rect 3675 -750 3685 -725
rect 3710 -750 3720 -725
rect 3675 -770 3720 -750
rect 3735 -585 3780 -575
rect 3735 -610 3745 -585
rect 3770 -610 3780 -585
rect 3735 -630 3780 -610
rect 3735 -655 3745 -630
rect 3770 -655 3780 -630
rect 3735 -675 3780 -655
rect 3735 -700 3745 -675
rect 3770 -700 3780 -675
rect 3735 -725 3780 -700
rect 3735 -750 3745 -725
rect 3770 -750 3780 -725
rect 3735 -770 3780 -750
rect 3795 -585 3840 -575
rect 3795 -610 3805 -585
rect 3830 -610 3840 -585
rect 3795 -630 3840 -610
rect 3795 -655 3805 -630
rect 3830 -655 3840 -630
rect 3795 -675 3840 -655
rect 3795 -700 3805 -675
rect 3830 -700 3840 -675
rect 3795 -725 3840 -700
rect 3795 -750 3805 -725
rect 3830 -750 3840 -725
rect 3795 -770 3840 -750
rect 3855 -585 3900 -575
rect 3855 -610 3865 -585
rect 3890 -610 3900 -585
rect 3855 -630 3900 -610
rect 3855 -655 3865 -630
rect 3890 -655 3900 -630
rect 3855 -675 3900 -655
rect 3855 -700 3865 -675
rect 3890 -700 3900 -675
rect 3855 -725 3900 -700
rect 3855 -750 3865 -725
rect 3890 -750 3900 -725
rect 3855 -770 3900 -750
rect 3915 -585 3960 -575
rect 3915 -610 3925 -585
rect 3950 -610 3960 -585
rect 3915 -630 3960 -610
rect 3915 -655 3925 -630
rect 3950 -655 3960 -630
rect 3915 -675 3960 -655
rect 3915 -700 3925 -675
rect 3950 -700 3960 -675
rect 3915 -725 3960 -700
rect 3915 -750 3925 -725
rect 3950 -750 3960 -725
rect 3915 -770 3960 -750
rect 3975 -585 4020 -575
rect 3975 -610 3985 -585
rect 4010 -610 4020 -585
rect 3975 -630 4020 -610
rect 3975 -655 3985 -630
rect 4010 -655 4020 -630
rect 3975 -675 4020 -655
rect 3975 -700 3985 -675
rect 4010 -700 4020 -675
rect 3975 -725 4020 -700
rect 3975 -750 3985 -725
rect 4010 -750 4020 -725
rect 3975 -770 4020 -750
rect 4035 -585 4080 -575
rect 4035 -610 4045 -585
rect 4070 -610 4080 -585
rect 4035 -630 4080 -610
rect 4035 -655 4045 -630
rect 4070 -655 4080 -630
rect 4035 -675 4080 -655
rect 4035 -700 4045 -675
rect 4070 -700 4080 -675
rect 4035 -725 4080 -700
rect 4035 -750 4045 -725
rect 4070 -750 4080 -725
rect 4035 -770 4080 -750
rect 4095 -585 4140 -575
rect 4095 -610 4105 -585
rect 4130 -610 4140 -585
rect 4095 -630 4140 -610
rect 4095 -655 4105 -630
rect 4130 -655 4140 -630
rect 4095 -675 4140 -655
rect 4095 -700 4105 -675
rect 4130 -700 4140 -675
rect 4095 -725 4140 -700
rect 4095 -750 4105 -725
rect 4130 -750 4140 -725
rect 4095 -770 4140 -750
rect 4155 -585 4200 -575
rect 4155 -610 4165 -585
rect 4190 -610 4200 -585
rect 4155 -630 4200 -610
rect 4155 -655 4165 -630
rect 4190 -655 4200 -630
rect 4155 -675 4200 -655
rect 4155 -700 4165 -675
rect 4190 -700 4200 -675
rect 4155 -725 4200 -700
rect 4155 -750 4165 -725
rect 4190 -750 4200 -725
rect 4155 -770 4200 -750
rect 4215 -585 4260 -575
rect 4215 -610 4225 -585
rect 4250 -610 4260 -585
rect 4215 -630 4260 -610
rect 4215 -655 4225 -630
rect 4250 -655 4260 -630
rect 4215 -675 4260 -655
rect 4215 -700 4225 -675
rect 4250 -700 4260 -675
rect 4215 -725 4260 -700
rect 4215 -750 4225 -725
rect 4250 -750 4260 -725
rect 4215 -770 4260 -750
rect 4275 -585 4320 -575
rect 4275 -610 4285 -585
rect 4310 -610 4320 -585
rect 4275 -630 4320 -610
rect 4275 -655 4285 -630
rect 4310 -655 4320 -630
rect 4275 -675 4320 -655
rect 4275 -700 4285 -675
rect 4310 -700 4320 -675
rect 4275 -725 4320 -700
rect 4275 -750 4285 -725
rect 4310 -750 4320 -725
rect 4275 -770 4320 -750
rect 4335 -585 4380 -575
rect 4335 -610 4345 -585
rect 4370 -610 4380 -585
rect 4335 -630 4380 -610
rect 4335 -655 4345 -630
rect 4370 -655 4380 -630
rect 4335 -675 4380 -655
rect 4335 -700 4345 -675
rect 4370 -700 4380 -675
rect 4335 -725 4380 -700
rect 4335 -750 4345 -725
rect 4370 -750 4380 -725
rect 4335 -770 4380 -750
rect 4395 -585 4440 -575
rect 4395 -610 4405 -585
rect 4430 -610 4440 -585
rect 4395 -630 4440 -610
rect 4395 -655 4405 -630
rect 4430 -655 4440 -630
rect 4395 -675 4440 -655
rect 4395 -700 4405 -675
rect 4430 -700 4440 -675
rect 4395 -725 4440 -700
rect 4395 -750 4405 -725
rect 4430 -750 4440 -725
rect 4395 -770 4440 -750
rect 4455 -585 4500 -575
rect 4455 -610 4465 -585
rect 4490 -610 4500 -585
rect 4455 -630 4500 -610
rect 4455 -655 4465 -630
rect 4490 -655 4500 -630
rect 4455 -675 4500 -655
rect 4455 -700 4465 -675
rect 4490 -700 4500 -675
rect 4455 -725 4500 -700
rect 4455 -750 4465 -725
rect 4490 -750 4500 -725
rect 4455 -770 4500 -750
rect 4515 -585 4560 -575
rect 4515 -610 4525 -585
rect 4550 -610 4560 -585
rect 4515 -630 4560 -610
rect 4515 -655 4525 -630
rect 4550 -655 4560 -630
rect 4515 -675 4560 -655
rect 4515 -700 4525 -675
rect 4550 -700 4560 -675
rect 4515 -725 4560 -700
rect 4515 -750 4525 -725
rect 4550 -750 4560 -725
rect 4515 -770 4560 -750
rect 4575 -585 4620 -575
rect 4575 -610 4585 -585
rect 4610 -610 4620 -585
rect 4575 -630 4620 -610
rect 4575 -655 4585 -630
rect 4610 -655 4620 -630
rect 4575 -675 4620 -655
rect 4575 -700 4585 -675
rect 4610 -700 4620 -675
rect 4575 -725 4620 -700
rect 4575 -750 4585 -725
rect 4610 -750 4620 -725
rect 4575 -770 4620 -750
rect 4635 -585 4680 -575
rect 4635 -610 4645 -585
rect 4670 -610 4680 -585
rect 4635 -630 4680 -610
rect 4635 -655 4645 -630
rect 4670 -655 4680 -630
rect 4635 -675 4680 -655
rect 4635 -700 4645 -675
rect 4670 -700 4680 -675
rect 4635 -725 4680 -700
rect 4635 -750 4645 -725
rect 4670 -750 4680 -725
rect 4635 -770 4680 -750
rect 4695 -585 4740 -575
rect 4695 -610 4705 -585
rect 4730 -610 4740 -585
rect 4695 -630 4740 -610
rect 4695 -655 4705 -630
rect 4730 -655 4740 -630
rect 4695 -675 4740 -655
rect 4695 -700 4705 -675
rect 4730 -700 4740 -675
rect 4695 -725 4740 -700
rect 4695 -750 4705 -725
rect 4730 -750 4740 -725
rect 4695 -770 4740 -750
rect 4755 -585 4800 -575
rect 4755 -610 4765 -585
rect 4790 -610 4800 -585
rect 4755 -630 4800 -610
rect 4755 -655 4765 -630
rect 4790 -655 4800 -630
rect 4755 -675 4800 -655
rect 4755 -700 4765 -675
rect 4790 -700 4800 -675
rect 4755 -725 4800 -700
rect 4755 -750 4765 -725
rect 4790 -750 4800 -725
rect 4755 -770 4800 -750
rect 4815 -585 4860 -575
rect 4815 -610 4825 -585
rect 4850 -610 4860 -585
rect 4815 -630 4860 -610
rect 4815 -655 4825 -630
rect 4850 -655 4860 -630
rect 4815 -675 4860 -655
rect 4815 -700 4825 -675
rect 4850 -700 4860 -675
rect 4815 -725 4860 -700
rect 4815 -750 4825 -725
rect 4850 -750 4860 -725
rect 4815 -770 4860 -750
rect 4875 -585 4920 -575
rect 4875 -610 4885 -585
rect 4910 -610 4920 -585
rect 4875 -630 4920 -610
rect 4875 -655 4885 -630
rect 4910 -655 4920 -630
rect 4875 -675 4920 -655
rect 4875 -700 4885 -675
rect 4910 -700 4920 -675
rect 4875 -725 4920 -700
rect 4875 -750 4885 -725
rect 4910 -750 4920 -725
rect 4875 -770 4920 -750
rect 4935 -585 4980 -575
rect 4935 -610 4945 -585
rect 4970 -610 4980 -585
rect 4935 -630 4980 -610
rect 4935 -655 4945 -630
rect 4970 -655 4980 -630
rect 4935 -675 4980 -655
rect 4935 -700 4945 -675
rect 4970 -700 4980 -675
rect 4935 -725 4980 -700
rect 4935 -750 4945 -725
rect 4970 -750 4980 -725
rect 4935 -770 4980 -750
rect 4995 -585 5040 -575
rect 4995 -610 5005 -585
rect 5030 -610 5040 -585
rect 4995 -630 5040 -610
rect 4995 -655 5005 -630
rect 5030 -655 5040 -630
rect 4995 -675 5040 -655
rect 4995 -700 5005 -675
rect 5030 -700 5040 -675
rect 4995 -725 5040 -700
rect 4995 -750 5005 -725
rect 5030 -750 5040 -725
rect 4995 -770 5040 -750
rect 5055 -585 5100 -575
rect 5055 -610 5065 -585
rect 5090 -610 5100 -585
rect 5055 -630 5100 -610
rect 5055 -655 5065 -630
rect 5090 -655 5100 -630
rect 5055 -675 5100 -655
rect 5055 -700 5065 -675
rect 5090 -700 5100 -675
rect 5055 -725 5100 -700
rect 5055 -750 5065 -725
rect 5090 -750 5100 -725
rect 5055 -770 5100 -750
rect 5115 -585 5160 -575
rect 5115 -610 5125 -585
rect 5150 -610 5160 -585
rect 5115 -630 5160 -610
rect 5115 -655 5125 -630
rect 5150 -655 5160 -630
rect 5115 -675 5160 -655
rect 5115 -700 5125 -675
rect 5150 -700 5160 -675
rect 5115 -725 5160 -700
rect 5115 -750 5125 -725
rect 5150 -750 5160 -725
rect 5115 -770 5160 -750
rect 5175 -585 5220 -575
rect 5175 -610 5185 -585
rect 5210 -610 5220 -585
rect 5175 -630 5220 -610
rect 5175 -655 5185 -630
rect 5210 -655 5220 -630
rect 5175 -675 5220 -655
rect 5175 -700 5185 -675
rect 5210 -700 5220 -675
rect 5175 -725 5220 -700
rect 5175 -750 5185 -725
rect 5210 -750 5220 -725
rect 5175 -770 5220 -750
rect 5235 -585 5280 -575
rect 5235 -610 5245 -585
rect 5270 -610 5280 -585
rect 5235 -630 5280 -610
rect 5235 -655 5245 -630
rect 5270 -655 5280 -630
rect 5235 -675 5280 -655
rect 5235 -700 5245 -675
rect 5270 -700 5280 -675
rect 5235 -725 5280 -700
rect 5235 -750 5245 -725
rect 5270 -750 5280 -725
rect 5235 -770 5280 -750
rect 5295 -585 5340 -575
rect 5295 -610 5305 -585
rect 5330 -610 5340 -585
rect 5295 -630 5340 -610
rect 5295 -655 5305 -630
rect 5330 -655 5340 -630
rect 5295 -675 5340 -655
rect 5295 -700 5305 -675
rect 5330 -700 5340 -675
rect 5295 -725 5340 -700
rect 5295 -750 5305 -725
rect 5330 -750 5340 -725
rect 5295 -770 5340 -750
rect 5355 -585 5400 -575
rect 5355 -610 5365 -585
rect 5390 -610 5400 -585
rect 5355 -630 5400 -610
rect 5355 -655 5365 -630
rect 5390 -655 5400 -630
rect 5355 -675 5400 -655
rect 5355 -700 5365 -675
rect 5390 -700 5400 -675
rect 5355 -725 5400 -700
rect 5355 -750 5365 -725
rect 5390 -750 5400 -725
rect 5355 -770 5400 -750
rect 5415 -585 5460 -575
rect 5415 -610 5425 -585
rect 5450 -610 5460 -585
rect 5415 -630 5460 -610
rect 5415 -655 5425 -630
rect 5450 -655 5460 -630
rect 5415 -675 5460 -655
rect 5415 -700 5425 -675
rect 5450 -700 5460 -675
rect 5415 -725 5460 -700
rect 5415 -750 5425 -725
rect 5450 -750 5460 -725
rect 5415 -770 5460 -750
rect 5475 -585 5520 -575
rect 5475 -610 5485 -585
rect 5510 -610 5520 -585
rect 5475 -630 5520 -610
rect 5475 -655 5485 -630
rect 5510 -655 5520 -630
rect 5475 -675 5520 -655
rect 5475 -700 5485 -675
rect 5510 -700 5520 -675
rect 5475 -725 5520 -700
rect 5475 -750 5485 -725
rect 5510 -750 5520 -725
rect 5475 -770 5520 -750
rect 5535 -585 5580 -575
rect 5535 -610 5545 -585
rect 5570 -610 5580 -585
rect 5535 -630 5580 -610
rect 5535 -655 5545 -630
rect 5570 -655 5580 -630
rect 5535 -675 5580 -655
rect 5535 -700 5545 -675
rect 5570 -700 5580 -675
rect 5535 -725 5580 -700
rect 5535 -750 5545 -725
rect 5570 -750 5580 -725
rect 5535 -770 5580 -750
rect 5595 -585 5640 -575
rect 5595 -610 5605 -585
rect 5630 -610 5640 -585
rect 5595 -630 5640 -610
rect 5595 -655 5605 -630
rect 5630 -655 5640 -630
rect 5595 -675 5640 -655
rect 5595 -700 5605 -675
rect 5630 -700 5640 -675
rect 5595 -725 5640 -700
rect 5595 -750 5605 -725
rect 5630 -750 5640 -725
rect 5595 -770 5640 -750
rect 5655 -585 5700 -575
rect 5655 -610 5665 -585
rect 5690 -610 5700 -585
rect 5655 -630 5700 -610
rect 5655 -655 5665 -630
rect 5690 -655 5700 -630
rect 5655 -675 5700 -655
rect 5655 -700 5665 -675
rect 5690 -700 5700 -675
rect 5655 -725 5700 -700
rect 5655 -750 5665 -725
rect 5690 -750 5700 -725
rect 5655 -770 5700 -750
rect 5715 -585 5760 -575
rect 5715 -610 5725 -585
rect 5750 -610 5760 -585
rect 5715 -630 5760 -610
rect 5715 -655 5725 -630
rect 5750 -655 5760 -630
rect 5715 -675 5760 -655
rect 5715 -700 5725 -675
rect 5750 -700 5760 -675
rect 5715 -725 5760 -700
rect 5715 -750 5725 -725
rect 5750 -750 5760 -725
rect 5715 -770 5760 -750
rect 5775 -585 5820 -575
rect 5775 -610 5785 -585
rect 5810 -610 5820 -585
rect 5775 -630 5820 -610
rect 5775 -655 5785 -630
rect 5810 -655 5820 -630
rect 5775 -675 5820 -655
rect 5775 -700 5785 -675
rect 5810 -700 5820 -675
rect 5775 -725 5820 -700
rect 5775 -750 5785 -725
rect 5810 -750 5820 -725
rect 5775 -770 5820 -750
rect 5835 -585 5880 -575
rect 5835 -610 5845 -585
rect 5870 -610 5880 -585
rect 5835 -630 5880 -610
rect 5835 -655 5845 -630
rect 5870 -655 5880 -630
rect 5835 -675 5880 -655
rect 5835 -700 5845 -675
rect 5870 -700 5880 -675
rect 5835 -725 5880 -700
rect 5835 -750 5845 -725
rect 5870 -750 5880 -725
rect 5835 -770 5880 -750
rect 5895 -585 5940 -575
rect 5895 -610 5905 -585
rect 5930 -610 5940 -585
rect 5895 -630 5940 -610
rect 5895 -655 5905 -630
rect 5930 -655 5940 -630
rect 5895 -675 5940 -655
rect 5895 -700 5905 -675
rect 5930 -700 5940 -675
rect 5895 -725 5940 -700
rect 5895 -750 5905 -725
rect 5930 -750 5940 -725
rect 5895 -770 5940 -750
rect 5955 -585 6000 -575
rect 5955 -610 5965 -585
rect 5990 -610 6000 -585
rect 5955 -630 6000 -610
rect 5955 -655 5965 -630
rect 5990 -655 6000 -630
rect 5955 -675 6000 -655
rect 5955 -700 5965 -675
rect 5990 -700 6000 -675
rect 5955 -725 6000 -700
rect 5955 -750 5965 -725
rect 5990 -750 6000 -725
rect 5955 -770 6000 -750
rect 6015 -585 6060 -575
rect 6015 -610 6025 -585
rect 6050 -610 6060 -585
rect 6015 -630 6060 -610
rect 6015 -655 6025 -630
rect 6050 -655 6060 -630
rect 6015 -675 6060 -655
rect 6015 -700 6025 -675
rect 6050 -700 6060 -675
rect 6015 -725 6060 -700
rect 6015 -750 6025 -725
rect 6050 -750 6060 -725
rect 6015 -770 6060 -750
rect 6075 -585 6120 -575
rect 6075 -610 6085 -585
rect 6110 -610 6120 -585
rect 6075 -630 6120 -610
rect 6075 -655 6085 -630
rect 6110 -655 6120 -630
rect 6075 -675 6120 -655
rect 6075 -700 6085 -675
rect 6110 -700 6120 -675
rect 6075 -725 6120 -700
rect 6075 -750 6085 -725
rect 6110 -750 6120 -725
rect 6075 -770 6120 -750
rect 6135 -585 6180 -575
rect 6135 -610 6145 -585
rect 6170 -610 6180 -585
rect 6135 -630 6180 -610
rect 6135 -655 6145 -630
rect 6170 -655 6180 -630
rect 6135 -675 6180 -655
rect 6135 -700 6145 -675
rect 6170 -700 6180 -675
rect 6135 -725 6180 -700
rect 6135 -750 6145 -725
rect 6170 -750 6180 -725
rect 6135 -770 6180 -750
rect 6195 -585 6240 -575
rect 6195 -610 6205 -585
rect 6230 -610 6240 -585
rect 6195 -630 6240 -610
rect 6195 -655 6205 -630
rect 6230 -655 6240 -630
rect 6195 -675 6240 -655
rect 6195 -700 6205 -675
rect 6230 -700 6240 -675
rect 6195 -725 6240 -700
rect 6195 -750 6205 -725
rect 6230 -750 6240 -725
rect 6195 -770 6240 -750
rect 6255 -585 6300 -575
rect 6255 -610 6265 -585
rect 6290 -610 6300 -585
rect 6255 -630 6300 -610
rect 6255 -655 6265 -630
rect 6290 -655 6300 -630
rect 6255 -675 6300 -655
rect 6255 -700 6265 -675
rect 6290 -700 6300 -675
rect 6255 -725 6300 -700
rect 6255 -750 6265 -725
rect 6290 -750 6300 -725
rect 6255 -770 6300 -750
rect 6315 -585 6360 -575
rect 6315 -610 6325 -585
rect 6350 -610 6360 -585
rect 6315 -630 6360 -610
rect 6315 -655 6325 -630
rect 6350 -655 6360 -630
rect 6315 -675 6360 -655
rect 6315 -700 6325 -675
rect 6350 -700 6360 -675
rect 6315 -725 6360 -700
rect 6315 -750 6325 -725
rect 6350 -750 6360 -725
rect 6315 -770 6360 -750
rect 6375 -585 6420 -575
rect 6375 -610 6385 -585
rect 6410 -610 6420 -585
rect 6375 -630 6420 -610
rect 6375 -655 6385 -630
rect 6410 -655 6420 -630
rect 6375 -675 6420 -655
rect 6375 -700 6385 -675
rect 6410 -700 6420 -675
rect 6375 -725 6420 -700
rect 6375 -750 6385 -725
rect 6410 -750 6420 -725
rect 6375 -770 6420 -750
rect 6435 -585 6480 -575
rect 6435 -610 6445 -585
rect 6470 -610 6480 -585
rect 6435 -630 6480 -610
rect 6435 -655 6445 -630
rect 6470 -655 6480 -630
rect 6435 -675 6480 -655
rect 6435 -700 6445 -675
rect 6470 -700 6480 -675
rect 6435 -725 6480 -700
rect 6435 -750 6445 -725
rect 6470 -750 6480 -725
rect 6435 -770 6480 -750
rect 6495 -585 6540 -575
rect 6495 -610 6505 -585
rect 6530 -610 6540 -585
rect 6495 -630 6540 -610
rect 6495 -655 6505 -630
rect 6530 -655 6540 -630
rect 6495 -675 6540 -655
rect 6495 -700 6505 -675
rect 6530 -700 6540 -675
rect 6495 -725 6540 -700
rect 6495 -750 6505 -725
rect 6530 -750 6540 -725
rect 6495 -770 6540 -750
rect 6555 -585 6600 -575
rect 6555 -610 6565 -585
rect 6590 -610 6600 -585
rect 6555 -630 6600 -610
rect 6555 -655 6565 -630
rect 6590 -655 6600 -630
rect 6555 -675 6600 -655
rect 6555 -700 6565 -675
rect 6590 -700 6600 -675
rect 6555 -725 6600 -700
rect 6555 -750 6565 -725
rect 6590 -750 6600 -725
rect 6555 -770 6600 -750
rect 6615 -585 6660 -575
rect 6615 -610 6625 -585
rect 6650 -610 6660 -585
rect 6615 -630 6660 -610
rect 6615 -655 6625 -630
rect 6650 -655 6660 -630
rect 6615 -675 6660 -655
rect 6615 -700 6625 -675
rect 6650 -700 6660 -675
rect 6615 -725 6660 -700
rect 6615 -750 6625 -725
rect 6650 -750 6660 -725
rect 6615 -770 6660 -750
rect 6675 -585 6720 -575
rect 6675 -610 6685 -585
rect 6710 -610 6720 -585
rect 6675 -630 6720 -610
rect 6675 -655 6685 -630
rect 6710 -655 6720 -630
rect 6675 -675 6720 -655
rect 6675 -700 6685 -675
rect 6710 -700 6720 -675
rect 6675 -725 6720 -700
rect 6675 -750 6685 -725
rect 6710 -750 6720 -725
rect 6675 -770 6720 -750
rect 6735 -585 6780 -575
rect 6735 -610 6745 -585
rect 6770 -610 6780 -585
rect 6735 -630 6780 -610
rect 6735 -655 6745 -630
rect 6770 -655 6780 -630
rect 6735 -675 6780 -655
rect 6735 -700 6745 -675
rect 6770 -700 6780 -675
rect 6735 -725 6780 -700
rect 6735 -750 6745 -725
rect 6770 -750 6780 -725
rect 6735 -770 6780 -750
rect 6795 -585 6840 -575
rect 6795 -610 6805 -585
rect 6830 -610 6840 -585
rect 6795 -630 6840 -610
rect 6795 -655 6805 -630
rect 6830 -655 6840 -630
rect 6795 -675 6840 -655
rect 6795 -700 6805 -675
rect 6830 -700 6840 -675
rect 6795 -725 6840 -700
rect 6795 -750 6805 -725
rect 6830 -750 6840 -725
rect 6795 -770 6840 -750
rect 6855 -585 6900 -575
rect 6855 -610 6865 -585
rect 6890 -610 6900 -585
rect 6855 -630 6900 -610
rect 6855 -655 6865 -630
rect 6890 -655 6900 -630
rect 6855 -675 6900 -655
rect 6855 -700 6865 -675
rect 6890 -700 6900 -675
rect 6855 -725 6900 -700
rect 6855 -750 6865 -725
rect 6890 -750 6900 -725
rect 6855 -770 6900 -750
rect 6915 -585 6960 -575
rect 6915 -610 6925 -585
rect 6950 -610 6960 -585
rect 6915 -630 6960 -610
rect 6915 -655 6925 -630
rect 6950 -655 6960 -630
rect 6915 -675 6960 -655
rect 6915 -700 6925 -675
rect 6950 -700 6960 -675
rect 6915 -725 6960 -700
rect 6915 -750 6925 -725
rect 6950 -750 6960 -725
rect 6915 -770 6960 -750
rect 6975 -585 7020 -575
rect 6975 -610 6985 -585
rect 7010 -610 7020 -585
rect 6975 -630 7020 -610
rect 6975 -655 6985 -630
rect 7010 -655 7020 -630
rect 6975 -675 7020 -655
rect 6975 -700 6985 -675
rect 7010 -700 7020 -675
rect 6975 -725 7020 -700
rect 6975 -750 6985 -725
rect 7010 -750 7020 -725
rect 6975 -770 7020 -750
rect 7035 -585 7080 -575
rect 7035 -610 7045 -585
rect 7070 -610 7080 -585
rect 7035 -630 7080 -610
rect 7035 -655 7045 -630
rect 7070 -655 7080 -630
rect 7035 -675 7080 -655
rect 7035 -700 7045 -675
rect 7070 -700 7080 -675
rect 7035 -725 7080 -700
rect 7035 -750 7045 -725
rect 7070 -750 7080 -725
rect 7035 -770 7080 -750
rect 7095 -585 7140 -575
rect 7095 -610 7105 -585
rect 7130 -610 7140 -585
rect 7095 -630 7140 -610
rect 7095 -655 7105 -630
rect 7130 -655 7140 -630
rect 7095 -675 7140 -655
rect 7095 -700 7105 -675
rect 7130 -700 7140 -675
rect 7095 -725 7140 -700
rect 7095 -750 7105 -725
rect 7130 -750 7140 -725
rect 7095 -770 7140 -750
rect 7155 -585 7200 -575
rect 7155 -610 7165 -585
rect 7190 -610 7200 -585
rect 7155 -630 7200 -610
rect 7155 -655 7165 -630
rect 7190 -655 7200 -630
rect 7155 -675 7200 -655
rect 7155 -700 7165 -675
rect 7190 -700 7200 -675
rect 7155 -725 7200 -700
rect 7155 -750 7165 -725
rect 7190 -750 7200 -725
rect 7155 -770 7200 -750
rect 7215 -585 7260 -575
rect 7215 -610 7225 -585
rect 7250 -610 7260 -585
rect 7215 -630 7260 -610
rect 7215 -655 7225 -630
rect 7250 -655 7260 -630
rect 7215 -675 7260 -655
rect 7215 -700 7225 -675
rect 7250 -700 7260 -675
rect 7215 -725 7260 -700
rect 7215 -750 7225 -725
rect 7250 -750 7260 -725
rect 7215 -770 7260 -750
rect 7275 -585 7320 -575
rect 7275 -610 7285 -585
rect 7310 -610 7320 -585
rect 7275 -630 7320 -610
rect 7275 -655 7285 -630
rect 7310 -655 7320 -630
rect 7275 -675 7320 -655
rect 7275 -700 7285 -675
rect 7310 -700 7320 -675
rect 7275 -725 7320 -700
rect 7275 -750 7285 -725
rect 7310 -750 7320 -725
rect 7275 -770 7320 -750
rect 7335 -585 7380 -575
rect 7335 -610 7345 -585
rect 7370 -610 7380 -585
rect 7335 -630 7380 -610
rect 7335 -655 7345 -630
rect 7370 -655 7380 -630
rect 7335 -675 7380 -655
rect 7335 -700 7345 -675
rect 7370 -700 7380 -675
rect 7335 -725 7380 -700
rect 7335 -750 7345 -725
rect 7370 -750 7380 -725
rect 7335 -770 7380 -750
rect 7395 -585 7440 -575
rect 7395 -610 7405 -585
rect 7430 -610 7440 -585
rect 7395 -630 7440 -610
rect 7395 -655 7405 -630
rect 7430 -655 7440 -630
rect 7395 -675 7440 -655
rect 7395 -700 7405 -675
rect 7430 -700 7440 -675
rect 7395 -725 7440 -700
rect 7395 -750 7405 -725
rect 7430 -750 7440 -725
rect 7395 -770 7440 -750
rect 7455 -585 7500 -575
rect 7455 -610 7465 -585
rect 7490 -610 7500 -585
rect 7455 -630 7500 -610
rect 7455 -655 7465 -630
rect 7490 -655 7500 -630
rect 7455 -675 7500 -655
rect 7455 -700 7465 -675
rect 7490 -700 7500 -675
rect 7455 -725 7500 -700
rect 7455 -750 7465 -725
rect 7490 -750 7500 -725
rect 7455 -770 7500 -750
rect 7515 -585 7560 -575
rect 7515 -610 7525 -585
rect 7550 -610 7560 -585
rect 7515 -630 7560 -610
rect 7515 -655 7525 -630
rect 7550 -655 7560 -630
rect 7515 -675 7560 -655
rect 7515 -700 7525 -675
rect 7550 -700 7560 -675
rect 7515 -725 7560 -700
rect 7515 -750 7525 -725
rect 7550 -750 7560 -725
rect 7515 -770 7560 -750
rect 7575 -585 7620 -575
rect 7575 -610 7585 -585
rect 7610 -610 7620 -585
rect 7575 -630 7620 -610
rect 7575 -655 7585 -630
rect 7610 -655 7620 -630
rect 7575 -675 7620 -655
rect 7575 -700 7585 -675
rect 7610 -700 7620 -675
rect 7575 -725 7620 -700
rect 7575 -750 7585 -725
rect 7610 -750 7620 -725
rect 7575 -770 7620 -750
rect 7635 -585 7680 -575
rect 7635 -610 7645 -585
rect 7670 -610 7680 -585
rect 7635 -630 7680 -610
rect 7635 -655 7645 -630
rect 7670 -655 7680 -630
rect 7635 -675 7680 -655
rect 7635 -700 7645 -675
rect 7670 -700 7680 -675
rect 7635 -725 7680 -700
rect 7635 -750 7645 -725
rect 7670 -750 7680 -725
rect 7635 -770 7680 -750
rect 7695 -585 7740 -575
rect 7695 -610 7705 -585
rect 7730 -610 7740 -585
rect 7695 -630 7740 -610
rect 7695 -655 7705 -630
rect 7730 -655 7740 -630
rect 7695 -675 7740 -655
rect 7695 -700 7705 -675
rect 7730 -700 7740 -675
rect 7695 -725 7740 -700
rect 7695 -750 7705 -725
rect 7730 -750 7740 -725
rect 7695 -770 7740 -750
rect 7755 -585 7800 -575
rect 7755 -610 7765 -585
rect 7790 -610 7800 -585
rect 7755 -630 7800 -610
rect 7755 -655 7765 -630
rect 7790 -655 7800 -630
rect 7755 -675 7800 -655
rect 7755 -700 7765 -675
rect 7790 -700 7800 -675
rect 7755 -725 7800 -700
rect 7755 -750 7765 -725
rect 7790 -750 7800 -725
rect 7755 -770 7800 -750
rect 7815 -585 7860 -575
rect 7815 -610 7825 -585
rect 7850 -610 7860 -585
rect 7815 -630 7860 -610
rect 7815 -655 7825 -630
rect 7850 -655 7860 -630
rect 7815 -675 7860 -655
rect 7815 -700 7825 -675
rect 7850 -700 7860 -675
rect 7815 -725 7860 -700
rect 7815 -750 7825 -725
rect 7850 -750 7860 -725
rect 7815 -770 7860 -750
rect 7875 -585 7920 -575
rect 7875 -610 7885 -585
rect 7910 -610 7920 -585
rect 7875 -630 7920 -610
rect 7875 -655 7885 -630
rect 7910 -655 7920 -630
rect 7875 -675 7920 -655
rect 7875 -700 7885 -675
rect 7910 -700 7920 -675
rect 7875 -725 7920 -700
rect 7875 -750 7885 -725
rect 7910 -750 7920 -725
rect 7875 -770 7920 -750
rect 7935 -585 7980 -575
rect 7935 -610 7945 -585
rect 7970 -610 7980 -585
rect 7935 -630 7980 -610
rect 7935 -655 7945 -630
rect 7970 -655 7980 -630
rect 7935 -675 7980 -655
rect 7935 -700 7945 -675
rect 7970 -700 7980 -675
rect 7935 -725 7980 -700
rect 7935 -750 7945 -725
rect 7970 -750 7980 -725
rect 7935 -770 7980 -750
rect 7995 -585 8040 -575
rect 7995 -610 8005 -585
rect 8030 -610 8040 -585
rect 7995 -630 8040 -610
rect 7995 -655 8005 -630
rect 8030 -655 8040 -630
rect 7995 -675 8040 -655
rect 7995 -700 8005 -675
rect 8030 -700 8040 -675
rect 7995 -725 8040 -700
rect 7995 -750 8005 -725
rect 8030 -750 8040 -725
rect 7995 -770 8040 -750
rect 8055 -585 8100 -575
rect 8055 -610 8065 -585
rect 8090 -610 8100 -585
rect 8055 -630 8100 -610
rect 8055 -655 8065 -630
rect 8090 -655 8100 -630
rect 8055 -675 8100 -655
rect 8055 -700 8065 -675
rect 8090 -700 8100 -675
rect 8055 -725 8100 -700
rect 8055 -750 8065 -725
rect 8090 -750 8100 -725
rect 8055 -770 8100 -750
rect 8115 -585 8160 -575
rect 8115 -610 8125 -585
rect 8150 -610 8160 -585
rect 8115 -630 8160 -610
rect 8115 -655 8125 -630
rect 8150 -655 8160 -630
rect 8115 -675 8160 -655
rect 8115 -700 8125 -675
rect 8150 -700 8160 -675
rect 8115 -725 8160 -700
rect 8115 -750 8125 -725
rect 8150 -750 8160 -725
rect 8115 -770 8160 -750
rect 8175 -585 8220 -575
rect 8175 -610 8185 -585
rect 8210 -610 8220 -585
rect 8175 -630 8220 -610
rect 8175 -655 8185 -630
rect 8210 -655 8220 -630
rect 8175 -675 8220 -655
rect 8175 -700 8185 -675
rect 8210 -700 8220 -675
rect 8175 -725 8220 -700
rect 8175 -750 8185 -725
rect 8210 -750 8220 -725
rect 8175 -770 8220 -750
rect 8235 -585 8280 -575
rect 8235 -610 8245 -585
rect 8270 -610 8280 -585
rect 8235 -630 8280 -610
rect 8235 -655 8245 -630
rect 8270 -655 8280 -630
rect 8235 -675 8280 -655
rect 8235 -700 8245 -675
rect 8270 -700 8280 -675
rect 8235 -725 8280 -700
rect 8235 -750 8245 -725
rect 8270 -750 8280 -725
rect 8235 -770 8280 -750
rect 8295 -585 8340 -575
rect 8295 -610 8305 -585
rect 8330 -610 8340 -585
rect 8295 -630 8340 -610
rect 8295 -655 8305 -630
rect 8330 -655 8340 -630
rect 8295 -675 8340 -655
rect 8295 -700 8305 -675
rect 8330 -700 8340 -675
rect 8295 -725 8340 -700
rect 8295 -750 8305 -725
rect 8330 -750 8340 -725
rect 8295 -770 8340 -750
rect 8355 -585 8400 -575
rect 8355 -610 8365 -585
rect 8390 -610 8400 -585
rect 8355 -630 8400 -610
rect 8355 -655 8365 -630
rect 8390 -655 8400 -630
rect 8355 -675 8400 -655
rect 8355 -700 8365 -675
rect 8390 -700 8400 -675
rect 8355 -725 8400 -700
rect 8355 -750 8365 -725
rect 8390 -750 8400 -725
rect 8355 -770 8400 -750
rect 8415 -585 8460 -575
rect 8415 -610 8425 -585
rect 8450 -610 8460 -585
rect 8415 -630 8460 -610
rect 8415 -655 8425 -630
rect 8450 -655 8460 -630
rect 8415 -675 8460 -655
rect 8415 -700 8425 -675
rect 8450 -700 8460 -675
rect 8415 -725 8460 -700
rect 8415 -750 8425 -725
rect 8450 -750 8460 -725
rect 8415 -770 8460 -750
rect 8475 -585 8520 -575
rect 8475 -610 8485 -585
rect 8510 -610 8520 -585
rect 8475 -630 8520 -610
rect 8475 -655 8485 -630
rect 8510 -655 8520 -630
rect 8475 -675 8520 -655
rect 8475 -700 8485 -675
rect 8510 -700 8520 -675
rect 8475 -725 8520 -700
rect 8475 -750 8485 -725
rect 8510 -750 8520 -725
rect 8475 -770 8520 -750
rect 8535 -585 8580 -575
rect 8535 -610 8545 -585
rect 8570 -610 8580 -585
rect 8535 -630 8580 -610
rect 8535 -655 8545 -630
rect 8570 -655 8580 -630
rect 8535 -675 8580 -655
rect 8535 -700 8545 -675
rect 8570 -700 8580 -675
rect 8535 -725 8580 -700
rect 8535 -750 8545 -725
rect 8570 -750 8580 -725
rect 8535 -770 8580 -750
rect 8595 -585 8640 -575
rect 8595 -610 8605 -585
rect 8630 -610 8640 -585
rect 8595 -630 8640 -610
rect 8595 -655 8605 -630
rect 8630 -655 8640 -630
rect 8595 -675 8640 -655
rect 8595 -700 8605 -675
rect 8630 -700 8640 -675
rect 8595 -725 8640 -700
rect 8595 -750 8605 -725
rect 8630 -750 8640 -725
rect 8595 -770 8640 -750
rect 8655 -585 8700 -575
rect 8655 -610 8665 -585
rect 8690 -610 8700 -585
rect 8655 -630 8700 -610
rect 8655 -655 8665 -630
rect 8690 -655 8700 -630
rect 8655 -675 8700 -655
rect 8655 -700 8665 -675
rect 8690 -700 8700 -675
rect 8655 -725 8700 -700
rect 8655 -750 8665 -725
rect 8690 -750 8700 -725
rect 8655 -770 8700 -750
rect 8715 -585 8760 -575
rect 8715 -610 8725 -585
rect 8750 -610 8760 -585
rect 8715 -630 8760 -610
rect 8715 -655 8725 -630
rect 8750 -655 8760 -630
rect 8715 -675 8760 -655
rect 8715 -700 8725 -675
rect 8750 -700 8760 -675
rect 8715 -725 8760 -700
rect 8715 -750 8725 -725
rect 8750 -750 8760 -725
rect 8715 -770 8760 -750
rect 8775 -585 8820 -575
rect 8775 -610 8785 -585
rect 8810 -610 8820 -585
rect 8775 -630 8820 -610
rect 8775 -655 8785 -630
rect 8810 -655 8820 -630
rect 8775 -675 8820 -655
rect 8775 -700 8785 -675
rect 8810 -700 8820 -675
rect 8775 -725 8820 -700
rect 8775 -750 8785 -725
rect 8810 -750 8820 -725
rect 8775 -770 8820 -750
rect 8835 -585 8880 -575
rect 8835 -610 8845 -585
rect 8870 -610 8880 -585
rect 8835 -630 8880 -610
rect 8835 -655 8845 -630
rect 8870 -655 8880 -630
rect 8835 -675 8880 -655
rect 8835 -700 8845 -675
rect 8870 -700 8880 -675
rect 8835 -725 8880 -700
rect 8835 -750 8845 -725
rect 8870 -750 8880 -725
rect 8835 -770 8880 -750
rect 8895 -585 8940 -575
rect 8895 -610 8905 -585
rect 8930 -610 8940 -585
rect 8895 -630 8940 -610
rect 8895 -655 8905 -630
rect 8930 -655 8940 -630
rect 8895 -675 8940 -655
rect 8895 -700 8905 -675
rect 8930 -700 8940 -675
rect 8895 -725 8940 -700
rect 8895 -750 8905 -725
rect 8930 -750 8940 -725
rect 8895 -770 8940 -750
rect 8955 -585 9000 -575
rect 8955 -610 8965 -585
rect 8990 -610 9000 -585
rect 8955 -630 9000 -610
rect 8955 -655 8965 -630
rect 8990 -655 9000 -630
rect 8955 -675 9000 -655
rect 8955 -700 8965 -675
rect 8990 -700 9000 -675
rect 8955 -725 9000 -700
rect 8955 -750 8965 -725
rect 8990 -750 9000 -725
rect 8955 -770 9000 -750
rect 9015 -585 9060 -575
rect 9015 -610 9025 -585
rect 9050 -610 9060 -585
rect 9015 -630 9060 -610
rect 9015 -655 9025 -630
rect 9050 -655 9060 -630
rect 9015 -675 9060 -655
rect 9015 -700 9025 -675
rect 9050 -700 9060 -675
rect 9015 -725 9060 -700
rect 9015 -750 9025 -725
rect 9050 -750 9060 -725
rect 9015 -770 9060 -750
rect 9075 -585 9120 -575
rect 9075 -610 9085 -585
rect 9110 -610 9120 -585
rect 9075 -630 9120 -610
rect 9075 -655 9085 -630
rect 9110 -655 9120 -630
rect 9075 -675 9120 -655
rect 9075 -700 9085 -675
rect 9110 -700 9120 -675
rect 9075 -725 9120 -700
rect 9075 -750 9085 -725
rect 9110 -750 9120 -725
rect 9075 -770 9120 -750
rect 9135 -585 9180 -575
rect 9135 -610 9145 -585
rect 9170 -610 9180 -585
rect 9135 -630 9180 -610
rect 9135 -655 9145 -630
rect 9170 -655 9180 -630
rect 9135 -675 9180 -655
rect 9135 -700 9145 -675
rect 9170 -700 9180 -675
rect 9135 -725 9180 -700
rect 9135 -750 9145 -725
rect 9170 -750 9180 -725
rect 9135 -770 9180 -750
rect 9195 -585 9240 -575
rect 9195 -610 9205 -585
rect 9230 -610 9240 -585
rect 9195 -630 9240 -610
rect 9195 -655 9205 -630
rect 9230 -655 9240 -630
rect 9195 -675 9240 -655
rect 9195 -700 9205 -675
rect 9230 -700 9240 -675
rect 9195 -725 9240 -700
rect 9195 -750 9205 -725
rect 9230 -750 9240 -725
rect 9195 -770 9240 -750
rect 9255 -585 9300 -575
rect 9255 -610 9265 -585
rect 9290 -610 9300 -585
rect 9255 -630 9300 -610
rect 9255 -655 9265 -630
rect 9290 -655 9300 -630
rect 9255 -675 9300 -655
rect 9255 -700 9265 -675
rect 9290 -700 9300 -675
rect 9255 -725 9300 -700
rect 9255 -750 9265 -725
rect 9290 -750 9300 -725
rect 9255 -770 9300 -750
rect 9315 -585 9360 -575
rect 9315 -610 9325 -585
rect 9350 -610 9360 -585
rect 9315 -630 9360 -610
rect 9315 -655 9325 -630
rect 9350 -655 9360 -630
rect 9315 -675 9360 -655
rect 9315 -700 9325 -675
rect 9350 -700 9360 -675
rect 9315 -725 9360 -700
rect 9315 -750 9325 -725
rect 9350 -750 9360 -725
rect 9315 -770 9360 -750
rect 9375 -585 9420 -575
rect 9375 -610 9385 -585
rect 9410 -610 9420 -585
rect 9375 -630 9420 -610
rect 9375 -655 9385 -630
rect 9410 -655 9420 -630
rect 9375 -675 9420 -655
rect 9375 -700 9385 -675
rect 9410 -700 9420 -675
rect 9375 -725 9420 -700
rect 9375 -750 9385 -725
rect 9410 -750 9420 -725
rect 9375 -770 9420 -750
rect 9435 -585 9480 -575
rect 9435 -610 9445 -585
rect 9470 -610 9480 -585
rect 9435 -630 9480 -610
rect 9435 -655 9445 -630
rect 9470 -655 9480 -630
rect 9435 -675 9480 -655
rect 9435 -700 9445 -675
rect 9470 -700 9480 -675
rect 9435 -725 9480 -700
rect 9435 -750 9445 -725
rect 9470 -750 9480 -725
rect 9435 -770 9480 -750
rect 9495 -585 9540 -575
rect 9495 -610 9505 -585
rect 9530 -610 9540 -585
rect 9495 -630 9540 -610
rect 9495 -655 9505 -630
rect 9530 -655 9540 -630
rect 9495 -675 9540 -655
rect 9495 -700 9505 -675
rect 9530 -700 9540 -675
rect 9495 -725 9540 -700
rect 9495 -750 9505 -725
rect 9530 -750 9540 -725
rect 9495 -770 9540 -750
rect 9555 -585 9600 -575
rect 9555 -610 9565 -585
rect 9590 -610 9600 -585
rect 9555 -630 9600 -610
rect 9555 -655 9565 -630
rect 9590 -655 9600 -630
rect 9555 -675 9600 -655
rect 9555 -700 9565 -675
rect 9590 -700 9600 -675
rect 9555 -725 9600 -700
rect 9555 -750 9565 -725
rect 9590 -750 9600 -725
rect 9555 -770 9600 -750
rect 9615 -585 9660 -575
rect 9615 -610 9625 -585
rect 9650 -610 9660 -585
rect 9615 -630 9660 -610
rect 9615 -655 9625 -630
rect 9650 -655 9660 -630
rect 9615 -675 9660 -655
rect 9615 -700 9625 -675
rect 9650 -700 9660 -675
rect 9615 -725 9660 -700
rect 9615 -750 9625 -725
rect 9650 -750 9660 -725
rect 9615 -770 9660 -750
rect 9675 -585 9720 -575
rect 9675 -610 9685 -585
rect 9710 -610 9720 -585
rect 9675 -630 9720 -610
rect 9675 -655 9685 -630
rect 9710 -655 9720 -630
rect 9675 -675 9720 -655
rect 9675 -700 9685 -675
rect 9710 -700 9720 -675
rect 9675 -725 9720 -700
rect 9675 -750 9685 -725
rect 9710 -750 9720 -725
rect 9675 -770 9720 -750
rect 9735 -585 9780 -575
rect 9735 -610 9745 -585
rect 9770 -610 9780 -585
rect 9735 -630 9780 -610
rect 9735 -655 9745 -630
rect 9770 -655 9780 -630
rect 9735 -675 9780 -655
rect 9735 -700 9745 -675
rect 9770 -700 9780 -675
rect 9735 -725 9780 -700
rect 9735 -750 9745 -725
rect 9770 -750 9780 -725
rect 9735 -770 9780 -750
rect 9795 -585 9840 -575
rect 9795 -610 9805 -585
rect 9830 -610 9840 -585
rect 9795 -630 9840 -610
rect 9795 -655 9805 -630
rect 9830 -655 9840 -630
rect 9795 -675 9840 -655
rect 9795 -700 9805 -675
rect 9830 -700 9840 -675
rect 9795 -725 9840 -700
rect 9795 -750 9805 -725
rect 9830 -750 9840 -725
rect 9795 -770 9840 -750
rect 9855 -585 9900 -575
rect 9855 -610 9865 -585
rect 9890 -610 9900 -585
rect 9855 -630 9900 -610
rect 9855 -655 9865 -630
rect 9890 -655 9900 -630
rect 9855 -675 9900 -655
rect 9855 -700 9865 -675
rect 9890 -700 9900 -675
rect 9855 -725 9900 -700
rect 9855 -750 9865 -725
rect 9890 -750 9900 -725
rect 9855 -770 9900 -750
rect 9915 -585 9960 -575
rect 9915 -610 9925 -585
rect 9950 -610 9960 -585
rect 9915 -630 9960 -610
rect 9915 -655 9925 -630
rect 9950 -655 9960 -630
rect 9915 -675 9960 -655
rect 9915 -700 9925 -675
rect 9950 -700 9960 -675
rect 9915 -725 9960 -700
rect 9915 -750 9925 -725
rect 9950 -750 9960 -725
rect 9915 -770 9960 -750
rect 9975 -585 10020 -575
rect 9975 -610 9985 -585
rect 10010 -610 10020 -585
rect 9975 -630 10020 -610
rect 9975 -655 9985 -630
rect 10010 -655 10020 -630
rect 9975 -675 10020 -655
rect 9975 -700 9985 -675
rect 10010 -700 10020 -675
rect 9975 -725 10020 -700
rect 9975 -750 9985 -725
rect 10010 -750 10020 -725
rect 9975 -770 10020 -750
rect 10035 -585 10080 -575
rect 10035 -610 10045 -585
rect 10070 -610 10080 -585
rect 10035 -630 10080 -610
rect 10035 -655 10045 -630
rect 10070 -655 10080 -630
rect 10035 -675 10080 -655
rect 10035 -700 10045 -675
rect 10070 -700 10080 -675
rect 10035 -725 10080 -700
rect 10035 -750 10045 -725
rect 10070 -750 10080 -725
rect 10035 -770 10080 -750
rect 10095 -585 10140 -575
rect 10095 -610 10105 -585
rect 10130 -610 10140 -585
rect 10095 -630 10140 -610
rect 10095 -655 10105 -630
rect 10130 -655 10140 -630
rect 10095 -675 10140 -655
rect 10095 -700 10105 -675
rect 10130 -700 10140 -675
rect 10095 -725 10140 -700
rect 10095 -750 10105 -725
rect 10130 -750 10140 -725
rect 10095 -770 10140 -750
rect 10155 -585 10200 -575
rect 10155 -610 10165 -585
rect 10190 -610 10200 -585
rect 10155 -630 10200 -610
rect 10155 -655 10165 -630
rect 10190 -655 10200 -630
rect 10155 -675 10200 -655
rect 10155 -700 10165 -675
rect 10190 -700 10200 -675
rect 10155 -725 10200 -700
rect 10155 -750 10165 -725
rect 10190 -750 10200 -725
rect 10155 -770 10200 -750
rect 10215 -585 10260 -575
rect 10215 -610 10225 -585
rect 10250 -610 10260 -585
rect 10215 -630 10260 -610
rect 10215 -655 10225 -630
rect 10250 -655 10260 -630
rect 10215 -675 10260 -655
rect 10215 -700 10225 -675
rect 10250 -700 10260 -675
rect 10215 -725 10260 -700
rect 10215 -750 10225 -725
rect 10250 -750 10260 -725
rect 10215 -770 10260 -750
rect 10275 -585 10320 -575
rect 10275 -610 10285 -585
rect 10310 -610 10320 -585
rect 10275 -630 10320 -610
rect 10275 -655 10285 -630
rect 10310 -655 10320 -630
rect 10275 -675 10320 -655
rect 10275 -700 10285 -675
rect 10310 -700 10320 -675
rect 10275 -725 10320 -700
rect 10275 -750 10285 -725
rect 10310 -750 10320 -725
rect 10275 -770 10320 -750
rect 10335 -585 10380 -575
rect 10335 -610 10345 -585
rect 10370 -610 10380 -585
rect 10335 -630 10380 -610
rect 10335 -655 10345 -630
rect 10370 -655 10380 -630
rect 10335 -675 10380 -655
rect 10335 -700 10345 -675
rect 10370 -700 10380 -675
rect 10335 -725 10380 -700
rect 10335 -750 10345 -725
rect 10370 -750 10380 -725
rect 10335 -770 10380 -750
rect 10395 -585 10440 -575
rect 10395 -610 10405 -585
rect 10430 -610 10440 -585
rect 10395 -630 10440 -610
rect 10395 -655 10405 -630
rect 10430 -655 10440 -630
rect 10395 -675 10440 -655
rect 10395 -700 10405 -675
rect 10430 -700 10440 -675
rect 10395 -725 10440 -700
rect 10395 -750 10405 -725
rect 10430 -750 10440 -725
rect 10395 -770 10440 -750
rect 10455 -585 10500 -575
rect 10455 -610 10465 -585
rect 10490 -610 10500 -585
rect 10455 -630 10500 -610
rect 10455 -655 10465 -630
rect 10490 -655 10500 -630
rect 10455 -675 10500 -655
rect 10455 -700 10465 -675
rect 10490 -700 10500 -675
rect 10455 -725 10500 -700
rect 10455 -750 10465 -725
rect 10490 -750 10500 -725
rect 10455 -770 10500 -750
rect 10515 -585 10560 -575
rect 10515 -610 10525 -585
rect 10550 -610 10560 -585
rect 10515 -630 10560 -610
rect 10515 -655 10525 -630
rect 10550 -655 10560 -630
rect 10515 -675 10560 -655
rect 10515 -700 10525 -675
rect 10550 -700 10560 -675
rect 10515 -725 10560 -700
rect 10515 -750 10525 -725
rect 10550 -750 10560 -725
rect 10515 -770 10560 -750
rect 10575 -585 10620 -575
rect 10575 -610 10585 -585
rect 10610 -610 10620 -585
rect 10575 -630 10620 -610
rect 10575 -655 10585 -630
rect 10610 -655 10620 -630
rect 10575 -675 10620 -655
rect 10575 -700 10585 -675
rect 10610 -700 10620 -675
rect 10575 -725 10620 -700
rect 10575 -750 10585 -725
rect 10610 -750 10620 -725
rect 10575 -770 10620 -750
rect 10635 -585 10680 -575
rect 10635 -610 10645 -585
rect 10670 -610 10680 -585
rect 10635 -630 10680 -610
rect 10635 -655 10645 -630
rect 10670 -655 10680 -630
rect 10635 -675 10680 -655
rect 10635 -700 10645 -675
rect 10670 -700 10680 -675
rect 10635 -725 10680 -700
rect 10635 -750 10645 -725
rect 10670 -750 10680 -725
rect 10635 -770 10680 -750
rect 10695 -585 10740 -575
rect 10695 -610 10705 -585
rect 10730 -610 10740 -585
rect 10695 -630 10740 -610
rect 10695 -655 10705 -630
rect 10730 -655 10740 -630
rect 10695 -675 10740 -655
rect 10695 -700 10705 -675
rect 10730 -700 10740 -675
rect 10695 -725 10740 -700
rect 10695 -750 10705 -725
rect 10730 -750 10740 -725
rect 10695 -770 10740 -750
rect 10755 -585 10800 -575
rect 10755 -610 10765 -585
rect 10790 -610 10800 -585
rect 10755 -630 10800 -610
rect 10755 -655 10765 -630
rect 10790 -655 10800 -630
rect 10755 -675 10800 -655
rect 10755 -700 10765 -675
rect 10790 -700 10800 -675
rect 10755 -725 10800 -700
rect 10755 -750 10765 -725
rect 10790 -750 10800 -725
rect 10755 -770 10800 -750
rect 10815 -585 10860 -575
rect 10815 -610 10825 -585
rect 10850 -610 10860 -585
rect 10815 -630 10860 -610
rect 10815 -655 10825 -630
rect 10850 -655 10860 -630
rect 10815 -675 10860 -655
rect 10815 -700 10825 -675
rect 10850 -700 10860 -675
rect 10815 -725 10860 -700
rect 10815 -750 10825 -725
rect 10850 -750 10860 -725
rect 10815 -770 10860 -750
rect 10875 -585 10920 -575
rect 10875 -610 10885 -585
rect 10910 -610 10920 -585
rect 10875 -630 10920 -610
rect 10875 -655 10885 -630
rect 10910 -655 10920 -630
rect 10875 -675 10920 -655
rect 10875 -700 10885 -675
rect 10910 -700 10920 -675
rect 10875 -725 10920 -700
rect 10875 -750 10885 -725
rect 10910 -750 10920 -725
rect 10875 -770 10920 -750
rect 10935 -585 10980 -575
rect 10935 -610 10945 -585
rect 10970 -610 10980 -585
rect 10935 -630 10980 -610
rect 10935 -655 10945 -630
rect 10970 -655 10980 -630
rect 10935 -675 10980 -655
rect 10935 -700 10945 -675
rect 10970 -700 10980 -675
rect 10935 -725 10980 -700
rect 10935 -750 10945 -725
rect 10970 -750 10980 -725
rect 10935 -770 10980 -750
rect 10995 -585 11040 -575
rect 10995 -610 11005 -585
rect 11030 -610 11040 -585
rect 10995 -630 11040 -610
rect 10995 -655 11005 -630
rect 11030 -655 11040 -630
rect 10995 -675 11040 -655
rect 10995 -700 11005 -675
rect 11030 -700 11040 -675
rect 10995 -725 11040 -700
rect 10995 -750 11005 -725
rect 11030 -750 11040 -725
rect 10995 -770 11040 -750
rect 11055 -585 11100 -575
rect 11055 -610 11065 -585
rect 11090 -610 11100 -585
rect 11055 -630 11100 -610
rect 11055 -655 11065 -630
rect 11090 -655 11100 -630
rect 11055 -675 11100 -655
rect 11055 -700 11065 -675
rect 11090 -700 11100 -675
rect 11055 -725 11100 -700
rect 11055 -750 11065 -725
rect 11090 -750 11100 -725
rect 11055 -770 11100 -750
rect 11115 -585 11160 -575
rect 11115 -610 11125 -585
rect 11150 -610 11160 -585
rect 11115 -630 11160 -610
rect 11115 -655 11125 -630
rect 11150 -655 11160 -630
rect 11115 -675 11160 -655
rect 11115 -700 11125 -675
rect 11150 -700 11160 -675
rect 11115 -725 11160 -700
rect 11115 -750 11125 -725
rect 11150 -750 11160 -725
rect 11115 -770 11160 -750
rect 11175 -585 11220 -575
rect 11175 -610 11185 -585
rect 11210 -610 11220 -585
rect 11175 -630 11220 -610
rect 11175 -655 11185 -630
rect 11210 -655 11220 -630
rect 11175 -675 11220 -655
rect 11175 -700 11185 -675
rect 11210 -700 11220 -675
rect 11175 -725 11220 -700
rect 11175 -750 11185 -725
rect 11210 -750 11220 -725
rect 11175 -770 11220 -750
rect 11235 -585 11280 -575
rect 11235 -610 11245 -585
rect 11270 -610 11280 -585
rect 11235 -630 11280 -610
rect 11235 -655 11245 -630
rect 11270 -655 11280 -630
rect 11235 -675 11280 -655
rect 11235 -700 11245 -675
rect 11270 -700 11280 -675
rect 11235 -725 11280 -700
rect 11235 -750 11245 -725
rect 11270 -750 11280 -725
rect 11235 -770 11280 -750
rect 11295 -585 11340 -575
rect 11295 -610 11305 -585
rect 11330 -610 11340 -585
rect 11295 -630 11340 -610
rect 11295 -655 11305 -630
rect 11330 -655 11340 -630
rect 11295 -675 11340 -655
rect 11295 -700 11305 -675
rect 11330 -700 11340 -675
rect 11295 -725 11340 -700
rect 11295 -750 11305 -725
rect 11330 -750 11340 -725
rect 11295 -770 11340 -750
rect 11355 -585 11400 -575
rect 11355 -610 11365 -585
rect 11390 -610 11400 -585
rect 11355 -630 11400 -610
rect 11355 -655 11365 -630
rect 11390 -655 11400 -630
rect 11355 -675 11400 -655
rect 11355 -700 11365 -675
rect 11390 -700 11400 -675
rect 11355 -725 11400 -700
rect 11355 -750 11365 -725
rect 11390 -750 11400 -725
rect 11355 -770 11400 -750
rect 11415 -585 11460 -575
rect 11415 -610 11425 -585
rect 11450 -610 11460 -585
rect 11415 -630 11460 -610
rect 11415 -655 11425 -630
rect 11450 -655 11460 -630
rect 11415 -675 11460 -655
rect 11415 -700 11425 -675
rect 11450 -700 11460 -675
rect 11415 -725 11460 -700
rect 11415 -750 11425 -725
rect 11450 -750 11460 -725
rect 11415 -770 11460 -750
rect 11475 -585 11520 -575
rect 11475 -610 11485 -585
rect 11510 -610 11520 -585
rect 11475 -630 11520 -610
rect 11475 -655 11485 -630
rect 11510 -655 11520 -630
rect 11475 -675 11520 -655
rect 11475 -700 11485 -675
rect 11510 -700 11520 -675
rect 11475 -725 11520 -700
rect 11475 -750 11485 -725
rect 11510 -750 11520 -725
rect 11475 -770 11520 -750
rect 11535 -585 11580 -575
rect 11535 -610 11545 -585
rect 11570 -610 11580 -585
rect 11535 -630 11580 -610
rect 11535 -655 11545 -630
rect 11570 -655 11580 -630
rect 11535 -675 11580 -655
rect 11535 -700 11545 -675
rect 11570 -700 11580 -675
rect 11535 -725 11580 -700
rect 11535 -750 11545 -725
rect 11570 -750 11580 -725
rect 11535 -770 11580 -750
rect 11595 -585 11640 -575
rect 11595 -610 11605 -585
rect 11630 -610 11640 -585
rect 11595 -630 11640 -610
rect 11595 -655 11605 -630
rect 11630 -655 11640 -630
rect 11595 -675 11640 -655
rect 11595 -700 11605 -675
rect 11630 -700 11640 -675
rect 11595 -725 11640 -700
rect 11595 -750 11605 -725
rect 11630 -750 11640 -725
rect 11595 -770 11640 -750
rect 11655 -585 11700 -575
rect 11655 -610 11665 -585
rect 11690 -610 11700 -585
rect 11655 -630 11700 -610
rect 11655 -655 11665 -630
rect 11690 -655 11700 -630
rect 11655 -675 11700 -655
rect 11655 -700 11665 -675
rect 11690 -700 11700 -675
rect 11655 -725 11700 -700
rect 11655 -750 11665 -725
rect 11690 -750 11700 -725
rect 11655 -770 11700 -750
rect 11715 -585 11760 -575
rect 11715 -610 11725 -585
rect 11750 -610 11760 -585
rect 11715 -630 11760 -610
rect 11715 -655 11725 -630
rect 11750 -655 11760 -630
rect 11715 -675 11760 -655
rect 11715 -700 11725 -675
rect 11750 -700 11760 -675
rect 11715 -725 11760 -700
rect 11715 -750 11725 -725
rect 11750 -750 11760 -725
rect 11715 -770 11760 -750
rect 11775 -585 11820 -575
rect 11775 -610 11785 -585
rect 11810 -610 11820 -585
rect 11775 -630 11820 -610
rect 11775 -655 11785 -630
rect 11810 -655 11820 -630
rect 11775 -675 11820 -655
rect 11775 -700 11785 -675
rect 11810 -700 11820 -675
rect 11775 -725 11820 -700
rect 11775 -750 11785 -725
rect 11810 -750 11820 -725
rect 11775 -770 11820 -750
rect 11835 -585 11880 -575
rect 11835 -610 11845 -585
rect 11870 -610 11880 -585
rect 11835 -630 11880 -610
rect 11835 -655 11845 -630
rect 11870 -655 11880 -630
rect 11835 -675 11880 -655
rect 11835 -700 11845 -675
rect 11870 -700 11880 -675
rect 11835 -725 11880 -700
rect 11835 -750 11845 -725
rect 11870 -750 11880 -725
rect 11835 -770 11880 -750
rect 11895 -585 11940 -575
rect 11895 -610 11905 -585
rect 11930 -610 11940 -585
rect 11895 -630 11940 -610
rect 11895 -655 11905 -630
rect 11930 -655 11940 -630
rect 11895 -675 11940 -655
rect 11895 -700 11905 -675
rect 11930 -700 11940 -675
rect 11895 -725 11940 -700
rect 11895 -750 11905 -725
rect 11930 -750 11940 -725
rect 11895 -770 11940 -750
rect 11955 -585 12000 -575
rect 11955 -610 11965 -585
rect 11990 -610 12000 -585
rect 11955 -630 12000 -610
rect 11955 -655 11965 -630
rect 11990 -655 12000 -630
rect 11955 -675 12000 -655
rect 11955 -700 11965 -675
rect 11990 -700 12000 -675
rect 11955 -725 12000 -700
rect 11955 -750 11965 -725
rect 11990 -750 12000 -725
rect 11955 -770 12000 -750
rect 12015 -585 12060 -575
rect 12015 -610 12025 -585
rect 12050 -610 12060 -585
rect 12015 -630 12060 -610
rect 12015 -655 12025 -630
rect 12050 -655 12060 -630
rect 12015 -675 12060 -655
rect 12015 -700 12025 -675
rect 12050 -700 12060 -675
rect 12015 -725 12060 -700
rect 12015 -750 12025 -725
rect 12050 -750 12060 -725
rect 12015 -770 12060 -750
rect 12075 -585 12120 -575
rect 12075 -610 12085 -585
rect 12110 -610 12120 -585
rect 12075 -630 12120 -610
rect 12075 -655 12085 -630
rect 12110 -655 12120 -630
rect 12075 -675 12120 -655
rect 12075 -700 12085 -675
rect 12110 -700 12120 -675
rect 12075 -725 12120 -700
rect 12075 -750 12085 -725
rect 12110 -750 12120 -725
rect 12075 -770 12120 -750
rect 12135 -585 12180 -575
rect 12135 -610 12145 -585
rect 12170 -610 12180 -585
rect 12135 -630 12180 -610
rect 12135 -655 12145 -630
rect 12170 -655 12180 -630
rect 12135 -675 12180 -655
rect 12135 -700 12145 -675
rect 12170 -700 12180 -675
rect 12135 -725 12180 -700
rect 12135 -750 12145 -725
rect 12170 -750 12180 -725
rect 12135 -770 12180 -750
rect 12195 -585 12240 -575
rect 12195 -610 12205 -585
rect 12230 -610 12240 -585
rect 12195 -630 12240 -610
rect 12195 -655 12205 -630
rect 12230 -655 12240 -630
rect 12195 -675 12240 -655
rect 12195 -700 12205 -675
rect 12230 -700 12240 -675
rect 12195 -725 12240 -700
rect 12195 -750 12205 -725
rect 12230 -750 12240 -725
rect 12195 -770 12240 -750
rect 12255 -585 12300 -575
rect 12255 -610 12265 -585
rect 12290 -610 12300 -585
rect 12255 -630 12300 -610
rect 12255 -655 12265 -630
rect 12290 -655 12300 -630
rect 12255 -675 12300 -655
rect 12255 -700 12265 -675
rect 12290 -700 12300 -675
rect 12255 -725 12300 -700
rect 12255 -750 12265 -725
rect 12290 -750 12300 -725
rect 12255 -770 12300 -750
rect 12315 -585 12360 -575
rect 12315 -610 12325 -585
rect 12350 -610 12360 -585
rect 12315 -630 12360 -610
rect 12315 -655 12325 -630
rect 12350 -655 12360 -630
rect 12315 -675 12360 -655
rect 12315 -700 12325 -675
rect 12350 -700 12360 -675
rect 12315 -725 12360 -700
rect 12315 -750 12325 -725
rect 12350 -750 12360 -725
rect 12315 -770 12360 -750
rect 12375 -585 12420 -575
rect 12375 -610 12385 -585
rect 12410 -610 12420 -585
rect 12375 -630 12420 -610
rect 12375 -655 12385 -630
rect 12410 -655 12420 -630
rect 12375 -675 12420 -655
rect 12375 -700 12385 -675
rect 12410 -700 12420 -675
rect 12375 -725 12420 -700
rect 12375 -750 12385 -725
rect 12410 -750 12420 -725
rect 12375 -770 12420 -750
rect 12435 -585 12480 -575
rect 12435 -610 12445 -585
rect 12470 -610 12480 -585
rect 12435 -630 12480 -610
rect 12435 -655 12445 -630
rect 12470 -655 12480 -630
rect 12435 -675 12480 -655
rect 12435 -700 12445 -675
rect 12470 -700 12480 -675
rect 12435 -725 12480 -700
rect 12435 -750 12445 -725
rect 12470 -750 12480 -725
rect 12435 -770 12480 -750
rect 12495 -585 12540 -575
rect 12495 -610 12505 -585
rect 12530 -610 12540 -585
rect 12495 -630 12540 -610
rect 12495 -655 12505 -630
rect 12530 -655 12540 -630
rect 12495 -675 12540 -655
rect 12495 -700 12505 -675
rect 12530 -700 12540 -675
rect 12495 -725 12540 -700
rect 12495 -750 12505 -725
rect 12530 -750 12540 -725
rect 12495 -770 12540 -750
rect 12555 -585 12600 -575
rect 12555 -610 12565 -585
rect 12590 -610 12600 -585
rect 12555 -630 12600 -610
rect 12555 -655 12565 -630
rect 12590 -655 12600 -630
rect 12555 -675 12600 -655
rect 12555 -700 12565 -675
rect 12590 -700 12600 -675
rect 12555 -725 12600 -700
rect 12555 -750 12565 -725
rect 12590 -750 12600 -725
rect 12555 -770 12600 -750
rect 12615 -585 12660 -575
rect 12615 -610 12625 -585
rect 12650 -610 12660 -585
rect 12615 -630 12660 -610
rect 12615 -655 12625 -630
rect 12650 -655 12660 -630
rect 12615 -675 12660 -655
rect 12615 -700 12625 -675
rect 12650 -700 12660 -675
rect 12615 -725 12660 -700
rect 12615 -750 12625 -725
rect 12650 -750 12660 -725
rect 12615 -770 12660 -750
rect 12675 -585 12720 -575
rect 12675 -610 12685 -585
rect 12710 -610 12720 -585
rect 12675 -630 12720 -610
rect 12675 -655 12685 -630
rect 12710 -655 12720 -630
rect 12675 -675 12720 -655
rect 12675 -700 12685 -675
rect 12710 -700 12720 -675
rect 12675 -725 12720 -700
rect 12675 -750 12685 -725
rect 12710 -750 12720 -725
rect 12675 -770 12720 -750
rect 12735 -585 12780 -575
rect 12735 -610 12745 -585
rect 12770 -610 12780 -585
rect 12735 -630 12780 -610
rect 12735 -655 12745 -630
rect 12770 -655 12780 -630
rect 12735 -675 12780 -655
rect 12735 -700 12745 -675
rect 12770 -700 12780 -675
rect 12735 -725 12780 -700
rect 12735 -750 12745 -725
rect 12770 -750 12780 -725
rect 12735 -770 12780 -750
rect 12795 -585 12840 -575
rect 12795 -610 12805 -585
rect 12830 -610 12840 -585
rect 12795 -630 12840 -610
rect 12795 -655 12805 -630
rect 12830 -655 12840 -630
rect 12795 -675 12840 -655
rect 12795 -700 12805 -675
rect 12830 -700 12840 -675
rect 12795 -725 12840 -700
rect 12795 -750 12805 -725
rect 12830 -750 12840 -725
rect 12795 -770 12840 -750
rect 12855 -585 12900 -575
rect 12855 -610 12865 -585
rect 12890 -610 12900 -585
rect 12855 -630 12900 -610
rect 12855 -655 12865 -630
rect 12890 -655 12900 -630
rect 12855 -675 12900 -655
rect 12855 -700 12865 -675
rect 12890 -700 12900 -675
rect 12855 -725 12900 -700
rect 12855 -750 12865 -725
rect 12890 -750 12900 -725
rect 12855 -770 12900 -750
rect 12915 -585 12960 -575
rect 12915 -610 12925 -585
rect 12950 -610 12960 -585
rect 12915 -630 12960 -610
rect 12915 -655 12925 -630
rect 12950 -655 12960 -630
rect 12915 -675 12960 -655
rect 12915 -700 12925 -675
rect 12950 -700 12960 -675
rect 12915 -725 12960 -700
rect 12915 -750 12925 -725
rect 12950 -750 12960 -725
rect 12915 -770 12960 -750
rect 12975 -585 13020 -575
rect 12975 -610 12985 -585
rect 13010 -610 13020 -585
rect 12975 -630 13020 -610
rect 12975 -655 12985 -630
rect 13010 -655 13020 -630
rect 12975 -675 13020 -655
rect 12975 -700 12985 -675
rect 13010 -700 13020 -675
rect 12975 -725 13020 -700
rect 12975 -750 12985 -725
rect 13010 -750 13020 -725
rect 12975 -770 13020 -750
rect 13035 -585 13080 -575
rect 13035 -610 13045 -585
rect 13070 -610 13080 -585
rect 13035 -630 13080 -610
rect 13035 -655 13045 -630
rect 13070 -655 13080 -630
rect 13035 -675 13080 -655
rect 13035 -700 13045 -675
rect 13070 -700 13080 -675
rect 13035 -725 13080 -700
rect 13035 -750 13045 -725
rect 13070 -750 13080 -725
rect 13035 -770 13080 -750
rect 13095 -585 13140 -575
rect 13095 -610 13105 -585
rect 13130 -610 13140 -585
rect 13095 -630 13140 -610
rect 13095 -655 13105 -630
rect 13130 -655 13140 -630
rect 13095 -675 13140 -655
rect 13095 -700 13105 -675
rect 13130 -700 13140 -675
rect 13095 -725 13140 -700
rect 13095 -750 13105 -725
rect 13130 -750 13140 -725
rect 13095 -770 13140 -750
rect 13155 -585 13200 -575
rect 13155 -610 13165 -585
rect 13190 -610 13200 -585
rect 13155 -630 13200 -610
rect 13155 -655 13165 -630
rect 13190 -655 13200 -630
rect 13155 -675 13200 -655
rect 13155 -700 13165 -675
rect 13190 -700 13200 -675
rect 13155 -725 13200 -700
rect 13155 -750 13165 -725
rect 13190 -750 13200 -725
rect 13155 -770 13200 -750
rect 13215 -585 13260 -575
rect 13215 -610 13225 -585
rect 13250 -610 13260 -585
rect 13215 -630 13260 -610
rect 13215 -655 13225 -630
rect 13250 -655 13260 -630
rect 13215 -675 13260 -655
rect 13215 -700 13225 -675
rect 13250 -700 13260 -675
rect 13215 -725 13260 -700
rect 13215 -750 13225 -725
rect 13250 -750 13260 -725
rect 13215 -770 13260 -750
rect 13275 -585 13320 -575
rect 13275 -610 13285 -585
rect 13310 -610 13320 -585
rect 13275 -630 13320 -610
rect 13275 -655 13285 -630
rect 13310 -655 13320 -630
rect 13275 -675 13320 -655
rect 13275 -700 13285 -675
rect 13310 -700 13320 -675
rect 13275 -725 13320 -700
rect 13275 -750 13285 -725
rect 13310 -750 13320 -725
rect 13275 -770 13320 -750
rect 13335 -585 13380 -575
rect 13335 -610 13345 -585
rect 13370 -610 13380 -585
rect 13335 -630 13380 -610
rect 13335 -655 13345 -630
rect 13370 -655 13380 -630
rect 13335 -675 13380 -655
rect 13335 -700 13345 -675
rect 13370 -700 13380 -675
rect 13335 -725 13380 -700
rect 13335 -750 13345 -725
rect 13370 -750 13380 -725
rect 13335 -770 13380 -750
rect 13395 -585 13440 -575
rect 13395 -610 13405 -585
rect 13430 -610 13440 -585
rect 13395 -630 13440 -610
rect 13395 -655 13405 -630
rect 13430 -655 13440 -630
rect 13395 -675 13440 -655
rect 13395 -700 13405 -675
rect 13430 -700 13440 -675
rect 13395 -725 13440 -700
rect 13395 -750 13405 -725
rect 13430 -750 13440 -725
rect 13395 -770 13440 -750
rect 13455 -585 13500 -575
rect 13455 -610 13465 -585
rect 13490 -610 13500 -585
rect 13455 -630 13500 -610
rect 13455 -655 13465 -630
rect 13490 -655 13500 -630
rect 13455 -675 13500 -655
rect 13455 -700 13465 -675
rect 13490 -700 13500 -675
rect 13455 -725 13500 -700
rect 13455 -750 13465 -725
rect 13490 -750 13500 -725
rect 13455 -770 13500 -750
rect 13515 -585 13560 -575
rect 13515 -610 13525 -585
rect 13550 -610 13560 -585
rect 13515 -630 13560 -610
rect 13515 -655 13525 -630
rect 13550 -655 13560 -630
rect 13515 -675 13560 -655
rect 13515 -700 13525 -675
rect 13550 -700 13560 -675
rect 13515 -725 13560 -700
rect 13515 -750 13525 -725
rect 13550 -750 13560 -725
rect 13515 -770 13560 -750
rect 13575 -585 13620 -575
rect 13575 -610 13585 -585
rect 13610 -610 13620 -585
rect 13575 -630 13620 -610
rect 13575 -655 13585 -630
rect 13610 -655 13620 -630
rect 13575 -675 13620 -655
rect 13575 -700 13585 -675
rect 13610 -700 13620 -675
rect 13575 -725 13620 -700
rect 13575 -750 13585 -725
rect 13610 -750 13620 -725
rect 13575 -770 13620 -750
rect 13635 -585 13680 -575
rect 13635 -610 13645 -585
rect 13670 -610 13680 -585
rect 13635 -630 13680 -610
rect 13635 -655 13645 -630
rect 13670 -655 13680 -630
rect 13635 -675 13680 -655
rect 13635 -700 13645 -675
rect 13670 -700 13680 -675
rect 13635 -725 13680 -700
rect 13635 -750 13645 -725
rect 13670 -750 13680 -725
rect 13635 -770 13680 -750
rect 13695 -585 13740 -575
rect 13695 -610 13705 -585
rect 13730 -610 13740 -585
rect 13695 -630 13740 -610
rect 13695 -655 13705 -630
rect 13730 -655 13740 -630
rect 13695 -675 13740 -655
rect 13695 -700 13705 -675
rect 13730 -700 13740 -675
rect 13695 -725 13740 -700
rect 13695 -750 13705 -725
rect 13730 -750 13740 -725
rect 13695 -770 13740 -750
rect 13755 -585 13800 -575
rect 13755 -610 13765 -585
rect 13790 -610 13800 -585
rect 13755 -630 13800 -610
rect 13755 -655 13765 -630
rect 13790 -655 13800 -630
rect 13755 -675 13800 -655
rect 13755 -700 13765 -675
rect 13790 -700 13800 -675
rect 13755 -725 13800 -700
rect 13755 -750 13765 -725
rect 13790 -750 13800 -725
rect 13755 -770 13800 -750
rect 13815 -585 13860 -575
rect 13815 -610 13825 -585
rect 13850 -610 13860 -585
rect 13815 -630 13860 -610
rect 13815 -655 13825 -630
rect 13850 -655 13860 -630
rect 13815 -675 13860 -655
rect 13815 -700 13825 -675
rect 13850 -700 13860 -675
rect 13815 -725 13860 -700
rect 13815 -750 13825 -725
rect 13850 -750 13860 -725
rect 13815 -770 13860 -750
rect 13875 -585 13920 -575
rect 13875 -610 13885 -585
rect 13910 -610 13920 -585
rect 13875 -630 13920 -610
rect 13875 -655 13885 -630
rect 13910 -655 13920 -630
rect 13875 -675 13920 -655
rect 13875 -700 13885 -675
rect 13910 -700 13920 -675
rect 13875 -725 13920 -700
rect 13875 -750 13885 -725
rect 13910 -750 13920 -725
rect 13875 -770 13920 -750
rect 13935 -585 13980 -575
rect 13935 -610 13945 -585
rect 13970 -610 13980 -585
rect 13935 -630 13980 -610
rect 13935 -655 13945 -630
rect 13970 -655 13980 -630
rect 13935 -675 13980 -655
rect 13935 -700 13945 -675
rect 13970 -700 13980 -675
rect 13935 -725 13980 -700
rect 13935 -750 13945 -725
rect 13970 -750 13980 -725
rect 13935 -770 13980 -750
rect 13995 -585 14040 -575
rect 13995 -610 14005 -585
rect 14030 -610 14040 -585
rect 13995 -630 14040 -610
rect 13995 -655 14005 -630
rect 14030 -655 14040 -630
rect 13995 -675 14040 -655
rect 13995 -700 14005 -675
rect 14030 -700 14040 -675
rect 13995 -725 14040 -700
rect 13995 -750 14005 -725
rect 14030 -750 14040 -725
rect 13995 -770 14040 -750
rect 14055 -585 14100 -575
rect 14055 -610 14065 -585
rect 14090 -610 14100 -585
rect 14055 -630 14100 -610
rect 14055 -655 14065 -630
rect 14090 -655 14100 -630
rect 14055 -675 14100 -655
rect 14055 -700 14065 -675
rect 14090 -700 14100 -675
rect 14055 -725 14100 -700
rect 14055 -750 14065 -725
rect 14090 -750 14100 -725
rect 14055 -770 14100 -750
rect 14115 -585 14160 -575
rect 14115 -610 14125 -585
rect 14150 -610 14160 -585
rect 14115 -630 14160 -610
rect 14115 -655 14125 -630
rect 14150 -655 14160 -630
rect 14115 -675 14160 -655
rect 14115 -700 14125 -675
rect 14150 -700 14160 -675
rect 14115 -725 14160 -700
rect 14115 -750 14125 -725
rect 14150 -750 14160 -725
rect 14115 -770 14160 -750
rect 14175 -585 14220 -575
rect 14175 -610 14185 -585
rect 14210 -610 14220 -585
rect 14175 -630 14220 -610
rect 14175 -655 14185 -630
rect 14210 -655 14220 -630
rect 14175 -675 14220 -655
rect 14175 -700 14185 -675
rect 14210 -700 14220 -675
rect 14175 -725 14220 -700
rect 14175 -750 14185 -725
rect 14210 -750 14220 -725
rect 14175 -770 14220 -750
rect 14235 -585 14280 -575
rect 14235 -610 14245 -585
rect 14270 -610 14280 -585
rect 14235 -630 14280 -610
rect 14235 -655 14245 -630
rect 14270 -655 14280 -630
rect 14235 -675 14280 -655
rect 14235 -700 14245 -675
rect 14270 -700 14280 -675
rect 14235 -725 14280 -700
rect 14235 -750 14245 -725
rect 14270 -750 14280 -725
rect 14235 -770 14280 -750
rect 14295 -585 14340 -575
rect 14295 -610 14305 -585
rect 14330 -610 14340 -585
rect 14295 -630 14340 -610
rect 14295 -655 14305 -630
rect 14330 -655 14340 -630
rect 14295 -675 14340 -655
rect 14295 -700 14305 -675
rect 14330 -700 14340 -675
rect 14295 -725 14340 -700
rect 14295 -750 14305 -725
rect 14330 -750 14340 -725
rect 14295 -770 14340 -750
rect 14355 -585 14400 -575
rect 14355 -610 14365 -585
rect 14390 -610 14400 -585
rect 14355 -630 14400 -610
rect 14355 -655 14365 -630
rect 14390 -655 14400 -630
rect 14355 -675 14400 -655
rect 14355 -700 14365 -675
rect 14390 -700 14400 -675
rect 14355 -725 14400 -700
rect 14355 -750 14365 -725
rect 14390 -750 14400 -725
rect 14355 -770 14400 -750
rect 14415 -585 14460 -575
rect 14415 -610 14425 -585
rect 14450 -610 14460 -585
rect 14415 -630 14460 -610
rect 14415 -655 14425 -630
rect 14450 -655 14460 -630
rect 14415 -675 14460 -655
rect 14415 -700 14425 -675
rect 14450 -700 14460 -675
rect 14415 -725 14460 -700
rect 14415 -750 14425 -725
rect 14450 -750 14460 -725
rect 14415 -770 14460 -750
rect 14475 -585 14520 -575
rect 14475 -610 14485 -585
rect 14510 -610 14520 -585
rect 14475 -630 14520 -610
rect 14475 -655 14485 -630
rect 14510 -655 14520 -630
rect 14475 -675 14520 -655
rect 14475 -700 14485 -675
rect 14510 -700 14520 -675
rect 14475 -725 14520 -700
rect 14475 -750 14485 -725
rect 14510 -750 14520 -725
rect 14475 -770 14520 -750
rect 14535 -585 14580 -575
rect 14535 -610 14545 -585
rect 14570 -610 14580 -585
rect 14535 -630 14580 -610
rect 14535 -655 14545 -630
rect 14570 -655 14580 -630
rect 14535 -675 14580 -655
rect 14535 -700 14545 -675
rect 14570 -700 14580 -675
rect 14535 -725 14580 -700
rect 14535 -750 14545 -725
rect 14570 -750 14580 -725
rect 14535 -770 14580 -750
rect 14595 -585 14640 -575
rect 14595 -610 14605 -585
rect 14630 -610 14640 -585
rect 14595 -630 14640 -610
rect 14595 -655 14605 -630
rect 14630 -655 14640 -630
rect 14595 -675 14640 -655
rect 14595 -700 14605 -675
rect 14630 -700 14640 -675
rect 14595 -725 14640 -700
rect 14595 -750 14605 -725
rect 14630 -750 14640 -725
rect 14595 -770 14640 -750
rect 14655 -585 14700 -575
rect 14655 -610 14665 -585
rect 14690 -610 14700 -585
rect 14655 -630 14700 -610
rect 14655 -655 14665 -630
rect 14690 -655 14700 -630
rect 14655 -675 14700 -655
rect 14655 -700 14665 -675
rect 14690 -700 14700 -675
rect 14655 -725 14700 -700
rect 14655 -750 14665 -725
rect 14690 -750 14700 -725
rect 14655 -770 14700 -750
rect 14715 -585 14760 -575
rect 14715 -610 14725 -585
rect 14750 -610 14760 -585
rect 14715 -630 14760 -610
rect 14715 -655 14725 -630
rect 14750 -655 14760 -630
rect 14715 -675 14760 -655
rect 14715 -700 14725 -675
rect 14750 -700 14760 -675
rect 14715 -725 14760 -700
rect 14715 -750 14725 -725
rect 14750 -750 14760 -725
rect 14715 -770 14760 -750
rect 14775 -585 14820 -575
rect 14775 -610 14785 -585
rect 14810 -610 14820 -585
rect 14775 -630 14820 -610
rect 14775 -655 14785 -630
rect 14810 -655 14820 -630
rect 14775 -675 14820 -655
rect 14775 -700 14785 -675
rect 14810 -700 14820 -675
rect 14775 -725 14820 -700
rect 14775 -750 14785 -725
rect 14810 -750 14820 -725
rect 14775 -770 14820 -750
rect 14835 -585 14880 -575
rect 14835 -610 14845 -585
rect 14870 -610 14880 -585
rect 14835 -630 14880 -610
rect 14835 -655 14845 -630
rect 14870 -655 14880 -630
rect 14835 -675 14880 -655
rect 14835 -700 14845 -675
rect 14870 -700 14880 -675
rect 14835 -725 14880 -700
rect 14835 -750 14845 -725
rect 14870 -750 14880 -725
rect 14835 -770 14880 -750
rect 14895 -585 14940 -575
rect 14895 -610 14905 -585
rect 14930 -610 14940 -585
rect 14895 -630 14940 -610
rect 14895 -655 14905 -630
rect 14930 -655 14940 -630
rect 14895 -675 14940 -655
rect 14895 -700 14905 -675
rect 14930 -700 14940 -675
rect 14895 -725 14940 -700
rect 14895 -750 14905 -725
rect 14930 -750 14940 -725
rect 14895 -770 14940 -750
rect 14955 -585 15000 -575
rect 14955 -610 14965 -585
rect 14990 -610 15000 -585
rect 14955 -630 15000 -610
rect 14955 -655 14965 -630
rect 14990 -655 15000 -630
rect 14955 -675 15000 -655
rect 14955 -700 14965 -675
rect 14990 -700 15000 -675
rect 14955 -725 15000 -700
rect 14955 -750 14965 -725
rect 14990 -750 15000 -725
rect 14955 -770 15000 -750
rect 15015 -585 15060 -575
rect 15015 -610 15025 -585
rect 15050 -610 15060 -585
rect 15015 -630 15060 -610
rect 15015 -655 15025 -630
rect 15050 -655 15060 -630
rect 15015 -675 15060 -655
rect 15015 -700 15025 -675
rect 15050 -700 15060 -675
rect 15015 -725 15060 -700
rect 15015 -750 15025 -725
rect 15050 -750 15060 -725
rect 15015 -770 15060 -750
rect 15075 -585 15120 -575
rect 15075 -610 15085 -585
rect 15110 -610 15120 -585
rect 15075 -630 15120 -610
rect 15075 -655 15085 -630
rect 15110 -655 15120 -630
rect 15075 -675 15120 -655
rect 15075 -700 15085 -675
rect 15110 -700 15120 -675
rect 15075 -725 15120 -700
rect 15075 -750 15085 -725
rect 15110 -750 15120 -725
rect 15075 -770 15120 -750
rect 15135 -585 15180 -575
rect 15135 -610 15145 -585
rect 15170 -610 15180 -585
rect 15135 -630 15180 -610
rect 15135 -655 15145 -630
rect 15170 -655 15180 -630
rect 15135 -675 15180 -655
rect 15135 -700 15145 -675
rect 15170 -700 15180 -675
rect 15135 -725 15180 -700
rect 15135 -750 15145 -725
rect 15170 -750 15180 -725
rect 15135 -770 15180 -750
rect 15195 -585 15240 -575
rect 15195 -610 15205 -585
rect 15230 -610 15240 -585
rect 15195 -630 15240 -610
rect 15195 -655 15205 -630
rect 15230 -655 15240 -630
rect 15195 -675 15240 -655
rect 15195 -700 15205 -675
rect 15230 -700 15240 -675
rect 15195 -725 15240 -700
rect 15195 -750 15205 -725
rect 15230 -750 15240 -725
rect 15195 -770 15240 -750
rect 15255 -585 15300 -575
rect 15255 -610 15265 -585
rect 15290 -610 15300 -585
rect 15255 -630 15300 -610
rect 15255 -655 15265 -630
rect 15290 -655 15300 -630
rect 15255 -675 15300 -655
rect 15255 -700 15265 -675
rect 15290 -700 15300 -675
rect 15255 -725 15300 -700
rect 15255 -750 15265 -725
rect 15290 -750 15300 -725
rect 15255 -770 15300 -750
rect 15315 -585 15360 -575
rect 15315 -610 15325 -585
rect 15350 -610 15360 -585
rect 15315 -630 15360 -610
rect 15315 -655 15325 -630
rect 15350 -655 15360 -630
rect 15315 -675 15360 -655
rect 15315 -700 15325 -675
rect 15350 -700 15360 -675
rect 15315 -725 15360 -700
rect 15315 -750 15325 -725
rect 15350 -750 15360 -725
rect 15315 -770 15360 -750
rect 15375 -585 15420 -575
rect 15375 -610 15385 -585
rect 15410 -610 15420 -585
rect 15375 -630 15420 -610
rect 15375 -655 15385 -630
rect 15410 -655 15420 -630
rect 15375 -675 15420 -655
rect 15375 -700 15385 -675
rect 15410 -700 15420 -675
rect 15375 -725 15420 -700
rect 15375 -750 15385 -725
rect 15410 -750 15420 -725
rect 15375 -770 15420 -750
rect 15435 -585 15480 -575
rect 15435 -610 15445 -585
rect 15470 -610 15480 -585
rect 15435 -630 15480 -610
rect 15435 -655 15445 -630
rect 15470 -655 15480 -630
rect 15435 -675 15480 -655
rect 15435 -700 15445 -675
rect 15470 -700 15480 -675
rect 15435 -725 15480 -700
rect 15435 -750 15445 -725
rect 15470 -750 15480 -725
rect 15435 -770 15480 -750
rect 15495 -585 15540 -575
rect 15495 -610 15505 -585
rect 15530 -610 15540 -585
rect 15495 -630 15540 -610
rect 15495 -655 15505 -630
rect 15530 -655 15540 -630
rect 15495 -675 15540 -655
rect 15495 -700 15505 -675
rect 15530 -700 15540 -675
rect 15495 -725 15540 -700
rect 15495 -750 15505 -725
rect 15530 -750 15540 -725
rect 15495 -770 15540 -750
rect 15555 -585 15600 -575
rect 15555 -610 15565 -585
rect 15590 -610 15600 -585
rect 15555 -630 15600 -610
rect 15555 -655 15565 -630
rect 15590 -655 15600 -630
rect 15555 -675 15600 -655
rect 15555 -700 15565 -675
rect 15590 -700 15600 -675
rect 15555 -725 15600 -700
rect 15555 -750 15565 -725
rect 15590 -750 15600 -725
rect 15555 -770 15600 -750
rect 15615 -585 15660 -575
rect 15615 -610 15625 -585
rect 15650 -610 15660 -585
rect 15615 -630 15660 -610
rect 15615 -655 15625 -630
rect 15650 -655 15660 -630
rect 15615 -675 15660 -655
rect 15615 -700 15625 -675
rect 15650 -700 15660 -675
rect 15615 -725 15660 -700
rect 15615 -750 15625 -725
rect 15650 -750 15660 -725
rect 15615 -770 15660 -750
rect 15675 -585 15720 -575
rect 15675 -610 15685 -585
rect 15710 -610 15720 -585
rect 15675 -630 15720 -610
rect 15675 -655 15685 -630
rect 15710 -655 15720 -630
rect 15675 -675 15720 -655
rect 15675 -700 15685 -675
rect 15710 -700 15720 -675
rect 15675 -725 15720 -700
rect 15675 -750 15685 -725
rect 15710 -750 15720 -725
rect 15675 -770 15720 -750
rect 15735 -585 15780 -575
rect 15735 -610 15745 -585
rect 15770 -610 15780 -585
rect 15735 -630 15780 -610
rect 15735 -655 15745 -630
rect 15770 -655 15780 -630
rect 15735 -675 15780 -655
rect 15735 -700 15745 -675
rect 15770 -700 15780 -675
rect 15735 -725 15780 -700
rect 15735 -750 15745 -725
rect 15770 -750 15780 -725
rect 15735 -770 15780 -750
rect 15795 -585 15840 -575
rect 15795 -610 15805 -585
rect 15830 -610 15840 -585
rect 15795 -630 15840 -610
rect 15795 -655 15805 -630
rect 15830 -655 15840 -630
rect 15795 -675 15840 -655
rect 15795 -700 15805 -675
rect 15830 -700 15840 -675
rect 15795 -725 15840 -700
rect 15795 -750 15805 -725
rect 15830 -750 15840 -725
rect 15795 -770 15840 -750
rect 15855 -585 15900 -575
rect 15855 -610 15865 -585
rect 15890 -610 15900 -585
rect 15855 -630 15900 -610
rect 15855 -655 15865 -630
rect 15890 -655 15900 -630
rect 15855 -675 15900 -655
rect 15855 -700 15865 -675
rect 15890 -700 15900 -675
rect 15855 -725 15900 -700
rect 15855 -750 15865 -725
rect 15890 -750 15900 -725
rect 15855 -770 15900 -750
rect 15915 -585 15960 -575
rect 15915 -610 15925 -585
rect 15950 -610 15960 -585
rect 15915 -630 15960 -610
rect 15915 -655 15925 -630
rect 15950 -655 15960 -630
rect 15915 -675 15960 -655
rect 15915 -700 15925 -675
rect 15950 -700 15960 -675
rect 15915 -725 15960 -700
rect 15915 -750 15925 -725
rect 15950 -750 15960 -725
rect 15915 -770 15960 -750
rect 15975 -585 16020 -575
rect 15975 -610 15985 -585
rect 16010 -610 16020 -585
rect 15975 -630 16020 -610
rect 15975 -655 15985 -630
rect 16010 -655 16020 -630
rect 15975 -675 16020 -655
rect 15975 -700 15985 -675
rect 16010 -700 16020 -675
rect 15975 -725 16020 -700
rect 15975 -750 15985 -725
rect 16010 -750 16020 -725
rect 15975 -770 16020 -750
rect 16035 -585 16080 -575
rect 16035 -610 16045 -585
rect 16070 -610 16080 -585
rect 16035 -630 16080 -610
rect 16035 -655 16045 -630
rect 16070 -655 16080 -630
rect 16035 -675 16080 -655
rect 16035 -700 16045 -675
rect 16070 -700 16080 -675
rect 16035 -725 16080 -700
rect 16035 -750 16045 -725
rect 16070 -750 16080 -725
rect 16035 -770 16080 -750
rect 16095 -585 16140 -575
rect 16095 -610 16105 -585
rect 16130 -610 16140 -585
rect 16095 -630 16140 -610
rect 16095 -655 16105 -630
rect 16130 -655 16140 -630
rect 16095 -675 16140 -655
rect 16095 -700 16105 -675
rect 16130 -700 16140 -675
rect 16095 -725 16140 -700
rect 16095 -750 16105 -725
rect 16130 -750 16140 -725
rect 16095 -770 16140 -750
rect 16155 -585 16200 -575
rect 16155 -610 16165 -585
rect 16190 -610 16200 -585
rect 16155 -630 16200 -610
rect 16155 -655 16165 -630
rect 16190 -655 16200 -630
rect 16155 -675 16200 -655
rect 16155 -700 16165 -675
rect 16190 -700 16200 -675
rect 16155 -725 16200 -700
rect 16155 -750 16165 -725
rect 16190 -750 16200 -725
rect 16155 -770 16200 -750
rect 16215 -585 16260 -575
rect 16215 -610 16225 -585
rect 16250 -610 16260 -585
rect 16215 -630 16260 -610
rect 16215 -655 16225 -630
rect 16250 -655 16260 -630
rect 16215 -675 16260 -655
rect 16215 -700 16225 -675
rect 16250 -700 16260 -675
rect 16215 -725 16260 -700
rect 16215 -750 16225 -725
rect 16250 -750 16260 -725
rect 16215 -770 16260 -750
rect 16275 -585 16320 -575
rect 16275 -610 16285 -585
rect 16310 -610 16320 -585
rect 16275 -630 16320 -610
rect 16275 -655 16285 -630
rect 16310 -655 16320 -630
rect 16275 -675 16320 -655
rect 16275 -700 16285 -675
rect 16310 -700 16320 -675
rect 16275 -725 16320 -700
rect 16275 -750 16285 -725
rect 16310 -750 16320 -725
rect 16275 -770 16320 -750
rect 16335 -585 16380 -575
rect 16335 -610 16345 -585
rect 16370 -610 16380 -585
rect 16335 -630 16380 -610
rect 16335 -655 16345 -630
rect 16370 -655 16380 -630
rect 16335 -675 16380 -655
rect 16335 -700 16345 -675
rect 16370 -700 16380 -675
rect 16335 -725 16380 -700
rect 16335 -750 16345 -725
rect 16370 -750 16380 -725
rect 16335 -770 16380 -750
rect 16395 -585 16440 -575
rect 16395 -610 16405 -585
rect 16430 -610 16440 -585
rect 16395 -630 16440 -610
rect 16395 -655 16405 -630
rect 16430 -655 16440 -630
rect 16395 -675 16440 -655
rect 16395 -700 16405 -675
rect 16430 -700 16440 -675
rect 16395 -725 16440 -700
rect 16395 -750 16405 -725
rect 16430 -750 16440 -725
rect 16395 -770 16440 -750
rect 16455 -585 16500 -575
rect 16455 -610 16465 -585
rect 16490 -610 16500 -585
rect 16455 -630 16500 -610
rect 16455 -655 16465 -630
rect 16490 -655 16500 -630
rect 16455 -675 16500 -655
rect 16455 -700 16465 -675
rect 16490 -700 16500 -675
rect 16455 -725 16500 -700
rect 16455 -750 16465 -725
rect 16490 -750 16500 -725
rect 16455 -770 16500 -750
rect 16515 -585 16560 -575
rect 16515 -610 16525 -585
rect 16550 -610 16560 -585
rect 16515 -630 16560 -610
rect 16515 -655 16525 -630
rect 16550 -655 16560 -630
rect 16515 -675 16560 -655
rect 16515 -700 16525 -675
rect 16550 -700 16560 -675
rect 16515 -725 16560 -700
rect 16515 -750 16525 -725
rect 16550 -750 16560 -725
rect 16515 -770 16560 -750
rect 16575 -585 16620 -575
rect 16575 -610 16585 -585
rect 16610 -610 16620 -585
rect 16575 -630 16620 -610
rect 16575 -655 16585 -630
rect 16610 -655 16620 -630
rect 16575 -675 16620 -655
rect 16575 -700 16585 -675
rect 16610 -700 16620 -675
rect 16575 -725 16620 -700
rect 16575 -750 16585 -725
rect 16610 -750 16620 -725
rect 16575 -770 16620 -750
rect 16635 -585 16680 -575
rect 16635 -610 16645 -585
rect 16670 -610 16680 -585
rect 16635 -630 16680 -610
rect 16635 -655 16645 -630
rect 16670 -655 16680 -630
rect 16635 -675 16680 -655
rect 16635 -700 16645 -675
rect 16670 -700 16680 -675
rect 16635 -725 16680 -700
rect 16635 -750 16645 -725
rect 16670 -750 16680 -725
rect 16635 -770 16680 -750
rect 16695 -585 16740 -575
rect 16695 -610 16705 -585
rect 16730 -610 16740 -585
rect 16695 -630 16740 -610
rect 16695 -655 16705 -630
rect 16730 -655 16740 -630
rect 16695 -675 16740 -655
rect 16695 -700 16705 -675
rect 16730 -700 16740 -675
rect 16695 -725 16740 -700
rect 16695 -750 16705 -725
rect 16730 -750 16740 -725
rect 16695 -770 16740 -750
rect 16755 -585 16800 -575
rect 16755 -610 16765 -585
rect 16790 -610 16800 -585
rect 16755 -630 16800 -610
rect 16755 -655 16765 -630
rect 16790 -655 16800 -630
rect 16755 -675 16800 -655
rect 16755 -700 16765 -675
rect 16790 -700 16800 -675
rect 16755 -725 16800 -700
rect 16755 -750 16765 -725
rect 16790 -750 16800 -725
rect 16755 -770 16800 -750
rect 16815 -585 16860 -575
rect 16815 -610 16825 -585
rect 16850 -610 16860 -585
rect 16815 -630 16860 -610
rect 16815 -655 16825 -630
rect 16850 -655 16860 -630
rect 16815 -675 16860 -655
rect 16815 -700 16825 -675
rect 16850 -700 16860 -675
rect 16815 -725 16860 -700
rect 16815 -750 16825 -725
rect 16850 -750 16860 -725
rect 16815 -770 16860 -750
rect 16875 -585 16920 -575
rect 16875 -610 16885 -585
rect 16910 -610 16920 -585
rect 16875 -630 16920 -610
rect 16875 -655 16885 -630
rect 16910 -655 16920 -630
rect 16875 -675 16920 -655
rect 16875 -700 16885 -675
rect 16910 -700 16920 -675
rect 16875 -725 16920 -700
rect 16875 -750 16885 -725
rect 16910 -750 16920 -725
rect 16875 -770 16920 -750
rect 16935 -585 16980 -575
rect 16935 -610 16945 -585
rect 16970 -610 16980 -585
rect 16935 -630 16980 -610
rect 16935 -655 16945 -630
rect 16970 -655 16980 -630
rect 16935 -675 16980 -655
rect 16935 -700 16945 -675
rect 16970 -700 16980 -675
rect 16935 -725 16980 -700
rect 16935 -750 16945 -725
rect 16970 -750 16980 -725
rect 16935 -770 16980 -750
rect 16995 -585 17040 -575
rect 16995 -610 17005 -585
rect 17030 -610 17040 -585
rect 16995 -630 17040 -610
rect 16995 -655 17005 -630
rect 17030 -655 17040 -630
rect 16995 -675 17040 -655
rect 16995 -700 17005 -675
rect 17030 -700 17040 -675
rect 16995 -725 17040 -700
rect 16995 -750 17005 -725
rect 17030 -750 17040 -725
rect 16995 -770 17040 -750
rect 17055 -585 17100 -575
rect 17055 -610 17065 -585
rect 17090 -610 17100 -585
rect 17055 -630 17100 -610
rect 17055 -655 17065 -630
rect 17090 -655 17100 -630
rect 17055 -675 17100 -655
rect 17055 -700 17065 -675
rect 17090 -700 17100 -675
rect 17055 -725 17100 -700
rect 17055 -750 17065 -725
rect 17090 -750 17100 -725
rect 17055 -770 17100 -750
rect 17115 -585 17160 -575
rect 17115 -610 17125 -585
rect 17150 -610 17160 -585
rect 17115 -630 17160 -610
rect 17115 -655 17125 -630
rect 17150 -655 17160 -630
rect 17115 -675 17160 -655
rect 17115 -700 17125 -675
rect 17150 -700 17160 -675
rect 17115 -725 17160 -700
rect 17115 -750 17125 -725
rect 17150 -750 17160 -725
rect 17115 -770 17160 -750
rect 17175 -585 17220 -575
rect 17175 -610 17185 -585
rect 17210 -610 17220 -585
rect 17175 -630 17220 -610
rect 17175 -655 17185 -630
rect 17210 -655 17220 -630
rect 17175 -675 17220 -655
rect 17175 -700 17185 -675
rect 17210 -700 17220 -675
rect 17175 -725 17220 -700
rect 17175 -750 17185 -725
rect 17210 -750 17220 -725
rect 17175 -770 17220 -750
rect 17235 -585 17280 -575
rect 17235 -610 17245 -585
rect 17270 -610 17280 -585
rect 17235 -630 17280 -610
rect 17235 -655 17245 -630
rect 17270 -655 17280 -630
rect 17235 -675 17280 -655
rect 17235 -700 17245 -675
rect 17270 -700 17280 -675
rect 17235 -725 17280 -700
rect 17235 -750 17245 -725
rect 17270 -750 17280 -725
rect 17235 -770 17280 -750
rect 17295 -585 17340 -575
rect 17295 -610 17305 -585
rect 17330 -610 17340 -585
rect 17295 -630 17340 -610
rect 17295 -655 17305 -630
rect 17330 -655 17340 -630
rect 17295 -675 17340 -655
rect 17295 -700 17305 -675
rect 17330 -700 17340 -675
rect 17295 -725 17340 -700
rect 17295 -750 17305 -725
rect 17330 -750 17340 -725
rect 17295 -770 17340 -750
rect 17355 -585 17400 -575
rect 17355 -610 17365 -585
rect 17390 -610 17400 -585
rect 17355 -630 17400 -610
rect 17355 -655 17365 -630
rect 17390 -655 17400 -630
rect 17355 -675 17400 -655
rect 17355 -700 17365 -675
rect 17390 -700 17400 -675
rect 17355 -725 17400 -700
rect 17355 -750 17365 -725
rect 17390 -750 17400 -725
rect 17355 -770 17400 -750
rect 17415 -585 17460 -575
rect 17415 -610 17425 -585
rect 17450 -610 17460 -585
rect 17415 -630 17460 -610
rect 17415 -655 17425 -630
rect 17450 -655 17460 -630
rect 17415 -675 17460 -655
rect 17415 -700 17425 -675
rect 17450 -700 17460 -675
rect 17415 -725 17460 -700
rect 17415 -750 17425 -725
rect 17450 -750 17460 -725
rect 17415 -770 17460 -750
rect 17475 -585 17520 -575
rect 17475 -610 17485 -585
rect 17510 -610 17520 -585
rect 17475 -630 17520 -610
rect 17475 -655 17485 -630
rect 17510 -655 17520 -630
rect 17475 -675 17520 -655
rect 17475 -700 17485 -675
rect 17510 -700 17520 -675
rect 17475 -725 17520 -700
rect 17475 -750 17485 -725
rect 17510 -750 17520 -725
rect 17475 -770 17520 -750
rect 17535 -585 17580 -575
rect 17535 -610 17545 -585
rect 17570 -610 17580 -585
rect 17535 -630 17580 -610
rect 17535 -655 17545 -630
rect 17570 -655 17580 -630
rect 17535 -675 17580 -655
rect 17535 -700 17545 -675
rect 17570 -700 17580 -675
rect 17535 -725 17580 -700
rect 17535 -750 17545 -725
rect 17570 -750 17580 -725
rect 17535 -770 17580 -750
rect 17595 -585 17640 -575
rect 17595 -610 17605 -585
rect 17630 -610 17640 -585
rect 17595 -630 17640 -610
rect 17595 -655 17605 -630
rect 17630 -655 17640 -630
rect 17595 -675 17640 -655
rect 17595 -700 17605 -675
rect 17630 -700 17640 -675
rect 17595 -725 17640 -700
rect 17595 -750 17605 -725
rect 17630 -750 17640 -725
rect 17595 -770 17640 -750
rect 17655 -585 17700 -575
rect 17655 -610 17665 -585
rect 17690 -610 17700 -585
rect 17655 -630 17700 -610
rect 17655 -655 17665 -630
rect 17690 -655 17700 -630
rect 17655 -675 17700 -655
rect 17655 -700 17665 -675
rect 17690 -700 17700 -675
rect 17655 -725 17700 -700
rect 17655 -750 17665 -725
rect 17690 -750 17700 -725
rect 17655 -770 17700 -750
rect 17715 -585 17760 -575
rect 17715 -610 17725 -585
rect 17750 -610 17760 -585
rect 17715 -630 17760 -610
rect 17715 -655 17725 -630
rect 17750 -655 17760 -630
rect 17715 -675 17760 -655
rect 17715 -700 17725 -675
rect 17750 -700 17760 -675
rect 17715 -725 17760 -700
rect 17715 -750 17725 -725
rect 17750 -750 17760 -725
rect 17715 -770 17760 -750
rect 17775 -585 17820 -575
rect 17775 -610 17785 -585
rect 17810 -610 17820 -585
rect 17775 -630 17820 -610
rect 17775 -655 17785 -630
rect 17810 -655 17820 -630
rect 17775 -675 17820 -655
rect 17775 -700 17785 -675
rect 17810 -700 17820 -675
rect 17775 -725 17820 -700
rect 17775 -750 17785 -725
rect 17810 -750 17820 -725
rect 17775 -770 17820 -750
rect 17835 -585 17880 -575
rect 17835 -610 17845 -585
rect 17870 -610 17880 -585
rect 17835 -630 17880 -610
rect 17835 -655 17845 -630
rect 17870 -655 17880 -630
rect 17835 -675 17880 -655
rect 17835 -700 17845 -675
rect 17870 -700 17880 -675
rect 17835 -725 17880 -700
rect 17835 -750 17845 -725
rect 17870 -750 17880 -725
rect 17835 -770 17880 -750
rect 17895 -585 17940 -575
rect 17895 -610 17905 -585
rect 17930 -610 17940 -585
rect 17895 -630 17940 -610
rect 17895 -655 17905 -630
rect 17930 -655 17940 -630
rect 17895 -675 17940 -655
rect 17895 -700 17905 -675
rect 17930 -700 17940 -675
rect 17895 -725 17940 -700
rect 17895 -750 17905 -725
rect 17930 -750 17940 -725
rect 17895 -770 17940 -750
rect 17955 -585 18000 -575
rect 17955 -610 17965 -585
rect 17990 -610 18000 -585
rect 17955 -630 18000 -610
rect 17955 -655 17965 -630
rect 17990 -655 18000 -630
rect 17955 -675 18000 -655
rect 17955 -700 17965 -675
rect 17990 -700 18000 -675
rect 17955 -725 18000 -700
rect 17955 -750 17965 -725
rect 17990 -750 18000 -725
rect 17955 -770 18000 -750
rect 18015 -585 18060 -575
rect 18015 -610 18025 -585
rect 18050 -610 18060 -585
rect 18015 -630 18060 -610
rect 18015 -655 18025 -630
rect 18050 -655 18060 -630
rect 18015 -675 18060 -655
rect 18015 -700 18025 -675
rect 18050 -700 18060 -675
rect 18015 -725 18060 -700
rect 18015 -750 18025 -725
rect 18050 -750 18060 -725
rect 18015 -770 18060 -750
rect 18075 -585 18120 -575
rect 18075 -610 18085 -585
rect 18110 -610 18120 -585
rect 18075 -630 18120 -610
rect 18075 -655 18085 -630
rect 18110 -655 18120 -630
rect 18075 -675 18120 -655
rect 18075 -700 18085 -675
rect 18110 -700 18120 -675
rect 18075 -725 18120 -700
rect 18075 -750 18085 -725
rect 18110 -750 18120 -725
rect 18075 -770 18120 -750
rect 18135 -585 18180 -575
rect 18135 -610 18145 -585
rect 18170 -610 18180 -585
rect 18135 -630 18180 -610
rect 18135 -655 18145 -630
rect 18170 -655 18180 -630
rect 18135 -675 18180 -655
rect 18135 -700 18145 -675
rect 18170 -700 18180 -675
rect 18135 -725 18180 -700
rect 18135 -750 18145 -725
rect 18170 -750 18180 -725
rect 18135 -770 18180 -750
rect 18195 -585 18240 -575
rect 18195 -610 18205 -585
rect 18230 -610 18240 -585
rect 18195 -630 18240 -610
rect 18195 -655 18205 -630
rect 18230 -655 18240 -630
rect 18195 -675 18240 -655
rect 18195 -700 18205 -675
rect 18230 -700 18240 -675
rect 18195 -725 18240 -700
rect 18195 -750 18205 -725
rect 18230 -750 18240 -725
rect 18195 -770 18240 -750
rect 18255 -585 18300 -575
rect 18255 -610 18265 -585
rect 18290 -610 18300 -585
rect 18255 -630 18300 -610
rect 18255 -655 18265 -630
rect 18290 -655 18300 -630
rect 18255 -675 18300 -655
rect 18255 -700 18265 -675
rect 18290 -700 18300 -675
rect 18255 -725 18300 -700
rect 18255 -750 18265 -725
rect 18290 -750 18300 -725
rect 18255 -770 18300 -750
rect 18315 -585 18360 -575
rect 18315 -610 18325 -585
rect 18350 -610 18360 -585
rect 18315 -630 18360 -610
rect 18315 -655 18325 -630
rect 18350 -655 18360 -630
rect 18315 -675 18360 -655
rect 18315 -700 18325 -675
rect 18350 -700 18360 -675
rect 18315 -725 18360 -700
rect 18315 -750 18325 -725
rect 18350 -750 18360 -725
rect 18315 -770 18360 -750
rect 18375 -585 18420 -575
rect 18375 -610 18385 -585
rect 18410 -610 18420 -585
rect 18375 -630 18420 -610
rect 18375 -655 18385 -630
rect 18410 -655 18420 -630
rect 18375 -675 18420 -655
rect 18375 -700 18385 -675
rect 18410 -700 18420 -675
rect 18375 -725 18420 -700
rect 18375 -750 18385 -725
rect 18410 -750 18420 -725
rect 18375 -770 18420 -750
rect 18435 -585 18480 -575
rect 18435 -610 18445 -585
rect 18470 -610 18480 -585
rect 18435 -630 18480 -610
rect 18435 -655 18445 -630
rect 18470 -655 18480 -630
rect 18435 -675 18480 -655
rect 18435 -700 18445 -675
rect 18470 -700 18480 -675
rect 18435 -725 18480 -700
rect 18435 -750 18445 -725
rect 18470 -750 18480 -725
rect 18435 -770 18480 -750
rect 18495 -585 18540 -575
rect 18495 -610 18505 -585
rect 18530 -610 18540 -585
rect 18495 -630 18540 -610
rect 18495 -655 18505 -630
rect 18530 -655 18540 -630
rect 18495 -675 18540 -655
rect 18495 -700 18505 -675
rect 18530 -700 18540 -675
rect 18495 -725 18540 -700
rect 18495 -750 18505 -725
rect 18530 -750 18540 -725
rect 18495 -770 18540 -750
rect 18555 -585 18600 -575
rect 18555 -610 18565 -585
rect 18590 -610 18600 -585
rect 18555 -630 18600 -610
rect 18555 -655 18565 -630
rect 18590 -655 18600 -630
rect 18555 -675 18600 -655
rect 18555 -700 18565 -675
rect 18590 -700 18600 -675
rect 18555 -725 18600 -700
rect 18555 -750 18565 -725
rect 18590 -750 18600 -725
rect 18555 -770 18600 -750
rect 18615 -585 18660 -575
rect 18615 -610 18625 -585
rect 18650 -610 18660 -585
rect 18615 -630 18660 -610
rect 18615 -655 18625 -630
rect 18650 -655 18660 -630
rect 18615 -675 18660 -655
rect 18615 -700 18625 -675
rect 18650 -700 18660 -675
rect 18615 -725 18660 -700
rect 18615 -750 18625 -725
rect 18650 -750 18660 -725
rect 18615 -770 18660 -750
rect 18675 -585 18720 -575
rect 18675 -610 18685 -585
rect 18710 -610 18720 -585
rect 18675 -630 18720 -610
rect 18675 -655 18685 -630
rect 18710 -655 18720 -630
rect 18675 -675 18720 -655
rect 18675 -700 18685 -675
rect 18710 -700 18720 -675
rect 18675 -725 18720 -700
rect 18675 -750 18685 -725
rect 18710 -750 18720 -725
rect 18675 -770 18720 -750
rect 18735 -585 18780 -575
rect 18735 -610 18745 -585
rect 18770 -610 18780 -585
rect 18735 -630 18780 -610
rect 18735 -655 18745 -630
rect 18770 -655 18780 -630
rect 18735 -675 18780 -655
rect 18735 -700 18745 -675
rect 18770 -700 18780 -675
rect 18735 -725 18780 -700
rect 18735 -750 18745 -725
rect 18770 -750 18780 -725
rect 18735 -770 18780 -750
rect 18795 -585 18840 -575
rect 18795 -610 18805 -585
rect 18830 -610 18840 -585
rect 18795 -630 18840 -610
rect 18795 -655 18805 -630
rect 18830 -655 18840 -630
rect 18795 -675 18840 -655
rect 18795 -700 18805 -675
rect 18830 -700 18840 -675
rect 18795 -725 18840 -700
rect 18795 -750 18805 -725
rect 18830 -750 18840 -725
rect 18795 -770 18840 -750
rect 18855 -585 18900 -575
rect 18855 -610 18865 -585
rect 18890 -610 18900 -585
rect 18855 -630 18900 -610
rect 18855 -655 18865 -630
rect 18890 -655 18900 -630
rect 18855 -675 18900 -655
rect 18855 -700 18865 -675
rect 18890 -700 18900 -675
rect 18855 -725 18900 -700
rect 18855 -750 18865 -725
rect 18890 -750 18900 -725
rect 18855 -770 18900 -750
rect 18915 -585 18960 -575
rect 18915 -610 18925 -585
rect 18950 -610 18960 -585
rect 18915 -630 18960 -610
rect 18915 -655 18925 -630
rect 18950 -655 18960 -630
rect 18915 -675 18960 -655
rect 18915 -700 18925 -675
rect 18950 -700 18960 -675
rect 18915 -725 18960 -700
rect 18915 -750 18925 -725
rect 18950 -750 18960 -725
rect 18915 -770 18960 -750
rect 18975 -585 19020 -575
rect 18975 -610 18985 -585
rect 19010 -610 19020 -585
rect 18975 -630 19020 -610
rect 18975 -655 18985 -630
rect 19010 -655 19020 -630
rect 18975 -675 19020 -655
rect 18975 -700 18985 -675
rect 19010 -700 19020 -675
rect 18975 -725 19020 -700
rect 18975 -750 18985 -725
rect 19010 -750 19020 -725
rect 18975 -770 19020 -750
rect 19035 -585 19080 -575
rect 19035 -610 19045 -585
rect 19070 -610 19080 -585
rect 19035 -630 19080 -610
rect 19035 -655 19045 -630
rect 19070 -655 19080 -630
rect 19035 -675 19080 -655
rect 19035 -700 19045 -675
rect 19070 -700 19080 -675
rect 19035 -725 19080 -700
rect 19035 -750 19045 -725
rect 19070 -750 19080 -725
rect 19035 -770 19080 -750
rect 19095 -585 19140 -575
rect 19095 -610 19105 -585
rect 19130 -610 19140 -585
rect 19095 -630 19140 -610
rect 19095 -655 19105 -630
rect 19130 -655 19140 -630
rect 19095 -675 19140 -655
rect 19095 -700 19105 -675
rect 19130 -700 19140 -675
rect 19095 -725 19140 -700
rect 19095 -750 19105 -725
rect 19130 -750 19140 -725
rect 19095 -770 19140 -750
rect 19155 -585 19200 -575
rect 19155 -610 19165 -585
rect 19190 -610 19200 -585
rect 19155 -630 19200 -610
rect 19155 -655 19165 -630
rect 19190 -655 19200 -630
rect 19155 -675 19200 -655
rect 19155 -700 19165 -675
rect 19190 -700 19200 -675
rect 19155 -725 19200 -700
rect 19155 -750 19165 -725
rect 19190 -750 19200 -725
rect 19155 -770 19200 -750
rect 19215 -585 19260 -575
rect 19215 -610 19225 -585
rect 19250 -610 19260 -585
rect 19215 -630 19260 -610
rect 19215 -655 19225 -630
rect 19250 -655 19260 -630
rect 19215 -675 19260 -655
rect 19215 -700 19225 -675
rect 19250 -700 19260 -675
rect 19215 -725 19260 -700
rect 19215 -750 19225 -725
rect 19250 -750 19260 -725
rect 19215 -770 19260 -750
rect 19275 -585 19320 -575
rect 19275 -610 19285 -585
rect 19310 -610 19320 -585
rect 19275 -630 19320 -610
rect 19275 -655 19285 -630
rect 19310 -655 19320 -630
rect 19275 -675 19320 -655
rect 19275 -700 19285 -675
rect 19310 -700 19320 -675
rect 19275 -725 19320 -700
rect 19275 -750 19285 -725
rect 19310 -750 19320 -725
rect 19275 -770 19320 -750
rect 19335 -585 19380 -575
rect 19335 -610 19345 -585
rect 19370 -610 19380 -585
rect 19335 -630 19380 -610
rect 19335 -655 19345 -630
rect 19370 -655 19380 -630
rect 19335 -675 19380 -655
rect 19335 -700 19345 -675
rect 19370 -700 19380 -675
rect 19335 -725 19380 -700
rect 19335 -750 19345 -725
rect 19370 -750 19380 -725
rect 19335 -770 19380 -750
rect 19395 -585 19440 -575
rect 19395 -610 19405 -585
rect 19430 -610 19440 -585
rect 19395 -630 19440 -610
rect 19395 -655 19405 -630
rect 19430 -655 19440 -630
rect 19395 -675 19440 -655
rect 19395 -700 19405 -675
rect 19430 -700 19440 -675
rect 19395 -725 19440 -700
rect 19395 -750 19405 -725
rect 19430 -750 19440 -725
rect 19395 -770 19440 -750
rect 19455 -585 19500 -575
rect 19455 -610 19465 -585
rect 19490 -610 19500 -585
rect 19455 -630 19500 -610
rect 19455 -655 19465 -630
rect 19490 -655 19500 -630
rect 19455 -675 19500 -655
rect 19455 -700 19465 -675
rect 19490 -700 19500 -675
rect 19455 -725 19500 -700
rect 19455 -750 19465 -725
rect 19490 -750 19500 -725
rect 19455 -770 19500 -750
rect 19515 -585 19560 -575
rect 19515 -610 19525 -585
rect 19550 -610 19560 -585
rect 19515 -630 19560 -610
rect 19515 -655 19525 -630
rect 19550 -655 19560 -630
rect 19515 -675 19560 -655
rect 19515 -700 19525 -675
rect 19550 -700 19560 -675
rect 19515 -725 19560 -700
rect 19515 -750 19525 -725
rect 19550 -750 19560 -725
rect 19515 -770 19560 -750
rect 19575 -585 19620 -575
rect 19575 -610 19585 -585
rect 19610 -610 19620 -585
rect 19575 -630 19620 -610
rect 19575 -655 19585 -630
rect 19610 -655 19620 -630
rect 19575 -675 19620 -655
rect 19575 -700 19585 -675
rect 19610 -700 19620 -675
rect 19575 -725 19620 -700
rect 19575 -750 19585 -725
rect 19610 -750 19620 -725
rect 19575 -770 19620 -750
rect 19635 -585 19680 -575
rect 19635 -610 19645 -585
rect 19670 -610 19680 -585
rect 19635 -630 19680 -610
rect 19635 -655 19645 -630
rect 19670 -655 19680 -630
rect 19635 -675 19680 -655
rect 19635 -700 19645 -675
rect 19670 -700 19680 -675
rect 19635 -725 19680 -700
rect 19635 -750 19645 -725
rect 19670 -750 19680 -725
rect 19635 -770 19680 -750
rect 19695 -585 19740 -575
rect 19695 -610 19705 -585
rect 19730 -610 19740 -585
rect 19695 -630 19740 -610
rect 19695 -655 19705 -630
rect 19730 -655 19740 -630
rect 19695 -675 19740 -655
rect 19695 -700 19705 -675
rect 19730 -700 19740 -675
rect 19695 -725 19740 -700
rect 19695 -750 19705 -725
rect 19730 -750 19740 -725
rect 19695 -770 19740 -750
rect 19755 -585 19800 -575
rect 19755 -610 19765 -585
rect 19790 -610 19800 -585
rect 19755 -630 19800 -610
rect 19755 -655 19765 -630
rect 19790 -655 19800 -630
rect 19755 -675 19800 -655
rect 19755 -700 19765 -675
rect 19790 -700 19800 -675
rect 19755 -725 19800 -700
rect 19755 -750 19765 -725
rect 19790 -750 19800 -725
rect 19755 -770 19800 -750
rect 19815 -585 19860 -575
rect 19815 -610 19825 -585
rect 19850 -610 19860 -585
rect 19815 -630 19860 -610
rect 19815 -655 19825 -630
rect 19850 -655 19860 -630
rect 19815 -675 19860 -655
rect 19815 -700 19825 -675
rect 19850 -700 19860 -675
rect 19815 -725 19860 -700
rect 19815 -750 19825 -725
rect 19850 -750 19860 -725
rect 19815 -770 19860 -750
rect 19875 -585 19920 -575
rect 19875 -610 19885 -585
rect 19910 -610 19920 -585
rect 19875 -630 19920 -610
rect 19875 -655 19885 -630
rect 19910 -655 19920 -630
rect 19875 -675 19920 -655
rect 19875 -700 19885 -675
rect 19910 -700 19920 -675
rect 19875 -725 19920 -700
rect 19875 -750 19885 -725
rect 19910 -750 19920 -725
rect 19875 -770 19920 -750
rect 19935 -585 19980 -575
rect 19935 -610 19945 -585
rect 19970 -610 19980 -585
rect 19935 -630 19980 -610
rect 19935 -655 19945 -630
rect 19970 -655 19980 -630
rect 19935 -675 19980 -655
rect 19935 -700 19945 -675
rect 19970 -700 19980 -675
rect 19935 -725 19980 -700
rect 19935 -750 19945 -725
rect 19970 -750 19980 -725
rect 19935 -770 19980 -750
rect 19995 -585 20040 -575
rect 19995 -610 20005 -585
rect 20030 -610 20040 -585
rect 19995 -630 20040 -610
rect 19995 -655 20005 -630
rect 20030 -655 20040 -630
rect 19995 -675 20040 -655
rect 19995 -700 20005 -675
rect 20030 -700 20040 -675
rect 19995 -725 20040 -700
rect 19995 -750 20005 -725
rect 20030 -750 20040 -725
rect 19995 -770 20040 -750
rect 20055 -585 20100 -575
rect 20055 -610 20065 -585
rect 20090 -610 20100 -585
rect 20055 -630 20100 -610
rect 20055 -655 20065 -630
rect 20090 -655 20100 -630
rect 20055 -675 20100 -655
rect 20055 -700 20065 -675
rect 20090 -700 20100 -675
rect 20055 -725 20100 -700
rect 20055 -750 20065 -725
rect 20090 -750 20100 -725
rect 20055 -770 20100 -750
rect 20115 -585 20160 -575
rect 20115 -610 20125 -585
rect 20150 -610 20160 -585
rect 20115 -630 20160 -610
rect 20115 -655 20125 -630
rect 20150 -655 20160 -630
rect 20115 -675 20160 -655
rect 20115 -700 20125 -675
rect 20150 -700 20160 -675
rect 20115 -725 20160 -700
rect 20115 -750 20125 -725
rect 20150 -750 20160 -725
rect 20115 -770 20160 -750
rect 20175 -585 20220 -575
rect 20175 -610 20185 -585
rect 20210 -610 20220 -585
rect 20175 -630 20220 -610
rect 20175 -655 20185 -630
rect 20210 -655 20220 -630
rect 20175 -675 20220 -655
rect 20175 -700 20185 -675
rect 20210 -700 20220 -675
rect 20175 -725 20220 -700
rect 20175 -750 20185 -725
rect 20210 -750 20220 -725
rect 20175 -770 20220 -750
rect 20235 -585 20280 -575
rect 20235 -610 20245 -585
rect 20270 -610 20280 -585
rect 20235 -630 20280 -610
rect 20235 -655 20245 -630
rect 20270 -655 20280 -630
rect 20235 -675 20280 -655
rect 20235 -700 20245 -675
rect 20270 -700 20280 -675
rect 20235 -725 20280 -700
rect 20235 -750 20245 -725
rect 20270 -750 20280 -725
rect 20235 -770 20280 -750
rect 20295 -585 20340 -575
rect 20295 -610 20305 -585
rect 20330 -610 20340 -585
rect 20295 -630 20340 -610
rect 20295 -655 20305 -630
rect 20330 -655 20340 -630
rect 20295 -675 20340 -655
rect 20295 -700 20305 -675
rect 20330 -700 20340 -675
rect 20295 -725 20340 -700
rect 20295 -750 20305 -725
rect 20330 -750 20340 -725
rect 20295 -770 20340 -750
rect 20355 -585 20400 -575
rect 20355 -610 20365 -585
rect 20390 -610 20400 -585
rect 20355 -630 20400 -610
rect 20355 -655 20365 -630
rect 20390 -655 20400 -630
rect 20355 -675 20400 -655
rect 20355 -700 20365 -675
rect 20390 -700 20400 -675
rect 20355 -725 20400 -700
rect 20355 -750 20365 -725
rect 20390 -750 20400 -725
rect 20355 -770 20400 -750
rect 20415 -585 20460 -575
rect 20415 -610 20425 -585
rect 20450 -610 20460 -585
rect 20415 -630 20460 -610
rect 20415 -655 20425 -630
rect 20450 -655 20460 -630
rect 20415 -675 20460 -655
rect 20415 -700 20425 -675
rect 20450 -700 20460 -675
rect 20415 -725 20460 -700
rect 20415 -750 20425 -725
rect 20450 -750 20460 -725
rect 20415 -770 20460 -750
rect 20475 -585 20520 -575
rect 20475 -610 20485 -585
rect 20510 -610 20520 -585
rect 20475 -630 20520 -610
rect 20475 -655 20485 -630
rect 20510 -655 20520 -630
rect 20475 -675 20520 -655
rect 20475 -700 20485 -675
rect 20510 -700 20520 -675
rect 20475 -725 20520 -700
rect 20475 -750 20485 -725
rect 20510 -750 20520 -725
rect 20475 -770 20520 -750
rect 20535 -585 20580 -575
rect 20535 -610 20545 -585
rect 20570 -610 20580 -585
rect 20535 -630 20580 -610
rect 20535 -655 20545 -630
rect 20570 -655 20580 -630
rect 20535 -675 20580 -655
rect 20535 -700 20545 -675
rect 20570 -700 20580 -675
rect 20535 -725 20580 -700
rect 20535 -750 20545 -725
rect 20570 -750 20580 -725
rect 20535 -770 20580 -750
rect 20595 -585 20640 -575
rect 20595 -610 20605 -585
rect 20630 -610 20640 -585
rect 20595 -630 20640 -610
rect 20595 -655 20605 -630
rect 20630 -655 20640 -630
rect 20595 -675 20640 -655
rect 20595 -700 20605 -675
rect 20630 -700 20640 -675
rect 20595 -725 20640 -700
rect 20595 -750 20605 -725
rect 20630 -750 20640 -725
rect 20595 -770 20640 -750
rect 20655 -585 20700 -575
rect 20655 -610 20665 -585
rect 20690 -610 20700 -585
rect 20655 -630 20700 -610
rect 20655 -655 20665 -630
rect 20690 -655 20700 -630
rect 20655 -675 20700 -655
rect 20655 -700 20665 -675
rect 20690 -700 20700 -675
rect 20655 -725 20700 -700
rect 20655 -750 20665 -725
rect 20690 -750 20700 -725
rect 20655 -770 20700 -750
rect 20715 -585 20760 -575
rect 20715 -610 20725 -585
rect 20750 -610 20760 -585
rect 20715 -630 20760 -610
rect 20715 -655 20725 -630
rect 20750 -655 20760 -630
rect 20715 -675 20760 -655
rect 20715 -700 20725 -675
rect 20750 -700 20760 -675
rect 20715 -725 20760 -700
rect 20715 -750 20725 -725
rect 20750 -750 20760 -725
rect 20715 -770 20760 -750
rect 20775 -585 20820 -575
rect 20775 -610 20785 -585
rect 20810 -610 20820 -585
rect 20775 -630 20820 -610
rect 20775 -655 20785 -630
rect 20810 -655 20820 -630
rect 20775 -675 20820 -655
rect 20775 -700 20785 -675
rect 20810 -700 20820 -675
rect 20775 -725 20820 -700
rect 20775 -750 20785 -725
rect 20810 -750 20820 -725
rect 20775 -770 20820 -750
rect 20835 -585 20880 -575
rect 20835 -610 20845 -585
rect 20870 -610 20880 -585
rect 20835 -630 20880 -610
rect 20835 -655 20845 -630
rect 20870 -655 20880 -630
rect 20835 -675 20880 -655
rect 20835 -700 20845 -675
rect 20870 -700 20880 -675
rect 20835 -725 20880 -700
rect 20835 -750 20845 -725
rect 20870 -750 20880 -725
rect 20835 -770 20880 -750
rect 20895 -585 20940 -575
rect 20895 -610 20905 -585
rect 20930 -610 20940 -585
rect 20895 -630 20940 -610
rect 20895 -655 20905 -630
rect 20930 -655 20940 -630
rect 20895 -675 20940 -655
rect 20895 -700 20905 -675
rect 20930 -700 20940 -675
rect 20895 -725 20940 -700
rect 20895 -750 20905 -725
rect 20930 -750 20940 -725
rect 20895 -770 20940 -750
rect 20955 -585 21000 -575
rect 20955 -610 20965 -585
rect 20990 -610 21000 -585
rect 20955 -630 21000 -610
rect 20955 -655 20965 -630
rect 20990 -655 21000 -630
rect 20955 -675 21000 -655
rect 20955 -700 20965 -675
rect 20990 -700 21000 -675
rect 20955 -725 21000 -700
rect 20955 -750 20965 -725
rect 20990 -750 21000 -725
rect 20955 -770 21000 -750
rect 21015 -585 21060 -575
rect 21015 -610 21025 -585
rect 21050 -610 21060 -585
rect 21015 -630 21060 -610
rect 21015 -655 21025 -630
rect 21050 -655 21060 -630
rect 21015 -675 21060 -655
rect 21015 -700 21025 -675
rect 21050 -700 21060 -675
rect 21015 -725 21060 -700
rect 21015 -750 21025 -725
rect 21050 -750 21060 -725
rect 21015 -770 21060 -750
rect 21075 -585 21120 -575
rect 21075 -610 21085 -585
rect 21110 -610 21120 -585
rect 21075 -630 21120 -610
rect 21075 -655 21085 -630
rect 21110 -655 21120 -630
rect 21075 -675 21120 -655
rect 21075 -700 21085 -675
rect 21110 -700 21120 -675
rect 21075 -725 21120 -700
rect 21075 -750 21085 -725
rect 21110 -750 21120 -725
rect 21075 -770 21120 -750
rect 21135 -585 21180 -575
rect 21135 -610 21145 -585
rect 21170 -610 21180 -585
rect 21135 -630 21180 -610
rect 21135 -655 21145 -630
rect 21170 -655 21180 -630
rect 21135 -675 21180 -655
rect 21135 -700 21145 -675
rect 21170 -700 21180 -675
rect 21135 -725 21180 -700
rect 21135 -750 21145 -725
rect 21170 -750 21180 -725
rect 21135 -770 21180 -750
rect 21195 -585 21240 -575
rect 21195 -610 21205 -585
rect 21230 -610 21240 -585
rect 21195 -630 21240 -610
rect 21195 -655 21205 -630
rect 21230 -655 21240 -630
rect 21195 -675 21240 -655
rect 21195 -700 21205 -675
rect 21230 -700 21240 -675
rect 21195 -725 21240 -700
rect 21195 -750 21205 -725
rect 21230 -750 21240 -725
rect 21195 -770 21240 -750
rect 21255 -585 21300 -575
rect 21255 -610 21265 -585
rect 21290 -610 21300 -585
rect 21255 -630 21300 -610
rect 21255 -655 21265 -630
rect 21290 -655 21300 -630
rect 21255 -675 21300 -655
rect 21255 -700 21265 -675
rect 21290 -700 21300 -675
rect 21255 -725 21300 -700
rect 21255 -750 21265 -725
rect 21290 -750 21300 -725
rect 21255 -770 21300 -750
rect 21315 -585 21360 -575
rect 21315 -610 21325 -585
rect 21350 -610 21360 -585
rect 21315 -630 21360 -610
rect 21315 -655 21325 -630
rect 21350 -655 21360 -630
rect 21315 -675 21360 -655
rect 21315 -700 21325 -675
rect 21350 -700 21360 -675
rect 21315 -725 21360 -700
rect 21315 -750 21325 -725
rect 21350 -750 21360 -725
rect 21315 -770 21360 -750
rect 21375 -585 21420 -575
rect 21375 -610 21385 -585
rect 21410 -610 21420 -585
rect 21375 -630 21420 -610
rect 21375 -655 21385 -630
rect 21410 -655 21420 -630
rect 21375 -675 21420 -655
rect 21375 -700 21385 -675
rect 21410 -700 21420 -675
rect 21375 -725 21420 -700
rect 21375 -750 21385 -725
rect 21410 -750 21420 -725
rect 21375 -770 21420 -750
rect 21435 -585 21480 -575
rect 21435 -610 21445 -585
rect 21470 -610 21480 -585
rect 21435 -630 21480 -610
rect 21435 -655 21445 -630
rect 21470 -655 21480 -630
rect 21435 -675 21480 -655
rect 21435 -700 21445 -675
rect 21470 -700 21480 -675
rect 21435 -725 21480 -700
rect 21435 -750 21445 -725
rect 21470 -750 21480 -725
rect 21435 -770 21480 -750
rect 21495 -585 21540 -575
rect 21495 -610 21505 -585
rect 21530 -610 21540 -585
rect 21495 -630 21540 -610
rect 21495 -655 21505 -630
rect 21530 -655 21540 -630
rect 21495 -675 21540 -655
rect 21495 -700 21505 -675
rect 21530 -700 21540 -675
rect 21495 -725 21540 -700
rect 21495 -750 21505 -725
rect 21530 -750 21540 -725
rect 21495 -770 21540 -750
rect 21555 -585 21600 -575
rect 21555 -610 21565 -585
rect 21590 -610 21600 -585
rect 21555 -630 21600 -610
rect 21555 -655 21565 -630
rect 21590 -655 21600 -630
rect 21555 -675 21600 -655
rect 21555 -700 21565 -675
rect 21590 -700 21600 -675
rect 21555 -725 21600 -700
rect 21555 -750 21565 -725
rect 21590 -750 21600 -725
rect 21555 -770 21600 -750
rect 21615 -585 21660 -575
rect 21615 -610 21625 -585
rect 21650 -610 21660 -585
rect 21615 -630 21660 -610
rect 21615 -655 21625 -630
rect 21650 -655 21660 -630
rect 21615 -675 21660 -655
rect 21615 -700 21625 -675
rect 21650 -700 21660 -675
rect 21615 -725 21660 -700
rect 21615 -750 21625 -725
rect 21650 -750 21660 -725
rect 21615 -770 21660 -750
rect 21675 -585 21720 -575
rect 21675 -610 21685 -585
rect 21710 -610 21720 -585
rect 21675 -630 21720 -610
rect 21675 -655 21685 -630
rect 21710 -655 21720 -630
rect 21675 -675 21720 -655
rect 21675 -700 21685 -675
rect 21710 -700 21720 -675
rect 21675 -725 21720 -700
rect 21675 -750 21685 -725
rect 21710 -750 21720 -725
rect 21675 -770 21720 -750
rect 21735 -585 21780 -575
rect 21735 -610 21745 -585
rect 21770 -610 21780 -585
rect 21735 -630 21780 -610
rect 21735 -655 21745 -630
rect 21770 -655 21780 -630
rect 21735 -675 21780 -655
rect 21735 -700 21745 -675
rect 21770 -700 21780 -675
rect 21735 -725 21780 -700
rect 21735 -750 21745 -725
rect 21770 -750 21780 -725
rect 21735 -770 21780 -750
rect 21795 -585 21840 -575
rect 21795 -610 21805 -585
rect 21830 -610 21840 -585
rect 21795 -630 21840 -610
rect 21795 -655 21805 -630
rect 21830 -655 21840 -630
rect 21795 -675 21840 -655
rect 21795 -700 21805 -675
rect 21830 -700 21840 -675
rect 21795 -725 21840 -700
rect 21795 -750 21805 -725
rect 21830 -750 21840 -725
rect 21795 -770 21840 -750
rect 21855 -585 21900 -575
rect 21855 -610 21865 -585
rect 21890 -610 21900 -585
rect 21855 -630 21900 -610
rect 21855 -655 21865 -630
rect 21890 -655 21900 -630
rect 21855 -675 21900 -655
rect 21855 -700 21865 -675
rect 21890 -700 21900 -675
rect 21855 -725 21900 -700
rect 21855 -750 21865 -725
rect 21890 -750 21900 -725
rect 21855 -770 21900 -750
rect 21915 -585 21960 -575
rect 21915 -610 21925 -585
rect 21950 -610 21960 -585
rect 21915 -630 21960 -610
rect 21915 -655 21925 -630
rect 21950 -655 21960 -630
rect 21915 -675 21960 -655
rect 21915 -700 21925 -675
rect 21950 -700 21960 -675
rect 21915 -725 21960 -700
rect 21915 -750 21925 -725
rect 21950 -750 21960 -725
rect 21915 -770 21960 -750
rect 21975 -585 22020 -575
rect 21975 -610 21985 -585
rect 22010 -610 22020 -585
rect 21975 -630 22020 -610
rect 21975 -655 21985 -630
rect 22010 -655 22020 -630
rect 21975 -675 22020 -655
rect 21975 -700 21985 -675
rect 22010 -700 22020 -675
rect 21975 -725 22020 -700
rect 21975 -750 21985 -725
rect 22010 -750 22020 -725
rect 21975 -770 22020 -750
rect 22035 -585 22080 -575
rect 22035 -610 22045 -585
rect 22070 -610 22080 -585
rect 22035 -630 22080 -610
rect 22035 -655 22045 -630
rect 22070 -655 22080 -630
rect 22035 -675 22080 -655
rect 22035 -700 22045 -675
rect 22070 -700 22080 -675
rect 22035 -725 22080 -700
rect 22035 -750 22045 -725
rect 22070 -750 22080 -725
rect 22035 -770 22080 -750
rect 22095 -585 22140 -575
rect 22095 -610 22105 -585
rect 22130 -610 22140 -585
rect 22095 -630 22140 -610
rect 22095 -655 22105 -630
rect 22130 -655 22140 -630
rect 22095 -675 22140 -655
rect 22095 -700 22105 -675
rect 22130 -700 22140 -675
rect 22095 -725 22140 -700
rect 22095 -750 22105 -725
rect 22130 -750 22140 -725
rect 22095 -770 22140 -750
rect 22155 -585 22200 -575
rect 22155 -610 22165 -585
rect 22190 -610 22200 -585
rect 22155 -630 22200 -610
rect 22155 -655 22165 -630
rect 22190 -655 22200 -630
rect 22155 -675 22200 -655
rect 22155 -700 22165 -675
rect 22190 -700 22200 -675
rect 22155 -725 22200 -700
rect 22155 -750 22165 -725
rect 22190 -750 22200 -725
rect 22155 -770 22200 -750
rect 22215 -585 22260 -575
rect 22215 -610 22225 -585
rect 22250 -610 22260 -585
rect 22215 -630 22260 -610
rect 22215 -655 22225 -630
rect 22250 -655 22260 -630
rect 22215 -675 22260 -655
rect 22215 -700 22225 -675
rect 22250 -700 22260 -675
rect 22215 -725 22260 -700
rect 22215 -750 22225 -725
rect 22250 -750 22260 -725
rect 22215 -770 22260 -750
rect 22275 -585 22320 -575
rect 22275 -610 22285 -585
rect 22310 -610 22320 -585
rect 22275 -630 22320 -610
rect 22275 -655 22285 -630
rect 22310 -655 22320 -630
rect 22275 -675 22320 -655
rect 22275 -700 22285 -675
rect 22310 -700 22320 -675
rect 22275 -725 22320 -700
rect 22275 -750 22285 -725
rect 22310 -750 22320 -725
rect 22275 -770 22320 -750
rect 22335 -585 22380 -575
rect 22335 -610 22345 -585
rect 22370 -610 22380 -585
rect 22335 -630 22380 -610
rect 22335 -655 22345 -630
rect 22370 -655 22380 -630
rect 22335 -675 22380 -655
rect 22335 -700 22345 -675
rect 22370 -700 22380 -675
rect 22335 -725 22380 -700
rect 22335 -750 22345 -725
rect 22370 -750 22380 -725
rect 22335 -770 22380 -750
rect 22395 -585 22440 -575
rect 22395 -610 22405 -585
rect 22430 -610 22440 -585
rect 22395 -630 22440 -610
rect 22395 -655 22405 -630
rect 22430 -655 22440 -630
rect 22395 -675 22440 -655
rect 22395 -700 22405 -675
rect 22430 -700 22440 -675
rect 22395 -725 22440 -700
rect 22395 -750 22405 -725
rect 22430 -750 22440 -725
rect 22395 -770 22440 -750
rect 22455 -585 22500 -575
rect 22455 -610 22465 -585
rect 22490 -610 22500 -585
rect 22455 -630 22500 -610
rect 22455 -655 22465 -630
rect 22490 -655 22500 -630
rect 22455 -675 22500 -655
rect 22455 -700 22465 -675
rect 22490 -700 22500 -675
rect 22455 -725 22500 -700
rect 22455 -750 22465 -725
rect 22490 -750 22500 -725
rect 22455 -770 22500 -750
rect 22515 -585 22560 -575
rect 22515 -610 22525 -585
rect 22550 -610 22560 -585
rect 22515 -630 22560 -610
rect 22515 -655 22525 -630
rect 22550 -655 22560 -630
rect 22515 -675 22560 -655
rect 22515 -700 22525 -675
rect 22550 -700 22560 -675
rect 22515 -725 22560 -700
rect 22515 -750 22525 -725
rect 22550 -750 22560 -725
rect 22515 -770 22560 -750
rect 22575 -585 22620 -575
rect 22575 -610 22585 -585
rect 22610 -610 22620 -585
rect 22575 -630 22620 -610
rect 22575 -655 22585 -630
rect 22610 -655 22620 -630
rect 22575 -675 22620 -655
rect 22575 -700 22585 -675
rect 22610 -700 22620 -675
rect 22575 -725 22620 -700
rect 22575 -750 22585 -725
rect 22610 -750 22620 -725
rect 22575 -770 22620 -750
rect 22635 -585 22680 -575
rect 22635 -610 22645 -585
rect 22670 -610 22680 -585
rect 22635 -630 22680 -610
rect 22635 -655 22645 -630
rect 22670 -655 22680 -630
rect 22635 -675 22680 -655
rect 22635 -700 22645 -675
rect 22670 -700 22680 -675
rect 22635 -725 22680 -700
rect 22635 -750 22645 -725
rect 22670 -750 22680 -725
rect 22635 -770 22680 -750
rect 22695 -585 22740 -575
rect 22695 -610 22705 -585
rect 22730 -610 22740 -585
rect 22695 -630 22740 -610
rect 22695 -655 22705 -630
rect 22730 -655 22740 -630
rect 22695 -675 22740 -655
rect 22695 -700 22705 -675
rect 22730 -700 22740 -675
rect 22695 -725 22740 -700
rect 22695 -750 22705 -725
rect 22730 -750 22740 -725
rect 22695 -770 22740 -750
rect 22755 -585 22800 -575
rect 22755 -610 22765 -585
rect 22790 -610 22800 -585
rect 22755 -630 22800 -610
rect 22755 -655 22765 -630
rect 22790 -655 22800 -630
rect 22755 -675 22800 -655
rect 22755 -700 22765 -675
rect 22790 -700 22800 -675
rect 22755 -725 22800 -700
rect 22755 -750 22765 -725
rect 22790 -750 22800 -725
rect 22755 -770 22800 -750
rect 22815 -585 22860 -575
rect 22815 -610 22825 -585
rect 22850 -610 22860 -585
rect 22815 -630 22860 -610
rect 22815 -655 22825 -630
rect 22850 -655 22860 -630
rect 22815 -675 22860 -655
rect 22815 -700 22825 -675
rect 22850 -700 22860 -675
rect 22815 -725 22860 -700
rect 22815 -750 22825 -725
rect 22850 -750 22860 -725
rect 22815 -770 22860 -750
rect 22875 -585 22920 -575
rect 22875 -610 22885 -585
rect 22910 -610 22920 -585
rect 22875 -630 22920 -610
rect 22875 -655 22885 -630
rect 22910 -655 22920 -630
rect 22875 -675 22920 -655
rect 22875 -700 22885 -675
rect 22910 -700 22920 -675
rect 22875 -725 22920 -700
rect 22875 -750 22885 -725
rect 22910 -750 22920 -725
rect 22875 -770 22920 -750
rect 22935 -585 22980 -575
rect 22935 -610 22945 -585
rect 22970 -610 22980 -585
rect 22935 -630 22980 -610
rect 22935 -655 22945 -630
rect 22970 -655 22980 -630
rect 22935 -675 22980 -655
rect 22935 -700 22945 -675
rect 22970 -700 22980 -675
rect 22935 -725 22980 -700
rect 22935 -750 22945 -725
rect 22970 -750 22980 -725
rect 22935 -770 22980 -750
rect 22995 -585 23040 -575
rect 22995 -610 23005 -585
rect 23030 -610 23040 -585
rect 22995 -630 23040 -610
rect 22995 -655 23005 -630
rect 23030 -655 23040 -630
rect 22995 -675 23040 -655
rect 22995 -700 23005 -675
rect 23030 -700 23040 -675
rect 22995 -725 23040 -700
rect 22995 -750 23005 -725
rect 23030 -750 23040 -725
rect 22995 -770 23040 -750
rect 23055 -585 23100 -575
rect 23055 -610 23065 -585
rect 23090 -610 23100 -585
rect 23055 -630 23100 -610
rect 23055 -655 23065 -630
rect 23090 -655 23100 -630
rect 23055 -675 23100 -655
rect 23055 -700 23065 -675
rect 23090 -700 23100 -675
rect 23055 -725 23100 -700
rect 23055 -750 23065 -725
rect 23090 -750 23100 -725
rect 23055 -770 23100 -750
rect 23115 -585 23160 -575
rect 23115 -610 23125 -585
rect 23150 -610 23160 -585
rect 23115 -630 23160 -610
rect 23115 -655 23125 -630
rect 23150 -655 23160 -630
rect 23115 -675 23160 -655
rect 23115 -700 23125 -675
rect 23150 -700 23160 -675
rect 23115 -725 23160 -700
rect 23115 -750 23125 -725
rect 23150 -750 23160 -725
rect 23115 -770 23160 -750
rect 23175 -585 23220 -575
rect 23175 -610 23185 -585
rect 23210 -610 23220 -585
rect 23175 -630 23220 -610
rect 23175 -655 23185 -630
rect 23210 -655 23220 -630
rect 23175 -675 23220 -655
rect 23175 -700 23185 -675
rect 23210 -700 23220 -675
rect 23175 -725 23220 -700
rect 23175 -750 23185 -725
rect 23210 -750 23220 -725
rect 23175 -770 23220 -750
rect 23235 -585 23280 -575
rect 23235 -610 23245 -585
rect 23270 -610 23280 -585
rect 23235 -630 23280 -610
rect 23235 -655 23245 -630
rect 23270 -655 23280 -630
rect 23235 -675 23280 -655
rect 23235 -700 23245 -675
rect 23270 -700 23280 -675
rect 23235 -725 23280 -700
rect 23235 -750 23245 -725
rect 23270 -750 23280 -725
rect 23235 -770 23280 -750
rect 23295 -585 23340 -575
rect 23295 -610 23305 -585
rect 23330 -610 23340 -585
rect 23295 -630 23340 -610
rect 23295 -655 23305 -630
rect 23330 -655 23340 -630
rect 23295 -675 23340 -655
rect 23295 -700 23305 -675
rect 23330 -700 23340 -675
rect 23295 -725 23340 -700
rect 23295 -750 23305 -725
rect 23330 -750 23340 -725
rect 23295 -770 23340 -750
rect 23355 -585 23400 -575
rect 23355 -610 23365 -585
rect 23390 -610 23400 -585
rect 23355 -630 23400 -610
rect 23355 -655 23365 -630
rect 23390 -655 23400 -630
rect 23355 -675 23400 -655
rect 23355 -700 23365 -675
rect 23390 -700 23400 -675
rect 23355 -725 23400 -700
rect 23355 -750 23365 -725
rect 23390 -750 23400 -725
rect 23355 -770 23400 -750
rect 23415 -585 23460 -575
rect 23415 -610 23425 -585
rect 23450 -610 23460 -585
rect 23415 -630 23460 -610
rect 23415 -655 23425 -630
rect 23450 -655 23460 -630
rect 23415 -675 23460 -655
rect 23415 -700 23425 -675
rect 23450 -700 23460 -675
rect 23415 -725 23460 -700
rect 23415 -750 23425 -725
rect 23450 -750 23460 -725
rect 23415 -770 23460 -750
rect 23475 -585 23520 -575
rect 23475 -610 23485 -585
rect 23510 -610 23520 -585
rect 23475 -630 23520 -610
rect 23475 -655 23485 -630
rect 23510 -655 23520 -630
rect 23475 -675 23520 -655
rect 23475 -700 23485 -675
rect 23510 -700 23520 -675
rect 23475 -725 23520 -700
rect 23475 -750 23485 -725
rect 23510 -750 23520 -725
rect 23475 -770 23520 -750
rect 23535 -585 23580 -575
rect 23535 -610 23545 -585
rect 23570 -610 23580 -585
rect 23535 -630 23580 -610
rect 23535 -655 23545 -630
rect 23570 -655 23580 -630
rect 23535 -675 23580 -655
rect 23535 -700 23545 -675
rect 23570 -700 23580 -675
rect 23535 -725 23580 -700
rect 23535 -750 23545 -725
rect 23570 -750 23580 -725
rect 23535 -770 23580 -750
rect 23595 -585 23640 -575
rect 23595 -610 23605 -585
rect 23630 -610 23640 -585
rect 23595 -630 23640 -610
rect 23595 -655 23605 -630
rect 23630 -655 23640 -630
rect 23595 -675 23640 -655
rect 23595 -700 23605 -675
rect 23630 -700 23640 -675
rect 23595 -725 23640 -700
rect 23595 -750 23605 -725
rect 23630 -750 23640 -725
rect 23595 -770 23640 -750
rect 23655 -585 23700 -575
rect 23655 -610 23665 -585
rect 23690 -610 23700 -585
rect 23655 -630 23700 -610
rect 23655 -655 23665 -630
rect 23690 -655 23700 -630
rect 23655 -675 23700 -655
rect 23655 -700 23665 -675
rect 23690 -700 23700 -675
rect 23655 -725 23700 -700
rect 23655 -750 23665 -725
rect 23690 -750 23700 -725
rect 23655 -770 23700 -750
rect 23715 -585 23760 -575
rect 23715 -610 23725 -585
rect 23750 -610 23760 -585
rect 23715 -630 23760 -610
rect 23715 -655 23725 -630
rect 23750 -655 23760 -630
rect 23715 -675 23760 -655
rect 23715 -700 23725 -675
rect 23750 -700 23760 -675
rect 23715 -725 23760 -700
rect 23715 -750 23725 -725
rect 23750 -750 23760 -725
rect 23715 -770 23760 -750
rect 23775 -585 23820 -575
rect 23775 -610 23785 -585
rect 23810 -610 23820 -585
rect 23775 -630 23820 -610
rect 23775 -655 23785 -630
rect 23810 -655 23820 -630
rect 23775 -675 23820 -655
rect 23775 -700 23785 -675
rect 23810 -700 23820 -675
rect 23775 -725 23820 -700
rect 23775 -750 23785 -725
rect 23810 -750 23820 -725
rect 23775 -770 23820 -750
rect 23835 -585 23880 -575
rect 23835 -610 23845 -585
rect 23870 -610 23880 -585
rect 23835 -630 23880 -610
rect 23835 -655 23845 -630
rect 23870 -655 23880 -630
rect 23835 -675 23880 -655
rect 23835 -700 23845 -675
rect 23870 -700 23880 -675
rect 23835 -725 23880 -700
rect 23835 -750 23845 -725
rect 23870 -750 23880 -725
rect 23835 -770 23880 -750
rect 23895 -585 23940 -575
rect 23895 -610 23905 -585
rect 23930 -610 23940 -585
rect 23895 -630 23940 -610
rect 23895 -655 23905 -630
rect 23930 -655 23940 -630
rect 23895 -675 23940 -655
rect 23895 -700 23905 -675
rect 23930 -700 23940 -675
rect 23895 -725 23940 -700
rect 23895 -750 23905 -725
rect 23930 -750 23940 -725
rect 23895 -770 23940 -750
rect 23955 -585 24000 -575
rect 23955 -610 23965 -585
rect 23990 -610 24000 -585
rect 23955 -630 24000 -610
rect 23955 -655 23965 -630
rect 23990 -655 24000 -630
rect 23955 -675 24000 -655
rect 23955 -700 23965 -675
rect 23990 -700 24000 -675
rect 23955 -725 24000 -700
rect 23955 -750 23965 -725
rect 23990 -750 24000 -725
rect 23955 -770 24000 -750
rect 24015 -585 24060 -575
rect 24015 -610 24025 -585
rect 24050 -610 24060 -585
rect 24015 -630 24060 -610
rect 24015 -655 24025 -630
rect 24050 -655 24060 -630
rect 24015 -675 24060 -655
rect 24015 -700 24025 -675
rect 24050 -700 24060 -675
rect 24015 -725 24060 -700
rect 24015 -750 24025 -725
rect 24050 -750 24060 -725
rect 24015 -770 24060 -750
rect 24075 -585 24120 -575
rect 24075 -610 24085 -585
rect 24110 -610 24120 -585
rect 24075 -630 24120 -610
rect 24075 -655 24085 -630
rect 24110 -655 24120 -630
rect 24075 -675 24120 -655
rect 24075 -700 24085 -675
rect 24110 -700 24120 -675
rect 24075 -725 24120 -700
rect 24075 -750 24085 -725
rect 24110 -750 24120 -725
rect 24075 -770 24120 -750
rect 24135 -585 24180 -575
rect 24135 -610 24145 -585
rect 24170 -610 24180 -585
rect 24135 -630 24180 -610
rect 24135 -655 24145 -630
rect 24170 -655 24180 -630
rect 24135 -675 24180 -655
rect 24135 -700 24145 -675
rect 24170 -700 24180 -675
rect 24135 -725 24180 -700
rect 24135 -750 24145 -725
rect 24170 -750 24180 -725
rect 24135 -770 24180 -750
rect 24195 -585 24240 -575
rect 24195 -610 24205 -585
rect 24230 -610 24240 -585
rect 24195 -630 24240 -610
rect 24195 -655 24205 -630
rect 24230 -655 24240 -630
rect 24195 -675 24240 -655
rect 24195 -700 24205 -675
rect 24230 -700 24240 -675
rect 24195 -725 24240 -700
rect 24195 -750 24205 -725
rect 24230 -750 24240 -725
rect 24195 -770 24240 -750
rect 24255 -585 24300 -575
rect 24255 -610 24265 -585
rect 24290 -610 24300 -585
rect 24255 -630 24300 -610
rect 24255 -655 24265 -630
rect 24290 -655 24300 -630
rect 24255 -675 24300 -655
rect 24255 -700 24265 -675
rect 24290 -700 24300 -675
rect 24255 -725 24300 -700
rect 24255 -750 24265 -725
rect 24290 -750 24300 -725
rect 24255 -770 24300 -750
rect 24315 -585 24360 -575
rect 24315 -610 24325 -585
rect 24350 -610 24360 -585
rect 24315 -630 24360 -610
rect 24315 -655 24325 -630
rect 24350 -655 24360 -630
rect 24315 -675 24360 -655
rect 24315 -700 24325 -675
rect 24350 -700 24360 -675
rect 24315 -725 24360 -700
rect 24315 -750 24325 -725
rect 24350 -750 24360 -725
rect 24315 -770 24360 -750
rect 24375 -585 24420 -575
rect 24375 -610 24385 -585
rect 24410 -610 24420 -585
rect 24375 -630 24420 -610
rect 24375 -655 24385 -630
rect 24410 -655 24420 -630
rect 24375 -675 24420 -655
rect 24375 -700 24385 -675
rect 24410 -700 24420 -675
rect 24375 -725 24420 -700
rect 24375 -750 24385 -725
rect 24410 -750 24420 -725
rect 24375 -770 24420 -750
rect 24435 -585 24480 -575
rect 24435 -610 24445 -585
rect 24470 -610 24480 -585
rect 24435 -630 24480 -610
rect 24435 -655 24445 -630
rect 24470 -655 24480 -630
rect 24435 -675 24480 -655
rect 24435 -700 24445 -675
rect 24470 -700 24480 -675
rect 24435 -725 24480 -700
rect 24435 -750 24445 -725
rect 24470 -750 24480 -725
rect 24435 -770 24480 -750
rect 24495 -585 24540 -575
rect 24495 -610 24505 -585
rect 24530 -610 24540 -585
rect 24495 -630 24540 -610
rect 24495 -655 24505 -630
rect 24530 -655 24540 -630
rect 24495 -675 24540 -655
rect 24495 -700 24505 -675
rect 24530 -700 24540 -675
rect 24495 -725 24540 -700
rect 24495 -750 24505 -725
rect 24530 -750 24540 -725
rect 24495 -770 24540 -750
rect 24555 -585 24600 -575
rect 24555 -610 24565 -585
rect 24590 -610 24600 -585
rect 24555 -630 24600 -610
rect 24555 -655 24565 -630
rect 24590 -655 24600 -630
rect 24555 -675 24600 -655
rect 24555 -700 24565 -675
rect 24590 -700 24600 -675
rect 24555 -725 24600 -700
rect 24555 -750 24565 -725
rect 24590 -750 24600 -725
rect 24555 -770 24600 -750
rect 24615 -585 24660 -575
rect 24615 -610 24625 -585
rect 24650 -610 24660 -585
rect 24615 -630 24660 -610
rect 24615 -655 24625 -630
rect 24650 -655 24660 -630
rect 24615 -675 24660 -655
rect 24615 -700 24625 -675
rect 24650 -700 24660 -675
rect 24615 -725 24660 -700
rect 24615 -750 24625 -725
rect 24650 -750 24660 -725
rect 24615 -770 24660 -750
rect 24675 -585 24720 -575
rect 24675 -610 24685 -585
rect 24710 -610 24720 -585
rect 24675 -630 24720 -610
rect 24675 -655 24685 -630
rect 24710 -655 24720 -630
rect 24675 -675 24720 -655
rect 24675 -700 24685 -675
rect 24710 -700 24720 -675
rect 24675 -725 24720 -700
rect 24675 -750 24685 -725
rect 24710 -750 24720 -725
rect 24675 -770 24720 -750
rect 24735 -585 24780 -575
rect 24735 -610 24745 -585
rect 24770 -610 24780 -585
rect 24735 -630 24780 -610
rect 24735 -655 24745 -630
rect 24770 -655 24780 -630
rect 24735 -675 24780 -655
rect 24735 -700 24745 -675
rect 24770 -700 24780 -675
rect 24735 -725 24780 -700
rect 24735 -750 24745 -725
rect 24770 -750 24780 -725
rect 24735 -770 24780 -750
rect 24795 -585 24840 -575
rect 24795 -610 24805 -585
rect 24830 -610 24840 -585
rect 24795 -630 24840 -610
rect 24795 -655 24805 -630
rect 24830 -655 24840 -630
rect 24795 -675 24840 -655
rect 24795 -700 24805 -675
rect 24830 -700 24840 -675
rect 24795 -725 24840 -700
rect 24795 -750 24805 -725
rect 24830 -750 24840 -725
rect 24795 -770 24840 -750
rect 24855 -585 24900 -575
rect 24855 -610 24865 -585
rect 24890 -610 24900 -585
rect 24855 -630 24900 -610
rect 24855 -655 24865 -630
rect 24890 -655 24900 -630
rect 24855 -675 24900 -655
rect 24855 -700 24865 -675
rect 24890 -700 24900 -675
rect 24855 -725 24900 -700
rect 24855 -750 24865 -725
rect 24890 -750 24900 -725
rect 24855 -770 24900 -750
rect 24915 -585 24960 -575
rect 24915 -610 24925 -585
rect 24950 -610 24960 -585
rect 24915 -630 24960 -610
rect 24915 -655 24925 -630
rect 24950 -655 24960 -630
rect 24915 -675 24960 -655
rect 24915 -700 24925 -675
rect 24950 -700 24960 -675
rect 24915 -725 24960 -700
rect 24915 -750 24925 -725
rect 24950 -750 24960 -725
rect 24915 -770 24960 -750
rect 24975 -585 25020 -575
rect 24975 -610 24985 -585
rect 25010 -610 25020 -585
rect 24975 -630 25020 -610
rect 24975 -655 24985 -630
rect 25010 -655 25020 -630
rect 24975 -675 25020 -655
rect 24975 -700 24985 -675
rect 25010 -700 25020 -675
rect 24975 -725 25020 -700
rect 24975 -750 24985 -725
rect 25010 -750 25020 -725
rect 24975 -770 25020 -750
rect 25035 -585 25080 -575
rect 25035 -610 25045 -585
rect 25070 -610 25080 -585
rect 25035 -630 25080 -610
rect 25035 -655 25045 -630
rect 25070 -655 25080 -630
rect 25035 -675 25080 -655
rect 25035 -700 25045 -675
rect 25070 -700 25080 -675
rect 25035 -725 25080 -700
rect 25035 -750 25045 -725
rect 25070 -750 25080 -725
rect 25035 -770 25080 -750
rect 25095 -585 25140 -575
rect 25095 -610 25105 -585
rect 25130 -610 25140 -585
rect 25095 -630 25140 -610
rect 25095 -655 25105 -630
rect 25130 -655 25140 -630
rect 25095 -675 25140 -655
rect 25095 -700 25105 -675
rect 25130 -700 25140 -675
rect 25095 -725 25140 -700
rect 25095 -750 25105 -725
rect 25130 -750 25140 -725
rect 25095 -770 25140 -750
rect 25155 -585 25200 -575
rect 25155 -610 25165 -585
rect 25190 -610 25200 -585
rect 25155 -630 25200 -610
rect 25155 -655 25165 -630
rect 25190 -655 25200 -630
rect 25155 -675 25200 -655
rect 25155 -700 25165 -675
rect 25190 -700 25200 -675
rect 25155 -725 25200 -700
rect 25155 -750 25165 -725
rect 25190 -750 25200 -725
rect 25155 -770 25200 -750
rect 25215 -585 25260 -575
rect 25215 -610 25225 -585
rect 25250 -610 25260 -585
rect 25215 -630 25260 -610
rect 25215 -655 25225 -630
rect 25250 -655 25260 -630
rect 25215 -675 25260 -655
rect 25215 -700 25225 -675
rect 25250 -700 25260 -675
rect 25215 -725 25260 -700
rect 25215 -750 25225 -725
rect 25250 -750 25260 -725
rect 25215 -770 25260 -750
rect 25275 -585 25320 -575
rect 25275 -610 25285 -585
rect 25310 -610 25320 -585
rect 25275 -630 25320 -610
rect 25275 -655 25285 -630
rect 25310 -655 25320 -630
rect 25275 -675 25320 -655
rect 25275 -700 25285 -675
rect 25310 -700 25320 -675
rect 25275 -725 25320 -700
rect 25275 -750 25285 -725
rect 25310 -750 25320 -725
rect 25275 -770 25320 -750
rect 25335 -585 25380 -575
rect 25335 -610 25345 -585
rect 25370 -610 25380 -585
rect 25335 -630 25380 -610
rect 25335 -655 25345 -630
rect 25370 -655 25380 -630
rect 25335 -675 25380 -655
rect 25335 -700 25345 -675
rect 25370 -700 25380 -675
rect 25335 -725 25380 -700
rect 25335 -750 25345 -725
rect 25370 -750 25380 -725
rect 25335 -770 25380 -750
rect 25395 -585 25440 -575
rect 25395 -610 25405 -585
rect 25430 -610 25440 -585
rect 25395 -630 25440 -610
rect 25395 -655 25405 -630
rect 25430 -655 25440 -630
rect 25395 -675 25440 -655
rect 25395 -700 25405 -675
rect 25430 -700 25440 -675
rect 25395 -725 25440 -700
rect 25395 -750 25405 -725
rect 25430 -750 25440 -725
rect 25395 -770 25440 -750
rect 25455 -585 25500 -575
rect 25455 -610 25465 -585
rect 25490 -610 25500 -585
rect 25455 -630 25500 -610
rect 25455 -655 25465 -630
rect 25490 -655 25500 -630
rect 25455 -675 25500 -655
rect 25455 -700 25465 -675
rect 25490 -700 25500 -675
rect 25455 -725 25500 -700
rect 25455 -750 25465 -725
rect 25490 -750 25500 -725
rect 25455 -770 25500 -750
rect 25515 -585 25560 -575
rect 25515 -610 25525 -585
rect 25550 -610 25560 -585
rect 25515 -630 25560 -610
rect 25515 -655 25525 -630
rect 25550 -655 25560 -630
rect 25515 -675 25560 -655
rect 25515 -700 25525 -675
rect 25550 -700 25560 -675
rect 25515 -725 25560 -700
rect 25515 -750 25525 -725
rect 25550 -750 25560 -725
rect 25515 -770 25560 -750
rect 25575 -585 25620 -575
rect 25575 -610 25585 -585
rect 25610 -610 25620 -585
rect 25575 -630 25620 -610
rect 25575 -655 25585 -630
rect 25610 -655 25620 -630
rect 25575 -675 25620 -655
rect 25575 -700 25585 -675
rect 25610 -700 25620 -675
rect 25575 -725 25620 -700
rect 25575 -750 25585 -725
rect 25610 -750 25620 -725
rect 25575 -770 25620 -750
rect 25635 -585 25680 -575
rect 25635 -610 25645 -585
rect 25670 -610 25680 -585
rect 25635 -630 25680 -610
rect 25635 -655 25645 -630
rect 25670 -655 25680 -630
rect 25635 -675 25680 -655
rect 25635 -700 25645 -675
rect 25670 -700 25680 -675
rect 25635 -725 25680 -700
rect 25635 -750 25645 -725
rect 25670 -750 25680 -725
rect 25635 -770 25680 -750
rect 25695 -585 25740 -575
rect 25695 -610 25705 -585
rect 25730 -610 25740 -585
rect 25695 -630 25740 -610
rect 25695 -655 25705 -630
rect 25730 -655 25740 -630
rect 25695 -675 25740 -655
rect 25695 -700 25705 -675
rect 25730 -700 25740 -675
rect 25695 -725 25740 -700
rect 25695 -750 25705 -725
rect 25730 -750 25740 -725
rect 25695 -770 25740 -750
rect 25755 -585 25800 -575
rect 25755 -610 25765 -585
rect 25790 -610 25800 -585
rect 25755 -630 25800 -610
rect 25755 -655 25765 -630
rect 25790 -655 25800 -630
rect 25755 -675 25800 -655
rect 25755 -700 25765 -675
rect 25790 -700 25800 -675
rect 25755 -725 25800 -700
rect 25755 -750 25765 -725
rect 25790 -750 25800 -725
rect 25755 -770 25800 -750
rect 25815 -585 25860 -575
rect 25815 -610 25825 -585
rect 25850 -610 25860 -585
rect 25815 -630 25860 -610
rect 25815 -655 25825 -630
rect 25850 -655 25860 -630
rect 25815 -675 25860 -655
rect 25815 -700 25825 -675
rect 25850 -700 25860 -675
rect 25815 -725 25860 -700
rect 25815 -750 25825 -725
rect 25850 -750 25860 -725
rect 25815 -770 25860 -750
rect 25875 -585 25920 -575
rect 25875 -610 25885 -585
rect 25910 -610 25920 -585
rect 25875 -630 25920 -610
rect 25875 -655 25885 -630
rect 25910 -655 25920 -630
rect 25875 -675 25920 -655
rect 25875 -700 25885 -675
rect 25910 -700 25920 -675
rect 25875 -725 25920 -700
rect 25875 -750 25885 -725
rect 25910 -750 25920 -725
rect 25875 -770 25920 -750
rect 25935 -585 25980 -575
rect 25935 -610 25945 -585
rect 25970 -610 25980 -585
rect 25935 -630 25980 -610
rect 25935 -655 25945 -630
rect 25970 -655 25980 -630
rect 25935 -675 25980 -655
rect 25935 -700 25945 -675
rect 25970 -700 25980 -675
rect 25935 -725 25980 -700
rect 25935 -750 25945 -725
rect 25970 -750 25980 -725
rect 25935 -770 25980 -750
rect 25995 -585 26040 -575
rect 25995 -610 26005 -585
rect 26030 -610 26040 -585
rect 25995 -630 26040 -610
rect 25995 -655 26005 -630
rect 26030 -655 26040 -630
rect 25995 -675 26040 -655
rect 25995 -700 26005 -675
rect 26030 -700 26040 -675
rect 25995 -725 26040 -700
rect 25995 -750 26005 -725
rect 26030 -750 26040 -725
rect 25995 -770 26040 -750
rect 26055 -585 26100 -575
rect 26055 -610 26065 -585
rect 26090 -610 26100 -585
rect 26055 -630 26100 -610
rect 26055 -655 26065 -630
rect 26090 -655 26100 -630
rect 26055 -675 26100 -655
rect 26055 -700 26065 -675
rect 26090 -700 26100 -675
rect 26055 -725 26100 -700
rect 26055 -750 26065 -725
rect 26090 -750 26100 -725
rect 26055 -770 26100 -750
rect 26115 -585 26160 -575
rect 26115 -610 26125 -585
rect 26150 -610 26160 -585
rect 26115 -630 26160 -610
rect 26115 -655 26125 -630
rect 26150 -655 26160 -630
rect 26115 -675 26160 -655
rect 26115 -700 26125 -675
rect 26150 -700 26160 -675
rect 26115 -725 26160 -700
rect 26115 -750 26125 -725
rect 26150 -750 26160 -725
rect 26115 -770 26160 -750
rect 26175 -585 26220 -575
rect 26175 -610 26185 -585
rect 26210 -610 26220 -585
rect 26175 -630 26220 -610
rect 26175 -655 26185 -630
rect 26210 -655 26220 -630
rect 26175 -675 26220 -655
rect 26175 -700 26185 -675
rect 26210 -700 26220 -675
rect 26175 -725 26220 -700
rect 26175 -750 26185 -725
rect 26210 -750 26220 -725
rect 26175 -770 26220 -750
rect 26235 -585 26280 -575
rect 26235 -610 26245 -585
rect 26270 -610 26280 -585
rect 26235 -630 26280 -610
rect 26235 -655 26245 -630
rect 26270 -655 26280 -630
rect 26235 -675 26280 -655
rect 26235 -700 26245 -675
rect 26270 -700 26280 -675
rect 26235 -725 26280 -700
rect 26235 -750 26245 -725
rect 26270 -750 26280 -725
rect 26235 -770 26280 -750
rect 26295 -585 26340 -575
rect 26295 -610 26305 -585
rect 26330 -610 26340 -585
rect 26295 -630 26340 -610
rect 26295 -655 26305 -630
rect 26330 -655 26340 -630
rect 26295 -675 26340 -655
rect 26295 -700 26305 -675
rect 26330 -700 26340 -675
rect 26295 -725 26340 -700
rect 26295 -750 26305 -725
rect 26330 -750 26340 -725
rect 26295 -770 26340 -750
rect 26355 -585 26400 -575
rect 26355 -610 26365 -585
rect 26390 -610 26400 -585
rect 26355 -630 26400 -610
rect 26355 -655 26365 -630
rect 26390 -655 26400 -630
rect 26355 -675 26400 -655
rect 26355 -700 26365 -675
rect 26390 -700 26400 -675
rect 26355 -725 26400 -700
rect 26355 -750 26365 -725
rect 26390 -750 26400 -725
rect 26355 -770 26400 -750
rect 26415 -585 26460 -575
rect 26415 -610 26425 -585
rect 26450 -610 26460 -585
rect 26415 -630 26460 -610
rect 26415 -655 26425 -630
rect 26450 -655 26460 -630
rect 26415 -675 26460 -655
rect 26415 -700 26425 -675
rect 26450 -700 26460 -675
rect 26415 -725 26460 -700
rect 26415 -750 26425 -725
rect 26450 -750 26460 -725
rect 26415 -770 26460 -750
rect 26475 -585 26520 -575
rect 26475 -610 26485 -585
rect 26510 -610 26520 -585
rect 26475 -630 26520 -610
rect 26475 -655 26485 -630
rect 26510 -655 26520 -630
rect 26475 -675 26520 -655
rect 26475 -700 26485 -675
rect 26510 -700 26520 -675
rect 26475 -725 26520 -700
rect 26475 -750 26485 -725
rect 26510 -750 26520 -725
rect 26475 -770 26520 -750
rect 26535 -585 26580 -575
rect 26535 -610 26545 -585
rect 26570 -610 26580 -585
rect 26535 -630 26580 -610
rect 26535 -655 26545 -630
rect 26570 -655 26580 -630
rect 26535 -675 26580 -655
rect 26535 -700 26545 -675
rect 26570 -700 26580 -675
rect 26535 -725 26580 -700
rect 26535 -750 26545 -725
rect 26570 -750 26580 -725
rect 26535 -770 26580 -750
rect 26595 -585 26640 -575
rect 26595 -610 26605 -585
rect 26630 -610 26640 -585
rect 26595 -630 26640 -610
rect 26595 -655 26605 -630
rect 26630 -655 26640 -630
rect 26595 -675 26640 -655
rect 26595 -700 26605 -675
rect 26630 -700 26640 -675
rect 26595 -725 26640 -700
rect 26595 -750 26605 -725
rect 26630 -750 26640 -725
rect 26595 -770 26640 -750
rect 26655 -585 26700 -575
rect 26655 -610 26665 -585
rect 26690 -610 26700 -585
rect 26655 -630 26700 -610
rect 26655 -655 26665 -630
rect 26690 -655 26700 -630
rect 26655 -675 26700 -655
rect 26655 -700 26665 -675
rect 26690 -700 26700 -675
rect 26655 -725 26700 -700
rect 26655 -750 26665 -725
rect 26690 -750 26700 -725
rect 26655 -770 26700 -750
rect 26715 -585 26760 -575
rect 26715 -610 26725 -585
rect 26750 -610 26760 -585
rect 26715 -630 26760 -610
rect 26715 -655 26725 -630
rect 26750 -655 26760 -630
rect 26715 -675 26760 -655
rect 26715 -700 26725 -675
rect 26750 -700 26760 -675
rect 26715 -725 26760 -700
rect 26715 -750 26725 -725
rect 26750 -750 26760 -725
rect 26715 -770 26760 -750
rect 26775 -585 26820 -575
rect 26775 -610 26785 -585
rect 26810 -610 26820 -585
rect 26775 -630 26820 -610
rect 26775 -655 26785 -630
rect 26810 -655 26820 -630
rect 26775 -675 26820 -655
rect 26775 -700 26785 -675
rect 26810 -700 26820 -675
rect 26775 -725 26820 -700
rect 26775 -750 26785 -725
rect 26810 -750 26820 -725
rect 26775 -770 26820 -750
rect 26835 -585 26880 -575
rect 26835 -610 26845 -585
rect 26870 -610 26880 -585
rect 26835 -630 26880 -610
rect 26835 -655 26845 -630
rect 26870 -655 26880 -630
rect 26835 -675 26880 -655
rect 26835 -700 26845 -675
rect 26870 -700 26880 -675
rect 26835 -725 26880 -700
rect 26835 -750 26845 -725
rect 26870 -750 26880 -725
rect 26835 -770 26880 -750
rect 26895 -585 26940 -575
rect 26895 -610 26905 -585
rect 26930 -610 26940 -585
rect 26895 -630 26940 -610
rect 26895 -655 26905 -630
rect 26930 -655 26940 -630
rect 26895 -675 26940 -655
rect 26895 -700 26905 -675
rect 26930 -700 26940 -675
rect 26895 -725 26940 -700
rect 26895 -750 26905 -725
rect 26930 -750 26940 -725
rect 26895 -770 26940 -750
rect 26955 -585 27000 -575
rect 26955 -610 26965 -585
rect 26990 -610 27000 -585
rect 26955 -630 27000 -610
rect 26955 -655 26965 -630
rect 26990 -655 27000 -630
rect 26955 -675 27000 -655
rect 26955 -700 26965 -675
rect 26990 -700 27000 -675
rect 26955 -725 27000 -700
rect 26955 -750 26965 -725
rect 26990 -750 27000 -725
rect 26955 -770 27000 -750
rect 27015 -585 27060 -575
rect 27015 -610 27025 -585
rect 27050 -610 27060 -585
rect 27015 -630 27060 -610
rect 27015 -655 27025 -630
rect 27050 -655 27060 -630
rect 27015 -675 27060 -655
rect 27015 -700 27025 -675
rect 27050 -700 27060 -675
rect 27015 -725 27060 -700
rect 27015 -750 27025 -725
rect 27050 -750 27060 -725
rect 27015 -770 27060 -750
rect 27075 -585 27120 -575
rect 27075 -610 27085 -585
rect 27110 -610 27120 -585
rect 27075 -630 27120 -610
rect 27075 -655 27085 -630
rect 27110 -655 27120 -630
rect 27075 -675 27120 -655
rect 27075 -700 27085 -675
rect 27110 -700 27120 -675
rect 27075 -725 27120 -700
rect 27075 -750 27085 -725
rect 27110 -750 27120 -725
rect 27075 -770 27120 -750
rect 27135 -585 27180 -575
rect 27135 -610 27145 -585
rect 27170 -610 27180 -585
rect 27135 -630 27180 -610
rect 27135 -655 27145 -630
rect 27170 -655 27180 -630
rect 27135 -675 27180 -655
rect 27135 -700 27145 -675
rect 27170 -700 27180 -675
rect 27135 -725 27180 -700
rect 27135 -750 27145 -725
rect 27170 -750 27180 -725
rect 27135 -770 27180 -750
rect 27195 -585 27240 -575
rect 27195 -610 27205 -585
rect 27230 -610 27240 -585
rect 27195 -630 27240 -610
rect 27195 -655 27205 -630
rect 27230 -655 27240 -630
rect 27195 -675 27240 -655
rect 27195 -700 27205 -675
rect 27230 -700 27240 -675
rect 27195 -725 27240 -700
rect 27195 -750 27205 -725
rect 27230 -750 27240 -725
rect 27195 -770 27240 -750
rect 27255 -585 27300 -575
rect 27255 -610 27265 -585
rect 27290 -610 27300 -585
rect 27255 -630 27300 -610
rect 27255 -655 27265 -630
rect 27290 -655 27300 -630
rect 27255 -675 27300 -655
rect 27255 -700 27265 -675
rect 27290 -700 27300 -675
rect 27255 -725 27300 -700
rect 27255 -750 27265 -725
rect 27290 -750 27300 -725
rect 27255 -770 27300 -750
rect 27315 -585 27360 -575
rect 27315 -610 27325 -585
rect 27350 -610 27360 -585
rect 27315 -630 27360 -610
rect 27315 -655 27325 -630
rect 27350 -655 27360 -630
rect 27315 -675 27360 -655
rect 27315 -700 27325 -675
rect 27350 -700 27360 -675
rect 27315 -725 27360 -700
rect 27315 -750 27325 -725
rect 27350 -750 27360 -725
rect 27315 -770 27360 -750
rect 27375 -585 27420 -575
rect 27375 -610 27385 -585
rect 27410 -610 27420 -585
rect 27375 -630 27420 -610
rect 27375 -655 27385 -630
rect 27410 -655 27420 -630
rect 27375 -675 27420 -655
rect 27375 -700 27385 -675
rect 27410 -700 27420 -675
rect 27375 -725 27420 -700
rect 27375 -750 27385 -725
rect 27410 -750 27420 -725
rect 27375 -770 27420 -750
rect 27435 -585 27480 -575
rect 27435 -610 27445 -585
rect 27470 -610 27480 -585
rect 27435 -630 27480 -610
rect 27435 -655 27445 -630
rect 27470 -655 27480 -630
rect 27435 -675 27480 -655
rect 27435 -700 27445 -675
rect 27470 -700 27480 -675
rect 27435 -725 27480 -700
rect 27435 -750 27445 -725
rect 27470 -750 27480 -725
rect 27435 -770 27480 -750
rect 27495 -585 27540 -575
rect 27495 -610 27505 -585
rect 27530 -610 27540 -585
rect 27495 -630 27540 -610
rect 27495 -655 27505 -630
rect 27530 -655 27540 -630
rect 27495 -675 27540 -655
rect 27495 -700 27505 -675
rect 27530 -700 27540 -675
rect 27495 -725 27540 -700
rect 27495 -750 27505 -725
rect 27530 -750 27540 -725
rect 27495 -770 27540 -750
rect 27555 -585 27600 -575
rect 27555 -610 27565 -585
rect 27590 -610 27600 -585
rect 27555 -630 27600 -610
rect 27555 -655 27565 -630
rect 27590 -655 27600 -630
rect 27555 -675 27600 -655
rect 27555 -700 27565 -675
rect 27590 -700 27600 -675
rect 27555 -725 27600 -700
rect 27555 -750 27565 -725
rect 27590 -750 27600 -725
rect 27555 -770 27600 -750
rect 27615 -585 27660 -575
rect 27615 -610 27625 -585
rect 27650 -610 27660 -585
rect 27615 -630 27660 -610
rect 27615 -655 27625 -630
rect 27650 -655 27660 -630
rect 27615 -675 27660 -655
rect 27615 -700 27625 -675
rect 27650 -700 27660 -675
rect 27615 -725 27660 -700
rect 27615 -750 27625 -725
rect 27650 -750 27660 -725
rect 27615 -770 27660 -750
rect 27675 -585 27720 -575
rect 27675 -610 27685 -585
rect 27710 -610 27720 -585
rect 27675 -630 27720 -610
rect 27675 -655 27685 -630
rect 27710 -655 27720 -630
rect 27675 -675 27720 -655
rect 27675 -700 27685 -675
rect 27710 -700 27720 -675
rect 27675 -725 27720 -700
rect 27675 -750 27685 -725
rect 27710 -750 27720 -725
rect 27675 -770 27720 -750
rect 27735 -585 27780 -575
rect 27735 -610 27745 -585
rect 27770 -610 27780 -585
rect 27735 -630 27780 -610
rect 27735 -655 27745 -630
rect 27770 -655 27780 -630
rect 27735 -675 27780 -655
rect 27735 -700 27745 -675
rect 27770 -700 27780 -675
rect 27735 -725 27780 -700
rect 27735 -750 27745 -725
rect 27770 -750 27780 -725
rect 27735 -770 27780 -750
rect 27795 -585 27840 -575
rect 27795 -610 27805 -585
rect 27830 -610 27840 -585
rect 27795 -630 27840 -610
rect 27795 -655 27805 -630
rect 27830 -655 27840 -630
rect 27795 -675 27840 -655
rect 27795 -700 27805 -675
rect 27830 -700 27840 -675
rect 27795 -725 27840 -700
rect 27795 -750 27805 -725
rect 27830 -750 27840 -725
rect 27795 -770 27840 -750
rect 27855 -585 27900 -575
rect 27855 -610 27865 -585
rect 27890 -610 27900 -585
rect 27855 -630 27900 -610
rect 27855 -655 27865 -630
rect 27890 -655 27900 -630
rect 27855 -675 27900 -655
rect 27855 -700 27865 -675
rect 27890 -700 27900 -675
rect 27855 -725 27900 -700
rect 27855 -750 27865 -725
rect 27890 -750 27900 -725
rect 27855 -770 27900 -750
rect 27915 -585 27960 -575
rect 27915 -610 27925 -585
rect 27950 -610 27960 -585
rect 27915 -630 27960 -610
rect 27915 -655 27925 -630
rect 27950 -655 27960 -630
rect 27915 -675 27960 -655
rect 27915 -700 27925 -675
rect 27950 -700 27960 -675
rect 27915 -725 27960 -700
rect 27915 -750 27925 -725
rect 27950 -750 27960 -725
rect 27915 -770 27960 -750
rect 27975 -585 28020 -575
rect 27975 -610 27985 -585
rect 28010 -610 28020 -585
rect 27975 -630 28020 -610
rect 27975 -655 27985 -630
rect 28010 -655 28020 -630
rect 27975 -675 28020 -655
rect 27975 -700 27985 -675
rect 28010 -700 28020 -675
rect 27975 -725 28020 -700
rect 27975 -750 27985 -725
rect 28010 -750 28020 -725
rect 27975 -770 28020 -750
rect 28035 -585 28080 -575
rect 28035 -610 28045 -585
rect 28070 -610 28080 -585
rect 28035 -630 28080 -610
rect 28035 -655 28045 -630
rect 28070 -655 28080 -630
rect 28035 -675 28080 -655
rect 28035 -700 28045 -675
rect 28070 -700 28080 -675
rect 28035 -725 28080 -700
rect 28035 -750 28045 -725
rect 28070 -750 28080 -725
rect 28035 -770 28080 -750
rect 28095 -585 28140 -575
rect 28095 -610 28105 -585
rect 28130 -610 28140 -585
rect 28095 -630 28140 -610
rect 28095 -655 28105 -630
rect 28130 -655 28140 -630
rect 28095 -675 28140 -655
rect 28095 -700 28105 -675
rect 28130 -700 28140 -675
rect 28095 -725 28140 -700
rect 28095 -750 28105 -725
rect 28130 -750 28140 -725
rect 28095 -770 28140 -750
rect 28155 -585 28200 -575
rect 28155 -610 28165 -585
rect 28190 -610 28200 -585
rect 28155 -630 28200 -610
rect 28155 -655 28165 -630
rect 28190 -655 28200 -630
rect 28155 -675 28200 -655
rect 28155 -700 28165 -675
rect 28190 -700 28200 -675
rect 28155 -725 28200 -700
rect 28155 -750 28165 -725
rect 28190 -750 28200 -725
rect 28155 -770 28200 -750
rect 28215 -585 28260 -575
rect 28215 -610 28225 -585
rect 28250 -610 28260 -585
rect 28215 -630 28260 -610
rect 28215 -655 28225 -630
rect 28250 -655 28260 -630
rect 28215 -675 28260 -655
rect 28215 -700 28225 -675
rect 28250 -700 28260 -675
rect 28215 -725 28260 -700
rect 28215 -750 28225 -725
rect 28250 -750 28260 -725
rect 28215 -770 28260 -750
rect 28275 -585 28320 -575
rect 28275 -610 28285 -585
rect 28310 -610 28320 -585
rect 28275 -630 28320 -610
rect 28275 -655 28285 -630
rect 28310 -655 28320 -630
rect 28275 -675 28320 -655
rect 28275 -700 28285 -675
rect 28310 -700 28320 -675
rect 28275 -725 28320 -700
rect 28275 -750 28285 -725
rect 28310 -750 28320 -725
rect 28275 -770 28320 -750
rect 28335 -585 28380 -575
rect 28335 -610 28345 -585
rect 28370 -610 28380 -585
rect 28335 -630 28380 -610
rect 28335 -655 28345 -630
rect 28370 -655 28380 -630
rect 28335 -675 28380 -655
rect 28335 -700 28345 -675
rect 28370 -700 28380 -675
rect 28335 -725 28380 -700
rect 28335 -750 28345 -725
rect 28370 -750 28380 -725
rect 28335 -770 28380 -750
rect 28395 -585 28440 -575
rect 28395 -610 28405 -585
rect 28430 -610 28440 -585
rect 28395 -630 28440 -610
rect 28395 -655 28405 -630
rect 28430 -655 28440 -630
rect 28395 -675 28440 -655
rect 28395 -700 28405 -675
rect 28430 -700 28440 -675
rect 28395 -725 28440 -700
rect 28395 -750 28405 -725
rect 28430 -750 28440 -725
rect 28395 -770 28440 -750
rect 28455 -585 28500 -575
rect 28455 -610 28465 -585
rect 28490 -610 28500 -585
rect 28455 -630 28500 -610
rect 28455 -655 28465 -630
rect 28490 -655 28500 -630
rect 28455 -675 28500 -655
rect 28455 -700 28465 -675
rect 28490 -700 28500 -675
rect 28455 -725 28500 -700
rect 28455 -750 28465 -725
rect 28490 -750 28500 -725
rect 28455 -770 28500 -750
rect 28515 -585 28560 -575
rect 28515 -610 28525 -585
rect 28550 -610 28560 -585
rect 28515 -630 28560 -610
rect 28515 -655 28525 -630
rect 28550 -655 28560 -630
rect 28515 -675 28560 -655
rect 28515 -700 28525 -675
rect 28550 -700 28560 -675
rect 28515 -725 28560 -700
rect 28515 -750 28525 -725
rect 28550 -750 28560 -725
rect 28515 -770 28560 -750
rect 28575 -585 28620 -575
rect 28575 -610 28585 -585
rect 28610 -610 28620 -585
rect 28575 -630 28620 -610
rect 28575 -655 28585 -630
rect 28610 -655 28620 -630
rect 28575 -675 28620 -655
rect 28575 -700 28585 -675
rect 28610 -700 28620 -675
rect 28575 -725 28620 -700
rect 28575 -750 28585 -725
rect 28610 -750 28620 -725
rect 28575 -770 28620 -750
rect 28635 -585 28680 -575
rect 28635 -610 28645 -585
rect 28670 -610 28680 -585
rect 28635 -630 28680 -610
rect 28635 -655 28645 -630
rect 28670 -655 28680 -630
rect 28635 -675 28680 -655
rect 28635 -700 28645 -675
rect 28670 -700 28680 -675
rect 28635 -725 28680 -700
rect 28635 -750 28645 -725
rect 28670 -750 28680 -725
rect 28635 -770 28680 -750
rect 28695 -585 28740 -575
rect 28695 -610 28705 -585
rect 28730 -610 28740 -585
rect 28695 -630 28740 -610
rect 28695 -655 28705 -630
rect 28730 -655 28740 -630
rect 28695 -675 28740 -655
rect 28695 -700 28705 -675
rect 28730 -700 28740 -675
rect 28695 -725 28740 -700
rect 28695 -750 28705 -725
rect 28730 -750 28740 -725
rect 28695 -770 28740 -750
rect 28755 -585 28800 -575
rect 28755 -610 28765 -585
rect 28790 -610 28800 -585
rect 28755 -630 28800 -610
rect 28755 -655 28765 -630
rect 28790 -655 28800 -630
rect 28755 -675 28800 -655
rect 28755 -700 28765 -675
rect 28790 -700 28800 -675
rect 28755 -725 28800 -700
rect 28755 -750 28765 -725
rect 28790 -750 28800 -725
rect 28755 -770 28800 -750
rect 28815 -585 28860 -575
rect 28815 -610 28825 -585
rect 28850 -610 28860 -585
rect 28815 -630 28860 -610
rect 28815 -655 28825 -630
rect 28850 -655 28860 -630
rect 28815 -675 28860 -655
rect 28815 -700 28825 -675
rect 28850 -700 28860 -675
rect 28815 -725 28860 -700
rect 28815 -750 28825 -725
rect 28850 -750 28860 -725
rect 28815 -770 28860 -750
rect 28875 -585 28920 -575
rect 28875 -610 28885 -585
rect 28910 -610 28920 -585
rect 28875 -630 28920 -610
rect 28875 -655 28885 -630
rect 28910 -655 28920 -630
rect 28875 -675 28920 -655
rect 28875 -700 28885 -675
rect 28910 -700 28920 -675
rect 28875 -725 28920 -700
rect 28875 -750 28885 -725
rect 28910 -750 28920 -725
rect 28875 -770 28920 -750
rect 28935 -585 28980 -575
rect 28935 -610 28945 -585
rect 28970 -610 28980 -585
rect 28935 -630 28980 -610
rect 28935 -655 28945 -630
rect 28970 -655 28980 -630
rect 28935 -675 28980 -655
rect 28935 -700 28945 -675
rect 28970 -700 28980 -675
rect 28935 -725 28980 -700
rect 28935 -750 28945 -725
rect 28970 -750 28980 -725
rect 28935 -770 28980 -750
rect 28995 -585 29040 -575
rect 28995 -610 29005 -585
rect 29030 -610 29040 -585
rect 28995 -630 29040 -610
rect 28995 -655 29005 -630
rect 29030 -655 29040 -630
rect 28995 -675 29040 -655
rect 28995 -700 29005 -675
rect 29030 -700 29040 -675
rect 28995 -725 29040 -700
rect 28995 -750 29005 -725
rect 29030 -750 29040 -725
rect 28995 -770 29040 -750
rect 29055 -585 29100 -575
rect 29055 -610 29065 -585
rect 29090 -610 29100 -585
rect 29055 -630 29100 -610
rect 29055 -655 29065 -630
rect 29090 -655 29100 -630
rect 29055 -675 29100 -655
rect 29055 -700 29065 -675
rect 29090 -700 29100 -675
rect 29055 -725 29100 -700
rect 29055 -750 29065 -725
rect 29090 -750 29100 -725
rect 29055 -770 29100 -750
rect 29115 -585 29160 -575
rect 29115 -610 29125 -585
rect 29150 -610 29160 -585
rect 29115 -630 29160 -610
rect 29115 -655 29125 -630
rect 29150 -655 29160 -630
rect 29115 -675 29160 -655
rect 29115 -700 29125 -675
rect 29150 -700 29160 -675
rect 29115 -725 29160 -700
rect 29115 -750 29125 -725
rect 29150 -750 29160 -725
rect 29115 -770 29160 -750
rect 29175 -585 29220 -575
rect 29175 -610 29185 -585
rect 29210 -610 29220 -585
rect 29175 -630 29220 -610
rect 29175 -655 29185 -630
rect 29210 -655 29220 -630
rect 29175 -675 29220 -655
rect 29175 -700 29185 -675
rect 29210 -700 29220 -675
rect 29175 -725 29220 -700
rect 29175 -750 29185 -725
rect 29210 -750 29220 -725
rect 29175 -770 29220 -750
rect 29235 -585 29280 -575
rect 29235 -610 29245 -585
rect 29270 -610 29280 -585
rect 29235 -630 29280 -610
rect 29235 -655 29245 -630
rect 29270 -655 29280 -630
rect 29235 -675 29280 -655
rect 29235 -700 29245 -675
rect 29270 -700 29280 -675
rect 29235 -725 29280 -700
rect 29235 -750 29245 -725
rect 29270 -750 29280 -725
rect 29235 -770 29280 -750
rect 29295 -585 29340 -575
rect 29295 -610 29305 -585
rect 29330 -610 29340 -585
rect 29295 -630 29340 -610
rect 29295 -655 29305 -630
rect 29330 -655 29340 -630
rect 29295 -675 29340 -655
rect 29295 -700 29305 -675
rect 29330 -700 29340 -675
rect 29295 -725 29340 -700
rect 29295 -750 29305 -725
rect 29330 -750 29340 -725
rect 29295 -770 29340 -750
rect 29355 -585 29400 -575
rect 29355 -610 29365 -585
rect 29390 -610 29400 -585
rect 29355 -630 29400 -610
rect 29355 -655 29365 -630
rect 29390 -655 29400 -630
rect 29355 -675 29400 -655
rect 29355 -700 29365 -675
rect 29390 -700 29400 -675
rect 29355 -725 29400 -700
rect 29355 -750 29365 -725
rect 29390 -750 29400 -725
rect 29355 -770 29400 -750
rect 29415 -585 29460 -575
rect 29415 -610 29425 -585
rect 29450 -610 29460 -585
rect 29415 -630 29460 -610
rect 29415 -655 29425 -630
rect 29450 -655 29460 -630
rect 29415 -675 29460 -655
rect 29415 -700 29425 -675
rect 29450 -700 29460 -675
rect 29415 -725 29460 -700
rect 29415 -750 29425 -725
rect 29450 -750 29460 -725
rect 29415 -770 29460 -750
rect 29475 -585 29520 -575
rect 29475 -610 29485 -585
rect 29510 -610 29520 -585
rect 29475 -630 29520 -610
rect 29475 -655 29485 -630
rect 29510 -655 29520 -630
rect 29475 -675 29520 -655
rect 29475 -700 29485 -675
rect 29510 -700 29520 -675
rect 29475 -725 29520 -700
rect 29475 -750 29485 -725
rect 29510 -750 29520 -725
rect 29475 -770 29520 -750
rect 29535 -585 29580 -575
rect 29535 -610 29545 -585
rect 29570 -610 29580 -585
rect 29535 -630 29580 -610
rect 29535 -655 29545 -630
rect 29570 -655 29580 -630
rect 29535 -675 29580 -655
rect 29535 -700 29545 -675
rect 29570 -700 29580 -675
rect 29535 -725 29580 -700
rect 29535 -750 29545 -725
rect 29570 -750 29580 -725
rect 29535 -770 29580 -750
rect 29595 -585 29640 -575
rect 29595 -610 29605 -585
rect 29630 -610 29640 -585
rect 29595 -630 29640 -610
rect 29595 -655 29605 -630
rect 29630 -655 29640 -630
rect 29595 -675 29640 -655
rect 29595 -700 29605 -675
rect 29630 -700 29640 -675
rect 29595 -725 29640 -700
rect 29595 -750 29605 -725
rect 29630 -750 29640 -725
rect 29595 -770 29640 -750
rect 29655 -585 29700 -575
rect 29655 -610 29665 -585
rect 29690 -610 29700 -585
rect 29655 -630 29700 -610
rect 29655 -655 29665 -630
rect 29690 -655 29700 -630
rect 29655 -675 29700 -655
rect 29655 -700 29665 -675
rect 29690 -700 29700 -675
rect 29655 -725 29700 -700
rect 29655 -750 29665 -725
rect 29690 -750 29700 -725
rect 29655 -770 29700 -750
rect 29715 -585 29760 -575
rect 29715 -610 29725 -585
rect 29750 -610 29760 -585
rect 29715 -630 29760 -610
rect 29715 -655 29725 -630
rect 29750 -655 29760 -630
rect 29715 -675 29760 -655
rect 29715 -700 29725 -675
rect 29750 -700 29760 -675
rect 29715 -725 29760 -700
rect 29715 -750 29725 -725
rect 29750 -750 29760 -725
rect 29715 -770 29760 -750
rect 29775 -585 29820 -575
rect 29775 -610 29785 -585
rect 29810 -610 29820 -585
rect 29775 -630 29820 -610
rect 29775 -655 29785 -630
rect 29810 -655 29820 -630
rect 29775 -675 29820 -655
rect 29775 -700 29785 -675
rect 29810 -700 29820 -675
rect 29775 -725 29820 -700
rect 29775 -750 29785 -725
rect 29810 -750 29820 -725
rect 29775 -770 29820 -750
rect 29835 -585 29880 -575
rect 29835 -610 29845 -585
rect 29870 -610 29880 -585
rect 29835 -630 29880 -610
rect 29835 -655 29845 -630
rect 29870 -655 29880 -630
rect 29835 -675 29880 -655
rect 29835 -700 29845 -675
rect 29870 -700 29880 -675
rect 29835 -725 29880 -700
rect 29835 -750 29845 -725
rect 29870 -750 29880 -725
rect 29835 -770 29880 -750
rect 29895 -585 29940 -575
rect 29895 -610 29905 -585
rect 29930 -610 29940 -585
rect 29895 -630 29940 -610
rect 29895 -655 29905 -630
rect 29930 -655 29940 -630
rect 29895 -675 29940 -655
rect 29895 -700 29905 -675
rect 29930 -700 29940 -675
rect 29895 -725 29940 -700
rect 29895 -750 29905 -725
rect 29930 -750 29940 -725
rect 29895 -770 29940 -750
rect 29955 -585 30000 -575
rect 29955 -610 29965 -585
rect 29990 -610 30000 -585
rect 29955 -630 30000 -610
rect 29955 -655 29965 -630
rect 29990 -655 30000 -630
rect 29955 -675 30000 -655
rect 29955 -700 29965 -675
rect 29990 -700 30000 -675
rect 29955 -725 30000 -700
rect 29955 -750 29965 -725
rect 29990 -750 30000 -725
rect 29955 -770 30000 -750
rect 30015 -585 30060 -575
rect 30015 -610 30025 -585
rect 30050 -610 30060 -585
rect 30015 -630 30060 -610
rect 30015 -655 30025 -630
rect 30050 -655 30060 -630
rect 30015 -675 30060 -655
rect 30015 -700 30025 -675
rect 30050 -700 30060 -675
rect 30015 -725 30060 -700
rect 30015 -750 30025 -725
rect 30050 -750 30060 -725
rect 30015 -770 30060 -750
rect 30075 -585 30120 -575
rect 30075 -610 30085 -585
rect 30110 -610 30120 -585
rect 30075 -630 30120 -610
rect 30075 -655 30085 -630
rect 30110 -655 30120 -630
rect 30075 -675 30120 -655
rect 30075 -700 30085 -675
rect 30110 -700 30120 -675
rect 30075 -725 30120 -700
rect 30075 -750 30085 -725
rect 30110 -750 30120 -725
rect 30075 -770 30120 -750
rect 30135 -585 30180 -575
rect 30135 -610 30145 -585
rect 30170 -610 30180 -585
rect 30135 -630 30180 -610
rect 30135 -655 30145 -630
rect 30170 -655 30180 -630
rect 30135 -675 30180 -655
rect 30135 -700 30145 -675
rect 30170 -700 30180 -675
rect 30135 -725 30180 -700
rect 30135 -750 30145 -725
rect 30170 -750 30180 -725
rect 30135 -770 30180 -750
rect 30195 -585 30240 -575
rect 30195 -610 30205 -585
rect 30230 -610 30240 -585
rect 30195 -630 30240 -610
rect 30195 -655 30205 -630
rect 30230 -655 30240 -630
rect 30195 -675 30240 -655
rect 30195 -700 30205 -675
rect 30230 -700 30240 -675
rect 30195 -725 30240 -700
rect 30195 -750 30205 -725
rect 30230 -750 30240 -725
rect 30195 -770 30240 -750
rect 30255 -585 30300 -575
rect 30255 -610 30265 -585
rect 30290 -610 30300 -585
rect 30255 -630 30300 -610
rect 30255 -655 30265 -630
rect 30290 -655 30300 -630
rect 30255 -675 30300 -655
rect 30255 -700 30265 -675
rect 30290 -700 30300 -675
rect 30255 -725 30300 -700
rect 30255 -750 30265 -725
rect 30290 -750 30300 -725
rect 30255 -770 30300 -750
rect 30315 -585 30360 -575
rect 30315 -610 30325 -585
rect 30350 -610 30360 -585
rect 30315 -630 30360 -610
rect 30315 -655 30325 -630
rect 30350 -655 30360 -630
rect 30315 -675 30360 -655
rect 30315 -700 30325 -675
rect 30350 -700 30360 -675
rect 30315 -725 30360 -700
rect 30315 -750 30325 -725
rect 30350 -750 30360 -725
rect 30315 -770 30360 -750
rect 30375 -585 30420 -575
rect 30375 -610 30385 -585
rect 30410 -610 30420 -585
rect 30375 -630 30420 -610
rect 30375 -655 30385 -630
rect 30410 -655 30420 -630
rect 30375 -675 30420 -655
rect 30375 -700 30385 -675
rect 30410 -700 30420 -675
rect 30375 -725 30420 -700
rect 30375 -750 30385 -725
rect 30410 -750 30420 -725
rect 30375 -770 30420 -750
rect 30435 -585 30480 -575
rect 30435 -610 30445 -585
rect 30470 -610 30480 -585
rect 30435 -630 30480 -610
rect 30435 -655 30445 -630
rect 30470 -655 30480 -630
rect 30435 -675 30480 -655
rect 30435 -700 30445 -675
rect 30470 -700 30480 -675
rect 30435 -725 30480 -700
rect 30435 -750 30445 -725
rect 30470 -750 30480 -725
rect 30435 -770 30480 -750
rect 30495 -585 30540 -575
rect 30495 -610 30505 -585
rect 30530 -610 30540 -585
rect 30495 -630 30540 -610
rect 30495 -655 30505 -630
rect 30530 -655 30540 -630
rect 30495 -675 30540 -655
rect 30495 -700 30505 -675
rect 30530 -700 30540 -675
rect 30495 -725 30540 -700
rect 30495 -750 30505 -725
rect 30530 -750 30540 -725
rect 30495 -770 30540 -750
rect 30555 -585 30600 -575
rect 30555 -610 30565 -585
rect 30590 -610 30600 -585
rect 30555 -630 30600 -610
rect 30555 -655 30565 -630
rect 30590 -655 30600 -630
rect 30555 -675 30600 -655
rect 30555 -700 30565 -675
rect 30590 -700 30600 -675
rect 30555 -725 30600 -700
rect 30555 -750 30565 -725
rect 30590 -750 30600 -725
rect 30555 -770 30600 -750
rect 30615 -585 30660 -575
rect 30615 -610 30625 -585
rect 30650 -610 30660 -585
rect 30615 -630 30660 -610
rect 30615 -655 30625 -630
rect 30650 -655 30660 -630
rect 30615 -675 30660 -655
rect 30615 -700 30625 -675
rect 30650 -700 30660 -675
rect 30615 -725 30660 -700
rect 30615 -750 30625 -725
rect 30650 -750 30660 -725
rect 30615 -770 30660 -750
rect 30675 -585 30715 -575
rect 30675 -610 30685 -585
rect 30710 -610 30715 -585
rect 30675 -630 30715 -610
rect 30675 -655 30685 -630
rect 30710 -655 30715 -630
rect 30675 -675 30715 -655
rect 30675 -700 30685 -675
rect 30710 -700 30715 -675
rect 30675 -725 30715 -700
rect 30675 -750 30685 -725
rect 30710 -750 30715 -725
rect 30675 -770 30715 -750
rect 75 -825 115 -810
rect 75 -850 85 -825
rect 110 -850 115 -825
rect 75 -860 115 -850
rect 315 -825 355 -810
rect 315 -850 325 -825
rect 350 -850 355 -825
rect 315 -860 355 -850
rect 555 -825 595 -810
rect 555 -850 565 -825
rect 590 -850 595 -825
rect 555 -860 595 -850
rect 1035 -825 1075 -810
rect 1035 -850 1045 -825
rect 1070 -850 1075 -825
rect 1035 -860 1075 -850
rect 1275 -825 1315 -810
rect 1275 -850 1285 -825
rect 1310 -850 1315 -825
rect 1275 -860 1315 -850
rect 1515 -825 1555 -810
rect 1515 -850 1525 -825
rect 1550 -850 1555 -825
rect 1515 -860 1555 -850
rect 1755 -825 1795 -810
rect 1755 -850 1765 -825
rect 1790 -850 1795 -825
rect 1755 -860 1795 -850
rect 1995 -825 2035 -810
rect 1995 -850 2005 -825
rect 2030 -850 2035 -825
rect 1995 -860 2035 -850
rect 2235 -825 2275 -810
rect 2235 -850 2245 -825
rect 2270 -850 2275 -825
rect 2235 -860 2275 -850
rect 2475 -825 2515 -810
rect 2475 -850 2485 -825
rect 2510 -850 2515 -825
rect 2475 -860 2515 -850
rect 2715 -825 2755 -810
rect 2715 -850 2725 -825
rect 2750 -850 2755 -825
rect 2715 -860 2755 -850
rect 3195 -825 3235 -810
rect 3195 -850 3205 -825
rect 3230 -850 3235 -825
rect 3195 -860 3235 -850
rect 3435 -825 3475 -810
rect 3435 -850 3445 -825
rect 3470 -850 3475 -825
rect 3435 -860 3475 -850
rect 3675 -825 3715 -810
rect 3675 -850 3685 -825
rect 3710 -850 3715 -825
rect 3675 -860 3715 -850
rect 3915 -825 3955 -810
rect 3915 -850 3925 -825
rect 3950 -850 3955 -825
rect 3915 -860 3955 -850
rect 4155 -825 4195 -810
rect 4155 -850 4165 -825
rect 4190 -850 4195 -825
rect 4155 -860 4195 -850
rect 4395 -825 4435 -810
rect 4395 -850 4405 -825
rect 4430 -850 4435 -825
rect 4395 -860 4435 -850
rect 4635 -825 4675 -810
rect 4635 -850 4645 -825
rect 4670 -850 4675 -825
rect 4635 -860 4675 -850
rect 4875 -825 4915 -810
rect 4875 -850 4885 -825
rect 4910 -850 4915 -825
rect 4875 -860 4915 -850
rect 5355 -825 5395 -810
rect 5355 -850 5365 -825
rect 5390 -850 5395 -825
rect 5355 -860 5395 -850
rect 5595 -825 5635 -810
rect 5595 -850 5605 -825
rect 5630 -850 5635 -825
rect 5595 -860 5635 -850
rect 5835 -825 5875 -810
rect 5835 -850 5845 -825
rect 5870 -850 5875 -825
rect 5835 -860 5875 -850
rect 6075 -825 6115 -810
rect 6075 -850 6085 -825
rect 6110 -850 6115 -825
rect 6075 -860 6115 -850
rect 6315 -825 6355 -810
rect 6315 -850 6325 -825
rect 6350 -850 6355 -825
rect 6315 -860 6355 -850
rect 6555 -825 6595 -810
rect 6555 -850 6565 -825
rect 6590 -850 6595 -825
rect 6555 -860 6595 -850
rect 6795 -825 6835 -810
rect 6795 -850 6805 -825
rect 6830 -850 6835 -825
rect 6795 -860 6835 -850
rect 7035 -825 7075 -810
rect 7035 -850 7045 -825
rect 7070 -850 7075 -825
rect 7035 -860 7075 -850
rect 7515 -825 7555 -810
rect 7515 -850 7525 -825
rect 7550 -850 7555 -825
rect 7515 -860 7555 -850
rect 7755 -825 7795 -810
rect 7755 -850 7765 -825
rect 7790 -850 7795 -825
rect 7755 -860 7795 -850
rect 7995 -825 8035 -810
rect 7995 -850 8005 -825
rect 8030 -850 8035 -825
rect 7995 -860 8035 -850
rect 8235 -825 8275 -810
rect 8235 -850 8245 -825
rect 8270 -850 8275 -825
rect 8235 -860 8275 -850
rect 8475 -825 8515 -810
rect 8475 -850 8485 -825
rect 8510 -850 8515 -825
rect 8475 -860 8515 -850
rect 8715 -825 8755 -810
rect 8715 -850 8725 -825
rect 8750 -850 8755 -825
rect 8715 -860 8755 -850
rect 8955 -825 8995 -810
rect 8955 -850 8965 -825
rect 8990 -850 8995 -825
rect 8955 -860 8995 -850
rect 9195 -825 9235 -810
rect 9195 -850 9205 -825
rect 9230 -850 9235 -825
rect 9195 -860 9235 -850
rect 9675 -825 9715 -810
rect 9675 -850 9685 -825
rect 9710 -850 9715 -825
rect 9675 -860 9715 -850
rect 9915 -825 9955 -810
rect 9915 -850 9925 -825
rect 9950 -850 9955 -825
rect 9915 -860 9955 -850
rect 10155 -825 10195 -810
rect 10155 -850 10165 -825
rect 10190 -850 10195 -825
rect 10155 -860 10195 -850
rect 10395 -825 10435 -810
rect 10395 -850 10405 -825
rect 10430 -850 10435 -825
rect 10395 -860 10435 -850
rect 10635 -825 10675 -810
rect 10635 -850 10645 -825
rect 10670 -850 10675 -825
rect 10635 -860 10675 -850
rect 10875 -825 10915 -810
rect 10875 -850 10885 -825
rect 10910 -850 10915 -825
rect 10875 -860 10915 -850
rect 11115 -825 11155 -810
rect 11115 -850 11125 -825
rect 11150 -850 11155 -825
rect 11115 -860 11155 -850
rect 11355 -825 11395 -810
rect 11355 -850 11365 -825
rect 11390 -850 11395 -825
rect 11355 -860 11395 -850
rect 11835 -825 11875 -810
rect 11835 -850 11845 -825
rect 11870 -850 11875 -825
rect 11835 -860 11875 -850
rect 12075 -825 12115 -810
rect 12075 -850 12085 -825
rect 12110 -850 12115 -825
rect 12075 -860 12115 -850
rect 12315 -825 12355 -810
rect 12315 -850 12325 -825
rect 12350 -850 12355 -825
rect 12315 -860 12355 -850
rect 12555 -825 12595 -810
rect 12555 -850 12565 -825
rect 12590 -850 12595 -825
rect 12555 -860 12595 -850
rect 12795 -825 12835 -810
rect 12795 -850 12805 -825
rect 12830 -850 12835 -825
rect 12795 -860 12835 -850
rect 13035 -825 13075 -810
rect 13035 -850 13045 -825
rect 13070 -850 13075 -825
rect 13035 -860 13075 -850
rect 13275 -825 13315 -810
rect 13275 -850 13285 -825
rect 13310 -850 13315 -825
rect 13275 -860 13315 -850
rect 13515 -825 13555 -810
rect 13515 -850 13525 -825
rect 13550 -850 13555 -825
rect 13515 -860 13555 -850
rect 13995 -825 14035 -810
rect 13995 -850 14005 -825
rect 14030 -850 14035 -825
rect 13995 -860 14035 -850
rect 14235 -825 14275 -810
rect 14235 -850 14245 -825
rect 14270 -850 14275 -825
rect 14235 -860 14275 -850
rect 14475 -825 14515 -810
rect 14475 -850 14485 -825
rect 14510 -850 14515 -825
rect 14475 -860 14515 -850
rect 14715 -825 14755 -810
rect 14715 -850 14725 -825
rect 14750 -850 14755 -825
rect 14715 -860 14755 -850
rect 14955 -825 14995 -810
rect 14955 -850 14965 -825
rect 14990 -850 14995 -825
rect 14955 -860 14995 -850
rect 15195 -825 15235 -810
rect 15195 -850 15205 -825
rect 15230 -850 15235 -825
rect 15195 -860 15235 -850
rect 15435 -825 15475 -810
rect 15435 -850 15445 -825
rect 15470 -850 15475 -825
rect 15435 -860 15475 -850
rect 15675 -825 15715 -810
rect 15675 -850 15685 -825
rect 15710 -850 15715 -825
rect 15675 -860 15715 -850
rect 16155 -825 16195 -810
rect 16155 -850 16165 -825
rect 16190 -850 16195 -825
rect 16155 -860 16195 -850
rect 16395 -825 16435 -810
rect 16395 -850 16405 -825
rect 16430 -850 16435 -825
rect 16395 -860 16435 -850
rect 16635 -825 16675 -810
rect 16635 -850 16645 -825
rect 16670 -850 16675 -825
rect 16635 -860 16675 -850
rect 16875 -825 16915 -810
rect 16875 -850 16885 -825
rect 16910 -850 16915 -825
rect 16875 -860 16915 -850
rect 17115 -825 17155 -810
rect 17115 -850 17125 -825
rect 17150 -850 17155 -825
rect 17115 -860 17155 -850
rect 17355 -825 17395 -810
rect 17355 -850 17365 -825
rect 17390 -850 17395 -825
rect 17355 -860 17395 -850
rect 17595 -825 17635 -810
rect 17595 -850 17605 -825
rect 17630 -850 17635 -825
rect 17595 -860 17635 -850
rect 17835 -825 17875 -810
rect 17835 -850 17845 -825
rect 17870 -850 17875 -825
rect 17835 -860 17875 -850
rect 18315 -825 18355 -810
rect 18315 -850 18325 -825
rect 18350 -850 18355 -825
rect 18315 -860 18355 -850
rect 18555 -825 18595 -810
rect 18555 -850 18565 -825
rect 18590 -850 18595 -825
rect 18555 -860 18595 -850
rect 18795 -825 18835 -810
rect 18795 -850 18805 -825
rect 18830 -850 18835 -825
rect 18795 -860 18835 -850
rect 19035 -825 19075 -810
rect 19035 -850 19045 -825
rect 19070 -850 19075 -825
rect 19035 -860 19075 -850
rect 19275 -825 19315 -810
rect 19275 -850 19285 -825
rect 19310 -850 19315 -825
rect 19275 -860 19315 -850
rect 19515 -825 19555 -810
rect 19515 -850 19525 -825
rect 19550 -850 19555 -825
rect 19515 -860 19555 -850
rect 19755 -825 19795 -810
rect 19755 -850 19765 -825
rect 19790 -850 19795 -825
rect 19755 -860 19795 -850
rect 19995 -825 20035 -810
rect 19995 -850 20005 -825
rect 20030 -850 20035 -825
rect 19995 -860 20035 -850
rect 20475 -825 20515 -810
rect 20475 -850 20485 -825
rect 20510 -850 20515 -825
rect 20475 -860 20515 -850
rect 20715 -825 20755 -810
rect 20715 -850 20725 -825
rect 20750 -850 20755 -825
rect 20715 -860 20755 -850
rect 20955 -825 20995 -810
rect 20955 -850 20965 -825
rect 20990 -850 20995 -825
rect 20955 -860 20995 -850
rect 21195 -825 21235 -810
rect 21195 -850 21205 -825
rect 21230 -850 21235 -825
rect 21195 -860 21235 -850
rect 21435 -825 21475 -810
rect 21435 -850 21445 -825
rect 21470 -850 21475 -825
rect 21435 -860 21475 -850
rect 21675 -825 21715 -810
rect 21675 -850 21685 -825
rect 21710 -850 21715 -825
rect 21675 -860 21715 -850
rect 21915 -825 21955 -810
rect 21915 -850 21925 -825
rect 21950 -850 21955 -825
rect 21915 -860 21955 -850
rect 22155 -825 22195 -810
rect 22155 -850 22165 -825
rect 22190 -850 22195 -825
rect 22155 -860 22195 -850
rect 22635 -825 22675 -810
rect 22635 -850 22645 -825
rect 22670 -850 22675 -825
rect 22635 -860 22675 -850
rect 22875 -825 22915 -810
rect 22875 -850 22885 -825
rect 22910 -850 22915 -825
rect 22875 -860 22915 -850
rect 23115 -825 23155 -810
rect 23115 -850 23125 -825
rect 23150 -850 23155 -825
rect 23115 -860 23155 -850
rect 23355 -825 23395 -810
rect 23355 -850 23365 -825
rect 23390 -850 23395 -825
rect 23355 -860 23395 -850
rect 23595 -825 23635 -810
rect 23595 -850 23605 -825
rect 23630 -850 23635 -825
rect 23595 -860 23635 -850
rect 23835 -825 23875 -810
rect 23835 -850 23845 -825
rect 23870 -850 23875 -825
rect 23835 -860 23875 -850
rect 24075 -825 24115 -810
rect 24075 -850 24085 -825
rect 24110 -850 24115 -825
rect 24075 -860 24115 -850
rect 24555 -825 24595 -810
rect 24555 -850 24565 -825
rect 24590 -850 24595 -825
rect 24555 -860 24595 -850
rect 24795 -825 24835 -810
rect 24795 -850 24805 -825
rect 24830 -850 24835 -825
rect 24795 -860 24835 -850
rect 25035 -825 25075 -810
rect 25035 -850 25045 -825
rect 25070 -850 25075 -825
rect 25035 -860 25075 -850
rect 25275 -825 25315 -810
rect 25275 -850 25285 -825
rect 25310 -850 25315 -825
rect 25275 -860 25315 -850
rect 25515 -825 25555 -810
rect 25515 -850 25525 -825
rect 25550 -850 25555 -825
rect 25515 -860 25555 -850
rect 25755 -825 25795 -810
rect 25755 -850 25765 -825
rect 25790 -850 25795 -825
rect 25755 -860 25795 -850
rect 25995 -825 26035 -810
rect 25995 -850 26005 -825
rect 26030 -850 26035 -825
rect 25995 -860 26035 -850
rect 26475 -825 26515 -810
rect 26475 -850 26485 -825
rect 26510 -850 26515 -825
rect 26475 -860 26515 -850
rect 26715 -825 26755 -810
rect 26715 -850 26725 -825
rect 26750 -850 26755 -825
rect 26715 -860 26755 -850
rect 26955 -825 26995 -810
rect 26955 -850 26965 -825
rect 26990 -850 26995 -825
rect 26955 -860 26995 -850
rect 27195 -825 27235 -810
rect 27195 -850 27205 -825
rect 27230 -850 27235 -825
rect 27195 -860 27235 -850
rect 27435 -825 27475 -810
rect 27435 -850 27445 -825
rect 27470 -850 27475 -825
rect 27435 -860 27475 -850
rect 27675 -825 27715 -810
rect 27675 -850 27685 -825
rect 27710 -850 27715 -825
rect 27675 -860 27715 -850
rect 27915 -825 27955 -810
rect 27915 -850 27925 -825
rect 27950 -850 27955 -825
rect 27915 -860 27955 -850
rect 28395 -825 28435 -810
rect 28395 -850 28405 -825
rect 28430 -850 28435 -825
rect 28395 -860 28435 -850
rect 28635 -825 28675 -810
rect 28635 -850 28645 -825
rect 28670 -850 28675 -825
rect 28635 -860 28675 -850
rect 28875 -825 28915 -810
rect 28875 -850 28885 -825
rect 28910 -850 28915 -825
rect 28875 -860 28915 -850
rect 29115 -825 29155 -810
rect 29115 -850 29125 -825
rect 29150 -850 29155 -825
rect 29115 -860 29155 -850
rect 29355 -825 29395 -810
rect 29355 -850 29365 -825
rect 29390 -850 29395 -825
rect 29355 -860 29395 -850
rect 29595 -825 29635 -810
rect 29595 -850 29605 -825
rect 29630 -850 29635 -825
rect 29595 -860 29635 -850
rect 30075 -825 30115 -810
rect 30075 -850 30085 -825
rect 30110 -850 30115 -825
rect 30075 -860 30115 -850
rect 30315 -825 30355 -810
rect 30315 -850 30325 -825
rect 30350 -850 30355 -825
rect 30315 -860 30355 -850
rect 30555 -825 30595 -810
rect 30555 -850 30565 -825
rect 30590 -850 30595 -825
rect 30555 -860 30595 -850
<< ndiffc >>
rect 196 -110 221 -85
rect 256 -110 281 -85
rect 321 -110 346 -85
rect 381 -110 406 -85
rect 441 -110 466 -85
rect 501 -110 526 -85
rect 561 -110 586 -85
rect 626 -110 651 -85
rect 686 -110 711 -85
rect 746 -110 771 -85
rect 806 -110 831 -85
rect 871 -110 896 -85
rect 931 -110 956 -85
rect 991 -110 1016 -85
rect 1051 -110 1076 -85
rect 1111 -110 1136 -85
rect 1171 -110 1196 -85
rect 1231 -110 1256 -85
rect 1291 -110 1316 -85
rect 1356 -110 1381 -85
rect 1416 -110 1441 -85
rect 1476 -110 1501 -85
rect 1536 -110 1561 -85
rect 1596 -110 1621 -85
rect 1661 -110 1686 -85
rect 1721 -110 1746 -85
rect 1781 -110 1806 -85
rect 1841 -110 1866 -85
rect 1906 -110 1931 -85
rect 1966 -110 1991 -85
rect 2026 -110 2051 -85
rect 2086 -110 2111 -85
rect 2146 -110 2171 -85
rect 2206 -110 2231 -85
rect 2266 -110 2291 -85
rect 2326 -110 2351 -85
rect 2391 -110 2416 -85
rect 2451 -110 2476 -85
rect 2511 -110 2536 -85
rect 2571 -110 2596 -85
rect 2631 -110 2656 -85
rect 2691 -110 2716 -85
rect 2751 -110 2776 -85
rect 2811 -110 2836 -85
rect 2876 -110 2901 -85
rect 2936 -110 2961 -85
rect 2996 -110 3021 -85
rect 3056 -110 3081 -85
rect 3116 -110 3141 -85
rect 3176 -110 3201 -85
rect 3236 -110 3261 -85
rect 3296 -110 3321 -85
rect 3361 -110 3386 -85
rect 3421 -110 3446 -85
rect 3481 -110 3506 -85
rect 3541 -110 3566 -85
rect 3601 -110 3626 -85
rect 3661 -110 3686 -85
rect 3721 -110 3746 -85
rect 3781 -110 3806 -85
rect 3846 -110 3871 -85
rect 3906 -110 3931 -85
rect 3966 -110 3991 -85
rect 4026 -110 4051 -85
rect 4086 -110 4111 -85
rect 4146 -110 4171 -85
rect 4206 -110 4231 -85
rect 4266 -110 4291 -85
rect 4331 -110 4356 -85
rect 4391 -110 4416 -85
rect 4451 -110 4476 -85
rect 4511 -110 4536 -85
rect 4571 -110 4596 -85
rect 4631 -110 4656 -85
rect 4691 -110 4716 -85
rect 4751 -110 4776 -85
rect 4816 -110 4841 -85
rect 4876 -110 4901 -85
rect 4936 -110 4961 -85
rect 4996 -110 5021 -85
rect 5056 -110 5081 -85
rect 5116 -110 5141 -85
rect 5176 -110 5201 -85
rect 5236 -110 5261 -85
rect 5301 -110 5326 -85
rect 5361 -110 5386 -85
rect 5421 -110 5446 -85
rect 5481 -110 5506 -85
rect 5541 -110 5566 -85
rect 5606 -110 5631 -85
rect 5666 -110 5691 -85
rect 5726 -110 5751 -85
rect 5786 -110 5811 -85
rect 5851 -110 5876 -85
rect 5911 -110 5936 -85
rect 5971 -110 5996 -85
rect 6031 -110 6056 -85
rect 6091 -110 6116 -85
rect 6151 -110 6176 -85
rect 6211 -110 6236 -85
rect 6271 -110 6296 -85
rect 6336 -110 6361 -85
rect 6396 -110 6421 -85
rect 6456 -110 6481 -85
rect 6516 -110 6541 -85
rect 6576 -110 6601 -85
rect 6636 -110 6661 -85
rect 6696 -110 6721 -85
rect 6756 -110 6781 -85
rect 6821 -110 6846 -85
rect 6881 -110 6906 -85
rect 6941 -110 6966 -85
rect 7001 -110 7026 -85
rect 7061 -110 7086 -85
rect 7121 -110 7146 -85
rect 7181 -110 7206 -85
rect 7241 -110 7266 -85
rect 7301 -110 7326 -85
rect 7361 -110 7386 -85
rect 7421 -110 7446 -85
rect 7481 -110 7506 -85
rect 7541 -110 7566 -85
rect 7601 -110 7626 -85
rect 7661 -110 7686 -85
rect 7721 -110 7746 -85
rect 7786 -110 7811 -85
rect 7846 -110 7871 -85
rect 7906 -110 7931 -85
rect 7966 -110 7991 -85
rect 8026 -110 8051 -85
rect 8086 -110 8111 -85
rect 8146 -110 8171 -85
rect 8206 -110 8231 -85
rect 8271 -110 8296 -85
rect 8331 -110 8356 -85
rect 8391 -110 8416 -85
rect 8451 -110 8476 -85
rect 8511 -110 8536 -85
rect 8571 -110 8596 -85
rect 8631 -110 8656 -85
rect 8691 -110 8716 -85
rect 8756 -110 8781 -85
rect 8816 -110 8841 -85
rect 8876 -110 8901 -85
rect 8936 -110 8961 -85
rect 8996 -110 9021 -85
rect 9056 -110 9081 -85
rect 9116 -110 9141 -85
rect 9176 -110 9201 -85
rect 9241 -110 9266 -85
rect 9301 -110 9326 -85
rect 9361 -110 9386 -85
rect 9421 -110 9446 -85
rect 9486 -110 9511 -85
rect 9546 -110 9571 -85
rect 9606 -110 9631 -85
rect 9666 -110 9691 -85
rect 9731 -110 9756 -85
rect 9791 -110 9816 -85
rect 9851 -110 9876 -85
rect 9911 -110 9936 -85
rect 9971 -110 9996 -85
rect 10031 -110 10056 -85
rect 10091 -110 10116 -85
rect 10151 -110 10176 -85
rect 10216 -110 10241 -85
rect 10276 -110 10301 -85
rect 10336 -110 10361 -85
rect 10396 -110 10421 -85
rect 10456 -110 10481 -85
rect 10516 -110 10541 -85
rect 10576 -110 10601 -85
rect 10636 -110 10661 -85
rect 10701 -110 10726 -85
rect 10761 -110 10786 -85
rect 10821 -110 10846 -85
rect 10881 -110 10906 -85
rect 10941 -110 10966 -85
rect 11001 -110 11026 -85
rect 11061 -110 11086 -85
rect 11121 -110 11146 -85
rect 11186 -110 11211 -85
rect 11246 -110 11271 -85
rect 11306 -110 11331 -85
rect 11366 -110 11391 -85
rect 11426 -110 11451 -85
rect 11486 -110 11511 -85
rect 11546 -110 11571 -85
rect 11606 -110 11631 -85
rect 11671 -110 11696 -85
rect 11731 -110 11756 -85
rect 11791 -110 11816 -85
rect 11851 -110 11876 -85
rect 11911 -110 11936 -85
rect 11971 -110 11996 -85
rect 12031 -110 12056 -85
rect 12091 -110 12116 -85
rect 12156 -110 12181 -85
rect 12216 -110 12241 -85
rect 12276 -110 12301 -85
rect 12336 -110 12361 -85
rect 12396 -110 12421 -85
rect 12456 -110 12481 -85
rect 12516 -110 12541 -85
rect 12576 -110 12601 -85
rect 12641 -110 12666 -85
rect 12701 -110 12726 -85
rect 12761 -110 12786 -85
rect 12821 -110 12846 -85
rect 12881 -110 12906 -85
rect 12941 -110 12966 -85
rect 13001 -110 13026 -85
rect 13061 -110 13086 -85
rect 13126 -110 13151 -85
rect 13186 -110 13211 -85
rect 13246 -110 13271 -85
rect 13306 -110 13331 -85
rect 13366 -110 13391 -85
rect 13426 -110 13451 -85
rect 13486 -110 13511 -85
rect 13546 -110 13571 -85
rect 13611 -110 13636 -85
rect 13671 -110 13696 -85
rect 13731 -110 13756 -85
rect 13791 -110 13816 -85
rect 13851 -110 13876 -85
rect 13911 -110 13936 -85
rect 13971 -110 13996 -85
rect 14031 -110 14056 -85
rect 14096 -110 14121 -85
rect 14156 -110 14181 -85
rect 14216 -110 14241 -85
rect 14276 -110 14301 -85
rect 14336 -110 14361 -85
rect 14396 -110 14421 -85
rect 14456 -110 14481 -85
rect 14516 -110 14541 -85
rect 14581 -110 14606 -85
rect 14641 -110 14666 -85
rect 14701 -110 14726 -85
rect 14761 -110 14786 -85
rect 14821 -110 14846 -85
rect 14881 -110 14906 -85
rect 14941 -110 14966 -85
rect 15001 -110 15026 -85
rect 15066 -110 15091 -85
rect 15126 -110 15151 -85
rect 15186 -110 15211 -85
rect 15246 -110 15271 -85
rect 15306 -110 15331 -85
rect 15366 -110 15391 -85
rect 15426 -110 15451 -85
rect 15486 -110 15511 -85
rect 15551 -110 15576 -85
rect 15611 -110 15636 -85
rect 15671 -110 15696 -85
rect 15731 -110 15756 -85
rect 15791 -110 15816 -85
rect 15851 -110 15876 -85
rect 15911 -110 15936 -85
rect 15971 -110 15996 -85
rect 16036 -110 16061 -85
rect 16096 -110 16121 -85
rect 16156 -110 16181 -85
rect 16216 -110 16241 -85
rect 16276 -110 16301 -85
rect 16336 -110 16361 -85
rect 16396 -110 16421 -85
rect 16456 -110 16481 -85
rect 16521 -110 16546 -85
rect 16581 -110 16606 -85
rect 16641 -110 16666 -85
rect 16701 -110 16726 -85
rect 16761 -110 16786 -85
rect 16821 -110 16846 -85
rect 16881 -110 16906 -85
rect 16941 -110 16966 -85
rect 17006 -110 17031 -85
rect 17066 -110 17091 -85
rect 17126 -110 17151 -85
rect 17186 -110 17211 -85
rect 17246 -110 17271 -85
rect 17306 -110 17331 -85
rect 17366 -110 17391 -85
rect 17426 -110 17451 -85
rect 17491 -110 17516 -85
rect 17551 -110 17576 -85
rect 17611 -110 17636 -85
rect 17671 -110 17696 -85
rect 17731 -110 17756 -85
rect 17791 -110 17816 -85
rect 17851 -110 17876 -85
rect 17911 -110 17936 -85
rect 17976 -110 18001 -85
rect 18036 -110 18061 -85
rect 18096 -110 18121 -85
rect 18156 -110 18181 -85
rect 18216 -110 18241 -85
rect 18276 -110 18301 -85
rect 18336 -110 18361 -85
rect 18396 -110 18421 -85
rect 18461 -110 18486 -85
rect 18521 -110 18546 -85
rect 18581 -110 18606 -85
rect 18641 -110 18666 -85
rect 18701 -110 18726 -85
rect 18761 -110 18786 -85
rect 18821 -110 18846 -85
rect 18881 -110 18906 -85
rect 18946 -110 18971 -85
rect 19006 -110 19031 -85
rect 19066 -110 19091 -85
rect 19126 -110 19151 -85
rect 19186 -110 19211 -85
rect 19246 -110 19271 -85
rect 19306 -110 19331 -85
rect 19366 -110 19391 -85
rect 19431 -110 19456 -85
rect 19491 -110 19516 -85
rect 19551 -110 19576 -85
rect 19611 -110 19636 -85
rect 19671 -110 19696 -85
rect 19731 -110 19756 -85
rect 19791 -110 19816 -85
rect 19851 -110 19876 -85
rect 19916 -110 19941 -85
rect 19976 -110 20001 -85
rect 20036 -110 20061 -85
rect 20096 -110 20121 -85
rect 20156 -110 20181 -85
rect 20216 -110 20241 -85
rect 20276 -110 20301 -85
rect 20336 -110 20361 -85
rect 20401 -110 20426 -85
rect 20461 -110 20486 -85
rect 20521 -110 20546 -85
rect 20581 -110 20606 -85
rect 20641 -110 20666 -85
rect 20701 -110 20726 -85
rect 20761 -110 20786 -85
rect 20821 -110 20846 -85
rect 20886 -110 20911 -85
rect 20946 -110 20971 -85
rect 21006 -110 21031 -85
rect 21066 -110 21091 -85
rect 21126 -110 21151 -85
rect -35 -360 -10 -335
rect -35 -405 -10 -380
rect 25 -360 50 -335
rect 25 -405 50 -380
rect 85 -360 110 -335
rect 85 -405 110 -380
rect 145 -360 170 -335
rect 145 -405 170 -380
rect 205 -360 230 -335
rect 205 -405 230 -380
rect 265 -360 290 -335
rect 265 -405 290 -380
rect 325 -360 350 -335
rect 325 -405 350 -380
rect 385 -360 410 -335
rect 385 -405 410 -380
rect 445 -360 470 -335
rect 445 -405 470 -380
rect 505 -360 530 -335
rect 505 -405 530 -380
rect 565 -360 590 -335
rect 565 -405 590 -380
rect 625 -360 650 -335
rect 625 -405 650 -380
rect 685 -360 710 -335
rect 685 -405 710 -380
rect 745 -360 770 -335
rect 745 -405 770 -380
rect 805 -360 830 -335
rect 805 -405 830 -380
rect 865 -360 890 -335
rect 865 -405 890 -380
rect 925 -360 950 -335
rect 925 -405 950 -380
rect 985 -360 1010 -335
rect 985 -405 1010 -380
rect 1045 -360 1070 -335
rect 1045 -405 1070 -380
rect 1105 -360 1130 -335
rect 1105 -405 1130 -380
rect 1165 -360 1190 -335
rect 1165 -405 1190 -380
rect 1225 -360 1250 -335
rect 1225 -405 1250 -380
rect 1285 -360 1310 -335
rect 1285 -405 1310 -380
rect 1345 -360 1370 -335
rect 1345 -405 1370 -380
rect 1405 -360 1430 -335
rect 1405 -405 1430 -380
rect 1465 -360 1490 -335
rect 1465 -405 1490 -380
rect 1525 -360 1550 -335
rect 1525 -405 1550 -380
rect 1585 -360 1610 -335
rect 1585 -405 1610 -380
rect 1645 -360 1670 -335
rect 1645 -405 1670 -380
rect 1705 -360 1730 -335
rect 1705 -405 1730 -380
rect 1765 -360 1790 -335
rect 1765 -405 1790 -380
rect 1825 -360 1850 -335
rect 1825 -405 1850 -380
rect 1885 -360 1910 -335
rect 1885 -405 1910 -380
rect 1945 -360 1970 -335
rect 1945 -405 1970 -380
rect 2005 -360 2030 -335
rect 2005 -405 2030 -380
rect 2065 -360 2090 -335
rect 2065 -405 2090 -380
rect 2125 -360 2150 -335
rect 2125 -405 2150 -380
rect 2185 -360 2210 -335
rect 2185 -405 2210 -380
rect 2245 -360 2270 -335
rect 2245 -405 2270 -380
rect 2305 -360 2330 -335
rect 2305 -405 2330 -380
rect 2365 -360 2390 -335
rect 2365 -405 2390 -380
rect 2425 -360 2450 -335
rect 2425 -405 2450 -380
rect 2485 -360 2510 -335
rect 2485 -405 2510 -380
rect 2545 -360 2570 -335
rect 2545 -405 2570 -380
rect 2605 -360 2630 -335
rect 2605 -405 2630 -380
rect 2665 -360 2690 -335
rect 2665 -405 2690 -380
rect 2725 -360 2750 -335
rect 2725 -405 2750 -380
rect 2785 -360 2810 -335
rect 2785 -405 2810 -380
rect 2845 -360 2870 -335
rect 2845 -405 2870 -380
rect 2905 -360 2930 -335
rect 2905 -405 2930 -380
rect 2965 -360 2990 -335
rect 2965 -405 2990 -380
rect 3025 -360 3050 -335
rect 3025 -405 3050 -380
rect 3085 -360 3110 -335
rect 3085 -405 3110 -380
rect 3145 -360 3170 -335
rect 3145 -405 3170 -380
rect 3205 -360 3230 -335
rect 3205 -405 3230 -380
rect 3265 -360 3290 -335
rect 3265 -405 3290 -380
rect 3325 -360 3350 -335
rect 3325 -405 3350 -380
rect 3385 -360 3410 -335
rect 3385 -405 3410 -380
rect 3445 -360 3470 -335
rect 3445 -405 3470 -380
rect 3505 -360 3530 -335
rect 3505 -405 3530 -380
rect 3565 -360 3590 -335
rect 3565 -405 3590 -380
rect 3625 -360 3650 -335
rect 3625 -405 3650 -380
rect 3685 -360 3710 -335
rect 3685 -405 3710 -380
rect 3745 -360 3770 -335
rect 3745 -405 3770 -380
rect 3805 -360 3830 -335
rect 3805 -405 3830 -380
rect 3865 -360 3890 -335
rect 3865 -405 3890 -380
rect 3925 -360 3950 -335
rect 3925 -405 3950 -380
rect 3985 -360 4010 -335
rect 3985 -405 4010 -380
rect 4045 -360 4070 -335
rect 4045 -405 4070 -380
rect 4105 -360 4130 -335
rect 4105 -405 4130 -380
rect 4165 -360 4190 -335
rect 4165 -405 4190 -380
rect 4225 -360 4250 -335
rect 4225 -405 4250 -380
rect 4285 -360 4310 -335
rect 4285 -405 4310 -380
rect 4345 -360 4370 -335
rect 4345 -405 4370 -380
rect 4405 -360 4430 -335
rect 4405 -405 4430 -380
rect 4465 -360 4490 -335
rect 4465 -405 4490 -380
rect 4525 -360 4550 -335
rect 4525 -405 4550 -380
rect 4585 -360 4610 -335
rect 4585 -405 4610 -380
rect 4645 -360 4670 -335
rect 4645 -405 4670 -380
rect 4705 -360 4730 -335
rect 4705 -405 4730 -380
rect 4765 -360 4790 -335
rect 4765 -405 4790 -380
rect 4825 -360 4850 -335
rect 4825 -405 4850 -380
rect 4885 -360 4910 -335
rect 4885 -405 4910 -380
rect 4945 -360 4970 -335
rect 4945 -405 4970 -380
rect 5005 -360 5030 -335
rect 5005 -405 5030 -380
rect 5065 -360 5090 -335
rect 5065 -405 5090 -380
rect 5125 -360 5150 -335
rect 5125 -405 5150 -380
rect 5185 -360 5210 -335
rect 5185 -405 5210 -380
rect 5245 -360 5270 -335
rect 5245 -405 5270 -380
rect 5305 -360 5330 -335
rect 5305 -405 5330 -380
rect 5365 -360 5390 -335
rect 5365 -405 5390 -380
rect 5425 -360 5450 -335
rect 5425 -405 5450 -380
rect 5485 -360 5510 -335
rect 5485 -405 5510 -380
rect 5545 -360 5570 -335
rect 5545 -405 5570 -380
rect 5605 -360 5630 -335
rect 5605 -405 5630 -380
rect 5665 -360 5690 -335
rect 5665 -405 5690 -380
rect 5725 -360 5750 -335
rect 5725 -405 5750 -380
rect 5785 -360 5810 -335
rect 5785 -405 5810 -380
rect 5845 -360 5870 -335
rect 5845 -405 5870 -380
rect 5905 -360 5930 -335
rect 5905 -405 5930 -380
rect 5965 -360 5990 -335
rect 5965 -405 5990 -380
rect 6025 -360 6050 -335
rect 6025 -405 6050 -380
rect 6085 -360 6110 -335
rect 6085 -405 6110 -380
rect 6145 -360 6170 -335
rect 6145 -405 6170 -380
rect 6205 -360 6230 -335
rect 6205 -405 6230 -380
rect 6265 -360 6290 -335
rect 6265 -405 6290 -380
rect 6325 -360 6350 -335
rect 6325 -405 6350 -380
rect 6385 -360 6410 -335
rect 6385 -405 6410 -380
rect 6445 -360 6470 -335
rect 6445 -405 6470 -380
rect 6505 -360 6530 -335
rect 6505 -405 6530 -380
rect 6565 -360 6590 -335
rect 6565 -405 6590 -380
rect 6625 -360 6650 -335
rect 6625 -405 6650 -380
rect 6685 -360 6710 -335
rect 6685 -405 6710 -380
rect 6745 -360 6770 -335
rect 6745 -405 6770 -380
rect 6805 -360 6830 -335
rect 6805 -405 6830 -380
rect 6865 -360 6890 -335
rect 6865 -405 6890 -380
rect 6925 -360 6950 -335
rect 6925 -405 6950 -380
rect 6985 -360 7010 -335
rect 6985 -405 7010 -380
rect 7045 -360 7070 -335
rect 7045 -405 7070 -380
rect 7105 -360 7130 -335
rect 7105 -405 7130 -380
rect 7165 -360 7190 -335
rect 7165 -405 7190 -380
rect 7225 -360 7250 -335
rect 7225 -405 7250 -380
rect 7285 -360 7310 -335
rect 7285 -405 7310 -380
rect 7345 -360 7370 -335
rect 7345 -405 7370 -380
rect 7405 -360 7430 -335
rect 7405 -405 7430 -380
rect 7465 -360 7490 -335
rect 7465 -405 7490 -380
rect 7525 -360 7550 -335
rect 7525 -405 7550 -380
rect 7585 -360 7610 -335
rect 7585 -405 7610 -380
rect 7645 -360 7670 -335
rect 7645 -405 7670 -380
rect 7705 -360 7730 -335
rect 7705 -405 7730 -380
rect 7765 -360 7790 -335
rect 7765 -405 7790 -380
rect 7825 -360 7850 -335
rect 7825 -405 7850 -380
rect 7885 -360 7910 -335
rect 7885 -405 7910 -380
rect 7945 -360 7970 -335
rect 7945 -405 7970 -380
rect 8005 -360 8030 -335
rect 8005 -405 8030 -380
rect 8065 -360 8090 -335
rect 8065 -405 8090 -380
rect 8125 -360 8150 -335
rect 8125 -405 8150 -380
rect 8185 -360 8210 -335
rect 8185 -405 8210 -380
rect 8245 -360 8270 -335
rect 8245 -405 8270 -380
rect 8305 -360 8330 -335
rect 8305 -405 8330 -380
rect 8365 -360 8390 -335
rect 8365 -405 8390 -380
rect 8425 -360 8450 -335
rect 8425 -405 8450 -380
rect 8485 -360 8510 -335
rect 8485 -405 8510 -380
rect 8545 -360 8570 -335
rect 8545 -405 8570 -380
rect 8605 -360 8630 -335
rect 8605 -405 8630 -380
rect 8665 -360 8690 -335
rect 8665 -405 8690 -380
rect 8725 -360 8750 -335
rect 8725 -405 8750 -380
rect 8785 -360 8810 -335
rect 8785 -405 8810 -380
rect 8845 -360 8870 -335
rect 8845 -405 8870 -380
rect 8905 -360 8930 -335
rect 8905 -405 8930 -380
rect 8965 -360 8990 -335
rect 8965 -405 8990 -380
rect 9025 -360 9050 -335
rect 9025 -405 9050 -380
rect 9085 -360 9110 -335
rect 9085 -405 9110 -380
rect 9145 -360 9170 -335
rect 9145 -405 9170 -380
rect 9205 -360 9230 -335
rect 9205 -405 9230 -380
rect 9265 -360 9290 -335
rect 9265 -405 9290 -380
rect 9325 -360 9350 -335
rect 9325 -405 9350 -380
rect 9385 -360 9410 -335
rect 9385 -405 9410 -380
rect 9445 -360 9470 -335
rect 9445 -405 9470 -380
rect 9505 -360 9530 -335
rect 9505 -405 9530 -380
rect 9565 -360 9590 -335
rect 9565 -405 9590 -380
rect 9625 -360 9650 -335
rect 9625 -405 9650 -380
rect 9685 -360 9710 -335
rect 9685 -405 9710 -380
rect 9745 -360 9770 -335
rect 9745 -405 9770 -380
rect 9805 -360 9830 -335
rect 9805 -405 9830 -380
rect 9865 -360 9890 -335
rect 9865 -405 9890 -380
rect 9925 -360 9950 -335
rect 9925 -405 9950 -380
rect 9985 -360 10010 -335
rect 9985 -405 10010 -380
rect 10045 -360 10070 -335
rect 10045 -405 10070 -380
rect 10105 -360 10130 -335
rect 10105 -405 10130 -380
rect 10165 -360 10190 -335
rect 10165 -405 10190 -380
rect 10225 -360 10250 -335
rect 10225 -405 10250 -380
rect 10285 -360 10310 -335
rect 10285 -405 10310 -380
rect 10345 -360 10370 -335
rect 10345 -405 10370 -380
rect 10405 -360 10430 -335
rect 10405 -405 10430 -380
rect 10465 -360 10490 -335
rect 10465 -405 10490 -380
rect 10525 -360 10550 -335
rect 10525 -405 10550 -380
rect 10585 -360 10610 -335
rect 10585 -405 10610 -380
rect 10645 -360 10670 -335
rect 10645 -405 10670 -380
rect 10705 -360 10730 -335
rect 10705 -405 10730 -380
rect 10765 -360 10790 -335
rect 10765 -405 10790 -380
rect 10825 -360 10850 -335
rect 10825 -405 10850 -380
rect 10885 -360 10910 -335
rect 10885 -405 10910 -380
rect 10945 -360 10970 -335
rect 10945 -405 10970 -380
rect 11005 -360 11030 -335
rect 11005 -405 11030 -380
rect 11065 -360 11090 -335
rect 11065 -405 11090 -380
rect 11125 -360 11150 -335
rect 11125 -405 11150 -380
rect 11185 -360 11210 -335
rect 11185 -405 11210 -380
rect 11245 -360 11270 -335
rect 11245 -405 11270 -380
rect 11305 -360 11330 -335
rect 11305 -405 11330 -380
rect 11365 -360 11390 -335
rect 11365 -405 11390 -380
rect 11425 -360 11450 -335
rect 11425 -405 11450 -380
rect 11485 -360 11510 -335
rect 11485 -405 11510 -380
rect 11545 -360 11570 -335
rect 11545 -405 11570 -380
rect 11605 -360 11630 -335
rect 11605 -405 11630 -380
rect 11665 -360 11690 -335
rect 11665 -405 11690 -380
rect 11725 -360 11750 -335
rect 11725 -405 11750 -380
rect 11785 -360 11810 -335
rect 11785 -405 11810 -380
rect 11845 -360 11870 -335
rect 11845 -405 11870 -380
rect 11905 -360 11930 -335
rect 11905 -405 11930 -380
rect 11965 -360 11990 -335
rect 11965 -405 11990 -380
rect 12025 -360 12050 -335
rect 12025 -405 12050 -380
rect 12085 -360 12110 -335
rect 12085 -405 12110 -380
rect 12145 -360 12170 -335
rect 12145 -405 12170 -380
rect 12205 -360 12230 -335
rect 12205 -405 12230 -380
rect 12265 -360 12290 -335
rect 12265 -405 12290 -380
rect 12325 -360 12350 -335
rect 12325 -405 12350 -380
rect 12385 -360 12410 -335
rect 12385 -405 12410 -380
rect 12445 -360 12470 -335
rect 12445 -405 12470 -380
rect 12505 -360 12530 -335
rect 12505 -405 12530 -380
rect 12565 -360 12590 -335
rect 12565 -405 12590 -380
rect 12625 -360 12650 -335
rect 12625 -405 12650 -380
rect 12685 -360 12710 -335
rect 12685 -405 12710 -380
rect 12745 -360 12770 -335
rect 12745 -405 12770 -380
rect 12805 -360 12830 -335
rect 12805 -405 12830 -380
rect 12865 -360 12890 -335
rect 12865 -405 12890 -380
rect 12925 -360 12950 -335
rect 12925 -405 12950 -380
rect 12985 -360 13010 -335
rect 12985 -405 13010 -380
rect 13045 -360 13070 -335
rect 13045 -405 13070 -380
rect 13105 -360 13130 -335
rect 13105 -405 13130 -380
rect 13165 -360 13190 -335
rect 13165 -405 13190 -380
rect 13225 -360 13250 -335
rect 13225 -405 13250 -380
rect 13285 -360 13310 -335
rect 13285 -405 13310 -380
rect 13345 -360 13370 -335
rect 13345 -405 13370 -380
rect 13405 -360 13430 -335
rect 13405 -405 13430 -380
rect 13465 -360 13490 -335
rect 13465 -405 13490 -380
rect 13525 -360 13550 -335
rect 13525 -405 13550 -380
rect 13585 -360 13610 -335
rect 13585 -405 13610 -380
rect 13645 -360 13670 -335
rect 13645 -405 13670 -380
rect 13705 -360 13730 -335
rect 13705 -405 13730 -380
rect 13765 -360 13790 -335
rect 13765 -405 13790 -380
rect 13825 -360 13850 -335
rect 13825 -405 13850 -380
rect 13885 -360 13910 -335
rect 13885 -405 13910 -380
rect 13945 -360 13970 -335
rect 13945 -405 13970 -380
rect 14005 -360 14030 -335
rect 14005 -405 14030 -380
rect 14065 -360 14090 -335
rect 14065 -405 14090 -380
rect 14125 -360 14150 -335
rect 14125 -405 14150 -380
rect 14185 -360 14210 -335
rect 14185 -405 14210 -380
rect 14245 -360 14270 -335
rect 14245 -405 14270 -380
rect 14305 -360 14330 -335
rect 14305 -405 14330 -380
rect 14365 -360 14390 -335
rect 14365 -405 14390 -380
rect 14425 -360 14450 -335
rect 14425 -405 14450 -380
rect 14485 -360 14510 -335
rect 14485 -405 14510 -380
rect 14545 -360 14570 -335
rect 14545 -405 14570 -380
rect 14605 -360 14630 -335
rect 14605 -405 14630 -380
rect 14665 -360 14690 -335
rect 14665 -405 14690 -380
rect 14725 -360 14750 -335
rect 14725 -405 14750 -380
rect 14785 -360 14810 -335
rect 14785 -405 14810 -380
rect 14845 -360 14870 -335
rect 14845 -405 14870 -380
rect 14905 -360 14930 -335
rect 14905 -405 14930 -380
rect 14965 -360 14990 -335
rect 14965 -405 14990 -380
rect 15025 -360 15050 -335
rect 15025 -405 15050 -380
rect 15085 -360 15110 -335
rect 15085 -405 15110 -380
rect 15145 -360 15170 -335
rect 15145 -405 15170 -380
rect 15205 -360 15230 -335
rect 15205 -405 15230 -380
rect 15265 -360 15290 -335
rect 15265 -405 15290 -380
rect 15325 -360 15350 -335
rect 15325 -405 15350 -380
rect 15385 -360 15410 -335
rect 15385 -405 15410 -380
rect 15445 -360 15470 -335
rect 15445 -405 15470 -380
rect 15505 -360 15530 -335
rect 15505 -405 15530 -380
rect 15565 -360 15590 -335
rect 15565 -405 15590 -380
rect 15625 -360 15650 -335
rect 15625 -405 15650 -380
rect 15685 -360 15710 -335
rect 15685 -405 15710 -380
rect 15745 -360 15770 -335
rect 15745 -405 15770 -380
rect 15805 -360 15830 -335
rect 15805 -405 15830 -380
rect 15865 -360 15890 -335
rect 15865 -405 15890 -380
rect 15925 -360 15950 -335
rect 15925 -405 15950 -380
rect 15985 -360 16010 -335
rect 15985 -405 16010 -380
rect 16045 -360 16070 -335
rect 16045 -405 16070 -380
rect 16105 -360 16130 -335
rect 16105 -405 16130 -380
rect 16165 -360 16190 -335
rect 16165 -405 16190 -380
rect 16225 -360 16250 -335
rect 16225 -405 16250 -380
rect 16285 -360 16310 -335
rect 16285 -405 16310 -380
rect 16345 -360 16370 -335
rect 16345 -405 16370 -380
rect 16405 -360 16430 -335
rect 16405 -405 16430 -380
rect 16465 -360 16490 -335
rect 16465 -405 16490 -380
rect 16525 -360 16550 -335
rect 16525 -405 16550 -380
rect 16585 -360 16610 -335
rect 16585 -405 16610 -380
rect 16645 -360 16670 -335
rect 16645 -405 16670 -380
rect 16705 -360 16730 -335
rect 16705 -405 16730 -380
rect 16765 -360 16790 -335
rect 16765 -405 16790 -380
rect 16825 -360 16850 -335
rect 16825 -405 16850 -380
rect 16885 -360 16910 -335
rect 16885 -405 16910 -380
rect 16945 -360 16970 -335
rect 16945 -405 16970 -380
rect 17005 -360 17030 -335
rect 17005 -405 17030 -380
rect 17065 -360 17090 -335
rect 17065 -405 17090 -380
rect 17125 -360 17150 -335
rect 17125 -405 17150 -380
rect 17185 -360 17210 -335
rect 17185 -405 17210 -380
rect 17245 -360 17270 -335
rect 17245 -405 17270 -380
rect 17305 -360 17330 -335
rect 17305 -405 17330 -380
rect 17365 -360 17390 -335
rect 17365 -405 17390 -380
rect 17425 -360 17450 -335
rect 17425 -405 17450 -380
rect 17485 -360 17510 -335
rect 17485 -405 17510 -380
rect 17545 -360 17570 -335
rect 17545 -405 17570 -380
rect 17605 -360 17630 -335
rect 17605 -405 17630 -380
rect 17665 -360 17690 -335
rect 17665 -405 17690 -380
rect 17725 -360 17750 -335
rect 17725 -405 17750 -380
rect 17785 -360 17810 -335
rect 17785 -405 17810 -380
rect 17845 -360 17870 -335
rect 17845 -405 17870 -380
rect 17905 -360 17930 -335
rect 17905 -405 17930 -380
rect 17965 -360 17990 -335
rect 17965 -405 17990 -380
rect 18025 -360 18050 -335
rect 18025 -405 18050 -380
rect 18085 -360 18110 -335
rect 18085 -405 18110 -380
rect 18145 -360 18170 -335
rect 18145 -405 18170 -380
rect 18205 -360 18230 -335
rect 18205 -405 18230 -380
rect 18265 -360 18290 -335
rect 18265 -405 18290 -380
rect 18325 -360 18350 -335
rect 18325 -405 18350 -380
rect 18385 -360 18410 -335
rect 18385 -405 18410 -380
rect 18445 -360 18470 -335
rect 18445 -405 18470 -380
rect 18505 -360 18530 -335
rect 18505 -405 18530 -380
rect 18565 -360 18590 -335
rect 18565 -405 18590 -380
rect 18625 -360 18650 -335
rect 18625 -405 18650 -380
rect 18685 -360 18710 -335
rect 18685 -405 18710 -380
rect 18745 -360 18770 -335
rect 18745 -405 18770 -380
rect 18805 -360 18830 -335
rect 18805 -405 18830 -380
rect 18865 -360 18890 -335
rect 18865 -405 18890 -380
rect 18925 -360 18950 -335
rect 18925 -405 18950 -380
rect 18985 -360 19010 -335
rect 18985 -405 19010 -380
rect 19045 -360 19070 -335
rect 19045 -405 19070 -380
rect 19105 -360 19130 -335
rect 19105 -405 19130 -380
rect 19165 -360 19190 -335
rect 19165 -405 19190 -380
rect 19225 -360 19250 -335
rect 19225 -405 19250 -380
rect 19285 -360 19310 -335
rect 19285 -405 19310 -380
rect 19345 -360 19370 -335
rect 19345 -405 19370 -380
rect 19405 -360 19430 -335
rect 19405 -405 19430 -380
rect 19465 -360 19490 -335
rect 19465 -405 19490 -380
rect 19525 -360 19550 -335
rect 19525 -405 19550 -380
rect 19585 -360 19610 -335
rect 19585 -405 19610 -380
rect 19645 -360 19670 -335
rect 19645 -405 19670 -380
rect 19705 -360 19730 -335
rect 19705 -405 19730 -380
rect 19765 -360 19790 -335
rect 19765 -405 19790 -380
rect 19825 -360 19850 -335
rect 19825 -405 19850 -380
rect 19885 -360 19910 -335
rect 19885 -405 19910 -380
rect 19945 -360 19970 -335
rect 19945 -405 19970 -380
rect 20005 -360 20030 -335
rect 20005 -405 20030 -380
rect 20065 -360 20090 -335
rect 20065 -405 20090 -380
rect 20125 -360 20150 -335
rect 20125 -405 20150 -380
rect 20185 -360 20210 -335
rect 20185 -405 20210 -380
rect 20245 -360 20270 -335
rect 20245 -405 20270 -380
rect 20305 -360 20330 -335
rect 20305 -405 20330 -380
rect 20365 -360 20390 -335
rect 20365 -405 20390 -380
rect 20425 -360 20450 -335
rect 20425 -405 20450 -380
rect 20485 -360 20510 -335
rect 20485 -405 20510 -380
rect 20545 -360 20570 -335
rect 20545 -405 20570 -380
rect 20605 -360 20630 -335
rect 20605 -405 20630 -380
rect 20665 -360 20690 -335
rect 20665 -405 20690 -380
rect 20725 -360 20750 -335
rect 20725 -405 20750 -380
rect 20785 -360 20810 -335
rect 20785 -405 20810 -380
rect 20845 -360 20870 -335
rect 20845 -405 20870 -380
rect 20905 -360 20930 -335
rect 20905 -405 20930 -380
rect 20965 -360 20990 -335
rect 20965 -405 20990 -380
rect 21025 -360 21050 -335
rect 21025 -405 21050 -380
rect 21085 -360 21110 -335
rect 21085 -405 21110 -380
rect 21145 -360 21170 -335
rect 21145 -405 21170 -380
rect 21205 -360 21230 -335
rect 21205 -405 21230 -380
rect 21265 -360 21290 -335
rect 21265 -405 21290 -380
rect 21325 -360 21350 -335
rect 21325 -405 21350 -380
rect 21385 -360 21410 -335
rect 21385 -405 21410 -380
rect 21445 -360 21470 -335
rect 21445 -405 21470 -380
rect 21505 -360 21530 -335
rect 21505 -405 21530 -380
rect 21565 -360 21590 -335
rect 21565 -405 21590 -380
rect 21625 -360 21650 -335
rect 21625 -405 21650 -380
rect 21685 -360 21710 -335
rect 21685 -405 21710 -380
rect 21745 -360 21770 -335
rect 21745 -405 21770 -380
rect 21805 -360 21830 -335
rect 21805 -405 21830 -380
rect 21865 -360 21890 -335
rect 21865 -405 21890 -380
rect 21925 -360 21950 -335
rect 21925 -405 21950 -380
rect 21985 -360 22010 -335
rect 21985 -405 22010 -380
rect 22045 -360 22070 -335
rect 22045 -405 22070 -380
rect 22105 -360 22130 -335
rect 22105 -405 22130 -380
rect 22165 -360 22190 -335
rect 22165 -405 22190 -380
rect 22225 -360 22250 -335
rect 22225 -405 22250 -380
rect 22285 -360 22310 -335
rect 22285 -405 22310 -380
rect 22345 -360 22370 -335
rect 22345 -405 22370 -380
rect 22405 -360 22430 -335
rect 22405 -405 22430 -380
rect 22465 -360 22490 -335
rect 22465 -405 22490 -380
rect 22525 -360 22550 -335
rect 22525 -405 22550 -380
rect 22585 -360 22610 -335
rect 22585 -405 22610 -380
rect 22645 -360 22670 -335
rect 22645 -405 22670 -380
rect 22705 -360 22730 -335
rect 22705 -405 22730 -380
rect 22765 -360 22790 -335
rect 22765 -405 22790 -380
rect 22825 -360 22850 -335
rect 22825 -405 22850 -380
rect 22885 -360 22910 -335
rect 22885 -405 22910 -380
rect 22945 -360 22970 -335
rect 22945 -405 22970 -380
rect 23005 -360 23030 -335
rect 23005 -405 23030 -380
rect 23065 -360 23090 -335
rect 23065 -405 23090 -380
rect 23125 -360 23150 -335
rect 23125 -405 23150 -380
rect 23185 -360 23210 -335
rect 23185 -405 23210 -380
rect 23245 -360 23270 -335
rect 23245 -405 23270 -380
rect 23305 -360 23330 -335
rect 23305 -405 23330 -380
rect 23365 -360 23390 -335
rect 23365 -405 23390 -380
rect 23425 -360 23450 -335
rect 23425 -405 23450 -380
rect 23485 -360 23510 -335
rect 23485 -405 23510 -380
rect 23545 -360 23570 -335
rect 23545 -405 23570 -380
rect 23605 -360 23630 -335
rect 23605 -405 23630 -380
rect 23665 -360 23690 -335
rect 23665 -405 23690 -380
rect 23725 -360 23750 -335
rect 23725 -405 23750 -380
rect 23785 -360 23810 -335
rect 23785 -405 23810 -380
rect 23845 -360 23870 -335
rect 23845 -405 23870 -380
rect 23905 -360 23930 -335
rect 23905 -405 23930 -380
rect 23965 -360 23990 -335
rect 23965 -405 23990 -380
rect 24025 -360 24050 -335
rect 24025 -405 24050 -380
rect 24085 -360 24110 -335
rect 24085 -405 24110 -380
rect 24145 -360 24170 -335
rect 24145 -405 24170 -380
rect 24205 -360 24230 -335
rect 24205 -405 24230 -380
rect 24265 -360 24290 -335
rect 24265 -405 24290 -380
rect 24325 -360 24350 -335
rect 24325 -405 24350 -380
rect 24385 -360 24410 -335
rect 24385 -405 24410 -380
rect 24445 -360 24470 -335
rect 24445 -405 24470 -380
rect 24505 -360 24530 -335
rect 24505 -405 24530 -380
rect 24565 -360 24590 -335
rect 24565 -405 24590 -380
rect 24625 -360 24650 -335
rect 24625 -405 24650 -380
rect 24685 -360 24710 -335
rect 24685 -405 24710 -380
rect 24745 -360 24770 -335
rect 24745 -405 24770 -380
rect 24805 -360 24830 -335
rect 24805 -405 24830 -380
rect 24865 -360 24890 -335
rect 24865 -405 24890 -380
rect 24925 -360 24950 -335
rect 24925 -405 24950 -380
rect 24985 -360 25010 -335
rect 24985 -405 25010 -380
rect 25045 -360 25070 -335
rect 25045 -405 25070 -380
rect 25105 -360 25130 -335
rect 25105 -405 25130 -380
rect 25165 -360 25190 -335
rect 25165 -405 25190 -380
rect 25225 -360 25250 -335
rect 25225 -405 25250 -380
rect 25285 -360 25310 -335
rect 25285 -405 25310 -380
rect 25345 -360 25370 -335
rect 25345 -405 25370 -380
rect 25405 -360 25430 -335
rect 25405 -405 25430 -380
rect 25465 -360 25490 -335
rect 25465 -405 25490 -380
rect 25525 -360 25550 -335
rect 25525 -405 25550 -380
rect 25585 -360 25610 -335
rect 25585 -405 25610 -380
rect 25645 -360 25670 -335
rect 25645 -405 25670 -380
rect 25705 -360 25730 -335
rect 25705 -405 25730 -380
rect 25765 -360 25790 -335
rect 25765 -405 25790 -380
rect 25825 -360 25850 -335
rect 25825 -405 25850 -380
rect 25885 -360 25910 -335
rect 25885 -405 25910 -380
rect 25945 -360 25970 -335
rect 25945 -405 25970 -380
rect 26005 -360 26030 -335
rect 26005 -405 26030 -380
rect 26065 -360 26090 -335
rect 26065 -405 26090 -380
rect 26125 -360 26150 -335
rect 26125 -405 26150 -380
rect 26185 -360 26210 -335
rect 26185 -405 26210 -380
rect 26245 -360 26270 -335
rect 26245 -405 26270 -380
rect 26305 -360 26330 -335
rect 26305 -405 26330 -380
rect 26365 -360 26390 -335
rect 26365 -405 26390 -380
rect 26425 -360 26450 -335
rect 26425 -405 26450 -380
rect 26485 -360 26510 -335
rect 26485 -405 26510 -380
rect 26545 -360 26570 -335
rect 26545 -405 26570 -380
rect 26605 -360 26630 -335
rect 26605 -405 26630 -380
rect 26665 -360 26690 -335
rect 26665 -405 26690 -380
rect 26725 -360 26750 -335
rect 26725 -405 26750 -380
rect 26785 -360 26810 -335
rect 26785 -405 26810 -380
rect 26845 -360 26870 -335
rect 26845 -405 26870 -380
rect 26905 -360 26930 -335
rect 26905 -405 26930 -380
rect 26965 -360 26990 -335
rect 26965 -405 26990 -380
rect 27025 -360 27050 -335
rect 27025 -405 27050 -380
rect 27085 -360 27110 -335
rect 27085 -405 27110 -380
rect 27145 -360 27170 -335
rect 27145 -405 27170 -380
rect 27205 -360 27230 -335
rect 27205 -405 27230 -380
rect 27265 -360 27290 -335
rect 27265 -405 27290 -380
rect 27325 -360 27350 -335
rect 27325 -405 27350 -380
rect 27385 -360 27410 -335
rect 27385 -405 27410 -380
rect 27445 -360 27470 -335
rect 27445 -405 27470 -380
rect 27505 -360 27530 -335
rect 27505 -405 27530 -380
rect 27565 -360 27590 -335
rect 27565 -405 27590 -380
rect 27625 -360 27650 -335
rect 27625 -405 27650 -380
rect 27685 -360 27710 -335
rect 27685 -405 27710 -380
rect 27745 -360 27770 -335
rect 27745 -405 27770 -380
rect 27805 -360 27830 -335
rect 27805 -405 27830 -380
rect 27865 -360 27890 -335
rect 27865 -405 27890 -380
rect 27925 -360 27950 -335
rect 27925 -405 27950 -380
rect 27985 -360 28010 -335
rect 27985 -405 28010 -380
rect 28045 -360 28070 -335
rect 28045 -405 28070 -380
rect 28105 -360 28130 -335
rect 28105 -405 28130 -380
rect 28165 -360 28190 -335
rect 28165 -405 28190 -380
rect 28225 -360 28250 -335
rect 28225 -405 28250 -380
rect 28285 -360 28310 -335
rect 28285 -405 28310 -380
rect 28345 -360 28370 -335
rect 28345 -405 28370 -380
rect 28405 -360 28430 -335
rect 28405 -405 28430 -380
rect 28465 -360 28490 -335
rect 28465 -405 28490 -380
rect 28525 -360 28550 -335
rect 28525 -405 28550 -380
rect 28585 -360 28610 -335
rect 28585 -405 28610 -380
rect 28645 -360 28670 -335
rect 28645 -405 28670 -380
rect 28705 -360 28730 -335
rect 28705 -405 28730 -380
rect 28765 -360 28790 -335
rect 28765 -405 28790 -380
rect 28825 -360 28850 -335
rect 28825 -405 28850 -380
rect 28885 -360 28910 -335
rect 28885 -405 28910 -380
rect 28945 -360 28970 -335
rect 28945 -405 28970 -380
rect 29005 -360 29030 -335
rect 29005 -405 29030 -380
rect 29065 -360 29090 -335
rect 29065 -405 29090 -380
rect 29125 -360 29150 -335
rect 29125 -405 29150 -380
rect 29185 -360 29210 -335
rect 29185 -405 29210 -380
rect 29245 -360 29270 -335
rect 29245 -405 29270 -380
rect 29305 -360 29330 -335
rect 29305 -405 29330 -380
rect 29365 -360 29390 -335
rect 29365 -405 29390 -380
rect 29425 -360 29450 -335
rect 29425 -405 29450 -380
rect 29485 -360 29510 -335
rect 29485 -405 29510 -380
rect 29545 -360 29570 -335
rect 29545 -405 29570 -380
rect 29605 -360 29630 -335
rect 29605 -405 29630 -380
rect 29665 -360 29690 -335
rect 29665 -405 29690 -380
rect 29725 -360 29750 -335
rect 29725 -405 29750 -380
rect 29785 -360 29810 -335
rect 29785 -405 29810 -380
rect 29845 -360 29870 -335
rect 29845 -405 29870 -380
rect 29905 -360 29930 -335
rect 29905 -405 29930 -380
rect 29965 -360 29990 -335
rect 29965 -405 29990 -380
rect 30025 -360 30050 -335
rect 30025 -405 30050 -380
rect 30085 -360 30110 -335
rect 30085 -405 30110 -380
rect 30145 -360 30170 -335
rect 30145 -405 30170 -380
rect 30205 -360 30230 -335
rect 30205 -405 30230 -380
rect 30265 -360 30290 -335
rect 30265 -405 30290 -380
rect 30325 -360 30350 -335
rect 30325 -405 30350 -380
rect 30385 -360 30410 -335
rect 30385 -405 30410 -380
rect 30445 -360 30470 -335
rect 30445 -405 30470 -380
rect 30505 -360 30530 -335
rect 30505 -405 30530 -380
rect 30565 -360 30590 -335
rect 30565 -405 30590 -380
rect 30625 -360 30650 -335
rect 30625 -405 30650 -380
rect 30685 -360 30710 -335
rect 30685 -405 30710 -380
<< pdiffc >>
rect 441 240 466 265
rect 746 240 771 265
rect 991 240 1016 265
rect 1231 240 1256 265
rect 1476 240 1501 265
rect 1781 240 1806 265
rect 2026 240 2051 265
rect 2511 240 2536 265
rect 2751 240 2776 265
rect 2996 240 3021 265
rect 3236 240 3261 265
rect 3481 240 3506 265
rect 3721 240 3746 265
rect 3966 240 3991 265
rect 4451 240 4476 265
rect 4691 240 4716 265
rect 4936 240 4961 265
rect 5176 240 5201 265
rect 5421 240 5446 265
rect 5726 240 5751 265
rect 5971 240 5996 265
rect 6211 240 6236 265
rect 6696 240 6721 265
rect 6941 240 6966 265
rect 7181 240 7206 265
rect 7421 240 7446 265
rect 7661 240 7686 265
rect 7906 240 7931 265
rect 8146 240 8171 265
rect 8391 240 8416 265
rect 8631 240 8656 265
rect 8876 240 8901 265
rect 9116 240 9141 265
rect 9606 240 9631 265
rect 9851 240 9876 265
rect 10091 240 10116 265
rect 10336 240 10361 265
rect 10576 240 10601 265
rect 10821 240 10846 265
rect 11061 240 11086 265
rect 11546 240 11571 265
rect 11791 240 11816 265
rect 12031 240 12056 265
rect 12276 240 12301 265
rect 12516 240 12541 265
rect 12761 240 12786 265
rect 13246 240 13271 265
rect 13486 240 13511 265
rect 13731 240 13756 265
rect 13971 240 13996 265
rect 14216 240 14241 265
rect 14456 240 14481 265
rect 14701 240 14726 265
rect 14941 240 14966 265
rect 15426 240 15451 265
rect 15671 240 15696 265
rect 15911 240 15936 265
rect 16156 240 16181 265
rect 16396 240 16421 265
rect 16641 240 16666 265
rect 16881 240 16906 265
rect 17126 240 17151 265
rect 17611 240 17636 265
rect 17851 240 17876 265
rect 18096 240 18121 265
rect 18336 240 18361 265
rect 18581 240 18606 265
rect 18821 240 18846 265
rect 19066 240 19091 265
rect 19306 240 19331 265
rect 19791 240 19816 265
rect 20036 240 20061 265
rect 20276 240 20301 265
rect 20521 240 20546 265
rect 21006 240 21031 265
rect 196 140 221 165
rect 196 95 221 120
rect 256 140 281 165
rect 256 95 281 120
rect 321 140 346 165
rect 321 95 346 120
rect 381 140 406 165
rect 381 95 406 120
rect 441 140 466 165
rect 441 95 466 120
rect 501 140 526 165
rect 501 95 526 120
rect 561 140 586 165
rect 561 95 586 120
rect 626 140 651 165
rect 626 95 651 120
rect 686 140 711 165
rect 686 95 711 120
rect 746 140 771 165
rect 746 95 771 120
rect 806 140 831 165
rect 806 95 831 120
rect 871 140 896 165
rect 871 95 896 120
rect 931 140 956 165
rect 931 95 956 120
rect 991 140 1016 165
rect 991 95 1016 120
rect 1051 140 1076 165
rect 1051 95 1076 120
rect 1111 140 1136 165
rect 1111 95 1136 120
rect 1171 140 1196 165
rect 1171 95 1196 120
rect 1231 140 1256 165
rect 1231 95 1256 120
rect 1291 140 1316 165
rect 1291 95 1316 120
rect 1356 140 1381 165
rect 1356 95 1381 120
rect 1416 140 1441 165
rect 1416 95 1441 120
rect 1476 140 1501 165
rect 1476 95 1501 120
rect 1536 140 1561 165
rect 1536 95 1561 120
rect 1596 140 1621 165
rect 1596 95 1621 120
rect 1661 140 1686 165
rect 1661 95 1686 120
rect 1721 140 1746 165
rect 1721 95 1746 120
rect 1781 140 1806 165
rect 1781 95 1806 120
rect 1841 140 1866 165
rect 1841 95 1866 120
rect 1906 140 1931 165
rect 1906 95 1931 120
rect 1966 140 1991 165
rect 1966 95 1991 120
rect 2026 140 2051 165
rect 2026 95 2051 120
rect 2086 140 2111 165
rect 2086 95 2111 120
rect 2146 140 2171 165
rect 2146 95 2171 120
rect 2206 140 2231 165
rect 2206 95 2231 120
rect 2266 140 2291 165
rect 2266 95 2291 120
rect 2326 140 2351 165
rect 2326 95 2351 120
rect 2391 140 2416 165
rect 2391 95 2416 120
rect 2451 140 2476 165
rect 2451 95 2476 120
rect 2511 140 2536 165
rect 2511 95 2536 120
rect 2571 140 2596 165
rect 2571 95 2596 120
rect 2631 140 2656 165
rect 2631 95 2656 120
rect 2691 140 2716 165
rect 2691 95 2716 120
rect 2751 140 2776 165
rect 2751 95 2776 120
rect 2811 140 2836 165
rect 2811 95 2836 120
rect 2876 140 2901 165
rect 2876 95 2901 120
rect 2936 140 2961 165
rect 2936 95 2961 120
rect 2996 140 3021 165
rect 2996 95 3021 120
rect 3056 140 3081 165
rect 3056 95 3081 120
rect 3116 140 3141 165
rect 3116 95 3141 120
rect 3176 140 3201 165
rect 3176 95 3201 120
rect 3236 140 3261 165
rect 3236 95 3261 120
rect 3296 140 3321 165
rect 3296 95 3321 120
rect 3361 140 3386 165
rect 3361 95 3386 120
rect 3421 140 3446 165
rect 3421 95 3446 120
rect 3481 140 3506 165
rect 3481 95 3506 120
rect 3541 140 3566 165
rect 3541 95 3566 120
rect 3601 140 3626 165
rect 3601 95 3626 120
rect 3661 140 3686 165
rect 3661 95 3686 120
rect 3721 140 3746 165
rect 3721 95 3746 120
rect 3781 140 3806 165
rect 3781 95 3806 120
rect 3846 140 3871 165
rect 3846 95 3871 120
rect 3906 140 3931 165
rect 3906 95 3931 120
rect 3966 140 3991 165
rect 3966 95 3991 120
rect 4026 140 4051 165
rect 4026 95 4051 120
rect 4086 140 4111 165
rect 4086 95 4111 120
rect 4146 140 4171 165
rect 4146 95 4171 120
rect 4206 140 4231 165
rect 4206 95 4231 120
rect 4266 140 4291 165
rect 4266 95 4291 120
rect 4331 140 4356 165
rect 4331 95 4356 120
rect 4391 140 4416 165
rect 4391 95 4416 120
rect 4451 140 4476 165
rect 4451 95 4476 120
rect 4511 140 4536 165
rect 4511 95 4536 120
rect 4571 140 4596 165
rect 4571 95 4596 120
rect 4631 140 4656 165
rect 4631 95 4656 120
rect 4691 140 4716 165
rect 4691 95 4716 120
rect 4751 140 4776 165
rect 4751 95 4776 120
rect 4816 140 4841 165
rect 4816 95 4841 120
rect 4876 140 4901 165
rect 4876 95 4901 120
rect 4936 140 4961 165
rect 4936 95 4961 120
rect 4996 140 5021 165
rect 4996 95 5021 120
rect 5056 140 5081 165
rect 5056 95 5081 120
rect 5116 140 5141 165
rect 5116 95 5141 120
rect 5176 140 5201 165
rect 5176 95 5201 120
rect 5236 140 5261 165
rect 5236 95 5261 120
rect 5301 140 5326 165
rect 5301 95 5326 120
rect 5361 140 5386 165
rect 5361 95 5386 120
rect 5421 140 5446 165
rect 5421 95 5446 120
rect 5481 140 5506 165
rect 5481 95 5506 120
rect 5541 140 5566 165
rect 5541 95 5566 120
rect 5606 140 5631 165
rect 5606 95 5631 120
rect 5666 140 5691 165
rect 5666 95 5691 120
rect 5726 140 5751 165
rect 5726 95 5751 120
rect 5786 140 5811 165
rect 5786 95 5811 120
rect 5851 140 5876 165
rect 5851 95 5876 120
rect 5911 140 5936 165
rect 5911 95 5936 120
rect 5971 140 5996 165
rect 5971 95 5996 120
rect 6031 140 6056 165
rect 6031 95 6056 120
rect 6091 140 6116 165
rect 6091 95 6116 120
rect 6151 140 6176 165
rect 6151 95 6176 120
rect 6211 140 6236 165
rect 6211 95 6236 120
rect 6271 140 6296 165
rect 6271 95 6296 120
rect 6336 140 6361 165
rect 6336 95 6361 120
rect 6396 140 6421 165
rect 6396 95 6421 120
rect 6456 140 6481 165
rect 6456 95 6481 120
rect 6516 140 6541 165
rect 6516 95 6541 120
rect 6576 140 6601 165
rect 6576 95 6601 120
rect 6636 140 6661 165
rect 6636 95 6661 120
rect 6696 140 6721 165
rect 6696 95 6721 120
rect 6756 140 6781 165
rect 6756 95 6781 120
rect 6821 140 6846 165
rect 6821 95 6846 120
rect 6881 140 6906 165
rect 6881 95 6906 120
rect 6941 140 6966 165
rect 6941 95 6966 120
rect 7001 140 7026 165
rect 7001 95 7026 120
rect 7061 140 7086 165
rect 7061 95 7086 120
rect 7121 140 7146 165
rect 7121 95 7146 120
rect 7181 140 7206 165
rect 7181 95 7206 120
rect 7241 140 7266 165
rect 7241 95 7266 120
rect 7301 140 7326 165
rect 7301 95 7326 120
rect 7361 140 7386 165
rect 7361 95 7386 120
rect 7421 140 7446 165
rect 7421 95 7446 120
rect 7481 140 7506 165
rect 7481 95 7506 120
rect 7541 140 7566 165
rect 7541 95 7566 120
rect 7601 140 7626 165
rect 7601 95 7626 120
rect 7661 140 7686 165
rect 7661 95 7686 120
rect 7721 140 7746 165
rect 7721 95 7746 120
rect 7786 140 7811 165
rect 7786 95 7811 120
rect 7846 140 7871 165
rect 7846 95 7871 120
rect 7906 140 7931 165
rect 7906 95 7931 120
rect 7966 140 7991 165
rect 7966 95 7991 120
rect 8026 140 8051 165
rect 8026 95 8051 120
rect 8086 140 8111 165
rect 8086 95 8111 120
rect 8146 140 8171 165
rect 8146 95 8171 120
rect 8206 140 8231 165
rect 8206 95 8231 120
rect 8271 140 8296 165
rect 8271 95 8296 120
rect 8331 140 8356 165
rect 8331 95 8356 120
rect 8391 140 8416 165
rect 8391 95 8416 120
rect 8451 140 8476 165
rect 8451 95 8476 120
rect 8511 140 8536 165
rect 8511 95 8536 120
rect 8571 140 8596 165
rect 8571 95 8596 120
rect 8631 140 8656 165
rect 8631 95 8656 120
rect 8691 140 8716 165
rect 8691 95 8716 120
rect 8756 140 8781 165
rect 8756 95 8781 120
rect 8816 140 8841 165
rect 8816 95 8841 120
rect 8876 140 8901 165
rect 8876 95 8901 120
rect 8936 140 8961 165
rect 8936 95 8961 120
rect 8996 140 9021 165
rect 8996 95 9021 120
rect 9056 140 9081 165
rect 9056 95 9081 120
rect 9116 140 9141 165
rect 9116 95 9141 120
rect 9176 140 9201 165
rect 9176 95 9201 120
rect 9241 140 9266 165
rect 9241 95 9266 120
rect 9301 140 9326 165
rect 9301 95 9326 120
rect 9361 140 9386 165
rect 9361 95 9386 120
rect 9421 140 9446 165
rect 9421 95 9446 120
rect 9486 140 9511 165
rect 9486 95 9511 120
rect 9546 140 9571 165
rect 9546 95 9571 120
rect 9606 140 9631 165
rect 9606 95 9631 120
rect 9666 140 9691 165
rect 9666 95 9691 120
rect 9731 140 9756 165
rect 9731 95 9756 120
rect 9791 140 9816 165
rect 9791 95 9816 120
rect 9851 140 9876 165
rect 9851 95 9876 120
rect 9911 140 9936 165
rect 9911 95 9936 120
rect 9971 140 9996 165
rect 9971 95 9996 120
rect 10031 140 10056 165
rect 10031 95 10056 120
rect 10091 140 10116 165
rect 10091 95 10116 120
rect 10151 140 10176 165
rect 10151 95 10176 120
rect 10216 140 10241 165
rect 10216 95 10241 120
rect 10276 140 10301 165
rect 10276 95 10301 120
rect 10336 140 10361 165
rect 10336 95 10361 120
rect 10396 140 10421 165
rect 10396 95 10421 120
rect 10456 140 10481 165
rect 10456 95 10481 120
rect 10516 140 10541 165
rect 10516 95 10541 120
rect 10576 140 10601 165
rect 10576 95 10601 120
rect 10636 140 10661 165
rect 10636 95 10661 120
rect 10701 140 10726 165
rect 10701 95 10726 120
rect 10761 140 10786 165
rect 10761 95 10786 120
rect 10821 140 10846 165
rect 10821 95 10846 120
rect 10881 140 10906 165
rect 10881 95 10906 120
rect 10941 140 10966 165
rect 10941 95 10966 120
rect 11001 140 11026 165
rect 11001 95 11026 120
rect 11061 140 11086 165
rect 11061 95 11086 120
rect 11121 140 11146 165
rect 11121 95 11146 120
rect 11186 140 11211 165
rect 11186 95 11211 120
rect 11246 140 11271 165
rect 11246 95 11271 120
rect 11306 140 11331 165
rect 11306 95 11331 120
rect 11366 140 11391 165
rect 11366 95 11391 120
rect 11426 140 11451 165
rect 11426 95 11451 120
rect 11486 140 11511 165
rect 11486 95 11511 120
rect 11546 140 11571 165
rect 11546 95 11571 120
rect 11606 140 11631 165
rect 11606 95 11631 120
rect 11671 140 11696 165
rect 11671 95 11696 120
rect 11731 140 11756 165
rect 11731 95 11756 120
rect 11791 140 11816 165
rect 11791 95 11816 120
rect 11851 140 11876 165
rect 11851 95 11876 120
rect 11911 140 11936 165
rect 11911 95 11936 120
rect 11971 140 11996 165
rect 11971 95 11996 120
rect 12031 140 12056 165
rect 12031 95 12056 120
rect 12091 140 12116 165
rect 12091 95 12116 120
rect 12156 140 12181 165
rect 12156 95 12181 120
rect 12216 140 12241 165
rect 12216 95 12241 120
rect 12276 140 12301 165
rect 12276 95 12301 120
rect 12336 140 12361 165
rect 12336 95 12361 120
rect 12396 140 12421 165
rect 12396 95 12421 120
rect 12456 140 12481 165
rect 12456 95 12481 120
rect 12516 140 12541 165
rect 12516 95 12541 120
rect 12576 140 12601 165
rect 12576 95 12601 120
rect 12641 140 12666 165
rect 12641 95 12666 120
rect 12701 140 12726 165
rect 12701 95 12726 120
rect 12761 140 12786 165
rect 12761 95 12786 120
rect 12821 140 12846 165
rect 12821 95 12846 120
rect 12881 140 12906 165
rect 12881 95 12906 120
rect 12941 140 12966 165
rect 12941 95 12966 120
rect 13001 140 13026 165
rect 13001 95 13026 120
rect 13061 140 13086 165
rect 13061 95 13086 120
rect 13126 140 13151 165
rect 13126 95 13151 120
rect 13186 140 13211 165
rect 13186 95 13211 120
rect 13246 140 13271 165
rect 13246 95 13271 120
rect 13306 140 13331 165
rect 13306 95 13331 120
rect 13366 140 13391 165
rect 13366 95 13391 120
rect 13426 140 13451 165
rect 13426 95 13451 120
rect 13486 140 13511 165
rect 13486 95 13511 120
rect 13546 140 13571 165
rect 13546 95 13571 120
rect 13611 140 13636 165
rect 13611 95 13636 120
rect 13671 140 13696 165
rect 13671 95 13696 120
rect 13731 140 13756 165
rect 13731 95 13756 120
rect 13791 140 13816 165
rect 13791 95 13816 120
rect 13851 140 13876 165
rect 13851 95 13876 120
rect 13911 140 13936 165
rect 13911 95 13936 120
rect 13971 140 13996 165
rect 13971 95 13996 120
rect 14031 140 14056 165
rect 14031 95 14056 120
rect 14096 140 14121 165
rect 14096 95 14121 120
rect 14156 140 14181 165
rect 14156 95 14181 120
rect 14216 140 14241 165
rect 14216 95 14241 120
rect 14276 140 14301 165
rect 14276 95 14301 120
rect 14336 140 14361 165
rect 14336 95 14361 120
rect 14396 140 14421 165
rect 14396 95 14421 120
rect 14456 140 14481 165
rect 14456 95 14481 120
rect 14516 140 14541 165
rect 14516 95 14541 120
rect 14581 140 14606 165
rect 14581 95 14606 120
rect 14641 140 14666 165
rect 14641 95 14666 120
rect 14701 140 14726 165
rect 14701 95 14726 120
rect 14761 140 14786 165
rect 14761 95 14786 120
rect 14821 140 14846 165
rect 14821 95 14846 120
rect 14881 140 14906 165
rect 14881 95 14906 120
rect 14941 140 14966 165
rect 14941 95 14966 120
rect 15001 140 15026 165
rect 15001 95 15026 120
rect 15066 140 15091 165
rect 15066 95 15091 120
rect 15126 140 15151 165
rect 15126 95 15151 120
rect 15186 140 15211 165
rect 15186 95 15211 120
rect 15246 140 15271 165
rect 15246 95 15271 120
rect 15306 140 15331 165
rect 15306 95 15331 120
rect 15366 140 15391 165
rect 15366 95 15391 120
rect 15426 140 15451 165
rect 15426 95 15451 120
rect 15486 140 15511 165
rect 15486 95 15511 120
rect 15551 140 15576 165
rect 15551 95 15576 120
rect 15611 140 15636 165
rect 15611 95 15636 120
rect 15671 140 15696 165
rect 15671 95 15696 120
rect 15731 140 15756 165
rect 15731 95 15756 120
rect 15791 140 15816 165
rect 15791 95 15816 120
rect 15851 140 15876 165
rect 15851 95 15876 120
rect 15911 140 15936 165
rect 15911 95 15936 120
rect 15971 140 15996 165
rect 15971 95 15996 120
rect 16036 140 16061 165
rect 16036 95 16061 120
rect 16096 140 16121 165
rect 16096 95 16121 120
rect 16156 140 16181 165
rect 16156 95 16181 120
rect 16216 140 16241 165
rect 16216 95 16241 120
rect 16276 140 16301 165
rect 16276 95 16301 120
rect 16336 140 16361 165
rect 16336 95 16361 120
rect 16396 140 16421 165
rect 16396 95 16421 120
rect 16456 140 16481 165
rect 16456 95 16481 120
rect 16521 140 16546 165
rect 16521 95 16546 120
rect 16581 140 16606 165
rect 16581 95 16606 120
rect 16641 140 16666 165
rect 16641 95 16666 120
rect 16701 140 16726 165
rect 16701 95 16726 120
rect 16761 140 16786 165
rect 16761 95 16786 120
rect 16821 140 16846 165
rect 16821 95 16846 120
rect 16881 140 16906 165
rect 16881 95 16906 120
rect 16941 140 16966 165
rect 16941 95 16966 120
rect 17006 140 17031 165
rect 17006 95 17031 120
rect 17066 140 17091 165
rect 17066 95 17091 120
rect 17126 140 17151 165
rect 17126 95 17151 120
rect 17186 140 17211 165
rect 17186 95 17211 120
rect 17246 140 17271 165
rect 17246 95 17271 120
rect 17306 140 17331 165
rect 17306 95 17331 120
rect 17366 140 17391 165
rect 17366 95 17391 120
rect 17426 140 17451 165
rect 17426 95 17451 120
rect 17491 140 17516 165
rect 17491 95 17516 120
rect 17551 140 17576 165
rect 17551 95 17576 120
rect 17611 140 17636 165
rect 17611 95 17636 120
rect 17671 140 17696 165
rect 17671 95 17696 120
rect 17731 140 17756 165
rect 17731 95 17756 120
rect 17791 140 17816 165
rect 17791 95 17816 120
rect 17851 140 17876 165
rect 17851 95 17876 120
rect 17911 140 17936 165
rect 17911 95 17936 120
rect 17976 140 18001 165
rect 17976 95 18001 120
rect 18036 140 18061 165
rect 18036 95 18061 120
rect 18096 140 18121 165
rect 18096 95 18121 120
rect 18156 140 18181 165
rect 18156 95 18181 120
rect 18216 140 18241 165
rect 18216 95 18241 120
rect 18276 140 18301 165
rect 18276 95 18301 120
rect 18336 140 18361 165
rect 18336 95 18361 120
rect 18396 140 18421 165
rect 18396 95 18421 120
rect 18461 140 18486 165
rect 18461 95 18486 120
rect 18521 140 18546 165
rect 18521 95 18546 120
rect 18581 140 18606 165
rect 18581 95 18606 120
rect 18641 140 18666 165
rect 18641 95 18666 120
rect 18701 140 18726 165
rect 18701 95 18726 120
rect 18761 140 18786 165
rect 18761 95 18786 120
rect 18821 140 18846 165
rect 18821 95 18846 120
rect 18881 140 18906 165
rect 18881 95 18906 120
rect 18946 140 18971 165
rect 18946 95 18971 120
rect 19006 140 19031 165
rect 19006 95 19031 120
rect 19066 140 19091 165
rect 19066 95 19091 120
rect 19126 140 19151 165
rect 19126 95 19151 120
rect 19186 140 19211 165
rect 19186 95 19211 120
rect 19246 140 19271 165
rect 19246 95 19271 120
rect 19306 140 19331 165
rect 19306 95 19331 120
rect 19366 140 19391 165
rect 19366 95 19391 120
rect 19431 140 19456 165
rect 19431 95 19456 120
rect 19491 140 19516 165
rect 19491 95 19516 120
rect 19551 140 19576 165
rect 19551 95 19576 120
rect 19611 140 19636 165
rect 19611 95 19636 120
rect 19671 140 19696 165
rect 19671 95 19696 120
rect 19731 140 19756 165
rect 19731 95 19756 120
rect 19791 140 19816 165
rect 19791 95 19816 120
rect 19851 140 19876 165
rect 19851 95 19876 120
rect 19916 140 19941 165
rect 19916 95 19941 120
rect 19976 140 20001 165
rect 19976 95 20001 120
rect 20036 140 20061 165
rect 20036 95 20061 120
rect 20096 140 20121 165
rect 20096 95 20121 120
rect 20156 140 20181 165
rect 20156 95 20181 120
rect 20216 140 20241 165
rect 20216 95 20241 120
rect 20276 140 20301 165
rect 20276 95 20301 120
rect 20336 140 20361 165
rect 20336 95 20361 120
rect 20401 140 20426 165
rect 20401 95 20426 120
rect 20461 140 20486 165
rect 20461 95 20486 120
rect 20521 140 20546 165
rect 20521 95 20546 120
rect 20581 140 20606 165
rect 20581 95 20606 120
rect 20641 140 20666 165
rect 20641 95 20666 120
rect 20701 140 20726 165
rect 20701 95 20726 120
rect 20761 140 20786 165
rect 20761 95 20786 120
rect 20821 140 20846 165
rect 20821 95 20846 120
rect 20886 140 20911 165
rect 20886 95 20911 120
rect 20946 140 20971 165
rect 20946 95 20971 120
rect 21006 140 21031 165
rect 21006 95 21031 120
rect 21066 140 21091 165
rect 21066 95 21091 120
rect 21126 140 21151 165
rect 21126 95 21151 120
rect -35 -610 -10 -585
rect -35 -655 -10 -630
rect -35 -700 -10 -675
rect -35 -750 -10 -725
rect 25 -610 50 -585
rect 25 -655 50 -630
rect 25 -700 50 -675
rect 25 -750 50 -725
rect 85 -610 110 -585
rect 85 -655 110 -630
rect 85 -700 110 -675
rect 85 -750 110 -725
rect 145 -610 170 -585
rect 145 -655 170 -630
rect 145 -700 170 -675
rect 145 -750 170 -725
rect 205 -610 230 -585
rect 205 -655 230 -630
rect 205 -700 230 -675
rect 205 -750 230 -725
rect 265 -610 290 -585
rect 265 -655 290 -630
rect 265 -700 290 -675
rect 265 -750 290 -725
rect 325 -610 350 -585
rect 325 -655 350 -630
rect 325 -700 350 -675
rect 325 -750 350 -725
rect 385 -610 410 -585
rect 385 -655 410 -630
rect 385 -700 410 -675
rect 385 -750 410 -725
rect 445 -610 470 -585
rect 445 -655 470 -630
rect 445 -700 470 -675
rect 445 -750 470 -725
rect 505 -610 530 -585
rect 505 -655 530 -630
rect 505 -700 530 -675
rect 505 -750 530 -725
rect 565 -610 590 -585
rect 565 -655 590 -630
rect 565 -700 590 -675
rect 565 -750 590 -725
rect 625 -610 650 -585
rect 625 -655 650 -630
rect 625 -700 650 -675
rect 625 -750 650 -725
rect 685 -610 710 -585
rect 685 -655 710 -630
rect 685 -700 710 -675
rect 685 -750 710 -725
rect 745 -610 770 -585
rect 745 -655 770 -630
rect 745 -700 770 -675
rect 745 -750 770 -725
rect 805 -610 830 -585
rect 805 -655 830 -630
rect 805 -700 830 -675
rect 805 -750 830 -725
rect 865 -610 890 -585
rect 865 -655 890 -630
rect 865 -700 890 -675
rect 865 -750 890 -725
rect 925 -610 950 -585
rect 925 -655 950 -630
rect 925 -700 950 -675
rect 925 -750 950 -725
rect 985 -610 1010 -585
rect 985 -655 1010 -630
rect 985 -700 1010 -675
rect 985 -750 1010 -725
rect 1045 -610 1070 -585
rect 1045 -655 1070 -630
rect 1045 -700 1070 -675
rect 1045 -750 1070 -725
rect 1105 -610 1130 -585
rect 1105 -655 1130 -630
rect 1105 -700 1130 -675
rect 1105 -750 1130 -725
rect 1165 -610 1190 -585
rect 1165 -655 1190 -630
rect 1165 -700 1190 -675
rect 1165 -750 1190 -725
rect 1225 -610 1250 -585
rect 1225 -655 1250 -630
rect 1225 -700 1250 -675
rect 1225 -750 1250 -725
rect 1285 -610 1310 -585
rect 1285 -655 1310 -630
rect 1285 -700 1310 -675
rect 1285 -750 1310 -725
rect 1345 -610 1370 -585
rect 1345 -655 1370 -630
rect 1345 -700 1370 -675
rect 1345 -750 1370 -725
rect 1405 -610 1430 -585
rect 1405 -655 1430 -630
rect 1405 -700 1430 -675
rect 1405 -750 1430 -725
rect 1465 -610 1490 -585
rect 1465 -655 1490 -630
rect 1465 -700 1490 -675
rect 1465 -750 1490 -725
rect 1525 -610 1550 -585
rect 1525 -655 1550 -630
rect 1525 -700 1550 -675
rect 1525 -750 1550 -725
rect 1585 -610 1610 -585
rect 1585 -655 1610 -630
rect 1585 -700 1610 -675
rect 1585 -750 1610 -725
rect 1645 -610 1670 -585
rect 1645 -655 1670 -630
rect 1645 -700 1670 -675
rect 1645 -750 1670 -725
rect 1705 -610 1730 -585
rect 1705 -655 1730 -630
rect 1705 -700 1730 -675
rect 1705 -750 1730 -725
rect 1765 -610 1790 -585
rect 1765 -655 1790 -630
rect 1765 -700 1790 -675
rect 1765 -750 1790 -725
rect 1825 -610 1850 -585
rect 1825 -655 1850 -630
rect 1825 -700 1850 -675
rect 1825 -750 1850 -725
rect 1885 -610 1910 -585
rect 1885 -655 1910 -630
rect 1885 -700 1910 -675
rect 1885 -750 1910 -725
rect 1945 -610 1970 -585
rect 1945 -655 1970 -630
rect 1945 -700 1970 -675
rect 1945 -750 1970 -725
rect 2005 -610 2030 -585
rect 2005 -655 2030 -630
rect 2005 -700 2030 -675
rect 2005 -750 2030 -725
rect 2065 -610 2090 -585
rect 2065 -655 2090 -630
rect 2065 -700 2090 -675
rect 2065 -750 2090 -725
rect 2125 -610 2150 -585
rect 2125 -655 2150 -630
rect 2125 -700 2150 -675
rect 2125 -750 2150 -725
rect 2185 -610 2210 -585
rect 2185 -655 2210 -630
rect 2185 -700 2210 -675
rect 2185 -750 2210 -725
rect 2245 -610 2270 -585
rect 2245 -655 2270 -630
rect 2245 -700 2270 -675
rect 2245 -750 2270 -725
rect 2305 -610 2330 -585
rect 2305 -655 2330 -630
rect 2305 -700 2330 -675
rect 2305 -750 2330 -725
rect 2365 -610 2390 -585
rect 2365 -655 2390 -630
rect 2365 -700 2390 -675
rect 2365 -750 2390 -725
rect 2425 -610 2450 -585
rect 2425 -655 2450 -630
rect 2425 -700 2450 -675
rect 2425 -750 2450 -725
rect 2485 -610 2510 -585
rect 2485 -655 2510 -630
rect 2485 -700 2510 -675
rect 2485 -750 2510 -725
rect 2545 -610 2570 -585
rect 2545 -655 2570 -630
rect 2545 -700 2570 -675
rect 2545 -750 2570 -725
rect 2605 -610 2630 -585
rect 2605 -655 2630 -630
rect 2605 -700 2630 -675
rect 2605 -750 2630 -725
rect 2665 -610 2690 -585
rect 2665 -655 2690 -630
rect 2665 -700 2690 -675
rect 2665 -750 2690 -725
rect 2725 -610 2750 -585
rect 2725 -655 2750 -630
rect 2725 -700 2750 -675
rect 2725 -750 2750 -725
rect 2785 -610 2810 -585
rect 2785 -655 2810 -630
rect 2785 -700 2810 -675
rect 2785 -750 2810 -725
rect 2845 -610 2870 -585
rect 2845 -655 2870 -630
rect 2845 -700 2870 -675
rect 2845 -750 2870 -725
rect 2905 -610 2930 -585
rect 2905 -655 2930 -630
rect 2905 -700 2930 -675
rect 2905 -750 2930 -725
rect 2965 -610 2990 -585
rect 2965 -655 2990 -630
rect 2965 -700 2990 -675
rect 2965 -750 2990 -725
rect 3025 -610 3050 -585
rect 3025 -655 3050 -630
rect 3025 -700 3050 -675
rect 3025 -750 3050 -725
rect 3085 -610 3110 -585
rect 3085 -655 3110 -630
rect 3085 -700 3110 -675
rect 3085 -750 3110 -725
rect 3145 -610 3170 -585
rect 3145 -655 3170 -630
rect 3145 -700 3170 -675
rect 3145 -750 3170 -725
rect 3205 -610 3230 -585
rect 3205 -655 3230 -630
rect 3205 -700 3230 -675
rect 3205 -750 3230 -725
rect 3265 -610 3290 -585
rect 3265 -655 3290 -630
rect 3265 -700 3290 -675
rect 3265 -750 3290 -725
rect 3325 -610 3350 -585
rect 3325 -655 3350 -630
rect 3325 -700 3350 -675
rect 3325 -750 3350 -725
rect 3385 -610 3410 -585
rect 3385 -655 3410 -630
rect 3385 -700 3410 -675
rect 3385 -750 3410 -725
rect 3445 -610 3470 -585
rect 3445 -655 3470 -630
rect 3445 -700 3470 -675
rect 3445 -750 3470 -725
rect 3505 -610 3530 -585
rect 3505 -655 3530 -630
rect 3505 -700 3530 -675
rect 3505 -750 3530 -725
rect 3565 -610 3590 -585
rect 3565 -655 3590 -630
rect 3565 -700 3590 -675
rect 3565 -750 3590 -725
rect 3625 -610 3650 -585
rect 3625 -655 3650 -630
rect 3625 -700 3650 -675
rect 3625 -750 3650 -725
rect 3685 -610 3710 -585
rect 3685 -655 3710 -630
rect 3685 -700 3710 -675
rect 3685 -750 3710 -725
rect 3745 -610 3770 -585
rect 3745 -655 3770 -630
rect 3745 -700 3770 -675
rect 3745 -750 3770 -725
rect 3805 -610 3830 -585
rect 3805 -655 3830 -630
rect 3805 -700 3830 -675
rect 3805 -750 3830 -725
rect 3865 -610 3890 -585
rect 3865 -655 3890 -630
rect 3865 -700 3890 -675
rect 3865 -750 3890 -725
rect 3925 -610 3950 -585
rect 3925 -655 3950 -630
rect 3925 -700 3950 -675
rect 3925 -750 3950 -725
rect 3985 -610 4010 -585
rect 3985 -655 4010 -630
rect 3985 -700 4010 -675
rect 3985 -750 4010 -725
rect 4045 -610 4070 -585
rect 4045 -655 4070 -630
rect 4045 -700 4070 -675
rect 4045 -750 4070 -725
rect 4105 -610 4130 -585
rect 4105 -655 4130 -630
rect 4105 -700 4130 -675
rect 4105 -750 4130 -725
rect 4165 -610 4190 -585
rect 4165 -655 4190 -630
rect 4165 -700 4190 -675
rect 4165 -750 4190 -725
rect 4225 -610 4250 -585
rect 4225 -655 4250 -630
rect 4225 -700 4250 -675
rect 4225 -750 4250 -725
rect 4285 -610 4310 -585
rect 4285 -655 4310 -630
rect 4285 -700 4310 -675
rect 4285 -750 4310 -725
rect 4345 -610 4370 -585
rect 4345 -655 4370 -630
rect 4345 -700 4370 -675
rect 4345 -750 4370 -725
rect 4405 -610 4430 -585
rect 4405 -655 4430 -630
rect 4405 -700 4430 -675
rect 4405 -750 4430 -725
rect 4465 -610 4490 -585
rect 4465 -655 4490 -630
rect 4465 -700 4490 -675
rect 4465 -750 4490 -725
rect 4525 -610 4550 -585
rect 4525 -655 4550 -630
rect 4525 -700 4550 -675
rect 4525 -750 4550 -725
rect 4585 -610 4610 -585
rect 4585 -655 4610 -630
rect 4585 -700 4610 -675
rect 4585 -750 4610 -725
rect 4645 -610 4670 -585
rect 4645 -655 4670 -630
rect 4645 -700 4670 -675
rect 4645 -750 4670 -725
rect 4705 -610 4730 -585
rect 4705 -655 4730 -630
rect 4705 -700 4730 -675
rect 4705 -750 4730 -725
rect 4765 -610 4790 -585
rect 4765 -655 4790 -630
rect 4765 -700 4790 -675
rect 4765 -750 4790 -725
rect 4825 -610 4850 -585
rect 4825 -655 4850 -630
rect 4825 -700 4850 -675
rect 4825 -750 4850 -725
rect 4885 -610 4910 -585
rect 4885 -655 4910 -630
rect 4885 -700 4910 -675
rect 4885 -750 4910 -725
rect 4945 -610 4970 -585
rect 4945 -655 4970 -630
rect 4945 -700 4970 -675
rect 4945 -750 4970 -725
rect 5005 -610 5030 -585
rect 5005 -655 5030 -630
rect 5005 -700 5030 -675
rect 5005 -750 5030 -725
rect 5065 -610 5090 -585
rect 5065 -655 5090 -630
rect 5065 -700 5090 -675
rect 5065 -750 5090 -725
rect 5125 -610 5150 -585
rect 5125 -655 5150 -630
rect 5125 -700 5150 -675
rect 5125 -750 5150 -725
rect 5185 -610 5210 -585
rect 5185 -655 5210 -630
rect 5185 -700 5210 -675
rect 5185 -750 5210 -725
rect 5245 -610 5270 -585
rect 5245 -655 5270 -630
rect 5245 -700 5270 -675
rect 5245 -750 5270 -725
rect 5305 -610 5330 -585
rect 5305 -655 5330 -630
rect 5305 -700 5330 -675
rect 5305 -750 5330 -725
rect 5365 -610 5390 -585
rect 5365 -655 5390 -630
rect 5365 -700 5390 -675
rect 5365 -750 5390 -725
rect 5425 -610 5450 -585
rect 5425 -655 5450 -630
rect 5425 -700 5450 -675
rect 5425 -750 5450 -725
rect 5485 -610 5510 -585
rect 5485 -655 5510 -630
rect 5485 -700 5510 -675
rect 5485 -750 5510 -725
rect 5545 -610 5570 -585
rect 5545 -655 5570 -630
rect 5545 -700 5570 -675
rect 5545 -750 5570 -725
rect 5605 -610 5630 -585
rect 5605 -655 5630 -630
rect 5605 -700 5630 -675
rect 5605 -750 5630 -725
rect 5665 -610 5690 -585
rect 5665 -655 5690 -630
rect 5665 -700 5690 -675
rect 5665 -750 5690 -725
rect 5725 -610 5750 -585
rect 5725 -655 5750 -630
rect 5725 -700 5750 -675
rect 5725 -750 5750 -725
rect 5785 -610 5810 -585
rect 5785 -655 5810 -630
rect 5785 -700 5810 -675
rect 5785 -750 5810 -725
rect 5845 -610 5870 -585
rect 5845 -655 5870 -630
rect 5845 -700 5870 -675
rect 5845 -750 5870 -725
rect 5905 -610 5930 -585
rect 5905 -655 5930 -630
rect 5905 -700 5930 -675
rect 5905 -750 5930 -725
rect 5965 -610 5990 -585
rect 5965 -655 5990 -630
rect 5965 -700 5990 -675
rect 5965 -750 5990 -725
rect 6025 -610 6050 -585
rect 6025 -655 6050 -630
rect 6025 -700 6050 -675
rect 6025 -750 6050 -725
rect 6085 -610 6110 -585
rect 6085 -655 6110 -630
rect 6085 -700 6110 -675
rect 6085 -750 6110 -725
rect 6145 -610 6170 -585
rect 6145 -655 6170 -630
rect 6145 -700 6170 -675
rect 6145 -750 6170 -725
rect 6205 -610 6230 -585
rect 6205 -655 6230 -630
rect 6205 -700 6230 -675
rect 6205 -750 6230 -725
rect 6265 -610 6290 -585
rect 6265 -655 6290 -630
rect 6265 -700 6290 -675
rect 6265 -750 6290 -725
rect 6325 -610 6350 -585
rect 6325 -655 6350 -630
rect 6325 -700 6350 -675
rect 6325 -750 6350 -725
rect 6385 -610 6410 -585
rect 6385 -655 6410 -630
rect 6385 -700 6410 -675
rect 6385 -750 6410 -725
rect 6445 -610 6470 -585
rect 6445 -655 6470 -630
rect 6445 -700 6470 -675
rect 6445 -750 6470 -725
rect 6505 -610 6530 -585
rect 6505 -655 6530 -630
rect 6505 -700 6530 -675
rect 6505 -750 6530 -725
rect 6565 -610 6590 -585
rect 6565 -655 6590 -630
rect 6565 -700 6590 -675
rect 6565 -750 6590 -725
rect 6625 -610 6650 -585
rect 6625 -655 6650 -630
rect 6625 -700 6650 -675
rect 6625 -750 6650 -725
rect 6685 -610 6710 -585
rect 6685 -655 6710 -630
rect 6685 -700 6710 -675
rect 6685 -750 6710 -725
rect 6745 -610 6770 -585
rect 6745 -655 6770 -630
rect 6745 -700 6770 -675
rect 6745 -750 6770 -725
rect 6805 -610 6830 -585
rect 6805 -655 6830 -630
rect 6805 -700 6830 -675
rect 6805 -750 6830 -725
rect 6865 -610 6890 -585
rect 6865 -655 6890 -630
rect 6865 -700 6890 -675
rect 6865 -750 6890 -725
rect 6925 -610 6950 -585
rect 6925 -655 6950 -630
rect 6925 -700 6950 -675
rect 6925 -750 6950 -725
rect 6985 -610 7010 -585
rect 6985 -655 7010 -630
rect 6985 -700 7010 -675
rect 6985 -750 7010 -725
rect 7045 -610 7070 -585
rect 7045 -655 7070 -630
rect 7045 -700 7070 -675
rect 7045 -750 7070 -725
rect 7105 -610 7130 -585
rect 7105 -655 7130 -630
rect 7105 -700 7130 -675
rect 7105 -750 7130 -725
rect 7165 -610 7190 -585
rect 7165 -655 7190 -630
rect 7165 -700 7190 -675
rect 7165 -750 7190 -725
rect 7225 -610 7250 -585
rect 7225 -655 7250 -630
rect 7225 -700 7250 -675
rect 7225 -750 7250 -725
rect 7285 -610 7310 -585
rect 7285 -655 7310 -630
rect 7285 -700 7310 -675
rect 7285 -750 7310 -725
rect 7345 -610 7370 -585
rect 7345 -655 7370 -630
rect 7345 -700 7370 -675
rect 7345 -750 7370 -725
rect 7405 -610 7430 -585
rect 7405 -655 7430 -630
rect 7405 -700 7430 -675
rect 7405 -750 7430 -725
rect 7465 -610 7490 -585
rect 7465 -655 7490 -630
rect 7465 -700 7490 -675
rect 7465 -750 7490 -725
rect 7525 -610 7550 -585
rect 7525 -655 7550 -630
rect 7525 -700 7550 -675
rect 7525 -750 7550 -725
rect 7585 -610 7610 -585
rect 7585 -655 7610 -630
rect 7585 -700 7610 -675
rect 7585 -750 7610 -725
rect 7645 -610 7670 -585
rect 7645 -655 7670 -630
rect 7645 -700 7670 -675
rect 7645 -750 7670 -725
rect 7705 -610 7730 -585
rect 7705 -655 7730 -630
rect 7705 -700 7730 -675
rect 7705 -750 7730 -725
rect 7765 -610 7790 -585
rect 7765 -655 7790 -630
rect 7765 -700 7790 -675
rect 7765 -750 7790 -725
rect 7825 -610 7850 -585
rect 7825 -655 7850 -630
rect 7825 -700 7850 -675
rect 7825 -750 7850 -725
rect 7885 -610 7910 -585
rect 7885 -655 7910 -630
rect 7885 -700 7910 -675
rect 7885 -750 7910 -725
rect 7945 -610 7970 -585
rect 7945 -655 7970 -630
rect 7945 -700 7970 -675
rect 7945 -750 7970 -725
rect 8005 -610 8030 -585
rect 8005 -655 8030 -630
rect 8005 -700 8030 -675
rect 8005 -750 8030 -725
rect 8065 -610 8090 -585
rect 8065 -655 8090 -630
rect 8065 -700 8090 -675
rect 8065 -750 8090 -725
rect 8125 -610 8150 -585
rect 8125 -655 8150 -630
rect 8125 -700 8150 -675
rect 8125 -750 8150 -725
rect 8185 -610 8210 -585
rect 8185 -655 8210 -630
rect 8185 -700 8210 -675
rect 8185 -750 8210 -725
rect 8245 -610 8270 -585
rect 8245 -655 8270 -630
rect 8245 -700 8270 -675
rect 8245 -750 8270 -725
rect 8305 -610 8330 -585
rect 8305 -655 8330 -630
rect 8305 -700 8330 -675
rect 8305 -750 8330 -725
rect 8365 -610 8390 -585
rect 8365 -655 8390 -630
rect 8365 -700 8390 -675
rect 8365 -750 8390 -725
rect 8425 -610 8450 -585
rect 8425 -655 8450 -630
rect 8425 -700 8450 -675
rect 8425 -750 8450 -725
rect 8485 -610 8510 -585
rect 8485 -655 8510 -630
rect 8485 -700 8510 -675
rect 8485 -750 8510 -725
rect 8545 -610 8570 -585
rect 8545 -655 8570 -630
rect 8545 -700 8570 -675
rect 8545 -750 8570 -725
rect 8605 -610 8630 -585
rect 8605 -655 8630 -630
rect 8605 -700 8630 -675
rect 8605 -750 8630 -725
rect 8665 -610 8690 -585
rect 8665 -655 8690 -630
rect 8665 -700 8690 -675
rect 8665 -750 8690 -725
rect 8725 -610 8750 -585
rect 8725 -655 8750 -630
rect 8725 -700 8750 -675
rect 8725 -750 8750 -725
rect 8785 -610 8810 -585
rect 8785 -655 8810 -630
rect 8785 -700 8810 -675
rect 8785 -750 8810 -725
rect 8845 -610 8870 -585
rect 8845 -655 8870 -630
rect 8845 -700 8870 -675
rect 8845 -750 8870 -725
rect 8905 -610 8930 -585
rect 8905 -655 8930 -630
rect 8905 -700 8930 -675
rect 8905 -750 8930 -725
rect 8965 -610 8990 -585
rect 8965 -655 8990 -630
rect 8965 -700 8990 -675
rect 8965 -750 8990 -725
rect 9025 -610 9050 -585
rect 9025 -655 9050 -630
rect 9025 -700 9050 -675
rect 9025 -750 9050 -725
rect 9085 -610 9110 -585
rect 9085 -655 9110 -630
rect 9085 -700 9110 -675
rect 9085 -750 9110 -725
rect 9145 -610 9170 -585
rect 9145 -655 9170 -630
rect 9145 -700 9170 -675
rect 9145 -750 9170 -725
rect 9205 -610 9230 -585
rect 9205 -655 9230 -630
rect 9205 -700 9230 -675
rect 9205 -750 9230 -725
rect 9265 -610 9290 -585
rect 9265 -655 9290 -630
rect 9265 -700 9290 -675
rect 9265 -750 9290 -725
rect 9325 -610 9350 -585
rect 9325 -655 9350 -630
rect 9325 -700 9350 -675
rect 9325 -750 9350 -725
rect 9385 -610 9410 -585
rect 9385 -655 9410 -630
rect 9385 -700 9410 -675
rect 9385 -750 9410 -725
rect 9445 -610 9470 -585
rect 9445 -655 9470 -630
rect 9445 -700 9470 -675
rect 9445 -750 9470 -725
rect 9505 -610 9530 -585
rect 9505 -655 9530 -630
rect 9505 -700 9530 -675
rect 9505 -750 9530 -725
rect 9565 -610 9590 -585
rect 9565 -655 9590 -630
rect 9565 -700 9590 -675
rect 9565 -750 9590 -725
rect 9625 -610 9650 -585
rect 9625 -655 9650 -630
rect 9625 -700 9650 -675
rect 9625 -750 9650 -725
rect 9685 -610 9710 -585
rect 9685 -655 9710 -630
rect 9685 -700 9710 -675
rect 9685 -750 9710 -725
rect 9745 -610 9770 -585
rect 9745 -655 9770 -630
rect 9745 -700 9770 -675
rect 9745 -750 9770 -725
rect 9805 -610 9830 -585
rect 9805 -655 9830 -630
rect 9805 -700 9830 -675
rect 9805 -750 9830 -725
rect 9865 -610 9890 -585
rect 9865 -655 9890 -630
rect 9865 -700 9890 -675
rect 9865 -750 9890 -725
rect 9925 -610 9950 -585
rect 9925 -655 9950 -630
rect 9925 -700 9950 -675
rect 9925 -750 9950 -725
rect 9985 -610 10010 -585
rect 9985 -655 10010 -630
rect 9985 -700 10010 -675
rect 9985 -750 10010 -725
rect 10045 -610 10070 -585
rect 10045 -655 10070 -630
rect 10045 -700 10070 -675
rect 10045 -750 10070 -725
rect 10105 -610 10130 -585
rect 10105 -655 10130 -630
rect 10105 -700 10130 -675
rect 10105 -750 10130 -725
rect 10165 -610 10190 -585
rect 10165 -655 10190 -630
rect 10165 -700 10190 -675
rect 10165 -750 10190 -725
rect 10225 -610 10250 -585
rect 10225 -655 10250 -630
rect 10225 -700 10250 -675
rect 10225 -750 10250 -725
rect 10285 -610 10310 -585
rect 10285 -655 10310 -630
rect 10285 -700 10310 -675
rect 10285 -750 10310 -725
rect 10345 -610 10370 -585
rect 10345 -655 10370 -630
rect 10345 -700 10370 -675
rect 10345 -750 10370 -725
rect 10405 -610 10430 -585
rect 10405 -655 10430 -630
rect 10405 -700 10430 -675
rect 10405 -750 10430 -725
rect 10465 -610 10490 -585
rect 10465 -655 10490 -630
rect 10465 -700 10490 -675
rect 10465 -750 10490 -725
rect 10525 -610 10550 -585
rect 10525 -655 10550 -630
rect 10525 -700 10550 -675
rect 10525 -750 10550 -725
rect 10585 -610 10610 -585
rect 10585 -655 10610 -630
rect 10585 -700 10610 -675
rect 10585 -750 10610 -725
rect 10645 -610 10670 -585
rect 10645 -655 10670 -630
rect 10645 -700 10670 -675
rect 10645 -750 10670 -725
rect 10705 -610 10730 -585
rect 10705 -655 10730 -630
rect 10705 -700 10730 -675
rect 10705 -750 10730 -725
rect 10765 -610 10790 -585
rect 10765 -655 10790 -630
rect 10765 -700 10790 -675
rect 10765 -750 10790 -725
rect 10825 -610 10850 -585
rect 10825 -655 10850 -630
rect 10825 -700 10850 -675
rect 10825 -750 10850 -725
rect 10885 -610 10910 -585
rect 10885 -655 10910 -630
rect 10885 -700 10910 -675
rect 10885 -750 10910 -725
rect 10945 -610 10970 -585
rect 10945 -655 10970 -630
rect 10945 -700 10970 -675
rect 10945 -750 10970 -725
rect 11005 -610 11030 -585
rect 11005 -655 11030 -630
rect 11005 -700 11030 -675
rect 11005 -750 11030 -725
rect 11065 -610 11090 -585
rect 11065 -655 11090 -630
rect 11065 -700 11090 -675
rect 11065 -750 11090 -725
rect 11125 -610 11150 -585
rect 11125 -655 11150 -630
rect 11125 -700 11150 -675
rect 11125 -750 11150 -725
rect 11185 -610 11210 -585
rect 11185 -655 11210 -630
rect 11185 -700 11210 -675
rect 11185 -750 11210 -725
rect 11245 -610 11270 -585
rect 11245 -655 11270 -630
rect 11245 -700 11270 -675
rect 11245 -750 11270 -725
rect 11305 -610 11330 -585
rect 11305 -655 11330 -630
rect 11305 -700 11330 -675
rect 11305 -750 11330 -725
rect 11365 -610 11390 -585
rect 11365 -655 11390 -630
rect 11365 -700 11390 -675
rect 11365 -750 11390 -725
rect 11425 -610 11450 -585
rect 11425 -655 11450 -630
rect 11425 -700 11450 -675
rect 11425 -750 11450 -725
rect 11485 -610 11510 -585
rect 11485 -655 11510 -630
rect 11485 -700 11510 -675
rect 11485 -750 11510 -725
rect 11545 -610 11570 -585
rect 11545 -655 11570 -630
rect 11545 -700 11570 -675
rect 11545 -750 11570 -725
rect 11605 -610 11630 -585
rect 11605 -655 11630 -630
rect 11605 -700 11630 -675
rect 11605 -750 11630 -725
rect 11665 -610 11690 -585
rect 11665 -655 11690 -630
rect 11665 -700 11690 -675
rect 11665 -750 11690 -725
rect 11725 -610 11750 -585
rect 11725 -655 11750 -630
rect 11725 -700 11750 -675
rect 11725 -750 11750 -725
rect 11785 -610 11810 -585
rect 11785 -655 11810 -630
rect 11785 -700 11810 -675
rect 11785 -750 11810 -725
rect 11845 -610 11870 -585
rect 11845 -655 11870 -630
rect 11845 -700 11870 -675
rect 11845 -750 11870 -725
rect 11905 -610 11930 -585
rect 11905 -655 11930 -630
rect 11905 -700 11930 -675
rect 11905 -750 11930 -725
rect 11965 -610 11990 -585
rect 11965 -655 11990 -630
rect 11965 -700 11990 -675
rect 11965 -750 11990 -725
rect 12025 -610 12050 -585
rect 12025 -655 12050 -630
rect 12025 -700 12050 -675
rect 12025 -750 12050 -725
rect 12085 -610 12110 -585
rect 12085 -655 12110 -630
rect 12085 -700 12110 -675
rect 12085 -750 12110 -725
rect 12145 -610 12170 -585
rect 12145 -655 12170 -630
rect 12145 -700 12170 -675
rect 12145 -750 12170 -725
rect 12205 -610 12230 -585
rect 12205 -655 12230 -630
rect 12205 -700 12230 -675
rect 12205 -750 12230 -725
rect 12265 -610 12290 -585
rect 12265 -655 12290 -630
rect 12265 -700 12290 -675
rect 12265 -750 12290 -725
rect 12325 -610 12350 -585
rect 12325 -655 12350 -630
rect 12325 -700 12350 -675
rect 12325 -750 12350 -725
rect 12385 -610 12410 -585
rect 12385 -655 12410 -630
rect 12385 -700 12410 -675
rect 12385 -750 12410 -725
rect 12445 -610 12470 -585
rect 12445 -655 12470 -630
rect 12445 -700 12470 -675
rect 12445 -750 12470 -725
rect 12505 -610 12530 -585
rect 12505 -655 12530 -630
rect 12505 -700 12530 -675
rect 12505 -750 12530 -725
rect 12565 -610 12590 -585
rect 12565 -655 12590 -630
rect 12565 -700 12590 -675
rect 12565 -750 12590 -725
rect 12625 -610 12650 -585
rect 12625 -655 12650 -630
rect 12625 -700 12650 -675
rect 12625 -750 12650 -725
rect 12685 -610 12710 -585
rect 12685 -655 12710 -630
rect 12685 -700 12710 -675
rect 12685 -750 12710 -725
rect 12745 -610 12770 -585
rect 12745 -655 12770 -630
rect 12745 -700 12770 -675
rect 12745 -750 12770 -725
rect 12805 -610 12830 -585
rect 12805 -655 12830 -630
rect 12805 -700 12830 -675
rect 12805 -750 12830 -725
rect 12865 -610 12890 -585
rect 12865 -655 12890 -630
rect 12865 -700 12890 -675
rect 12865 -750 12890 -725
rect 12925 -610 12950 -585
rect 12925 -655 12950 -630
rect 12925 -700 12950 -675
rect 12925 -750 12950 -725
rect 12985 -610 13010 -585
rect 12985 -655 13010 -630
rect 12985 -700 13010 -675
rect 12985 -750 13010 -725
rect 13045 -610 13070 -585
rect 13045 -655 13070 -630
rect 13045 -700 13070 -675
rect 13045 -750 13070 -725
rect 13105 -610 13130 -585
rect 13105 -655 13130 -630
rect 13105 -700 13130 -675
rect 13105 -750 13130 -725
rect 13165 -610 13190 -585
rect 13165 -655 13190 -630
rect 13165 -700 13190 -675
rect 13165 -750 13190 -725
rect 13225 -610 13250 -585
rect 13225 -655 13250 -630
rect 13225 -700 13250 -675
rect 13225 -750 13250 -725
rect 13285 -610 13310 -585
rect 13285 -655 13310 -630
rect 13285 -700 13310 -675
rect 13285 -750 13310 -725
rect 13345 -610 13370 -585
rect 13345 -655 13370 -630
rect 13345 -700 13370 -675
rect 13345 -750 13370 -725
rect 13405 -610 13430 -585
rect 13405 -655 13430 -630
rect 13405 -700 13430 -675
rect 13405 -750 13430 -725
rect 13465 -610 13490 -585
rect 13465 -655 13490 -630
rect 13465 -700 13490 -675
rect 13465 -750 13490 -725
rect 13525 -610 13550 -585
rect 13525 -655 13550 -630
rect 13525 -700 13550 -675
rect 13525 -750 13550 -725
rect 13585 -610 13610 -585
rect 13585 -655 13610 -630
rect 13585 -700 13610 -675
rect 13585 -750 13610 -725
rect 13645 -610 13670 -585
rect 13645 -655 13670 -630
rect 13645 -700 13670 -675
rect 13645 -750 13670 -725
rect 13705 -610 13730 -585
rect 13705 -655 13730 -630
rect 13705 -700 13730 -675
rect 13705 -750 13730 -725
rect 13765 -610 13790 -585
rect 13765 -655 13790 -630
rect 13765 -700 13790 -675
rect 13765 -750 13790 -725
rect 13825 -610 13850 -585
rect 13825 -655 13850 -630
rect 13825 -700 13850 -675
rect 13825 -750 13850 -725
rect 13885 -610 13910 -585
rect 13885 -655 13910 -630
rect 13885 -700 13910 -675
rect 13885 -750 13910 -725
rect 13945 -610 13970 -585
rect 13945 -655 13970 -630
rect 13945 -700 13970 -675
rect 13945 -750 13970 -725
rect 14005 -610 14030 -585
rect 14005 -655 14030 -630
rect 14005 -700 14030 -675
rect 14005 -750 14030 -725
rect 14065 -610 14090 -585
rect 14065 -655 14090 -630
rect 14065 -700 14090 -675
rect 14065 -750 14090 -725
rect 14125 -610 14150 -585
rect 14125 -655 14150 -630
rect 14125 -700 14150 -675
rect 14125 -750 14150 -725
rect 14185 -610 14210 -585
rect 14185 -655 14210 -630
rect 14185 -700 14210 -675
rect 14185 -750 14210 -725
rect 14245 -610 14270 -585
rect 14245 -655 14270 -630
rect 14245 -700 14270 -675
rect 14245 -750 14270 -725
rect 14305 -610 14330 -585
rect 14305 -655 14330 -630
rect 14305 -700 14330 -675
rect 14305 -750 14330 -725
rect 14365 -610 14390 -585
rect 14365 -655 14390 -630
rect 14365 -700 14390 -675
rect 14365 -750 14390 -725
rect 14425 -610 14450 -585
rect 14425 -655 14450 -630
rect 14425 -700 14450 -675
rect 14425 -750 14450 -725
rect 14485 -610 14510 -585
rect 14485 -655 14510 -630
rect 14485 -700 14510 -675
rect 14485 -750 14510 -725
rect 14545 -610 14570 -585
rect 14545 -655 14570 -630
rect 14545 -700 14570 -675
rect 14545 -750 14570 -725
rect 14605 -610 14630 -585
rect 14605 -655 14630 -630
rect 14605 -700 14630 -675
rect 14605 -750 14630 -725
rect 14665 -610 14690 -585
rect 14665 -655 14690 -630
rect 14665 -700 14690 -675
rect 14665 -750 14690 -725
rect 14725 -610 14750 -585
rect 14725 -655 14750 -630
rect 14725 -700 14750 -675
rect 14725 -750 14750 -725
rect 14785 -610 14810 -585
rect 14785 -655 14810 -630
rect 14785 -700 14810 -675
rect 14785 -750 14810 -725
rect 14845 -610 14870 -585
rect 14845 -655 14870 -630
rect 14845 -700 14870 -675
rect 14845 -750 14870 -725
rect 14905 -610 14930 -585
rect 14905 -655 14930 -630
rect 14905 -700 14930 -675
rect 14905 -750 14930 -725
rect 14965 -610 14990 -585
rect 14965 -655 14990 -630
rect 14965 -700 14990 -675
rect 14965 -750 14990 -725
rect 15025 -610 15050 -585
rect 15025 -655 15050 -630
rect 15025 -700 15050 -675
rect 15025 -750 15050 -725
rect 15085 -610 15110 -585
rect 15085 -655 15110 -630
rect 15085 -700 15110 -675
rect 15085 -750 15110 -725
rect 15145 -610 15170 -585
rect 15145 -655 15170 -630
rect 15145 -700 15170 -675
rect 15145 -750 15170 -725
rect 15205 -610 15230 -585
rect 15205 -655 15230 -630
rect 15205 -700 15230 -675
rect 15205 -750 15230 -725
rect 15265 -610 15290 -585
rect 15265 -655 15290 -630
rect 15265 -700 15290 -675
rect 15265 -750 15290 -725
rect 15325 -610 15350 -585
rect 15325 -655 15350 -630
rect 15325 -700 15350 -675
rect 15325 -750 15350 -725
rect 15385 -610 15410 -585
rect 15385 -655 15410 -630
rect 15385 -700 15410 -675
rect 15385 -750 15410 -725
rect 15445 -610 15470 -585
rect 15445 -655 15470 -630
rect 15445 -700 15470 -675
rect 15445 -750 15470 -725
rect 15505 -610 15530 -585
rect 15505 -655 15530 -630
rect 15505 -700 15530 -675
rect 15505 -750 15530 -725
rect 15565 -610 15590 -585
rect 15565 -655 15590 -630
rect 15565 -700 15590 -675
rect 15565 -750 15590 -725
rect 15625 -610 15650 -585
rect 15625 -655 15650 -630
rect 15625 -700 15650 -675
rect 15625 -750 15650 -725
rect 15685 -610 15710 -585
rect 15685 -655 15710 -630
rect 15685 -700 15710 -675
rect 15685 -750 15710 -725
rect 15745 -610 15770 -585
rect 15745 -655 15770 -630
rect 15745 -700 15770 -675
rect 15745 -750 15770 -725
rect 15805 -610 15830 -585
rect 15805 -655 15830 -630
rect 15805 -700 15830 -675
rect 15805 -750 15830 -725
rect 15865 -610 15890 -585
rect 15865 -655 15890 -630
rect 15865 -700 15890 -675
rect 15865 -750 15890 -725
rect 15925 -610 15950 -585
rect 15925 -655 15950 -630
rect 15925 -700 15950 -675
rect 15925 -750 15950 -725
rect 15985 -610 16010 -585
rect 15985 -655 16010 -630
rect 15985 -700 16010 -675
rect 15985 -750 16010 -725
rect 16045 -610 16070 -585
rect 16045 -655 16070 -630
rect 16045 -700 16070 -675
rect 16045 -750 16070 -725
rect 16105 -610 16130 -585
rect 16105 -655 16130 -630
rect 16105 -700 16130 -675
rect 16105 -750 16130 -725
rect 16165 -610 16190 -585
rect 16165 -655 16190 -630
rect 16165 -700 16190 -675
rect 16165 -750 16190 -725
rect 16225 -610 16250 -585
rect 16225 -655 16250 -630
rect 16225 -700 16250 -675
rect 16225 -750 16250 -725
rect 16285 -610 16310 -585
rect 16285 -655 16310 -630
rect 16285 -700 16310 -675
rect 16285 -750 16310 -725
rect 16345 -610 16370 -585
rect 16345 -655 16370 -630
rect 16345 -700 16370 -675
rect 16345 -750 16370 -725
rect 16405 -610 16430 -585
rect 16405 -655 16430 -630
rect 16405 -700 16430 -675
rect 16405 -750 16430 -725
rect 16465 -610 16490 -585
rect 16465 -655 16490 -630
rect 16465 -700 16490 -675
rect 16465 -750 16490 -725
rect 16525 -610 16550 -585
rect 16525 -655 16550 -630
rect 16525 -700 16550 -675
rect 16525 -750 16550 -725
rect 16585 -610 16610 -585
rect 16585 -655 16610 -630
rect 16585 -700 16610 -675
rect 16585 -750 16610 -725
rect 16645 -610 16670 -585
rect 16645 -655 16670 -630
rect 16645 -700 16670 -675
rect 16645 -750 16670 -725
rect 16705 -610 16730 -585
rect 16705 -655 16730 -630
rect 16705 -700 16730 -675
rect 16705 -750 16730 -725
rect 16765 -610 16790 -585
rect 16765 -655 16790 -630
rect 16765 -700 16790 -675
rect 16765 -750 16790 -725
rect 16825 -610 16850 -585
rect 16825 -655 16850 -630
rect 16825 -700 16850 -675
rect 16825 -750 16850 -725
rect 16885 -610 16910 -585
rect 16885 -655 16910 -630
rect 16885 -700 16910 -675
rect 16885 -750 16910 -725
rect 16945 -610 16970 -585
rect 16945 -655 16970 -630
rect 16945 -700 16970 -675
rect 16945 -750 16970 -725
rect 17005 -610 17030 -585
rect 17005 -655 17030 -630
rect 17005 -700 17030 -675
rect 17005 -750 17030 -725
rect 17065 -610 17090 -585
rect 17065 -655 17090 -630
rect 17065 -700 17090 -675
rect 17065 -750 17090 -725
rect 17125 -610 17150 -585
rect 17125 -655 17150 -630
rect 17125 -700 17150 -675
rect 17125 -750 17150 -725
rect 17185 -610 17210 -585
rect 17185 -655 17210 -630
rect 17185 -700 17210 -675
rect 17185 -750 17210 -725
rect 17245 -610 17270 -585
rect 17245 -655 17270 -630
rect 17245 -700 17270 -675
rect 17245 -750 17270 -725
rect 17305 -610 17330 -585
rect 17305 -655 17330 -630
rect 17305 -700 17330 -675
rect 17305 -750 17330 -725
rect 17365 -610 17390 -585
rect 17365 -655 17390 -630
rect 17365 -700 17390 -675
rect 17365 -750 17390 -725
rect 17425 -610 17450 -585
rect 17425 -655 17450 -630
rect 17425 -700 17450 -675
rect 17425 -750 17450 -725
rect 17485 -610 17510 -585
rect 17485 -655 17510 -630
rect 17485 -700 17510 -675
rect 17485 -750 17510 -725
rect 17545 -610 17570 -585
rect 17545 -655 17570 -630
rect 17545 -700 17570 -675
rect 17545 -750 17570 -725
rect 17605 -610 17630 -585
rect 17605 -655 17630 -630
rect 17605 -700 17630 -675
rect 17605 -750 17630 -725
rect 17665 -610 17690 -585
rect 17665 -655 17690 -630
rect 17665 -700 17690 -675
rect 17665 -750 17690 -725
rect 17725 -610 17750 -585
rect 17725 -655 17750 -630
rect 17725 -700 17750 -675
rect 17725 -750 17750 -725
rect 17785 -610 17810 -585
rect 17785 -655 17810 -630
rect 17785 -700 17810 -675
rect 17785 -750 17810 -725
rect 17845 -610 17870 -585
rect 17845 -655 17870 -630
rect 17845 -700 17870 -675
rect 17845 -750 17870 -725
rect 17905 -610 17930 -585
rect 17905 -655 17930 -630
rect 17905 -700 17930 -675
rect 17905 -750 17930 -725
rect 17965 -610 17990 -585
rect 17965 -655 17990 -630
rect 17965 -700 17990 -675
rect 17965 -750 17990 -725
rect 18025 -610 18050 -585
rect 18025 -655 18050 -630
rect 18025 -700 18050 -675
rect 18025 -750 18050 -725
rect 18085 -610 18110 -585
rect 18085 -655 18110 -630
rect 18085 -700 18110 -675
rect 18085 -750 18110 -725
rect 18145 -610 18170 -585
rect 18145 -655 18170 -630
rect 18145 -700 18170 -675
rect 18145 -750 18170 -725
rect 18205 -610 18230 -585
rect 18205 -655 18230 -630
rect 18205 -700 18230 -675
rect 18205 -750 18230 -725
rect 18265 -610 18290 -585
rect 18265 -655 18290 -630
rect 18265 -700 18290 -675
rect 18265 -750 18290 -725
rect 18325 -610 18350 -585
rect 18325 -655 18350 -630
rect 18325 -700 18350 -675
rect 18325 -750 18350 -725
rect 18385 -610 18410 -585
rect 18385 -655 18410 -630
rect 18385 -700 18410 -675
rect 18385 -750 18410 -725
rect 18445 -610 18470 -585
rect 18445 -655 18470 -630
rect 18445 -700 18470 -675
rect 18445 -750 18470 -725
rect 18505 -610 18530 -585
rect 18505 -655 18530 -630
rect 18505 -700 18530 -675
rect 18505 -750 18530 -725
rect 18565 -610 18590 -585
rect 18565 -655 18590 -630
rect 18565 -700 18590 -675
rect 18565 -750 18590 -725
rect 18625 -610 18650 -585
rect 18625 -655 18650 -630
rect 18625 -700 18650 -675
rect 18625 -750 18650 -725
rect 18685 -610 18710 -585
rect 18685 -655 18710 -630
rect 18685 -700 18710 -675
rect 18685 -750 18710 -725
rect 18745 -610 18770 -585
rect 18745 -655 18770 -630
rect 18745 -700 18770 -675
rect 18745 -750 18770 -725
rect 18805 -610 18830 -585
rect 18805 -655 18830 -630
rect 18805 -700 18830 -675
rect 18805 -750 18830 -725
rect 18865 -610 18890 -585
rect 18865 -655 18890 -630
rect 18865 -700 18890 -675
rect 18865 -750 18890 -725
rect 18925 -610 18950 -585
rect 18925 -655 18950 -630
rect 18925 -700 18950 -675
rect 18925 -750 18950 -725
rect 18985 -610 19010 -585
rect 18985 -655 19010 -630
rect 18985 -700 19010 -675
rect 18985 -750 19010 -725
rect 19045 -610 19070 -585
rect 19045 -655 19070 -630
rect 19045 -700 19070 -675
rect 19045 -750 19070 -725
rect 19105 -610 19130 -585
rect 19105 -655 19130 -630
rect 19105 -700 19130 -675
rect 19105 -750 19130 -725
rect 19165 -610 19190 -585
rect 19165 -655 19190 -630
rect 19165 -700 19190 -675
rect 19165 -750 19190 -725
rect 19225 -610 19250 -585
rect 19225 -655 19250 -630
rect 19225 -700 19250 -675
rect 19225 -750 19250 -725
rect 19285 -610 19310 -585
rect 19285 -655 19310 -630
rect 19285 -700 19310 -675
rect 19285 -750 19310 -725
rect 19345 -610 19370 -585
rect 19345 -655 19370 -630
rect 19345 -700 19370 -675
rect 19345 -750 19370 -725
rect 19405 -610 19430 -585
rect 19405 -655 19430 -630
rect 19405 -700 19430 -675
rect 19405 -750 19430 -725
rect 19465 -610 19490 -585
rect 19465 -655 19490 -630
rect 19465 -700 19490 -675
rect 19465 -750 19490 -725
rect 19525 -610 19550 -585
rect 19525 -655 19550 -630
rect 19525 -700 19550 -675
rect 19525 -750 19550 -725
rect 19585 -610 19610 -585
rect 19585 -655 19610 -630
rect 19585 -700 19610 -675
rect 19585 -750 19610 -725
rect 19645 -610 19670 -585
rect 19645 -655 19670 -630
rect 19645 -700 19670 -675
rect 19645 -750 19670 -725
rect 19705 -610 19730 -585
rect 19705 -655 19730 -630
rect 19705 -700 19730 -675
rect 19705 -750 19730 -725
rect 19765 -610 19790 -585
rect 19765 -655 19790 -630
rect 19765 -700 19790 -675
rect 19765 -750 19790 -725
rect 19825 -610 19850 -585
rect 19825 -655 19850 -630
rect 19825 -700 19850 -675
rect 19825 -750 19850 -725
rect 19885 -610 19910 -585
rect 19885 -655 19910 -630
rect 19885 -700 19910 -675
rect 19885 -750 19910 -725
rect 19945 -610 19970 -585
rect 19945 -655 19970 -630
rect 19945 -700 19970 -675
rect 19945 -750 19970 -725
rect 20005 -610 20030 -585
rect 20005 -655 20030 -630
rect 20005 -700 20030 -675
rect 20005 -750 20030 -725
rect 20065 -610 20090 -585
rect 20065 -655 20090 -630
rect 20065 -700 20090 -675
rect 20065 -750 20090 -725
rect 20125 -610 20150 -585
rect 20125 -655 20150 -630
rect 20125 -700 20150 -675
rect 20125 -750 20150 -725
rect 20185 -610 20210 -585
rect 20185 -655 20210 -630
rect 20185 -700 20210 -675
rect 20185 -750 20210 -725
rect 20245 -610 20270 -585
rect 20245 -655 20270 -630
rect 20245 -700 20270 -675
rect 20245 -750 20270 -725
rect 20305 -610 20330 -585
rect 20305 -655 20330 -630
rect 20305 -700 20330 -675
rect 20305 -750 20330 -725
rect 20365 -610 20390 -585
rect 20365 -655 20390 -630
rect 20365 -700 20390 -675
rect 20365 -750 20390 -725
rect 20425 -610 20450 -585
rect 20425 -655 20450 -630
rect 20425 -700 20450 -675
rect 20425 -750 20450 -725
rect 20485 -610 20510 -585
rect 20485 -655 20510 -630
rect 20485 -700 20510 -675
rect 20485 -750 20510 -725
rect 20545 -610 20570 -585
rect 20545 -655 20570 -630
rect 20545 -700 20570 -675
rect 20545 -750 20570 -725
rect 20605 -610 20630 -585
rect 20605 -655 20630 -630
rect 20605 -700 20630 -675
rect 20605 -750 20630 -725
rect 20665 -610 20690 -585
rect 20665 -655 20690 -630
rect 20665 -700 20690 -675
rect 20665 -750 20690 -725
rect 20725 -610 20750 -585
rect 20725 -655 20750 -630
rect 20725 -700 20750 -675
rect 20725 -750 20750 -725
rect 20785 -610 20810 -585
rect 20785 -655 20810 -630
rect 20785 -700 20810 -675
rect 20785 -750 20810 -725
rect 20845 -610 20870 -585
rect 20845 -655 20870 -630
rect 20845 -700 20870 -675
rect 20845 -750 20870 -725
rect 20905 -610 20930 -585
rect 20905 -655 20930 -630
rect 20905 -700 20930 -675
rect 20905 -750 20930 -725
rect 20965 -610 20990 -585
rect 20965 -655 20990 -630
rect 20965 -700 20990 -675
rect 20965 -750 20990 -725
rect 21025 -610 21050 -585
rect 21025 -655 21050 -630
rect 21025 -700 21050 -675
rect 21025 -750 21050 -725
rect 21085 -610 21110 -585
rect 21085 -655 21110 -630
rect 21085 -700 21110 -675
rect 21085 -750 21110 -725
rect 21145 -610 21170 -585
rect 21145 -655 21170 -630
rect 21145 -700 21170 -675
rect 21145 -750 21170 -725
rect 21205 -610 21230 -585
rect 21205 -655 21230 -630
rect 21205 -700 21230 -675
rect 21205 -750 21230 -725
rect 21265 -610 21290 -585
rect 21265 -655 21290 -630
rect 21265 -700 21290 -675
rect 21265 -750 21290 -725
rect 21325 -610 21350 -585
rect 21325 -655 21350 -630
rect 21325 -700 21350 -675
rect 21325 -750 21350 -725
rect 21385 -610 21410 -585
rect 21385 -655 21410 -630
rect 21385 -700 21410 -675
rect 21385 -750 21410 -725
rect 21445 -610 21470 -585
rect 21445 -655 21470 -630
rect 21445 -700 21470 -675
rect 21445 -750 21470 -725
rect 21505 -610 21530 -585
rect 21505 -655 21530 -630
rect 21505 -700 21530 -675
rect 21505 -750 21530 -725
rect 21565 -610 21590 -585
rect 21565 -655 21590 -630
rect 21565 -700 21590 -675
rect 21565 -750 21590 -725
rect 21625 -610 21650 -585
rect 21625 -655 21650 -630
rect 21625 -700 21650 -675
rect 21625 -750 21650 -725
rect 21685 -610 21710 -585
rect 21685 -655 21710 -630
rect 21685 -700 21710 -675
rect 21685 -750 21710 -725
rect 21745 -610 21770 -585
rect 21745 -655 21770 -630
rect 21745 -700 21770 -675
rect 21745 -750 21770 -725
rect 21805 -610 21830 -585
rect 21805 -655 21830 -630
rect 21805 -700 21830 -675
rect 21805 -750 21830 -725
rect 21865 -610 21890 -585
rect 21865 -655 21890 -630
rect 21865 -700 21890 -675
rect 21865 -750 21890 -725
rect 21925 -610 21950 -585
rect 21925 -655 21950 -630
rect 21925 -700 21950 -675
rect 21925 -750 21950 -725
rect 21985 -610 22010 -585
rect 21985 -655 22010 -630
rect 21985 -700 22010 -675
rect 21985 -750 22010 -725
rect 22045 -610 22070 -585
rect 22045 -655 22070 -630
rect 22045 -700 22070 -675
rect 22045 -750 22070 -725
rect 22105 -610 22130 -585
rect 22105 -655 22130 -630
rect 22105 -700 22130 -675
rect 22105 -750 22130 -725
rect 22165 -610 22190 -585
rect 22165 -655 22190 -630
rect 22165 -700 22190 -675
rect 22165 -750 22190 -725
rect 22225 -610 22250 -585
rect 22225 -655 22250 -630
rect 22225 -700 22250 -675
rect 22225 -750 22250 -725
rect 22285 -610 22310 -585
rect 22285 -655 22310 -630
rect 22285 -700 22310 -675
rect 22285 -750 22310 -725
rect 22345 -610 22370 -585
rect 22345 -655 22370 -630
rect 22345 -700 22370 -675
rect 22345 -750 22370 -725
rect 22405 -610 22430 -585
rect 22405 -655 22430 -630
rect 22405 -700 22430 -675
rect 22405 -750 22430 -725
rect 22465 -610 22490 -585
rect 22465 -655 22490 -630
rect 22465 -700 22490 -675
rect 22465 -750 22490 -725
rect 22525 -610 22550 -585
rect 22525 -655 22550 -630
rect 22525 -700 22550 -675
rect 22525 -750 22550 -725
rect 22585 -610 22610 -585
rect 22585 -655 22610 -630
rect 22585 -700 22610 -675
rect 22585 -750 22610 -725
rect 22645 -610 22670 -585
rect 22645 -655 22670 -630
rect 22645 -700 22670 -675
rect 22645 -750 22670 -725
rect 22705 -610 22730 -585
rect 22705 -655 22730 -630
rect 22705 -700 22730 -675
rect 22705 -750 22730 -725
rect 22765 -610 22790 -585
rect 22765 -655 22790 -630
rect 22765 -700 22790 -675
rect 22765 -750 22790 -725
rect 22825 -610 22850 -585
rect 22825 -655 22850 -630
rect 22825 -700 22850 -675
rect 22825 -750 22850 -725
rect 22885 -610 22910 -585
rect 22885 -655 22910 -630
rect 22885 -700 22910 -675
rect 22885 -750 22910 -725
rect 22945 -610 22970 -585
rect 22945 -655 22970 -630
rect 22945 -700 22970 -675
rect 22945 -750 22970 -725
rect 23005 -610 23030 -585
rect 23005 -655 23030 -630
rect 23005 -700 23030 -675
rect 23005 -750 23030 -725
rect 23065 -610 23090 -585
rect 23065 -655 23090 -630
rect 23065 -700 23090 -675
rect 23065 -750 23090 -725
rect 23125 -610 23150 -585
rect 23125 -655 23150 -630
rect 23125 -700 23150 -675
rect 23125 -750 23150 -725
rect 23185 -610 23210 -585
rect 23185 -655 23210 -630
rect 23185 -700 23210 -675
rect 23185 -750 23210 -725
rect 23245 -610 23270 -585
rect 23245 -655 23270 -630
rect 23245 -700 23270 -675
rect 23245 -750 23270 -725
rect 23305 -610 23330 -585
rect 23305 -655 23330 -630
rect 23305 -700 23330 -675
rect 23305 -750 23330 -725
rect 23365 -610 23390 -585
rect 23365 -655 23390 -630
rect 23365 -700 23390 -675
rect 23365 -750 23390 -725
rect 23425 -610 23450 -585
rect 23425 -655 23450 -630
rect 23425 -700 23450 -675
rect 23425 -750 23450 -725
rect 23485 -610 23510 -585
rect 23485 -655 23510 -630
rect 23485 -700 23510 -675
rect 23485 -750 23510 -725
rect 23545 -610 23570 -585
rect 23545 -655 23570 -630
rect 23545 -700 23570 -675
rect 23545 -750 23570 -725
rect 23605 -610 23630 -585
rect 23605 -655 23630 -630
rect 23605 -700 23630 -675
rect 23605 -750 23630 -725
rect 23665 -610 23690 -585
rect 23665 -655 23690 -630
rect 23665 -700 23690 -675
rect 23665 -750 23690 -725
rect 23725 -610 23750 -585
rect 23725 -655 23750 -630
rect 23725 -700 23750 -675
rect 23725 -750 23750 -725
rect 23785 -610 23810 -585
rect 23785 -655 23810 -630
rect 23785 -700 23810 -675
rect 23785 -750 23810 -725
rect 23845 -610 23870 -585
rect 23845 -655 23870 -630
rect 23845 -700 23870 -675
rect 23845 -750 23870 -725
rect 23905 -610 23930 -585
rect 23905 -655 23930 -630
rect 23905 -700 23930 -675
rect 23905 -750 23930 -725
rect 23965 -610 23990 -585
rect 23965 -655 23990 -630
rect 23965 -700 23990 -675
rect 23965 -750 23990 -725
rect 24025 -610 24050 -585
rect 24025 -655 24050 -630
rect 24025 -700 24050 -675
rect 24025 -750 24050 -725
rect 24085 -610 24110 -585
rect 24085 -655 24110 -630
rect 24085 -700 24110 -675
rect 24085 -750 24110 -725
rect 24145 -610 24170 -585
rect 24145 -655 24170 -630
rect 24145 -700 24170 -675
rect 24145 -750 24170 -725
rect 24205 -610 24230 -585
rect 24205 -655 24230 -630
rect 24205 -700 24230 -675
rect 24205 -750 24230 -725
rect 24265 -610 24290 -585
rect 24265 -655 24290 -630
rect 24265 -700 24290 -675
rect 24265 -750 24290 -725
rect 24325 -610 24350 -585
rect 24325 -655 24350 -630
rect 24325 -700 24350 -675
rect 24325 -750 24350 -725
rect 24385 -610 24410 -585
rect 24385 -655 24410 -630
rect 24385 -700 24410 -675
rect 24385 -750 24410 -725
rect 24445 -610 24470 -585
rect 24445 -655 24470 -630
rect 24445 -700 24470 -675
rect 24445 -750 24470 -725
rect 24505 -610 24530 -585
rect 24505 -655 24530 -630
rect 24505 -700 24530 -675
rect 24505 -750 24530 -725
rect 24565 -610 24590 -585
rect 24565 -655 24590 -630
rect 24565 -700 24590 -675
rect 24565 -750 24590 -725
rect 24625 -610 24650 -585
rect 24625 -655 24650 -630
rect 24625 -700 24650 -675
rect 24625 -750 24650 -725
rect 24685 -610 24710 -585
rect 24685 -655 24710 -630
rect 24685 -700 24710 -675
rect 24685 -750 24710 -725
rect 24745 -610 24770 -585
rect 24745 -655 24770 -630
rect 24745 -700 24770 -675
rect 24745 -750 24770 -725
rect 24805 -610 24830 -585
rect 24805 -655 24830 -630
rect 24805 -700 24830 -675
rect 24805 -750 24830 -725
rect 24865 -610 24890 -585
rect 24865 -655 24890 -630
rect 24865 -700 24890 -675
rect 24865 -750 24890 -725
rect 24925 -610 24950 -585
rect 24925 -655 24950 -630
rect 24925 -700 24950 -675
rect 24925 -750 24950 -725
rect 24985 -610 25010 -585
rect 24985 -655 25010 -630
rect 24985 -700 25010 -675
rect 24985 -750 25010 -725
rect 25045 -610 25070 -585
rect 25045 -655 25070 -630
rect 25045 -700 25070 -675
rect 25045 -750 25070 -725
rect 25105 -610 25130 -585
rect 25105 -655 25130 -630
rect 25105 -700 25130 -675
rect 25105 -750 25130 -725
rect 25165 -610 25190 -585
rect 25165 -655 25190 -630
rect 25165 -700 25190 -675
rect 25165 -750 25190 -725
rect 25225 -610 25250 -585
rect 25225 -655 25250 -630
rect 25225 -700 25250 -675
rect 25225 -750 25250 -725
rect 25285 -610 25310 -585
rect 25285 -655 25310 -630
rect 25285 -700 25310 -675
rect 25285 -750 25310 -725
rect 25345 -610 25370 -585
rect 25345 -655 25370 -630
rect 25345 -700 25370 -675
rect 25345 -750 25370 -725
rect 25405 -610 25430 -585
rect 25405 -655 25430 -630
rect 25405 -700 25430 -675
rect 25405 -750 25430 -725
rect 25465 -610 25490 -585
rect 25465 -655 25490 -630
rect 25465 -700 25490 -675
rect 25465 -750 25490 -725
rect 25525 -610 25550 -585
rect 25525 -655 25550 -630
rect 25525 -700 25550 -675
rect 25525 -750 25550 -725
rect 25585 -610 25610 -585
rect 25585 -655 25610 -630
rect 25585 -700 25610 -675
rect 25585 -750 25610 -725
rect 25645 -610 25670 -585
rect 25645 -655 25670 -630
rect 25645 -700 25670 -675
rect 25645 -750 25670 -725
rect 25705 -610 25730 -585
rect 25705 -655 25730 -630
rect 25705 -700 25730 -675
rect 25705 -750 25730 -725
rect 25765 -610 25790 -585
rect 25765 -655 25790 -630
rect 25765 -700 25790 -675
rect 25765 -750 25790 -725
rect 25825 -610 25850 -585
rect 25825 -655 25850 -630
rect 25825 -700 25850 -675
rect 25825 -750 25850 -725
rect 25885 -610 25910 -585
rect 25885 -655 25910 -630
rect 25885 -700 25910 -675
rect 25885 -750 25910 -725
rect 25945 -610 25970 -585
rect 25945 -655 25970 -630
rect 25945 -700 25970 -675
rect 25945 -750 25970 -725
rect 26005 -610 26030 -585
rect 26005 -655 26030 -630
rect 26005 -700 26030 -675
rect 26005 -750 26030 -725
rect 26065 -610 26090 -585
rect 26065 -655 26090 -630
rect 26065 -700 26090 -675
rect 26065 -750 26090 -725
rect 26125 -610 26150 -585
rect 26125 -655 26150 -630
rect 26125 -700 26150 -675
rect 26125 -750 26150 -725
rect 26185 -610 26210 -585
rect 26185 -655 26210 -630
rect 26185 -700 26210 -675
rect 26185 -750 26210 -725
rect 26245 -610 26270 -585
rect 26245 -655 26270 -630
rect 26245 -700 26270 -675
rect 26245 -750 26270 -725
rect 26305 -610 26330 -585
rect 26305 -655 26330 -630
rect 26305 -700 26330 -675
rect 26305 -750 26330 -725
rect 26365 -610 26390 -585
rect 26365 -655 26390 -630
rect 26365 -700 26390 -675
rect 26365 -750 26390 -725
rect 26425 -610 26450 -585
rect 26425 -655 26450 -630
rect 26425 -700 26450 -675
rect 26425 -750 26450 -725
rect 26485 -610 26510 -585
rect 26485 -655 26510 -630
rect 26485 -700 26510 -675
rect 26485 -750 26510 -725
rect 26545 -610 26570 -585
rect 26545 -655 26570 -630
rect 26545 -700 26570 -675
rect 26545 -750 26570 -725
rect 26605 -610 26630 -585
rect 26605 -655 26630 -630
rect 26605 -700 26630 -675
rect 26605 -750 26630 -725
rect 26665 -610 26690 -585
rect 26665 -655 26690 -630
rect 26665 -700 26690 -675
rect 26665 -750 26690 -725
rect 26725 -610 26750 -585
rect 26725 -655 26750 -630
rect 26725 -700 26750 -675
rect 26725 -750 26750 -725
rect 26785 -610 26810 -585
rect 26785 -655 26810 -630
rect 26785 -700 26810 -675
rect 26785 -750 26810 -725
rect 26845 -610 26870 -585
rect 26845 -655 26870 -630
rect 26845 -700 26870 -675
rect 26845 -750 26870 -725
rect 26905 -610 26930 -585
rect 26905 -655 26930 -630
rect 26905 -700 26930 -675
rect 26905 -750 26930 -725
rect 26965 -610 26990 -585
rect 26965 -655 26990 -630
rect 26965 -700 26990 -675
rect 26965 -750 26990 -725
rect 27025 -610 27050 -585
rect 27025 -655 27050 -630
rect 27025 -700 27050 -675
rect 27025 -750 27050 -725
rect 27085 -610 27110 -585
rect 27085 -655 27110 -630
rect 27085 -700 27110 -675
rect 27085 -750 27110 -725
rect 27145 -610 27170 -585
rect 27145 -655 27170 -630
rect 27145 -700 27170 -675
rect 27145 -750 27170 -725
rect 27205 -610 27230 -585
rect 27205 -655 27230 -630
rect 27205 -700 27230 -675
rect 27205 -750 27230 -725
rect 27265 -610 27290 -585
rect 27265 -655 27290 -630
rect 27265 -700 27290 -675
rect 27265 -750 27290 -725
rect 27325 -610 27350 -585
rect 27325 -655 27350 -630
rect 27325 -700 27350 -675
rect 27325 -750 27350 -725
rect 27385 -610 27410 -585
rect 27385 -655 27410 -630
rect 27385 -700 27410 -675
rect 27385 -750 27410 -725
rect 27445 -610 27470 -585
rect 27445 -655 27470 -630
rect 27445 -700 27470 -675
rect 27445 -750 27470 -725
rect 27505 -610 27530 -585
rect 27505 -655 27530 -630
rect 27505 -700 27530 -675
rect 27505 -750 27530 -725
rect 27565 -610 27590 -585
rect 27565 -655 27590 -630
rect 27565 -700 27590 -675
rect 27565 -750 27590 -725
rect 27625 -610 27650 -585
rect 27625 -655 27650 -630
rect 27625 -700 27650 -675
rect 27625 -750 27650 -725
rect 27685 -610 27710 -585
rect 27685 -655 27710 -630
rect 27685 -700 27710 -675
rect 27685 -750 27710 -725
rect 27745 -610 27770 -585
rect 27745 -655 27770 -630
rect 27745 -700 27770 -675
rect 27745 -750 27770 -725
rect 27805 -610 27830 -585
rect 27805 -655 27830 -630
rect 27805 -700 27830 -675
rect 27805 -750 27830 -725
rect 27865 -610 27890 -585
rect 27865 -655 27890 -630
rect 27865 -700 27890 -675
rect 27865 -750 27890 -725
rect 27925 -610 27950 -585
rect 27925 -655 27950 -630
rect 27925 -700 27950 -675
rect 27925 -750 27950 -725
rect 27985 -610 28010 -585
rect 27985 -655 28010 -630
rect 27985 -700 28010 -675
rect 27985 -750 28010 -725
rect 28045 -610 28070 -585
rect 28045 -655 28070 -630
rect 28045 -700 28070 -675
rect 28045 -750 28070 -725
rect 28105 -610 28130 -585
rect 28105 -655 28130 -630
rect 28105 -700 28130 -675
rect 28105 -750 28130 -725
rect 28165 -610 28190 -585
rect 28165 -655 28190 -630
rect 28165 -700 28190 -675
rect 28165 -750 28190 -725
rect 28225 -610 28250 -585
rect 28225 -655 28250 -630
rect 28225 -700 28250 -675
rect 28225 -750 28250 -725
rect 28285 -610 28310 -585
rect 28285 -655 28310 -630
rect 28285 -700 28310 -675
rect 28285 -750 28310 -725
rect 28345 -610 28370 -585
rect 28345 -655 28370 -630
rect 28345 -700 28370 -675
rect 28345 -750 28370 -725
rect 28405 -610 28430 -585
rect 28405 -655 28430 -630
rect 28405 -700 28430 -675
rect 28405 -750 28430 -725
rect 28465 -610 28490 -585
rect 28465 -655 28490 -630
rect 28465 -700 28490 -675
rect 28465 -750 28490 -725
rect 28525 -610 28550 -585
rect 28525 -655 28550 -630
rect 28525 -700 28550 -675
rect 28525 -750 28550 -725
rect 28585 -610 28610 -585
rect 28585 -655 28610 -630
rect 28585 -700 28610 -675
rect 28585 -750 28610 -725
rect 28645 -610 28670 -585
rect 28645 -655 28670 -630
rect 28645 -700 28670 -675
rect 28645 -750 28670 -725
rect 28705 -610 28730 -585
rect 28705 -655 28730 -630
rect 28705 -700 28730 -675
rect 28705 -750 28730 -725
rect 28765 -610 28790 -585
rect 28765 -655 28790 -630
rect 28765 -700 28790 -675
rect 28765 -750 28790 -725
rect 28825 -610 28850 -585
rect 28825 -655 28850 -630
rect 28825 -700 28850 -675
rect 28825 -750 28850 -725
rect 28885 -610 28910 -585
rect 28885 -655 28910 -630
rect 28885 -700 28910 -675
rect 28885 -750 28910 -725
rect 28945 -610 28970 -585
rect 28945 -655 28970 -630
rect 28945 -700 28970 -675
rect 28945 -750 28970 -725
rect 29005 -610 29030 -585
rect 29005 -655 29030 -630
rect 29005 -700 29030 -675
rect 29005 -750 29030 -725
rect 29065 -610 29090 -585
rect 29065 -655 29090 -630
rect 29065 -700 29090 -675
rect 29065 -750 29090 -725
rect 29125 -610 29150 -585
rect 29125 -655 29150 -630
rect 29125 -700 29150 -675
rect 29125 -750 29150 -725
rect 29185 -610 29210 -585
rect 29185 -655 29210 -630
rect 29185 -700 29210 -675
rect 29185 -750 29210 -725
rect 29245 -610 29270 -585
rect 29245 -655 29270 -630
rect 29245 -700 29270 -675
rect 29245 -750 29270 -725
rect 29305 -610 29330 -585
rect 29305 -655 29330 -630
rect 29305 -700 29330 -675
rect 29305 -750 29330 -725
rect 29365 -610 29390 -585
rect 29365 -655 29390 -630
rect 29365 -700 29390 -675
rect 29365 -750 29390 -725
rect 29425 -610 29450 -585
rect 29425 -655 29450 -630
rect 29425 -700 29450 -675
rect 29425 -750 29450 -725
rect 29485 -610 29510 -585
rect 29485 -655 29510 -630
rect 29485 -700 29510 -675
rect 29485 -750 29510 -725
rect 29545 -610 29570 -585
rect 29545 -655 29570 -630
rect 29545 -700 29570 -675
rect 29545 -750 29570 -725
rect 29605 -610 29630 -585
rect 29605 -655 29630 -630
rect 29605 -700 29630 -675
rect 29605 -750 29630 -725
rect 29665 -610 29690 -585
rect 29665 -655 29690 -630
rect 29665 -700 29690 -675
rect 29665 -750 29690 -725
rect 29725 -610 29750 -585
rect 29725 -655 29750 -630
rect 29725 -700 29750 -675
rect 29725 -750 29750 -725
rect 29785 -610 29810 -585
rect 29785 -655 29810 -630
rect 29785 -700 29810 -675
rect 29785 -750 29810 -725
rect 29845 -610 29870 -585
rect 29845 -655 29870 -630
rect 29845 -700 29870 -675
rect 29845 -750 29870 -725
rect 29905 -610 29930 -585
rect 29905 -655 29930 -630
rect 29905 -700 29930 -675
rect 29905 -750 29930 -725
rect 29965 -610 29990 -585
rect 29965 -655 29990 -630
rect 29965 -700 29990 -675
rect 29965 -750 29990 -725
rect 30025 -610 30050 -585
rect 30025 -655 30050 -630
rect 30025 -700 30050 -675
rect 30025 -750 30050 -725
rect 30085 -610 30110 -585
rect 30085 -655 30110 -630
rect 30085 -700 30110 -675
rect 30085 -750 30110 -725
rect 30145 -610 30170 -585
rect 30145 -655 30170 -630
rect 30145 -700 30170 -675
rect 30145 -750 30170 -725
rect 30205 -610 30230 -585
rect 30205 -655 30230 -630
rect 30205 -700 30230 -675
rect 30205 -750 30230 -725
rect 30265 -610 30290 -585
rect 30265 -655 30290 -630
rect 30265 -700 30290 -675
rect 30265 -750 30290 -725
rect 30325 -610 30350 -585
rect 30325 -655 30350 -630
rect 30325 -700 30350 -675
rect 30325 -750 30350 -725
rect 30385 -610 30410 -585
rect 30385 -655 30410 -630
rect 30385 -700 30410 -675
rect 30385 -750 30410 -725
rect 30445 -610 30470 -585
rect 30445 -655 30470 -630
rect 30445 -700 30470 -675
rect 30445 -750 30470 -725
rect 30505 -610 30530 -585
rect 30505 -655 30530 -630
rect 30505 -700 30530 -675
rect 30505 -750 30530 -725
rect 30565 -610 30590 -585
rect 30565 -655 30590 -630
rect 30565 -700 30590 -675
rect 30565 -750 30590 -725
rect 30625 -610 30650 -585
rect 30625 -655 30650 -630
rect 30625 -700 30650 -675
rect 30625 -750 30650 -725
rect 30685 -610 30710 -585
rect 30685 -655 30710 -630
rect 30685 -700 30710 -675
rect 30685 -750 30710 -725
rect 85 -850 110 -825
rect 325 -850 350 -825
rect 565 -850 590 -825
rect 1045 -850 1070 -825
rect 1285 -850 1310 -825
rect 1525 -850 1550 -825
rect 1765 -850 1790 -825
rect 2005 -850 2030 -825
rect 2245 -850 2270 -825
rect 2485 -850 2510 -825
rect 2725 -850 2750 -825
rect 3205 -850 3230 -825
rect 3445 -850 3470 -825
rect 3685 -850 3710 -825
rect 3925 -850 3950 -825
rect 4165 -850 4190 -825
rect 4405 -850 4430 -825
rect 4645 -850 4670 -825
rect 4885 -850 4910 -825
rect 5365 -850 5390 -825
rect 5605 -850 5630 -825
rect 5845 -850 5870 -825
rect 6085 -850 6110 -825
rect 6325 -850 6350 -825
rect 6565 -850 6590 -825
rect 6805 -850 6830 -825
rect 7045 -850 7070 -825
rect 7525 -850 7550 -825
rect 7765 -850 7790 -825
rect 8005 -850 8030 -825
rect 8245 -850 8270 -825
rect 8485 -850 8510 -825
rect 8725 -850 8750 -825
rect 8965 -850 8990 -825
rect 9205 -850 9230 -825
rect 9685 -850 9710 -825
rect 9925 -850 9950 -825
rect 10165 -850 10190 -825
rect 10405 -850 10430 -825
rect 10645 -850 10670 -825
rect 10885 -850 10910 -825
rect 11125 -850 11150 -825
rect 11365 -850 11390 -825
rect 11845 -850 11870 -825
rect 12085 -850 12110 -825
rect 12325 -850 12350 -825
rect 12565 -850 12590 -825
rect 12805 -850 12830 -825
rect 13045 -850 13070 -825
rect 13285 -850 13310 -825
rect 13525 -850 13550 -825
rect 14005 -850 14030 -825
rect 14245 -850 14270 -825
rect 14485 -850 14510 -825
rect 14725 -850 14750 -825
rect 14965 -850 14990 -825
rect 15205 -850 15230 -825
rect 15445 -850 15470 -825
rect 15685 -850 15710 -825
rect 16165 -850 16190 -825
rect 16405 -850 16430 -825
rect 16645 -850 16670 -825
rect 16885 -850 16910 -825
rect 17125 -850 17150 -825
rect 17365 -850 17390 -825
rect 17605 -850 17630 -825
rect 17845 -850 17870 -825
rect 18325 -850 18350 -825
rect 18565 -850 18590 -825
rect 18805 -850 18830 -825
rect 19045 -850 19070 -825
rect 19285 -850 19310 -825
rect 19525 -850 19550 -825
rect 19765 -850 19790 -825
rect 20005 -850 20030 -825
rect 20485 -850 20510 -825
rect 20725 -850 20750 -825
rect 20965 -850 20990 -825
rect 21205 -850 21230 -825
rect 21445 -850 21470 -825
rect 21685 -850 21710 -825
rect 21925 -850 21950 -825
rect 22165 -850 22190 -825
rect 22645 -850 22670 -825
rect 22885 -850 22910 -825
rect 23125 -850 23150 -825
rect 23365 -850 23390 -825
rect 23605 -850 23630 -825
rect 23845 -850 23870 -825
rect 24085 -850 24110 -825
rect 24565 -850 24590 -825
rect 24805 -850 24830 -825
rect 25045 -850 25070 -825
rect 25285 -850 25310 -825
rect 25525 -850 25550 -825
rect 25765 -850 25790 -825
rect 26005 -850 26030 -825
rect 26485 -850 26510 -825
rect 26725 -850 26750 -825
rect 26965 -850 26990 -825
rect 27205 -850 27230 -825
rect 27445 -850 27470 -825
rect 27685 -850 27710 -825
rect 27925 -850 27950 -825
rect 28405 -850 28430 -825
rect 28645 -850 28670 -825
rect 28885 -850 28910 -825
rect 29125 -850 29150 -825
rect 29365 -850 29390 -825
rect 29605 -850 29630 -825
rect 30085 -850 30110 -825
rect 30325 -850 30350 -825
rect 30565 -850 30590 -825
<< psubdiff >>
rect -250 475 -120 490
rect -250 375 -235 475
rect -135 375 -120 475
rect -250 360 -120 375
rect 300 475 430 490
rect 300 375 315 475
rect 415 375 430 475
rect 300 360 430 375
rect 850 475 980 490
rect 850 375 865 475
rect 965 375 980 475
rect 850 360 980 375
rect 1400 475 1530 490
rect 1400 375 1415 475
rect 1515 375 1530 475
rect 1400 360 1530 375
rect 1950 475 2080 490
rect 1950 375 1965 475
rect 2065 375 2080 475
rect 1950 360 2080 375
rect 2500 475 2630 490
rect 2500 375 2515 475
rect 2615 375 2630 475
rect 2500 360 2630 375
rect 3050 475 3180 490
rect 3050 375 3065 475
rect 3165 375 3180 475
rect 3050 360 3180 375
rect 3600 475 3730 490
rect 3600 375 3615 475
rect 3715 375 3730 475
rect 3600 360 3730 375
rect 4150 475 4280 490
rect 4150 375 4165 475
rect 4265 375 4280 475
rect 4150 360 4280 375
rect 4700 475 4830 490
rect 4700 375 4715 475
rect 4815 375 4830 475
rect 4700 360 4830 375
rect 5250 475 5380 490
rect 5250 375 5265 475
rect 5365 375 5380 475
rect 5250 360 5380 375
rect 5800 475 5930 490
rect 5800 375 5815 475
rect 5915 375 5930 475
rect 5800 360 5930 375
rect 6350 475 6480 490
rect 6350 375 6365 475
rect 6465 375 6480 475
rect 6350 360 6480 375
rect 6900 475 7030 490
rect 6900 375 6915 475
rect 7015 375 7030 475
rect 6900 360 7030 375
rect 7450 475 7580 490
rect 7450 375 7465 475
rect 7565 375 7580 475
rect 7450 360 7580 375
rect 8000 475 8130 490
rect 8000 375 8015 475
rect 8115 375 8130 475
rect 8000 360 8130 375
rect 8550 475 8680 490
rect 8550 375 8565 475
rect 8665 375 8680 475
rect 8550 360 8680 375
rect 9100 475 9230 490
rect 9100 375 9115 475
rect 9215 375 9230 475
rect 9100 360 9230 375
rect 9650 475 9780 490
rect 9650 375 9665 475
rect 9765 375 9780 475
rect 9650 360 9780 375
rect 10200 475 10330 490
rect 10200 375 10215 475
rect 10315 375 10330 475
rect 10200 360 10330 375
rect 10750 475 10880 490
rect 10750 375 10765 475
rect 10865 375 10880 475
rect 10750 360 10880 375
rect 11300 475 11430 490
rect 11300 375 11315 475
rect 11415 375 11430 475
rect 11300 360 11430 375
rect 11850 475 11980 490
rect 11850 375 11865 475
rect 11965 375 11980 475
rect 11850 360 11980 375
rect 12400 475 12530 490
rect 12400 375 12415 475
rect 12515 375 12530 475
rect 12400 360 12530 375
rect 12950 475 13080 490
rect 12950 375 12965 475
rect 13065 375 13080 475
rect 12950 360 13080 375
rect 13500 475 13630 490
rect 13500 375 13515 475
rect 13615 375 13630 475
rect 13500 360 13630 375
rect 14050 475 14180 490
rect 14050 375 14065 475
rect 14165 375 14180 475
rect 14050 360 14180 375
rect 14600 475 14730 490
rect 14600 375 14615 475
rect 14715 375 14730 475
rect 14600 360 14730 375
rect 15150 475 15280 490
rect 15150 375 15165 475
rect 15265 375 15280 475
rect 15150 360 15280 375
rect 15700 475 15830 490
rect 15700 375 15715 475
rect 15815 375 15830 475
rect 15700 360 15830 375
rect 16250 475 16380 490
rect 16250 375 16265 475
rect 16365 375 16380 475
rect 16250 360 16380 375
rect 16800 475 16930 490
rect 16800 375 16815 475
rect 16915 375 16930 475
rect 16800 360 16930 375
rect 17350 475 17480 490
rect 17350 375 17365 475
rect 17465 375 17480 475
rect 17350 360 17480 375
rect 17900 475 18030 490
rect 17900 375 17915 475
rect 18015 375 18030 475
rect 17900 360 18030 375
rect 18450 475 18580 490
rect 18450 375 18465 475
rect 18565 375 18580 475
rect 18450 360 18580 375
rect 19000 475 19130 490
rect 19000 375 19015 475
rect 19115 375 19130 475
rect 19000 360 19130 375
rect 19550 475 19680 490
rect 19550 375 19565 475
rect 19665 375 19680 475
rect 19550 360 19680 375
rect 20100 475 20230 490
rect 20100 375 20115 475
rect 20215 375 20230 475
rect 20100 360 20230 375
rect 20650 475 20780 490
rect 20650 375 20665 475
rect 20765 375 20780 475
rect 20650 360 20780 375
rect 21200 475 21330 490
rect 21200 375 21215 475
rect 21315 375 21330 475
rect 21200 360 21330 375
rect 21530 265 21660 280
rect 21530 165 21545 265
rect 21645 165 21660 265
rect 21530 150 21660 165
rect -455 -5 -325 10
rect -455 -105 -440 -5
rect -340 -105 -325 -5
rect 21750 -5 21880 10
rect -455 -120 -325 -105
rect 21750 -105 21765 -5
rect 21865 -105 21880 -5
rect 21750 -120 21880 -105
rect 22300 -5 22430 10
rect 22300 -105 22315 -5
rect 22415 -105 22430 -5
rect 22300 -120 22430 -105
rect 22850 -5 22980 10
rect 22850 -105 22865 -5
rect 22965 -105 22980 -5
rect 22850 -120 22980 -105
rect 23400 -5 23530 10
rect 23400 -105 23415 -5
rect 23515 -105 23530 -5
rect 23400 -120 23530 -105
rect 23950 -5 24080 10
rect 23950 -105 23965 -5
rect 24065 -105 24080 -5
rect 23950 -120 24080 -105
rect 24500 -5 24630 10
rect 24500 -105 24515 -5
rect 24615 -105 24630 -5
rect 24500 -120 24630 -105
rect 25050 -5 25180 10
rect 25050 -105 25065 -5
rect 25165 -105 25180 -5
rect 25050 -120 25180 -105
rect 25600 -5 25730 10
rect 25600 -105 25615 -5
rect 25715 -105 25730 -5
rect 25600 -120 25730 -105
rect 26150 -5 26280 10
rect 26150 -105 26165 -5
rect 26265 -105 26280 -5
rect 26150 -120 26280 -105
rect 26700 -5 26830 10
rect 26700 -105 26715 -5
rect 26815 -105 26830 -5
rect 26700 -120 26830 -105
rect 27250 -5 27380 10
rect 27250 -105 27265 -5
rect 27365 -105 27380 -5
rect 27250 -120 27380 -105
rect 27800 -5 27930 10
rect 27800 -105 27815 -5
rect 27915 -105 27930 -5
rect 27800 -120 27930 -105
rect 28350 -5 28480 10
rect 28350 -105 28365 -5
rect 28465 -105 28480 -5
rect 28350 -120 28480 -105
rect 28900 -5 29030 10
rect 28900 -105 28915 -5
rect 29015 -105 29030 -5
rect 28900 -120 29030 -105
rect 29450 -5 29580 10
rect 29450 -105 29465 -5
rect 29565 -105 29580 -5
rect 29450 -120 29580 -105
rect 30000 -5 30130 10
rect 30000 -105 30015 -5
rect 30115 -105 30130 -5
rect 30000 -120 30130 -105
rect 30550 -5 30680 10
rect 30550 -105 30565 -5
rect 30665 -105 30680 -5
rect 30550 -120 30680 -105
rect 1620 -200 1690 -185
rect 1620 -240 1635 -200
rect 1675 -240 1690 -200
rect 1620 -255 1690 -240
rect 4045 -195 4115 -180
rect 4045 -235 4060 -195
rect 4100 -235 4115 -195
rect 4045 -250 4115 -235
rect 6440 -220 6510 -205
rect 6440 -260 6455 -220
rect 6495 -260 6510 -220
rect 6440 -275 6510 -260
rect 7865 -220 7935 -205
rect 7865 -260 7880 -220
rect 7920 -260 7935 -220
rect 7865 -275 7935 -260
rect 9555 -210 9625 -195
rect 9555 -250 9570 -210
rect 9610 -250 9625 -210
rect 9555 -265 9625 -250
rect 11935 -220 12005 -205
rect 11935 -260 11950 -220
rect 11990 -260 12005 -220
rect 11935 -275 12005 -260
rect 13855 -220 13925 -205
rect 13855 -260 13870 -220
rect 13910 -260 13925 -220
rect 13855 -275 13925 -260
rect 15800 -220 15870 -205
rect 15800 -260 15815 -220
rect 15855 -260 15870 -220
rect 15800 -275 15870 -260
rect 17690 -210 17760 -195
rect 17690 -250 17705 -210
rect 17745 -250 17760 -210
rect 17690 -265 17760 -250
rect 19630 -210 19700 -195
rect 19630 -250 19645 -210
rect 19685 -250 19700 -210
rect 19630 -265 19700 -250
rect 31065 -220 31195 -205
rect 31065 -320 31080 -220
rect 31180 -320 31195 -220
rect 31065 -335 31195 -320
rect -455 -555 -325 -540
rect -455 -655 -440 -555
rect -340 -655 -325 -555
rect -455 -670 -325 -655
rect 31065 -770 31195 -755
rect 31065 -870 31080 -770
rect 31180 -870 31195 -770
rect 31065 -885 31195 -870
rect -290 -965 -160 -950
rect -290 -1065 -275 -965
rect -175 -1065 -160 -965
rect -290 -1080 -160 -1065
rect 260 -965 390 -950
rect 260 -1065 275 -965
rect 375 -1065 390 -965
rect 260 -1080 390 -1065
rect 810 -965 940 -950
rect 810 -1065 825 -965
rect 925 -1065 940 -965
rect 810 -1080 940 -1065
rect 1360 -965 1490 -950
rect 1360 -1065 1375 -965
rect 1475 -1065 1490 -965
rect 1360 -1080 1490 -1065
rect 1910 -965 2040 -950
rect 1910 -1065 1925 -965
rect 2025 -1065 2040 -965
rect 1910 -1080 2040 -1065
rect 2460 -965 2590 -950
rect 2460 -1065 2475 -965
rect 2575 -1065 2590 -965
rect 2460 -1080 2590 -1065
rect 3010 -965 3140 -950
rect 3010 -1065 3025 -965
rect 3125 -1065 3140 -965
rect 3010 -1080 3140 -1065
rect 3560 -965 3690 -950
rect 3560 -1065 3575 -965
rect 3675 -1065 3690 -965
rect 3560 -1080 3690 -1065
rect 4110 -965 4240 -950
rect 4110 -1065 4125 -965
rect 4225 -1065 4240 -965
rect 4110 -1080 4240 -1065
rect 4660 -965 4790 -950
rect 4660 -1065 4675 -965
rect 4775 -1065 4790 -965
rect 4660 -1080 4790 -1065
rect 5210 -965 5340 -950
rect 5210 -1065 5225 -965
rect 5325 -1065 5340 -965
rect 5210 -1080 5340 -1065
rect 5760 -965 5890 -950
rect 5760 -1065 5775 -965
rect 5875 -1065 5890 -965
rect 5760 -1080 5890 -1065
rect 6310 -965 6440 -950
rect 6310 -1065 6325 -965
rect 6425 -1065 6440 -965
rect 6310 -1080 6440 -1065
rect 6860 -965 6990 -950
rect 6860 -1065 6875 -965
rect 6975 -1065 6990 -965
rect 6860 -1080 6990 -1065
rect 7410 -965 7540 -950
rect 7410 -1065 7425 -965
rect 7525 -1065 7540 -965
rect 7410 -1080 7540 -1065
rect 7960 -965 8090 -950
rect 7960 -1065 7975 -965
rect 8075 -1065 8090 -965
rect 7960 -1080 8090 -1065
rect 8510 -965 8640 -950
rect 8510 -1065 8525 -965
rect 8625 -1065 8640 -965
rect 8510 -1080 8640 -1065
rect 9060 -965 9190 -950
rect 9060 -1065 9075 -965
rect 9175 -1065 9190 -965
rect 9060 -1080 9190 -1065
rect 9610 -965 9740 -950
rect 9610 -1065 9625 -965
rect 9725 -1065 9740 -965
rect 9610 -1080 9740 -1065
rect 10160 -965 10290 -950
rect 10160 -1065 10175 -965
rect 10275 -1065 10290 -965
rect 10160 -1080 10290 -1065
rect 10710 -965 10840 -950
rect 10710 -1065 10725 -965
rect 10825 -1065 10840 -965
rect 10710 -1080 10840 -1065
rect 11260 -965 11390 -950
rect 11260 -1065 11275 -965
rect 11375 -1065 11390 -965
rect 11260 -1080 11390 -1065
rect 11810 -965 11940 -950
rect 11810 -1065 11825 -965
rect 11925 -1065 11940 -965
rect 11810 -1080 11940 -1065
rect 12360 -965 12490 -950
rect 12360 -1065 12375 -965
rect 12475 -1065 12490 -965
rect 12360 -1080 12490 -1065
rect 12910 -965 13040 -950
rect 12910 -1065 12925 -965
rect 13025 -1065 13040 -965
rect 12910 -1080 13040 -1065
rect 13460 -965 13590 -950
rect 13460 -1065 13475 -965
rect 13575 -1065 13590 -965
rect 13460 -1080 13590 -1065
rect 14010 -965 14140 -950
rect 14010 -1065 14025 -965
rect 14125 -1065 14140 -965
rect 14010 -1080 14140 -1065
rect 14560 -965 14690 -950
rect 14560 -1065 14575 -965
rect 14675 -1065 14690 -965
rect 14560 -1080 14690 -1065
rect 15110 -965 15240 -950
rect 15110 -1065 15125 -965
rect 15225 -1065 15240 -965
rect 15110 -1080 15240 -1065
rect 15660 -965 15790 -950
rect 15660 -1065 15675 -965
rect 15775 -1065 15790 -965
rect 15660 -1080 15790 -1065
rect 16210 -965 16340 -950
rect 16210 -1065 16225 -965
rect 16325 -1065 16340 -965
rect 16210 -1080 16340 -1065
rect 16760 -965 16890 -950
rect 16760 -1065 16775 -965
rect 16875 -1065 16890 -965
rect 16760 -1080 16890 -1065
rect 17310 -965 17440 -950
rect 17310 -1065 17325 -965
rect 17425 -1065 17440 -965
rect 17310 -1080 17440 -1065
rect 17860 -965 17990 -950
rect 17860 -1065 17875 -965
rect 17975 -1065 17990 -965
rect 17860 -1080 17990 -1065
rect 18410 -965 18540 -950
rect 18410 -1065 18425 -965
rect 18525 -1065 18540 -965
rect 18410 -1080 18540 -1065
rect 18960 -965 19090 -950
rect 18960 -1065 18975 -965
rect 19075 -1065 19090 -965
rect 18960 -1080 19090 -1065
rect 19510 -965 19640 -950
rect 19510 -1065 19525 -965
rect 19625 -1065 19640 -965
rect 19510 -1080 19640 -1065
rect 20060 -965 20190 -950
rect 20060 -1065 20075 -965
rect 20175 -1065 20190 -965
rect 20060 -1080 20190 -1065
rect 20610 -965 20740 -950
rect 20610 -1065 20625 -965
rect 20725 -1065 20740 -965
rect 20610 -1080 20740 -1065
rect 21160 -965 21290 -950
rect 21160 -1065 21175 -965
rect 21275 -1065 21290 -965
rect 21160 -1080 21290 -1065
rect 22050 -965 22180 -950
rect 22050 -1065 22065 -965
rect 22165 -1065 22180 -965
rect 22050 -1080 22180 -1065
rect 22600 -965 22730 -950
rect 22600 -1065 22615 -965
rect 22715 -1065 22730 -965
rect 22600 -1080 22730 -1065
rect 23150 -965 23280 -950
rect 23150 -1065 23165 -965
rect 23265 -1065 23280 -965
rect 23150 -1080 23280 -1065
rect 23700 -965 23830 -950
rect 23700 -1065 23715 -965
rect 23815 -1065 23830 -965
rect 23700 -1080 23830 -1065
rect 24250 -965 24380 -950
rect 24250 -1065 24265 -965
rect 24365 -1065 24380 -965
rect 24250 -1080 24380 -1065
rect 24800 -965 24930 -950
rect 24800 -1065 24815 -965
rect 24915 -1065 24930 -965
rect 24800 -1080 24930 -1065
rect 25350 -965 25480 -950
rect 25350 -1065 25365 -965
rect 25465 -1065 25480 -965
rect 25350 -1080 25480 -1065
rect 25900 -965 26030 -950
rect 25900 -1065 25915 -965
rect 26015 -1065 26030 -965
rect 25900 -1080 26030 -1065
rect 26450 -965 26580 -950
rect 26450 -1065 26465 -965
rect 26565 -1065 26580 -965
rect 26450 -1080 26580 -1065
rect 27000 -965 27130 -950
rect 27000 -1065 27015 -965
rect 27115 -1065 27130 -965
rect 27000 -1080 27130 -1065
rect 27550 -965 27680 -950
rect 27550 -1065 27565 -965
rect 27665 -1065 27680 -965
rect 27550 -1080 27680 -1065
rect 28100 -965 28230 -950
rect 28100 -1065 28115 -965
rect 28215 -1065 28230 -965
rect 28100 -1080 28230 -1065
rect 28650 -965 28780 -950
rect 28650 -1065 28665 -965
rect 28765 -1065 28780 -965
rect 28650 -1080 28780 -1065
rect 29200 -965 29330 -950
rect 29200 -1065 29215 -965
rect 29315 -1065 29330 -965
rect 29200 -1080 29330 -1065
rect 29750 -965 29880 -950
rect 29750 -1065 29765 -965
rect 29865 -1065 29880 -965
rect 29750 -1080 29880 -1065
rect 30300 -965 30430 -950
rect 30300 -1065 30315 -965
rect 30415 -1065 30430 -965
rect 30300 -1080 30430 -1065
rect 30850 -965 30980 -950
rect 30850 -1065 30865 -965
rect 30965 -1065 30980 -965
rect 30850 -1080 30980 -1065
<< nsubdiff >>
rect 2250 305 2315 320
rect 180 275 245 290
rect 180 240 195 275
rect 230 240 245 275
rect 180 225 245 240
rect 2250 270 2265 305
rect 2300 270 2315 305
rect 4190 305 4255 320
rect 2250 255 2315 270
rect 4190 270 4205 305
rect 4240 270 4255 305
rect 6440 305 6505 320
rect 4190 255 4255 270
rect 6440 270 6455 305
rect 6490 270 6505 305
rect 9345 305 9410 320
rect 6440 255 6505 270
rect 9345 270 9360 305
rect 9395 270 9410 305
rect 11290 305 11355 320
rect 9345 255 9410 270
rect 11290 270 11305 305
rect 11340 270 11355 305
rect 12985 305 13050 320
rect 11290 255 11355 270
rect 12985 270 13000 305
rect 13035 270 13050 305
rect 15170 305 15235 320
rect 12985 255 13050 270
rect 15170 270 15185 305
rect 15220 270 15235 305
rect 17350 305 17415 320
rect 15170 255 15235 270
rect 17350 270 17365 305
rect 17400 270 17415 305
rect 19535 305 19600 320
rect 17350 255 17415 270
rect 19535 270 19550 305
rect 19585 270 19600 305
rect 20745 305 20810 320
rect 19535 255 19600 270
rect 20745 270 20760 305
rect 20795 270 20810 305
rect 20745 255 20810 270
rect 785 -835 850 -820
rect 785 -870 800 -835
rect 835 -870 850 -835
rect 2945 -835 3010 -820
rect 785 -885 850 -870
rect 2945 -870 2960 -835
rect 2995 -870 3010 -835
rect 5105 -835 5170 -820
rect 2945 -885 3010 -870
rect 5105 -870 5120 -835
rect 5155 -870 5170 -835
rect 7265 -835 7330 -820
rect 5105 -885 5170 -870
rect 7265 -870 7280 -835
rect 7315 -870 7330 -835
rect 9425 -835 9490 -820
rect 7265 -885 7330 -870
rect 9425 -870 9440 -835
rect 9475 -870 9490 -835
rect 11585 -835 11650 -820
rect 9425 -885 9490 -870
rect 11585 -870 11600 -835
rect 11635 -870 11650 -835
rect 13745 -835 13810 -820
rect 11585 -885 11650 -870
rect 13745 -870 13760 -835
rect 13795 -870 13810 -835
rect 15905 -835 15970 -820
rect 13745 -885 13810 -870
rect 15905 -870 15920 -835
rect 15955 -870 15970 -835
rect 18065 -835 18130 -820
rect 15905 -885 15970 -870
rect 18065 -870 18080 -835
rect 18115 -870 18130 -835
rect 20225 -835 20290 -820
rect 18065 -885 18130 -870
rect 20225 -870 20240 -835
rect 20275 -870 20290 -835
rect 22385 -835 22450 -820
rect 20225 -885 20290 -870
rect 22385 -870 22400 -835
rect 22435 -870 22450 -835
rect 24305 -835 24370 -820
rect 22385 -885 22450 -870
rect 24305 -870 24320 -835
rect 24355 -870 24370 -835
rect 26225 -835 26290 -820
rect 24305 -885 24370 -870
rect 26225 -870 26240 -835
rect 26275 -870 26290 -835
rect 28145 -835 28210 -820
rect 26225 -885 26290 -870
rect 28145 -870 28160 -835
rect 28195 -870 28210 -835
rect 29825 -835 29890 -820
rect 28145 -885 28210 -870
rect 29825 -870 29840 -835
rect 29875 -870 29890 -835
rect 29825 -885 29890 -870
<< psubdiffcont >>
rect -235 375 -135 475
rect 315 375 415 475
rect 865 375 965 475
rect 1415 375 1515 475
rect 1965 375 2065 475
rect 2515 375 2615 475
rect 3065 375 3165 475
rect 3615 375 3715 475
rect 4165 375 4265 475
rect 4715 375 4815 475
rect 5265 375 5365 475
rect 5815 375 5915 475
rect 6365 375 6465 475
rect 6915 375 7015 475
rect 7465 375 7565 475
rect 8015 375 8115 475
rect 8565 375 8665 475
rect 9115 375 9215 475
rect 9665 375 9765 475
rect 10215 375 10315 475
rect 10765 375 10865 475
rect 11315 375 11415 475
rect 11865 375 11965 475
rect 12415 375 12515 475
rect 12965 375 13065 475
rect 13515 375 13615 475
rect 14065 375 14165 475
rect 14615 375 14715 475
rect 15165 375 15265 475
rect 15715 375 15815 475
rect 16265 375 16365 475
rect 16815 375 16915 475
rect 17365 375 17465 475
rect 17915 375 18015 475
rect 18465 375 18565 475
rect 19015 375 19115 475
rect 19565 375 19665 475
rect 20115 375 20215 475
rect 20665 375 20765 475
rect 21215 375 21315 475
rect 21545 165 21645 265
rect -440 -105 -340 -5
rect 21765 -105 21865 -5
rect 22315 -105 22415 -5
rect 22865 -105 22965 -5
rect 23415 -105 23515 -5
rect 23965 -105 24065 -5
rect 24515 -105 24615 -5
rect 25065 -105 25165 -5
rect 25615 -105 25715 -5
rect 26165 -105 26265 -5
rect 26715 -105 26815 -5
rect 27265 -105 27365 -5
rect 27815 -105 27915 -5
rect 28365 -105 28465 -5
rect 28915 -105 29015 -5
rect 29465 -105 29565 -5
rect 30015 -105 30115 -5
rect 30565 -105 30665 -5
rect 1635 -240 1675 -200
rect 4060 -235 4100 -195
rect 6455 -260 6495 -220
rect 7880 -260 7920 -220
rect 9570 -250 9610 -210
rect 11950 -260 11990 -220
rect 13870 -260 13910 -220
rect 15815 -260 15855 -220
rect 17705 -250 17745 -210
rect 19645 -250 19685 -210
rect 31080 -320 31180 -220
rect -440 -655 -340 -555
rect 31080 -870 31180 -770
rect -275 -1065 -175 -965
rect 275 -1065 375 -965
rect 825 -1065 925 -965
rect 1375 -1065 1475 -965
rect 1925 -1065 2025 -965
rect 2475 -1065 2575 -965
rect 3025 -1065 3125 -965
rect 3575 -1065 3675 -965
rect 4125 -1065 4225 -965
rect 4675 -1065 4775 -965
rect 5225 -1065 5325 -965
rect 5775 -1065 5875 -965
rect 6325 -1065 6425 -965
rect 6875 -1065 6975 -965
rect 7425 -1065 7525 -965
rect 7975 -1065 8075 -965
rect 8525 -1065 8625 -965
rect 9075 -1065 9175 -965
rect 9625 -1065 9725 -965
rect 10175 -1065 10275 -965
rect 10725 -1065 10825 -965
rect 11275 -1065 11375 -965
rect 11825 -1065 11925 -965
rect 12375 -1065 12475 -965
rect 12925 -1065 13025 -965
rect 13475 -1065 13575 -965
rect 14025 -1065 14125 -965
rect 14575 -1065 14675 -965
rect 15125 -1065 15225 -965
rect 15675 -1065 15775 -965
rect 16225 -1065 16325 -965
rect 16775 -1065 16875 -965
rect 17325 -1065 17425 -965
rect 17875 -1065 17975 -965
rect 18425 -1065 18525 -965
rect 18975 -1065 19075 -965
rect 19525 -1065 19625 -965
rect 20075 -1065 20175 -965
rect 20625 -1065 20725 -965
rect 21175 -1065 21275 -965
rect 22065 -1065 22165 -965
rect 22615 -1065 22715 -965
rect 23165 -1065 23265 -965
rect 23715 -1065 23815 -965
rect 24265 -1065 24365 -965
rect 24815 -1065 24915 -965
rect 25365 -1065 25465 -965
rect 25915 -1065 26015 -965
rect 26465 -1065 26565 -965
rect 27015 -1065 27115 -965
rect 27565 -1065 27665 -965
rect 28115 -1065 28215 -965
rect 28665 -1065 28765 -965
rect 29215 -1065 29315 -965
rect 29765 -1065 29865 -965
rect 30315 -1065 30415 -965
rect 30865 -1065 30965 -965
<< nsubdiffcont >>
rect 195 240 230 275
rect 2265 270 2300 305
rect 4205 270 4240 305
rect 6455 270 6490 305
rect 9360 270 9395 305
rect 11305 270 11340 305
rect 13000 270 13035 305
rect 15185 270 15220 305
rect 17365 270 17400 305
rect 19550 270 19585 305
rect 20760 270 20795 305
rect 800 -870 835 -835
rect 2960 -870 2995 -835
rect 5120 -870 5155 -835
rect 7280 -870 7315 -835
rect 9440 -870 9475 -835
rect 11600 -870 11635 -835
rect 13760 -870 13795 -835
rect 15920 -870 15955 -835
rect 18080 -870 18115 -835
rect 20240 -870 20275 -835
rect 22400 -870 22435 -835
rect 24320 -870 24355 -835
rect 26240 -870 26275 -835
rect 28160 -870 28195 -835
rect 29840 -870 29875 -835
<< poly >>
rect 356 200 551 215
rect 231 185 246 200
rect 356 185 371 200
rect 416 185 431 200
rect 476 185 491 200
rect 536 185 551 200
rect 661 200 1586 215
rect 661 185 676 200
rect 721 185 736 200
rect 781 185 796 200
rect 841 185 856 200
rect 906 185 921 200
rect 966 185 981 200
rect 1026 185 1041 200
rect 1086 185 1101 200
rect 1146 185 1161 200
rect 1206 185 1221 200
rect 1266 185 1281 200
rect 1326 185 1341 200
rect 1391 185 1406 200
rect 1451 185 1466 200
rect 1511 185 1526 200
rect 1571 185 1586 200
rect 1696 200 5531 215
rect 1696 185 1711 200
rect 1756 185 1771 200
rect 1816 185 1831 200
rect 1876 185 1891 200
rect 1941 185 1956 200
rect 2001 185 2016 200
rect 2061 185 2076 200
rect 2121 185 2136 200
rect 2181 185 2196 200
rect 2241 185 2256 200
rect 2301 185 2316 200
rect 2361 185 2376 200
rect 2426 185 2441 200
rect 2486 185 2501 200
rect 2546 185 2561 200
rect 2606 185 2621 200
rect 2666 185 2681 200
rect 2726 185 2741 200
rect 2786 185 2801 200
rect 2846 185 2861 200
rect 2911 185 2926 200
rect 2971 185 2986 200
rect 3031 185 3046 200
rect 3091 185 3106 200
rect 3151 185 3166 200
rect 3211 185 3226 200
rect 3271 185 3286 200
rect 3331 185 3346 200
rect 3396 185 3411 200
rect 3456 185 3471 200
rect 3516 185 3531 200
rect 3576 185 3591 200
rect 3636 185 3651 200
rect 3696 185 3711 200
rect 3756 185 3771 200
rect 3816 185 3831 200
rect 3881 185 3896 200
rect 3941 185 3956 200
rect 4001 185 4016 200
rect 4061 185 4076 200
rect 4121 185 4136 200
rect 4181 185 4196 200
rect 4241 185 4256 200
rect 4301 185 4316 200
rect 4366 185 4381 200
rect 4426 185 4441 200
rect 4486 185 4501 200
rect 4546 185 4561 200
rect 4606 185 4621 200
rect 4666 185 4681 200
rect 4726 185 4741 200
rect 4786 185 4801 200
rect 4851 185 4866 200
rect 4911 185 4926 200
rect 4971 185 4986 200
rect 5031 185 5046 200
rect 5091 185 5106 200
rect 5151 185 5166 200
rect 5211 185 5226 200
rect 5271 185 5286 200
rect 5336 185 5351 200
rect 5396 185 5411 200
rect 5456 185 5471 200
rect 5516 185 5531 200
rect 5641 200 21116 215
rect 5641 185 5656 200
rect 5701 185 5716 200
rect 5761 185 5776 200
rect 5821 185 5836 200
rect 5886 185 5901 200
rect 5946 185 5961 200
rect 6006 185 6021 200
rect 6066 185 6081 200
rect 6126 185 6141 200
rect 6186 185 6201 200
rect 6246 185 6261 200
rect 6306 185 6321 200
rect 6371 185 6386 200
rect 6431 185 6446 200
rect 6491 185 6506 200
rect 6551 185 6566 200
rect 6611 185 6626 200
rect 6671 185 6686 200
rect 6731 185 6746 200
rect 6791 185 6806 200
rect 6856 185 6871 200
rect 6916 185 6931 200
rect 6976 185 6991 200
rect 7036 185 7051 200
rect 7096 185 7111 200
rect 7156 185 7171 200
rect 7216 185 7231 200
rect 7276 185 7291 200
rect 7336 185 7351 200
rect 7396 185 7411 200
rect 7456 185 7471 200
rect 7516 185 7531 200
rect 7576 185 7591 200
rect 7636 185 7651 200
rect 7696 185 7711 200
rect 7756 185 7771 200
rect 7821 185 7836 200
rect 7881 185 7896 200
rect 7941 185 7956 200
rect 8001 185 8016 200
rect 8061 185 8076 200
rect 8121 185 8136 200
rect 8181 185 8196 200
rect 8241 185 8256 200
rect 8306 185 8321 200
rect 8366 185 8381 200
rect 8426 185 8441 200
rect 8486 185 8501 200
rect 8546 185 8561 200
rect 8606 185 8621 200
rect 8666 185 8681 200
rect 8726 185 8741 200
rect 8791 185 8806 200
rect 8851 185 8866 200
rect 8911 185 8926 200
rect 8971 185 8986 200
rect 9031 185 9046 200
rect 9091 185 9106 200
rect 9151 185 9166 200
rect 9211 185 9226 200
rect 9276 185 9291 200
rect 9336 185 9351 200
rect 9396 185 9411 200
rect 9456 185 9471 200
rect 9521 185 9536 200
rect 9581 185 9596 200
rect 9641 185 9656 200
rect 9701 185 9716 200
rect 9766 185 9781 200
rect 9826 185 9841 200
rect 9886 185 9901 200
rect 9946 185 9961 200
rect 10006 185 10021 200
rect 10066 185 10081 200
rect 10126 185 10141 200
rect 10186 185 10201 200
rect 10251 185 10266 200
rect 10311 185 10326 200
rect 10371 185 10386 200
rect 10431 185 10446 200
rect 10491 185 10506 200
rect 10551 185 10566 200
rect 10611 185 10626 200
rect 10671 185 10686 200
rect 10736 185 10751 200
rect 10796 185 10811 200
rect 10856 185 10871 200
rect 10916 185 10931 200
rect 10976 185 10991 200
rect 11036 185 11051 200
rect 11096 185 11111 200
rect 11156 185 11171 200
rect 11221 185 11236 200
rect 11281 185 11296 200
rect 11341 185 11356 200
rect 11401 185 11416 200
rect 11461 185 11476 200
rect 11521 185 11536 200
rect 11581 185 11596 200
rect 11641 185 11656 200
rect 11706 185 11721 200
rect 11766 185 11781 200
rect 11826 185 11841 200
rect 11886 185 11901 200
rect 11946 185 11961 200
rect 12006 185 12021 200
rect 12066 185 12081 200
rect 12126 185 12141 200
rect 12191 185 12206 200
rect 12251 185 12266 200
rect 12311 185 12326 200
rect 12371 185 12386 200
rect 12431 185 12446 200
rect 12491 185 12506 200
rect 12551 185 12566 200
rect 12611 185 12626 200
rect 12676 185 12691 200
rect 12736 185 12751 200
rect 12796 185 12811 200
rect 12856 185 12871 200
rect 12916 185 12931 200
rect 12976 185 12991 200
rect 13036 185 13051 200
rect 13096 185 13111 200
rect 13161 185 13176 200
rect 13221 185 13236 200
rect 13281 185 13296 200
rect 13341 185 13356 200
rect 13401 185 13416 200
rect 13461 185 13476 200
rect 13521 185 13536 200
rect 13581 185 13596 200
rect 13646 185 13661 200
rect 13706 185 13721 200
rect 13766 185 13781 200
rect 13826 185 13841 200
rect 13886 185 13901 200
rect 13946 185 13961 200
rect 14006 185 14021 200
rect 14066 185 14081 200
rect 14131 185 14146 200
rect 14191 185 14206 200
rect 14251 185 14266 200
rect 14311 185 14326 200
rect 14371 185 14386 200
rect 14431 185 14446 200
rect 14491 185 14506 200
rect 14551 185 14566 200
rect 14616 185 14631 200
rect 14676 185 14691 200
rect 14736 185 14751 200
rect 14796 185 14811 200
rect 14856 185 14871 200
rect 14916 185 14931 200
rect 14976 185 14991 200
rect 15036 185 15051 200
rect 15101 185 15116 200
rect 15161 185 15176 200
rect 15221 185 15236 200
rect 15281 185 15296 200
rect 15341 185 15356 200
rect 15401 185 15416 200
rect 15461 185 15476 200
rect 15521 185 15536 200
rect 15586 185 15601 200
rect 15646 185 15661 200
rect 15706 185 15721 200
rect 15766 185 15781 200
rect 15826 185 15841 200
rect 15886 185 15901 200
rect 15946 185 15961 200
rect 16006 185 16021 200
rect 16071 185 16086 200
rect 16131 185 16146 200
rect 16191 185 16206 200
rect 16251 185 16266 200
rect 16311 185 16326 200
rect 16371 185 16386 200
rect 16431 185 16446 200
rect 16491 185 16506 200
rect 16556 185 16571 200
rect 16616 185 16631 200
rect 16676 185 16691 200
rect 16736 185 16751 200
rect 16796 185 16811 200
rect 16856 185 16871 200
rect 16916 185 16931 200
rect 16976 185 16991 200
rect 17041 185 17056 200
rect 17101 185 17116 200
rect 17161 185 17176 200
rect 17221 185 17236 200
rect 17281 185 17296 200
rect 17341 185 17356 200
rect 17401 185 17416 200
rect 17461 185 17476 200
rect 17526 185 17541 200
rect 17586 185 17601 200
rect 17646 185 17661 200
rect 17706 185 17721 200
rect 17766 185 17781 200
rect 17826 185 17841 200
rect 17886 185 17901 200
rect 17946 185 17961 200
rect 18011 185 18026 200
rect 18071 185 18086 200
rect 18131 185 18146 200
rect 18191 185 18206 200
rect 18251 185 18266 200
rect 18311 185 18326 200
rect 18371 185 18386 200
rect 18431 185 18446 200
rect 18496 185 18511 200
rect 18556 185 18571 200
rect 18616 185 18631 200
rect 18676 185 18691 200
rect 18736 185 18751 200
rect 18796 185 18811 200
rect 18856 185 18871 200
rect 18916 185 18931 200
rect 18981 185 18996 200
rect 19041 185 19056 200
rect 19101 185 19116 200
rect 19161 185 19176 200
rect 19221 185 19236 200
rect 19281 185 19296 200
rect 19341 185 19356 200
rect 19401 185 19416 200
rect 19466 185 19481 200
rect 19526 185 19541 200
rect 19586 185 19601 200
rect 19646 185 19661 200
rect 19706 185 19721 200
rect 19766 185 19781 200
rect 19826 185 19841 200
rect 19886 185 19901 200
rect 19951 185 19966 200
rect 20011 185 20026 200
rect 20071 185 20086 200
rect 20131 185 20146 200
rect 20191 185 20206 200
rect 20251 185 20266 200
rect 20311 185 20326 200
rect 20371 185 20386 200
rect 20436 185 20451 200
rect 20496 185 20511 200
rect 20556 185 20571 200
rect 20616 185 20631 200
rect 20676 185 20691 200
rect 20736 185 20751 200
rect 20796 185 20811 200
rect 20856 185 20871 200
rect 20921 185 20936 200
rect 20981 185 20996 200
rect 21041 185 21056 200
rect 21101 185 21116 200
rect 231 25 246 85
rect 356 25 371 85
rect 191 15 246 25
rect 191 -5 201 15
rect 221 -5 246 15
rect 191 -15 246 -5
rect 316 15 371 25
rect 316 -5 326 15
rect 346 -5 371 15
rect 316 -15 371 -5
rect 231 -70 246 -15
rect 356 -70 371 -15
rect 416 -70 431 85
rect 476 -70 491 85
rect 536 -70 551 85
rect 661 25 676 85
rect 621 15 676 25
rect 621 -5 631 15
rect 651 -5 676 15
rect 621 -15 676 -5
rect 661 -70 676 -15
rect 721 -70 736 85
rect 781 -70 796 85
rect 841 -70 856 85
rect 906 -70 921 85
rect 966 -70 981 85
rect 1026 -70 1041 85
rect 1086 -70 1101 85
rect 1146 -70 1161 85
rect 1206 -70 1221 85
rect 1266 -70 1281 85
rect 1326 -70 1341 85
rect 1391 -70 1406 85
rect 1451 -70 1466 85
rect 1511 -70 1526 85
rect 1571 -70 1586 85
rect 1696 25 1711 85
rect 1656 15 1711 25
rect 1656 -5 1666 15
rect 1686 -5 1711 15
rect 1656 -15 1711 -5
rect 1696 -70 1711 -15
rect 1756 -70 1771 85
rect 1816 -70 1831 85
rect 1876 -70 1891 85
rect 1941 -70 1956 85
rect 2001 -70 2016 85
rect 2061 -70 2076 85
rect 2121 -70 2136 85
rect 2181 -70 2196 85
rect 2241 -70 2256 85
rect 2301 -70 2316 85
rect 2361 -70 2376 85
rect 2426 -70 2441 85
rect 2486 -70 2501 85
rect 2546 -70 2561 85
rect 2606 -70 2621 85
rect 2666 -70 2681 85
rect 2726 -70 2741 85
rect 2786 -70 2801 85
rect 2846 -70 2861 85
rect 2911 -70 2926 85
rect 2971 -70 2986 85
rect 3031 -70 3046 85
rect 3091 -70 3106 85
rect 3151 -70 3166 85
rect 3211 -70 3226 85
rect 3271 -70 3286 85
rect 3331 -70 3346 85
rect 3396 -70 3411 85
rect 3456 -70 3471 85
rect 3516 -70 3531 85
rect 3576 -70 3591 85
rect 3636 -70 3651 85
rect 3696 -70 3711 85
rect 3756 -70 3771 85
rect 3816 -70 3831 85
rect 3881 -70 3896 85
rect 3941 -70 3956 85
rect 4001 -70 4016 85
rect 4061 -70 4076 85
rect 4121 -70 4136 85
rect 4181 -70 4196 85
rect 4241 -70 4256 85
rect 4301 -70 4316 85
rect 4366 -70 4381 85
rect 4426 -70 4441 85
rect 4486 -70 4501 85
rect 4546 -70 4561 85
rect 4606 -70 4621 85
rect 4666 -70 4681 85
rect 4726 -70 4741 85
rect 4786 -70 4801 85
rect 4851 -70 4866 85
rect 4911 -70 4926 85
rect 4971 -70 4986 85
rect 5031 -70 5046 85
rect 5091 -70 5106 85
rect 5151 -70 5166 85
rect 5211 -70 5226 85
rect 5271 -70 5286 85
rect 5336 -70 5351 85
rect 5396 -70 5411 85
rect 5456 -70 5471 85
rect 5516 -70 5531 85
rect 5641 25 5656 85
rect 5601 15 5656 25
rect 5601 -5 5611 15
rect 5631 -5 5656 15
rect 5601 -15 5656 -5
rect 5641 -70 5656 -15
rect 5701 -70 5716 85
rect 5761 -70 5776 85
rect 5821 -70 5836 85
rect 5886 -70 5901 85
rect 5946 -70 5961 85
rect 6006 -70 6021 85
rect 6066 -70 6081 85
rect 6126 -70 6141 85
rect 6186 -70 6201 85
rect 6246 -70 6261 85
rect 6306 -70 6321 85
rect 6371 -70 6386 85
rect 6431 -70 6446 85
rect 6491 -70 6506 85
rect 6551 -70 6566 85
rect 6611 -70 6626 85
rect 6671 -70 6686 85
rect 6731 -70 6746 85
rect 6791 -70 6806 85
rect 6856 -70 6871 85
rect 6916 -70 6931 85
rect 6976 -70 6991 85
rect 7036 -70 7051 85
rect 7096 -70 7111 85
rect 7156 -70 7171 85
rect 7216 -70 7231 85
rect 7276 -70 7291 85
rect 7336 -70 7351 85
rect 7396 -70 7411 85
rect 7456 -70 7471 85
rect 7516 -70 7531 85
rect 7576 -70 7591 85
rect 7636 -70 7651 85
rect 7696 -70 7711 85
rect 7756 -70 7771 85
rect 7821 -70 7836 85
rect 7881 -70 7896 85
rect 7941 -70 7956 85
rect 8001 -70 8016 85
rect 8061 -70 8076 85
rect 8121 -70 8136 85
rect 8181 -70 8196 85
rect 8241 -70 8256 85
rect 8306 -70 8321 85
rect 8366 -70 8381 85
rect 8426 -70 8441 85
rect 8486 -70 8501 85
rect 8546 -70 8561 85
rect 8606 -70 8621 85
rect 8666 -70 8681 85
rect 8726 -70 8741 85
rect 8791 -70 8806 85
rect 8851 -70 8866 85
rect 8911 -70 8926 85
rect 8971 -70 8986 85
rect 9031 -70 9046 85
rect 9091 -70 9106 85
rect 9151 -70 9166 85
rect 9211 -70 9226 85
rect 9276 -70 9291 85
rect 9336 -70 9351 85
rect 9396 -70 9411 85
rect 9456 -70 9471 85
rect 9521 -70 9536 85
rect 9581 -70 9596 85
rect 9641 -70 9656 85
rect 9701 -70 9716 85
rect 9766 -70 9781 85
rect 9826 -70 9841 85
rect 9886 -70 9901 85
rect 9946 -70 9961 85
rect 10006 -70 10021 85
rect 10066 -70 10081 85
rect 10126 -70 10141 85
rect 10186 -70 10201 85
rect 10251 -70 10266 85
rect 10311 -70 10326 85
rect 10371 -70 10386 85
rect 10431 -70 10446 85
rect 10491 -70 10506 85
rect 10551 -70 10566 85
rect 10611 -70 10626 85
rect 10671 -70 10686 85
rect 10736 -70 10751 85
rect 10796 -70 10811 85
rect 10856 -70 10871 85
rect 10916 -70 10931 85
rect 10976 -70 10991 85
rect 11036 -70 11051 85
rect 11096 -70 11111 85
rect 11156 -70 11171 85
rect 11221 -70 11236 85
rect 11281 -70 11296 85
rect 11341 -70 11356 85
rect 11401 -70 11416 85
rect 11461 -70 11476 85
rect 11521 -70 11536 85
rect 11581 -70 11596 85
rect 11641 -70 11656 85
rect 11706 -70 11721 85
rect 11766 -70 11781 85
rect 11826 -70 11841 85
rect 11886 -70 11901 85
rect 11946 -70 11961 85
rect 12006 -70 12021 85
rect 12066 -70 12081 85
rect 12126 -70 12141 85
rect 12191 -70 12206 85
rect 12251 -70 12266 85
rect 12311 -70 12326 85
rect 12371 -70 12386 85
rect 12431 -70 12446 85
rect 12491 -70 12506 85
rect 12551 -70 12566 85
rect 12611 -70 12626 85
rect 12676 -70 12691 85
rect 12736 -70 12751 85
rect 12796 -70 12811 85
rect 12856 -70 12871 85
rect 12916 -70 12931 85
rect 12976 -70 12991 85
rect 13036 -70 13051 85
rect 13096 -70 13111 85
rect 13161 -70 13176 85
rect 13221 -70 13236 85
rect 13281 -70 13296 85
rect 13341 -70 13356 85
rect 13401 -70 13416 85
rect 13461 -70 13476 85
rect 13521 -70 13536 85
rect 13581 -70 13596 85
rect 13646 -70 13661 85
rect 13706 -70 13721 85
rect 13766 -70 13781 85
rect 13826 -70 13841 85
rect 13886 -70 13901 85
rect 13946 -70 13961 85
rect 14006 -70 14021 85
rect 14066 -70 14081 85
rect 14131 -70 14146 85
rect 14191 -70 14206 85
rect 14251 -70 14266 85
rect 14311 -70 14326 85
rect 14371 -70 14386 85
rect 14431 -70 14446 85
rect 14491 -70 14506 85
rect 14551 -70 14566 85
rect 14616 -70 14631 85
rect 14676 -70 14691 85
rect 14736 -70 14751 85
rect 14796 -70 14811 85
rect 14856 -70 14871 85
rect 14916 -70 14931 85
rect 14976 -70 14991 85
rect 15036 -70 15051 85
rect 15101 -70 15116 85
rect 15161 -70 15176 85
rect 15221 -70 15236 85
rect 15281 -70 15296 85
rect 15341 -70 15356 85
rect 15401 -70 15416 85
rect 15461 -70 15476 85
rect 15521 -70 15536 85
rect 15586 -70 15601 85
rect 15646 -70 15661 85
rect 15706 -70 15721 85
rect 15766 -70 15781 85
rect 15826 -70 15841 85
rect 15886 -70 15901 85
rect 15946 -70 15961 85
rect 16006 -70 16021 85
rect 16071 -70 16086 85
rect 16131 -70 16146 85
rect 16191 -70 16206 85
rect 16251 -70 16266 85
rect 16311 -70 16326 85
rect 16371 -70 16386 85
rect 16431 -70 16446 85
rect 16491 -70 16506 85
rect 16556 -70 16571 85
rect 16616 -70 16631 85
rect 16676 -70 16691 85
rect 16736 -70 16751 85
rect 16796 -70 16811 85
rect 16856 -70 16871 85
rect 16916 -70 16931 85
rect 16976 -70 16991 85
rect 17041 -70 17056 85
rect 17101 -70 17116 85
rect 17161 -70 17176 85
rect 17221 -70 17236 85
rect 17281 -70 17296 85
rect 17341 -70 17356 85
rect 17401 -70 17416 85
rect 17461 -70 17476 85
rect 17526 -70 17541 85
rect 17586 -70 17601 85
rect 17646 -70 17661 85
rect 17706 -70 17721 85
rect 17766 -70 17781 85
rect 17826 -70 17841 85
rect 17886 -70 17901 85
rect 17946 -70 17961 85
rect 18011 -70 18026 85
rect 18071 -70 18086 85
rect 18131 -70 18146 85
rect 18191 -70 18206 85
rect 18251 -70 18266 85
rect 18311 -70 18326 85
rect 18371 -70 18386 85
rect 18431 -70 18446 85
rect 18496 -70 18511 85
rect 18556 -70 18571 85
rect 18616 -70 18631 85
rect 18676 -70 18691 85
rect 18736 -70 18751 85
rect 18796 -70 18811 85
rect 18856 -70 18871 85
rect 18916 -70 18931 85
rect 18981 -70 18996 85
rect 19041 -70 19056 85
rect 19101 -70 19116 85
rect 19161 -70 19176 85
rect 19221 -70 19236 85
rect 19281 -70 19296 85
rect 19341 -70 19356 85
rect 19401 -70 19416 85
rect 19466 -70 19481 85
rect 19526 -70 19541 85
rect 19586 -70 19601 85
rect 19646 -70 19661 85
rect 19706 -70 19721 85
rect 19766 -70 19781 85
rect 19826 -70 19841 85
rect 19886 -70 19901 85
rect 19951 -70 19966 85
rect 20011 -70 20026 85
rect 20071 -70 20086 85
rect 20131 -70 20146 85
rect 20191 -70 20206 85
rect 20251 -70 20266 85
rect 20311 -70 20326 85
rect 20371 -70 20386 85
rect 20436 -70 20451 85
rect 20496 -70 20511 85
rect 20556 -70 20571 85
rect 20616 -70 20631 85
rect 20676 -70 20691 85
rect 20736 -70 20751 85
rect 20796 -70 20811 85
rect 20856 -70 20871 85
rect 20921 -70 20936 85
rect 20981 -70 20996 85
rect 21041 -70 21056 85
rect 21101 -70 21116 85
rect 231 -135 246 -120
rect 356 -135 371 -120
rect 416 -135 431 -120
rect 476 -135 491 -120
rect 536 -135 551 -120
rect 661 -135 676 -120
rect 721 -135 736 -120
rect 781 -135 796 -120
rect 841 -135 856 -120
rect 906 -135 921 -120
rect 966 -135 981 -120
rect 1026 -135 1041 -120
rect 1086 -135 1101 -120
rect 1146 -135 1161 -120
rect 1206 -135 1221 -120
rect 1266 -135 1281 -120
rect 1326 -135 1341 -120
rect 1391 -135 1406 -120
rect 1451 -135 1466 -120
rect 1511 -135 1526 -120
rect 1571 -135 1586 -120
rect 1696 -135 1711 -120
rect 1756 -135 1771 -120
rect 1816 -135 1831 -120
rect 1876 -135 1891 -120
rect 1941 -135 1956 -120
rect 2001 -135 2016 -120
rect 2061 -135 2076 -120
rect 2121 -135 2136 -120
rect 2181 -135 2196 -120
rect 2241 -135 2256 -120
rect 2301 -135 2316 -120
rect 2361 -135 2376 -120
rect 2426 -135 2441 -120
rect 2486 -135 2501 -120
rect 2546 -135 2561 -120
rect 2606 -135 2621 -120
rect 2666 -135 2681 -120
rect 2726 -135 2741 -120
rect 2786 -135 2801 -120
rect 2846 -135 2861 -120
rect 2911 -135 2926 -120
rect 2971 -135 2986 -120
rect 3031 -135 3046 -120
rect 3091 -135 3106 -120
rect 3151 -135 3166 -120
rect 3211 -135 3226 -120
rect 3271 -135 3286 -120
rect 3331 -135 3346 -120
rect 3396 -135 3411 -120
rect 3456 -135 3471 -120
rect 3516 -135 3531 -120
rect 3576 -135 3591 -120
rect 3636 -135 3651 -120
rect 3696 -135 3711 -120
rect 3756 -135 3771 -120
rect 3816 -135 3831 -120
rect 3881 -135 3896 -120
rect 3941 -135 3956 -120
rect 4001 -135 4016 -120
rect 4061 -135 4076 -120
rect 4121 -135 4136 -120
rect 4181 -135 4196 -120
rect 4241 -135 4256 -120
rect 4301 -135 4316 -120
rect 4366 -135 4381 -120
rect 4426 -135 4441 -120
rect 4486 -135 4501 -120
rect 4546 -135 4561 -120
rect 4606 -135 4621 -120
rect 4666 -135 4681 -120
rect 4726 -135 4741 -120
rect 4786 -135 4801 -120
rect 4851 -135 4866 -120
rect 4911 -135 4926 -120
rect 4971 -135 4986 -120
rect 5031 -135 5046 -120
rect 5091 -135 5106 -120
rect 5151 -135 5166 -120
rect 5211 -135 5226 -120
rect 5271 -135 5286 -120
rect 5336 -135 5351 -120
rect 5396 -135 5411 -120
rect 5456 -135 5471 -120
rect 5516 -135 5531 -120
rect 5641 -135 5656 -120
rect 5701 -135 5716 -120
rect 5761 -135 5776 -120
rect 5821 -135 5836 -120
rect 5886 -135 5901 -120
rect 5946 -135 5961 -120
rect 6006 -135 6021 -120
rect 6066 -135 6081 -120
rect 6126 -135 6141 -120
rect 6186 -135 6201 -120
rect 6246 -135 6261 -120
rect 6306 -135 6321 -120
rect 6371 -135 6386 -120
rect 6431 -135 6446 -120
rect 6491 -135 6506 -120
rect 6551 -135 6566 -120
rect 6611 -135 6626 -120
rect 6671 -135 6686 -120
rect 6731 -135 6746 -120
rect 6791 -135 6806 -120
rect 6856 -135 6871 -120
rect 6916 -135 6931 -120
rect 6976 -135 6991 -120
rect 7036 -135 7051 -120
rect 7096 -135 7111 -120
rect 7156 -135 7171 -120
rect 7216 -135 7231 -120
rect 7276 -135 7291 -120
rect 7336 -135 7351 -120
rect 7396 -135 7411 -120
rect 7456 -135 7471 -120
rect 7516 -135 7531 -120
rect 7576 -135 7591 -120
rect 7636 -135 7651 -120
rect 7696 -135 7711 -120
rect 7756 -135 7771 -120
rect 7821 -135 7836 -120
rect 7881 -135 7896 -120
rect 7941 -135 7956 -120
rect 8001 -135 8016 -120
rect 8061 -135 8076 -120
rect 8121 -135 8136 -120
rect 8181 -135 8196 -120
rect 8241 -135 8256 -120
rect 8306 -135 8321 -120
rect 8366 -135 8381 -120
rect 8426 -135 8441 -120
rect 8486 -135 8501 -120
rect 8546 -135 8561 -120
rect 8606 -135 8621 -120
rect 8666 -135 8681 -120
rect 8726 -135 8741 -120
rect 8791 -135 8806 -120
rect 8851 -135 8866 -120
rect 8911 -135 8926 -120
rect 8971 -135 8986 -120
rect 9031 -135 9046 -120
rect 9091 -135 9106 -120
rect 9151 -135 9166 -120
rect 9211 -135 9226 -120
rect 9276 -135 9291 -120
rect 9336 -135 9351 -120
rect 9396 -135 9411 -120
rect 9456 -135 9471 -120
rect 9521 -135 9536 -120
rect 9581 -135 9596 -120
rect 9641 -135 9656 -120
rect 9701 -135 9716 -120
rect 9766 -135 9781 -120
rect 9826 -135 9841 -120
rect 9886 -135 9901 -120
rect 9946 -135 9961 -120
rect 10006 -135 10021 -120
rect 10066 -135 10081 -120
rect 10126 -135 10141 -120
rect 10186 -135 10201 -120
rect 10251 -135 10266 -120
rect 10311 -135 10326 -120
rect 10371 -135 10386 -120
rect 10431 -135 10446 -120
rect 10491 -135 10506 -120
rect 10551 -135 10566 -120
rect 10611 -135 10626 -120
rect 10671 -135 10686 -120
rect 10736 -135 10751 -120
rect 10796 -135 10811 -120
rect 10856 -135 10871 -120
rect 10916 -135 10931 -120
rect 10976 -135 10991 -120
rect 11036 -135 11051 -120
rect 11096 -135 11111 -120
rect 11156 -135 11171 -120
rect 11221 -135 11236 -120
rect 11281 -135 11296 -120
rect 11341 -135 11356 -120
rect 11401 -135 11416 -120
rect 11461 -135 11476 -120
rect 11521 -135 11536 -120
rect 11581 -135 11596 -120
rect 11641 -135 11656 -120
rect 11706 -135 11721 -120
rect 11766 -135 11781 -120
rect 11826 -135 11841 -120
rect 11886 -135 11901 -120
rect 11946 -135 11961 -120
rect 12006 -135 12021 -120
rect 12066 -135 12081 -120
rect 12126 -135 12141 -120
rect 12191 -135 12206 -120
rect 12251 -135 12266 -120
rect 12311 -135 12326 -120
rect 12371 -135 12386 -120
rect 12431 -135 12446 -120
rect 12491 -135 12506 -120
rect 12551 -135 12566 -120
rect 12611 -135 12626 -120
rect 12676 -135 12691 -120
rect 12736 -135 12751 -120
rect 12796 -135 12811 -120
rect 12856 -135 12871 -120
rect 12916 -135 12931 -120
rect 12976 -135 12991 -120
rect 13036 -135 13051 -120
rect 13096 -135 13111 -120
rect 13161 -135 13176 -120
rect 13221 -135 13236 -120
rect 13281 -135 13296 -120
rect 13341 -135 13356 -120
rect 13401 -135 13416 -120
rect 13461 -135 13476 -120
rect 13521 -135 13536 -120
rect 13581 -135 13596 -120
rect 13646 -135 13661 -120
rect 13706 -135 13721 -120
rect 13766 -135 13781 -120
rect 13826 -135 13841 -120
rect 13886 -135 13901 -120
rect 13946 -135 13961 -120
rect 14006 -135 14021 -120
rect 14066 -135 14081 -120
rect 14131 -135 14146 -120
rect 14191 -135 14206 -120
rect 14251 -135 14266 -120
rect 14311 -135 14326 -120
rect 14371 -135 14386 -120
rect 14431 -135 14446 -120
rect 14491 -135 14506 -120
rect 14551 -135 14566 -120
rect 14616 -135 14631 -120
rect 14676 -135 14691 -120
rect 14736 -135 14751 -120
rect 14796 -135 14811 -120
rect 14856 -135 14871 -120
rect 14916 -135 14931 -120
rect 14976 -135 14991 -120
rect 15036 -135 15051 -120
rect 15101 -135 15116 -120
rect 15161 -135 15176 -120
rect 15221 -135 15236 -120
rect 15281 -135 15296 -120
rect 15341 -135 15356 -120
rect 15401 -135 15416 -120
rect 15461 -135 15476 -120
rect 15521 -135 15536 -120
rect 15586 -135 15601 -120
rect 15646 -135 15661 -120
rect 15706 -135 15721 -120
rect 15766 -135 15781 -120
rect 15826 -135 15841 -120
rect 15886 -135 15901 -120
rect 15946 -135 15961 -120
rect 16006 -135 16021 -120
rect 16071 -135 16086 -120
rect 16131 -135 16146 -120
rect 16191 -135 16206 -120
rect 16251 -135 16266 -120
rect 16311 -135 16326 -120
rect 16371 -135 16386 -120
rect 16431 -135 16446 -120
rect 16491 -135 16506 -120
rect 16556 -135 16571 -120
rect 16616 -135 16631 -120
rect 16676 -135 16691 -120
rect 16736 -135 16751 -120
rect 16796 -135 16811 -120
rect 16856 -135 16871 -120
rect 16916 -135 16931 -120
rect 16976 -135 16991 -120
rect 17041 -135 17056 -120
rect 17101 -135 17116 -120
rect 17161 -135 17176 -120
rect 17221 -135 17236 -120
rect 17281 -135 17296 -120
rect 17341 -135 17356 -120
rect 17401 -135 17416 -120
rect 17461 -135 17476 -120
rect 17526 -135 17541 -120
rect 17586 -135 17601 -120
rect 17646 -135 17661 -120
rect 17706 -135 17721 -120
rect 17766 -135 17781 -120
rect 17826 -135 17841 -120
rect 17886 -135 17901 -120
rect 17946 -135 17961 -120
rect 18011 -135 18026 -120
rect 18071 -135 18086 -120
rect 18131 -135 18146 -120
rect 18191 -135 18206 -120
rect 18251 -135 18266 -120
rect 18311 -135 18326 -120
rect 18371 -135 18386 -120
rect 18431 -135 18446 -120
rect 18496 -135 18511 -120
rect 18556 -135 18571 -120
rect 18616 -135 18631 -120
rect 18676 -135 18691 -120
rect 18736 -135 18751 -120
rect 18796 -135 18811 -120
rect 18856 -135 18871 -120
rect 18916 -135 18931 -120
rect 18981 -135 18996 -120
rect 19041 -135 19056 -120
rect 19101 -135 19116 -120
rect 19161 -135 19176 -120
rect 19221 -135 19236 -120
rect 19281 -135 19296 -120
rect 19341 -135 19356 -120
rect 19401 -135 19416 -120
rect 19466 -135 19481 -120
rect 19526 -135 19541 -120
rect 19586 -135 19601 -120
rect 19646 -135 19661 -120
rect 19706 -135 19721 -120
rect 19766 -135 19781 -120
rect 19826 -135 19841 -120
rect 19886 -135 19901 -120
rect 19951 -135 19966 -120
rect 20011 -135 20026 -120
rect 20071 -135 20086 -120
rect 20131 -135 20146 -120
rect 20191 -135 20206 -120
rect 20251 -135 20266 -120
rect 20311 -135 20326 -120
rect 20371 -135 20386 -120
rect 20436 -135 20451 -120
rect 20496 -135 20511 -120
rect 20556 -135 20571 -120
rect 20616 -135 20631 -120
rect 20676 -135 20691 -120
rect 20736 -135 20751 -120
rect 20796 -135 20811 -120
rect 20856 -135 20871 -120
rect 20921 -135 20936 -120
rect 20981 -135 20996 -120
rect 21041 -135 21056 -120
rect 21101 -135 21116 -120
rect 0 -320 15 -305
rect 60 -320 75 -305
rect 120 -320 135 -305
rect 180 -320 195 -305
rect 240 -320 255 -305
rect 300 -320 315 -305
rect 360 -320 375 -305
rect 420 -320 435 -305
rect 480 -320 495 -305
rect 540 -320 555 -305
rect 600 -320 615 -305
rect 660 -320 675 -305
rect 720 -320 735 -305
rect 780 -320 795 -305
rect 840 -320 855 -305
rect 900 -320 915 -305
rect 960 -320 975 -305
rect 1020 -320 1035 -305
rect 1080 -320 1095 -305
rect 1140 -320 1155 -305
rect 1200 -320 1215 -305
rect 1260 -320 1275 -305
rect 1320 -320 1335 -305
rect 1380 -320 1395 -305
rect 1440 -320 1455 -305
rect 1500 -320 1515 -305
rect 1560 -320 1575 -305
rect 1620 -320 1635 -305
rect 1680 -320 1695 -305
rect 1740 -320 1755 -305
rect 1800 -320 1815 -305
rect 1860 -320 1875 -305
rect 1920 -320 1935 -305
rect 1980 -320 1995 -305
rect 2040 -320 2055 -305
rect 2100 -320 2115 -305
rect 2160 -320 2175 -305
rect 2220 -320 2235 -305
rect 2280 -320 2295 -305
rect 2340 -320 2355 -305
rect 2400 -320 2415 -305
rect 2460 -320 2475 -305
rect 2520 -320 2535 -305
rect 2580 -320 2595 -305
rect 2640 -320 2655 -305
rect 2700 -320 2715 -305
rect 2760 -320 2775 -305
rect 2820 -320 2835 -305
rect 2880 -320 2895 -305
rect 2940 -320 2955 -305
rect 3000 -320 3015 -305
rect 3060 -320 3075 -305
rect 3120 -320 3135 -305
rect 3180 -320 3195 -305
rect 3240 -320 3255 -305
rect 3300 -320 3315 -305
rect 3360 -320 3375 -305
rect 3420 -320 3435 -305
rect 3480 -320 3495 -305
rect 3540 -320 3555 -305
rect 3600 -320 3615 -305
rect 3660 -320 3675 -305
rect 3720 -320 3735 -305
rect 3780 -320 3795 -305
rect 3840 -320 3855 -305
rect 3900 -320 3915 -305
rect 3960 -320 3975 -305
rect 4020 -320 4035 -305
rect 4080 -320 4095 -305
rect 4140 -320 4155 -305
rect 4200 -320 4215 -305
rect 4260 -320 4275 -305
rect 4320 -320 4335 -305
rect 4380 -320 4395 -305
rect 4440 -320 4455 -305
rect 4500 -320 4515 -305
rect 4560 -320 4575 -305
rect 4620 -320 4635 -305
rect 4680 -320 4695 -305
rect 4740 -320 4755 -305
rect 4800 -320 4815 -305
rect 4860 -320 4875 -305
rect 4920 -320 4935 -305
rect 4980 -320 4995 -305
rect 5040 -320 5055 -305
rect 5100 -320 5115 -305
rect 5160 -320 5175 -305
rect 5220 -320 5235 -305
rect 5280 -320 5295 -305
rect 5340 -320 5355 -305
rect 5400 -320 5415 -305
rect 5460 -320 5475 -305
rect 5520 -320 5535 -305
rect 5580 -320 5595 -305
rect 5640 -320 5655 -305
rect 5700 -320 5715 -305
rect 5760 -320 5775 -305
rect 5820 -320 5835 -305
rect 5880 -320 5895 -305
rect 5940 -320 5955 -305
rect 6000 -320 6015 -305
rect 6060 -320 6075 -305
rect 6120 -320 6135 -305
rect 6180 -320 6195 -305
rect 6240 -320 6255 -305
rect 6300 -320 6315 -305
rect 6360 -320 6375 -305
rect 6420 -320 6435 -305
rect 6480 -320 6495 -305
rect 6540 -320 6555 -305
rect 6600 -320 6615 -305
rect 6660 -320 6675 -305
rect 6720 -320 6735 -305
rect 6780 -320 6795 -305
rect 6840 -320 6855 -305
rect 6900 -320 6915 -305
rect 6960 -320 6975 -305
rect 7020 -320 7035 -305
rect 7080 -320 7095 -305
rect 7140 -320 7155 -305
rect 7200 -320 7215 -305
rect 7260 -320 7275 -305
rect 7320 -320 7335 -305
rect 7380 -320 7395 -305
rect 7440 -320 7455 -305
rect 7500 -320 7515 -305
rect 7560 -320 7575 -305
rect 7620 -320 7635 -305
rect 7680 -320 7695 -305
rect 7740 -320 7755 -305
rect 7800 -320 7815 -305
rect 7860 -320 7875 -305
rect 7920 -320 7935 -305
rect 7980 -320 7995 -305
rect 8040 -320 8055 -305
rect 8100 -320 8115 -305
rect 8160 -320 8175 -305
rect 8220 -320 8235 -305
rect 8280 -320 8295 -305
rect 8340 -320 8355 -305
rect 8400 -320 8415 -305
rect 8460 -320 8475 -305
rect 8520 -320 8535 -305
rect 8580 -320 8595 -305
rect 8640 -320 8655 -305
rect 8700 -320 8715 -305
rect 8760 -320 8775 -305
rect 8820 -320 8835 -305
rect 8880 -320 8895 -305
rect 8940 -320 8955 -305
rect 9000 -320 9015 -305
rect 9060 -320 9075 -305
rect 9120 -320 9135 -305
rect 9180 -320 9195 -305
rect 9240 -320 9255 -305
rect 9300 -320 9315 -305
rect 9360 -320 9375 -305
rect 9420 -320 9435 -305
rect 9480 -320 9495 -305
rect 9540 -320 9555 -305
rect 9600 -320 9615 -305
rect 9660 -320 9675 -305
rect 9720 -320 9735 -305
rect 9780 -320 9795 -305
rect 9840 -320 9855 -305
rect 9900 -320 9915 -305
rect 9960 -320 9975 -305
rect 10020 -320 10035 -305
rect 10080 -320 10095 -305
rect 10140 -320 10155 -305
rect 10200 -320 10215 -305
rect 10260 -320 10275 -305
rect 10320 -320 10335 -305
rect 10380 -320 10395 -305
rect 10440 -320 10455 -305
rect 10500 -320 10515 -305
rect 10560 -320 10575 -305
rect 10620 -320 10635 -305
rect 10680 -320 10695 -305
rect 10740 -320 10755 -305
rect 10800 -320 10815 -305
rect 10860 -320 10875 -305
rect 10920 -320 10935 -305
rect 10980 -320 10995 -305
rect 11040 -320 11055 -305
rect 11100 -320 11115 -305
rect 11160 -320 11175 -305
rect 11220 -320 11235 -305
rect 11280 -320 11295 -305
rect 11340 -320 11355 -305
rect 11400 -320 11415 -305
rect 11460 -320 11475 -305
rect 11520 -320 11535 -305
rect 11580 -320 11595 -305
rect 11640 -320 11655 -305
rect 11700 -320 11715 -305
rect 11760 -320 11775 -305
rect 11820 -320 11835 -305
rect 11880 -320 11895 -305
rect 11940 -320 11955 -305
rect 12000 -320 12015 -305
rect 12060 -320 12075 -305
rect 12120 -320 12135 -305
rect 12180 -320 12195 -305
rect 12240 -320 12255 -305
rect 12300 -320 12315 -305
rect 12360 -320 12375 -305
rect 12420 -320 12435 -305
rect 12480 -320 12495 -305
rect 12540 -320 12555 -305
rect 12600 -320 12615 -305
rect 12660 -320 12675 -305
rect 12720 -320 12735 -305
rect 12780 -320 12795 -305
rect 12840 -320 12855 -305
rect 12900 -320 12915 -305
rect 12960 -320 12975 -305
rect 13020 -320 13035 -305
rect 13080 -320 13095 -305
rect 13140 -320 13155 -305
rect 13200 -320 13215 -305
rect 13260 -320 13275 -305
rect 13320 -320 13335 -305
rect 13380 -320 13395 -305
rect 13440 -320 13455 -305
rect 13500 -320 13515 -305
rect 13560 -320 13575 -305
rect 13620 -320 13635 -305
rect 13680 -320 13695 -305
rect 13740 -320 13755 -305
rect 13800 -320 13815 -305
rect 13860 -320 13875 -305
rect 13920 -320 13935 -305
rect 13980 -320 13995 -305
rect 14040 -320 14055 -305
rect 14100 -320 14115 -305
rect 14160 -320 14175 -305
rect 14220 -320 14235 -305
rect 14280 -320 14295 -305
rect 14340 -320 14355 -305
rect 14400 -320 14415 -305
rect 14460 -320 14475 -305
rect 14520 -320 14535 -305
rect 14580 -320 14595 -305
rect 14640 -320 14655 -305
rect 14700 -320 14715 -305
rect 14760 -320 14775 -305
rect 14820 -320 14835 -305
rect 14880 -320 14895 -305
rect 14940 -320 14955 -305
rect 15000 -320 15015 -305
rect 15060 -320 15075 -305
rect 15120 -320 15135 -305
rect 15180 -320 15195 -305
rect 15240 -320 15255 -305
rect 15300 -320 15315 -305
rect 15360 -320 15375 -305
rect 15420 -320 15435 -305
rect 15480 -320 15495 -305
rect 15540 -320 15555 -305
rect 15600 -320 15615 -305
rect 15660 -320 15675 -305
rect 15720 -320 15735 -305
rect 15780 -320 15795 -305
rect 15840 -320 15855 -305
rect 15900 -320 15915 -305
rect 15960 -320 15975 -305
rect 16020 -320 16035 -305
rect 16080 -320 16095 -305
rect 16140 -320 16155 -305
rect 16200 -320 16215 -305
rect 16260 -320 16275 -305
rect 16320 -320 16335 -305
rect 16380 -320 16395 -305
rect 16440 -320 16455 -305
rect 16500 -320 16515 -305
rect 16560 -320 16575 -305
rect 16620 -320 16635 -305
rect 16680 -320 16695 -305
rect 16740 -320 16755 -305
rect 16800 -320 16815 -305
rect 16860 -320 16875 -305
rect 16920 -320 16935 -305
rect 16980 -320 16995 -305
rect 17040 -320 17055 -305
rect 17100 -320 17115 -305
rect 17160 -320 17175 -305
rect 17220 -320 17235 -305
rect 17280 -320 17295 -305
rect 17340 -320 17355 -305
rect 17400 -320 17415 -305
rect 17460 -320 17475 -305
rect 17520 -320 17535 -305
rect 17580 -320 17595 -305
rect 17640 -320 17655 -305
rect 17700 -320 17715 -305
rect 17760 -320 17775 -305
rect 17820 -320 17835 -305
rect 17880 -320 17895 -305
rect 17940 -320 17955 -305
rect 18000 -320 18015 -305
rect 18060 -320 18075 -305
rect 18120 -320 18135 -305
rect 18180 -320 18195 -305
rect 18240 -320 18255 -305
rect 18300 -320 18315 -305
rect 18360 -320 18375 -305
rect 18420 -320 18435 -305
rect 18480 -320 18495 -305
rect 18540 -320 18555 -305
rect 18600 -320 18615 -305
rect 18660 -320 18675 -305
rect 18720 -320 18735 -305
rect 18780 -320 18795 -305
rect 18840 -320 18855 -305
rect 18900 -320 18915 -305
rect 18960 -320 18975 -305
rect 19020 -320 19035 -305
rect 19080 -320 19095 -305
rect 19140 -320 19155 -305
rect 19200 -320 19215 -305
rect 19260 -320 19275 -305
rect 19320 -320 19335 -305
rect 19380 -320 19395 -305
rect 19440 -320 19455 -305
rect 19500 -320 19515 -305
rect 19560 -320 19575 -305
rect 19620 -320 19635 -305
rect 19680 -320 19695 -305
rect 19740 -320 19755 -305
rect 19800 -320 19815 -305
rect 19860 -320 19875 -305
rect 19920 -320 19935 -305
rect 19980 -320 19995 -305
rect 20040 -320 20055 -305
rect 20100 -320 20115 -305
rect 20160 -320 20175 -305
rect 20220 -320 20235 -305
rect 20280 -320 20295 -305
rect 20340 -320 20355 -305
rect 20400 -320 20415 -305
rect 20460 -320 20475 -305
rect 20520 -320 20535 -305
rect 20580 -320 20595 -305
rect 20640 -320 20655 -305
rect 20700 -320 20715 -305
rect 20760 -320 20775 -305
rect 20820 -320 20835 -305
rect 20880 -320 20895 -305
rect 20940 -320 20955 -305
rect 21000 -320 21015 -305
rect 21060 -320 21075 -305
rect 21120 -320 21135 -305
rect 21180 -320 21195 -305
rect 21240 -320 21255 -305
rect 21300 -320 21315 -305
rect 21360 -320 21375 -305
rect 21420 -320 21435 -305
rect 21480 -320 21495 -305
rect 21540 -320 21555 -305
rect 21600 -320 21615 -305
rect 21660 -320 21675 -305
rect 21720 -320 21735 -305
rect 21780 -320 21795 -305
rect 21840 -320 21855 -305
rect 21900 -320 21915 -305
rect 21960 -320 21975 -305
rect 22020 -320 22035 -305
rect 22080 -320 22095 -305
rect 22140 -320 22155 -305
rect 22200 -320 22215 -305
rect 22260 -320 22275 -305
rect 22320 -320 22335 -305
rect 22380 -320 22395 -305
rect 22440 -320 22455 -305
rect 22500 -320 22515 -305
rect 22560 -320 22575 -305
rect 22620 -320 22635 -305
rect 22680 -320 22695 -305
rect 22740 -320 22755 -305
rect 22800 -320 22815 -305
rect 22860 -320 22875 -305
rect 22920 -320 22935 -305
rect 22980 -320 22995 -305
rect 23040 -320 23055 -305
rect 23100 -320 23115 -305
rect 23160 -320 23175 -305
rect 23220 -320 23235 -305
rect 23280 -320 23295 -305
rect 23340 -320 23355 -305
rect 23400 -320 23415 -305
rect 23460 -320 23475 -305
rect 23520 -320 23535 -305
rect 23580 -320 23595 -305
rect 23640 -320 23655 -305
rect 23700 -320 23715 -305
rect 23760 -320 23775 -305
rect 23820 -320 23835 -305
rect 23880 -320 23895 -305
rect 23940 -320 23955 -305
rect 24000 -320 24015 -305
rect 24060 -320 24075 -305
rect 24120 -320 24135 -305
rect 24180 -320 24195 -305
rect 24240 -320 24255 -305
rect 24300 -320 24315 -305
rect 24360 -320 24375 -305
rect 24420 -320 24435 -305
rect 24480 -320 24495 -305
rect 24540 -320 24555 -305
rect 24600 -320 24615 -305
rect 24660 -320 24675 -305
rect 24720 -320 24735 -305
rect 24780 -320 24795 -305
rect 24840 -320 24855 -305
rect 24900 -320 24915 -305
rect 24960 -320 24975 -305
rect 25020 -320 25035 -305
rect 25080 -320 25095 -305
rect 25140 -320 25155 -305
rect 25200 -320 25215 -305
rect 25260 -320 25275 -305
rect 25320 -320 25335 -305
rect 25380 -320 25395 -305
rect 25440 -320 25455 -305
rect 25500 -320 25515 -305
rect 25560 -320 25575 -305
rect 25620 -320 25635 -305
rect 25680 -320 25695 -305
rect 25740 -320 25755 -305
rect 25800 -320 25815 -305
rect 25860 -320 25875 -305
rect 25920 -320 25935 -305
rect 25980 -320 25995 -305
rect 26040 -320 26055 -305
rect 26100 -320 26115 -305
rect 26160 -320 26175 -305
rect 26220 -320 26235 -305
rect 26280 -320 26295 -305
rect 26340 -320 26355 -305
rect 26400 -320 26415 -305
rect 26460 -320 26475 -305
rect 26520 -320 26535 -305
rect 26580 -320 26595 -305
rect 26640 -320 26655 -305
rect 26700 -320 26715 -305
rect 26760 -320 26775 -305
rect 26820 -320 26835 -305
rect 26880 -320 26895 -305
rect 26940 -320 26955 -305
rect 27000 -320 27015 -305
rect 27060 -320 27075 -305
rect 27120 -320 27135 -305
rect 27180 -320 27195 -305
rect 27240 -320 27255 -305
rect 27300 -320 27315 -305
rect 27360 -320 27375 -305
rect 27420 -320 27435 -305
rect 27480 -320 27495 -305
rect 27540 -320 27555 -305
rect 27600 -320 27615 -305
rect 27660 -320 27675 -305
rect 27720 -320 27735 -305
rect 27780 -320 27795 -305
rect 27840 -320 27855 -305
rect 27900 -320 27915 -305
rect 27960 -320 27975 -305
rect 28020 -320 28035 -305
rect 28080 -320 28095 -305
rect 28140 -320 28155 -305
rect 28200 -320 28215 -305
rect 28260 -320 28275 -305
rect 28320 -320 28335 -305
rect 28380 -320 28395 -305
rect 28440 -320 28455 -305
rect 28500 -320 28515 -305
rect 28560 -320 28575 -305
rect 28620 -320 28635 -305
rect 28680 -320 28695 -305
rect 28740 -320 28755 -305
rect 28800 -320 28815 -305
rect 28860 -320 28875 -305
rect 28920 -320 28935 -305
rect 28980 -320 28995 -305
rect 29040 -320 29055 -305
rect 29100 -320 29115 -305
rect 29160 -320 29175 -305
rect 29220 -320 29235 -305
rect 29280 -320 29295 -305
rect 29340 -320 29355 -305
rect 29400 -320 29415 -305
rect 29460 -320 29475 -305
rect 29520 -320 29535 -305
rect 29580 -320 29595 -305
rect 29640 -320 29655 -305
rect 29700 -320 29715 -305
rect 29760 -320 29775 -305
rect 29820 -320 29835 -305
rect 29880 -320 29895 -305
rect 29940 -320 29955 -305
rect 30000 -320 30015 -305
rect 30060 -320 30075 -305
rect 30120 -320 30135 -305
rect 30180 -320 30195 -305
rect 30240 -320 30255 -305
rect 30300 -320 30315 -305
rect 30360 -320 30375 -305
rect 30420 -320 30435 -305
rect 30480 -320 30495 -305
rect 30540 -320 30555 -305
rect 30600 -320 30615 -305
rect 30660 -320 30675 -305
rect 0 -575 15 -420
rect 60 -575 75 -420
rect 120 -575 135 -420
rect 180 -575 195 -420
rect 240 -575 255 -420
rect 300 -575 315 -420
rect 360 -575 375 -420
rect 420 -575 435 -420
rect 480 -575 495 -420
rect 540 -575 555 -420
rect 600 -575 615 -420
rect 660 -575 675 -420
rect 720 -575 735 -420
rect 780 -575 795 -420
rect 840 -575 855 -420
rect 900 -575 915 -420
rect 960 -575 975 -420
rect 1020 -575 1035 -420
rect 1080 -575 1095 -420
rect 1140 -575 1155 -420
rect 1200 -575 1215 -420
rect 1260 -575 1275 -420
rect 1320 -575 1335 -420
rect 1380 -575 1395 -420
rect 1440 -575 1455 -420
rect 1500 -575 1515 -420
rect 1560 -575 1575 -420
rect 1620 -575 1635 -420
rect 1680 -575 1695 -420
rect 1740 -575 1755 -420
rect 1800 -575 1815 -420
rect 1860 -575 1875 -420
rect 1920 -575 1935 -420
rect 1980 -575 1995 -420
rect 2040 -575 2055 -420
rect 2100 -575 2115 -420
rect 2160 -575 2175 -420
rect 2220 -575 2235 -420
rect 2280 -575 2295 -420
rect 2340 -575 2355 -420
rect 2400 -575 2415 -420
rect 2460 -575 2475 -420
rect 2520 -575 2535 -420
rect 2580 -575 2595 -420
rect 2640 -575 2655 -420
rect 2700 -575 2715 -420
rect 2760 -575 2775 -420
rect 2820 -575 2835 -420
rect 2880 -575 2895 -420
rect 2940 -575 2955 -420
rect 3000 -575 3015 -420
rect 3060 -575 3075 -420
rect 3120 -575 3135 -420
rect 3180 -575 3195 -420
rect 3240 -575 3255 -420
rect 3300 -575 3315 -420
rect 3360 -575 3375 -420
rect 3420 -575 3435 -420
rect 3480 -575 3495 -420
rect 3540 -575 3555 -420
rect 3600 -575 3615 -420
rect 3660 -575 3675 -420
rect 3720 -575 3735 -420
rect 3780 -575 3795 -420
rect 3840 -575 3855 -420
rect 3900 -575 3915 -420
rect 3960 -575 3975 -420
rect 4020 -575 4035 -420
rect 4080 -575 4095 -420
rect 4140 -575 4155 -420
rect 4200 -575 4215 -420
rect 4260 -575 4275 -420
rect 4320 -575 4335 -420
rect 4380 -575 4395 -420
rect 4440 -575 4455 -420
rect 4500 -575 4515 -420
rect 4560 -575 4575 -420
rect 4620 -575 4635 -420
rect 4680 -575 4695 -420
rect 4740 -575 4755 -420
rect 4800 -575 4815 -420
rect 4860 -575 4875 -420
rect 4920 -575 4935 -420
rect 4980 -575 4995 -420
rect 5040 -575 5055 -420
rect 5100 -575 5115 -420
rect 5160 -575 5175 -420
rect 5220 -575 5235 -420
rect 5280 -575 5295 -420
rect 5340 -575 5355 -420
rect 5400 -575 5415 -420
rect 5460 -575 5475 -420
rect 5520 -575 5535 -420
rect 5580 -575 5595 -420
rect 5640 -575 5655 -420
rect 5700 -575 5715 -420
rect 5760 -575 5775 -420
rect 5820 -575 5835 -420
rect 5880 -575 5895 -420
rect 5940 -575 5955 -420
rect 6000 -575 6015 -420
rect 6060 -575 6075 -420
rect 6120 -575 6135 -420
rect 6180 -575 6195 -420
rect 6240 -575 6255 -420
rect 6300 -575 6315 -420
rect 6360 -575 6375 -420
rect 6420 -575 6435 -420
rect 6480 -575 6495 -420
rect 6540 -575 6555 -420
rect 6600 -575 6615 -420
rect 6660 -575 6675 -420
rect 6720 -575 6735 -420
rect 6780 -575 6795 -420
rect 6840 -575 6855 -420
rect 6900 -575 6915 -420
rect 6960 -575 6975 -420
rect 7020 -575 7035 -420
rect 7080 -575 7095 -420
rect 7140 -575 7155 -420
rect 7200 -575 7215 -420
rect 7260 -575 7275 -420
rect 7320 -575 7335 -420
rect 7380 -575 7395 -420
rect 7440 -575 7455 -420
rect 7500 -575 7515 -420
rect 7560 -575 7575 -420
rect 7620 -575 7635 -420
rect 7680 -575 7695 -420
rect 7740 -575 7755 -420
rect 7800 -575 7815 -420
rect 7860 -575 7875 -420
rect 7920 -575 7935 -420
rect 7980 -575 7995 -420
rect 8040 -575 8055 -420
rect 8100 -575 8115 -420
rect 8160 -575 8175 -420
rect 8220 -575 8235 -420
rect 8280 -575 8295 -420
rect 8340 -575 8355 -420
rect 8400 -575 8415 -420
rect 8460 -575 8475 -420
rect 8520 -575 8535 -420
rect 8580 -575 8595 -420
rect 8640 -575 8655 -420
rect 8700 -575 8715 -420
rect 8760 -575 8775 -420
rect 8820 -575 8835 -420
rect 8880 -575 8895 -420
rect 8940 -575 8955 -420
rect 9000 -575 9015 -420
rect 9060 -575 9075 -420
rect 9120 -575 9135 -420
rect 9180 -575 9195 -420
rect 9240 -575 9255 -420
rect 9300 -575 9315 -420
rect 9360 -575 9375 -420
rect 9420 -575 9435 -420
rect 9480 -575 9495 -420
rect 9540 -575 9555 -420
rect 9600 -575 9615 -420
rect 9660 -575 9675 -420
rect 9720 -575 9735 -420
rect 9780 -575 9795 -420
rect 9840 -575 9855 -420
rect 9900 -575 9915 -420
rect 9960 -575 9975 -420
rect 10020 -575 10035 -420
rect 10080 -575 10095 -420
rect 10140 -575 10155 -420
rect 10200 -575 10215 -420
rect 10260 -575 10275 -420
rect 10320 -575 10335 -420
rect 10380 -575 10395 -420
rect 10440 -575 10455 -420
rect 10500 -575 10515 -420
rect 10560 -575 10575 -420
rect 10620 -575 10635 -420
rect 10680 -575 10695 -420
rect 10740 -575 10755 -420
rect 10800 -575 10815 -420
rect 10860 -575 10875 -420
rect 10920 -575 10935 -420
rect 10980 -575 10995 -420
rect 11040 -575 11055 -420
rect 11100 -575 11115 -420
rect 11160 -575 11175 -420
rect 11220 -575 11235 -420
rect 11280 -575 11295 -420
rect 11340 -575 11355 -420
rect 11400 -575 11415 -420
rect 11460 -575 11475 -420
rect 11520 -575 11535 -420
rect 11580 -575 11595 -420
rect 11640 -575 11655 -420
rect 11700 -575 11715 -420
rect 11760 -575 11775 -420
rect 11820 -575 11835 -420
rect 11880 -575 11895 -420
rect 11940 -575 11955 -420
rect 12000 -575 12015 -420
rect 12060 -575 12075 -420
rect 12120 -575 12135 -420
rect 12180 -575 12195 -420
rect 12240 -575 12255 -420
rect 12300 -575 12315 -420
rect 12360 -575 12375 -420
rect 12420 -575 12435 -420
rect 12480 -575 12495 -420
rect 12540 -575 12555 -420
rect 12600 -575 12615 -420
rect 12660 -575 12675 -420
rect 12720 -575 12735 -420
rect 12780 -575 12795 -420
rect 12840 -575 12855 -420
rect 12900 -575 12915 -420
rect 12960 -575 12975 -420
rect 13020 -575 13035 -420
rect 13080 -575 13095 -420
rect 13140 -575 13155 -420
rect 13200 -575 13215 -420
rect 13260 -575 13275 -420
rect 13320 -575 13335 -420
rect 13380 -575 13395 -420
rect 13440 -575 13455 -420
rect 13500 -575 13515 -420
rect 13560 -575 13575 -420
rect 13620 -575 13635 -420
rect 13680 -575 13695 -420
rect 13740 -575 13755 -420
rect 13800 -575 13815 -420
rect 13860 -575 13875 -420
rect 13920 -575 13935 -420
rect 13980 -575 13995 -420
rect 14040 -575 14055 -420
rect 14100 -575 14115 -420
rect 14160 -575 14175 -420
rect 14220 -575 14235 -420
rect 14280 -575 14295 -420
rect 14340 -575 14355 -420
rect 14400 -575 14415 -420
rect 14460 -575 14475 -420
rect 14520 -575 14535 -420
rect 14580 -575 14595 -420
rect 14640 -575 14655 -420
rect 14700 -575 14715 -420
rect 14760 -575 14775 -420
rect 14820 -575 14835 -420
rect 14880 -575 14895 -420
rect 14940 -575 14955 -420
rect 15000 -575 15015 -420
rect 15060 -575 15075 -420
rect 15120 -575 15135 -420
rect 15180 -575 15195 -420
rect 15240 -575 15255 -420
rect 15300 -575 15315 -420
rect 15360 -575 15375 -420
rect 15420 -575 15435 -420
rect 15480 -575 15495 -420
rect 15540 -575 15555 -420
rect 15600 -575 15615 -420
rect 15660 -575 15675 -420
rect 15720 -575 15735 -420
rect 15780 -575 15795 -420
rect 15840 -575 15855 -420
rect 15900 -575 15915 -420
rect 15960 -575 15975 -420
rect 16020 -575 16035 -420
rect 16080 -575 16095 -420
rect 16140 -575 16155 -420
rect 16200 -575 16215 -420
rect 16260 -575 16275 -420
rect 16320 -575 16335 -420
rect 16380 -575 16395 -420
rect 16440 -575 16455 -420
rect 16500 -575 16515 -420
rect 16560 -575 16575 -420
rect 16620 -575 16635 -420
rect 16680 -575 16695 -420
rect 16740 -575 16755 -420
rect 16800 -575 16815 -420
rect 16860 -575 16875 -420
rect 16920 -575 16935 -420
rect 16980 -575 16995 -420
rect 17040 -575 17055 -420
rect 17100 -575 17115 -420
rect 17160 -575 17175 -420
rect 17220 -575 17235 -420
rect 17280 -575 17295 -420
rect 17340 -575 17355 -420
rect 17400 -575 17415 -420
rect 17460 -575 17475 -420
rect 17520 -575 17535 -420
rect 17580 -575 17595 -420
rect 17640 -575 17655 -420
rect 17700 -575 17715 -420
rect 17760 -575 17775 -420
rect 17820 -575 17835 -420
rect 17880 -575 17895 -420
rect 17940 -575 17955 -420
rect 18000 -575 18015 -420
rect 18060 -575 18075 -420
rect 18120 -575 18135 -420
rect 18180 -575 18195 -420
rect 18240 -575 18255 -420
rect 18300 -575 18315 -420
rect 18360 -575 18375 -420
rect 18420 -575 18435 -420
rect 18480 -575 18495 -420
rect 18540 -575 18555 -420
rect 18600 -575 18615 -420
rect 18660 -575 18675 -420
rect 18720 -575 18735 -420
rect 18780 -575 18795 -420
rect 18840 -575 18855 -420
rect 18900 -575 18915 -420
rect 18960 -575 18975 -420
rect 19020 -575 19035 -420
rect 19080 -575 19095 -420
rect 19140 -575 19155 -420
rect 19200 -575 19215 -420
rect 19260 -575 19275 -420
rect 19320 -575 19335 -420
rect 19380 -575 19395 -420
rect 19440 -575 19455 -420
rect 19500 -575 19515 -420
rect 19560 -575 19575 -420
rect 19620 -575 19635 -420
rect 19680 -575 19695 -420
rect 19740 -575 19755 -420
rect 19800 -575 19815 -420
rect 19860 -575 19875 -420
rect 19920 -575 19935 -420
rect 19980 -575 19995 -420
rect 20040 -575 20055 -420
rect 20100 -575 20115 -420
rect 20160 -575 20175 -420
rect 20220 -575 20235 -420
rect 20280 -575 20295 -420
rect 20340 -575 20355 -420
rect 20400 -575 20415 -420
rect 20460 -575 20475 -420
rect 20520 -575 20535 -420
rect 20580 -575 20595 -420
rect 20640 -575 20655 -420
rect 20700 -575 20715 -420
rect 20760 -575 20775 -420
rect 20820 -575 20835 -420
rect 20880 -575 20895 -420
rect 20940 -575 20955 -420
rect 21000 -575 21015 -420
rect 21060 -575 21075 -420
rect 21120 -575 21135 -420
rect 21180 -575 21195 -420
rect 21240 -575 21255 -420
rect 21300 -575 21315 -420
rect 21360 -575 21375 -420
rect 21420 -575 21435 -420
rect 21480 -575 21495 -420
rect 21540 -575 21555 -420
rect 21600 -575 21615 -420
rect 21660 -575 21675 -420
rect 21720 -575 21735 -420
rect 21780 -575 21795 -420
rect 21840 -575 21855 -420
rect 21900 -575 21915 -420
rect 21960 -575 21975 -420
rect 22020 -575 22035 -420
rect 22080 -575 22095 -420
rect 22140 -575 22155 -420
rect 22200 -575 22215 -420
rect 22260 -575 22275 -420
rect 22320 -575 22335 -420
rect 22380 -575 22395 -420
rect 22440 -575 22455 -420
rect 22500 -575 22515 -420
rect 22560 -575 22575 -420
rect 22620 -575 22635 -420
rect 22680 -575 22695 -420
rect 22740 -575 22755 -420
rect 22800 -575 22815 -420
rect 22860 -575 22875 -420
rect 22920 -575 22935 -420
rect 22980 -575 22995 -420
rect 23040 -575 23055 -420
rect 23100 -575 23115 -420
rect 23160 -575 23175 -420
rect 23220 -575 23235 -420
rect 23280 -575 23295 -420
rect 23340 -575 23355 -420
rect 23400 -575 23415 -420
rect 23460 -575 23475 -420
rect 23520 -575 23535 -420
rect 23580 -575 23595 -420
rect 23640 -575 23655 -420
rect 23700 -575 23715 -420
rect 23760 -575 23775 -420
rect 23820 -575 23835 -420
rect 23880 -575 23895 -420
rect 23940 -575 23955 -420
rect 24000 -575 24015 -420
rect 24060 -575 24075 -420
rect 24120 -575 24135 -420
rect 24180 -575 24195 -420
rect 24240 -575 24255 -420
rect 24300 -575 24315 -420
rect 24360 -575 24375 -420
rect 24420 -575 24435 -420
rect 24480 -575 24495 -420
rect 24540 -575 24555 -420
rect 24600 -575 24615 -420
rect 24660 -575 24675 -420
rect 24720 -575 24735 -420
rect 24780 -575 24795 -420
rect 24840 -575 24855 -420
rect 24900 -575 24915 -420
rect 24960 -575 24975 -420
rect 25020 -575 25035 -420
rect 25080 -575 25095 -420
rect 25140 -575 25155 -420
rect 25200 -575 25215 -420
rect 25260 -575 25275 -420
rect 25320 -575 25335 -420
rect 25380 -575 25395 -420
rect 25440 -575 25455 -420
rect 25500 -575 25515 -420
rect 25560 -575 25575 -420
rect 25620 -575 25635 -420
rect 25680 -575 25695 -420
rect 25740 -575 25755 -420
rect 25800 -575 25815 -420
rect 25860 -575 25875 -420
rect 25920 -575 25935 -420
rect 25980 -575 25995 -420
rect 26040 -575 26055 -420
rect 26100 -575 26115 -420
rect 26160 -575 26175 -420
rect 26220 -575 26235 -420
rect 26280 -575 26295 -420
rect 26340 -575 26355 -420
rect 26400 -575 26415 -420
rect 26460 -575 26475 -420
rect 26520 -575 26535 -420
rect 26580 -575 26595 -420
rect 26640 -575 26655 -420
rect 26700 -575 26715 -420
rect 26760 -575 26775 -420
rect 26820 -575 26835 -420
rect 26880 -575 26895 -420
rect 26940 -575 26955 -420
rect 27000 -575 27015 -420
rect 27060 -575 27075 -420
rect 27120 -575 27135 -420
rect 27180 -575 27195 -420
rect 27240 -575 27255 -420
rect 27300 -575 27315 -420
rect 27360 -575 27375 -420
rect 27420 -575 27435 -420
rect 27480 -575 27495 -420
rect 27540 -575 27555 -420
rect 27600 -575 27615 -420
rect 27660 -575 27675 -420
rect 27720 -575 27735 -420
rect 27780 -575 27795 -420
rect 27840 -575 27855 -420
rect 27900 -575 27915 -420
rect 27960 -575 27975 -420
rect 28020 -575 28035 -420
rect 28080 -575 28095 -420
rect 28140 -575 28155 -420
rect 28200 -575 28215 -420
rect 28260 -575 28275 -420
rect 28320 -575 28335 -420
rect 28380 -575 28395 -420
rect 28440 -575 28455 -420
rect 28500 -575 28515 -420
rect 28560 -575 28575 -420
rect 28620 -575 28635 -420
rect 28680 -575 28695 -420
rect 28740 -575 28755 -420
rect 28800 -575 28815 -420
rect 28860 -575 28875 -420
rect 28920 -575 28935 -420
rect 28980 -575 28995 -420
rect 29040 -575 29055 -420
rect 29100 -575 29115 -420
rect 29160 -575 29175 -420
rect 29220 -575 29235 -420
rect 29280 -575 29295 -420
rect 29340 -575 29355 -420
rect 29400 -575 29415 -420
rect 29460 -575 29475 -420
rect 29520 -575 29535 -420
rect 29580 -575 29595 -420
rect 29640 -575 29655 -420
rect 29700 -575 29715 -420
rect 29760 -575 29775 -420
rect 29820 -575 29835 -420
rect 29880 -575 29895 -420
rect 29940 -575 29955 -420
rect 30000 -575 30015 -420
rect 30060 -575 30075 -420
rect 30120 -575 30135 -420
rect 30180 -575 30195 -420
rect 30240 -575 30255 -420
rect 30300 -575 30315 -420
rect 30360 -575 30375 -420
rect 30420 -575 30435 -420
rect 30480 -575 30495 -420
rect 30540 -575 30555 -420
rect 30600 -575 30615 -420
rect 30660 -475 30675 -420
rect 30660 -485 30715 -475
rect 30660 -505 30685 -485
rect 30705 -505 30715 -485
rect 30660 -515 30715 -505
rect 30660 -575 30675 -515
rect 0 -785 15 -770
rect 60 -785 75 -770
rect 120 -785 135 -770
rect 180 -785 195 -770
rect 240 -785 255 -770
rect 300 -785 315 -770
rect 360 -785 375 -770
rect 420 -785 435 -770
rect 480 -785 495 -770
rect 540 -785 555 -770
rect 600 -785 615 -770
rect 660 -785 675 -770
rect 720 -785 735 -770
rect 780 -785 795 -770
rect 840 -785 855 -770
rect 900 -785 915 -770
rect 960 -785 975 -770
rect 1020 -785 1035 -770
rect 1080 -785 1095 -770
rect 1140 -785 1155 -770
rect 1200 -785 1215 -770
rect 1260 -785 1275 -770
rect 1320 -785 1335 -770
rect 1380 -785 1395 -770
rect 1440 -785 1455 -770
rect 1500 -785 1515 -770
rect 1560 -785 1575 -770
rect 1620 -785 1635 -770
rect 1680 -785 1695 -770
rect 1740 -785 1755 -770
rect 1800 -785 1815 -770
rect 1860 -785 1875 -770
rect 1920 -785 1935 -770
rect 1980 -785 1995 -770
rect 2040 -785 2055 -770
rect 2100 -785 2115 -770
rect 2160 -785 2175 -770
rect 2220 -785 2235 -770
rect 2280 -785 2295 -770
rect 2340 -785 2355 -770
rect 2400 -785 2415 -770
rect 2460 -785 2475 -770
rect 2520 -785 2535 -770
rect 2580 -785 2595 -770
rect 2640 -785 2655 -770
rect 2700 -785 2715 -770
rect 2760 -785 2775 -770
rect 2820 -785 2835 -770
rect 2880 -785 2895 -770
rect 2940 -785 2955 -770
rect 3000 -785 3015 -770
rect 3060 -785 3075 -770
rect 3120 -785 3135 -770
rect 3180 -785 3195 -770
rect 3240 -785 3255 -770
rect 3300 -785 3315 -770
rect 3360 -785 3375 -770
rect 3420 -785 3435 -770
rect 3480 -785 3495 -770
rect 3540 -785 3555 -770
rect 3600 -785 3615 -770
rect 3660 -785 3675 -770
rect 3720 -785 3735 -770
rect 3780 -785 3795 -770
rect 3840 -785 3855 -770
rect 3900 -785 3915 -770
rect 3960 -785 3975 -770
rect 4020 -785 4035 -770
rect 4080 -785 4095 -770
rect 4140 -785 4155 -770
rect 4200 -785 4215 -770
rect 4260 -785 4275 -770
rect 4320 -785 4335 -770
rect 4380 -785 4395 -770
rect 4440 -785 4455 -770
rect 4500 -785 4515 -770
rect 4560 -785 4575 -770
rect 4620 -785 4635 -770
rect 4680 -785 4695 -770
rect 4740 -785 4755 -770
rect 4800 -785 4815 -770
rect 4860 -785 4875 -770
rect 4920 -785 4935 -770
rect 4980 -785 4995 -770
rect 5040 -785 5055 -770
rect 5100 -785 5115 -770
rect 5160 -785 5175 -770
rect 5220 -785 5235 -770
rect 5280 -785 5295 -770
rect 5340 -785 5355 -770
rect 5400 -785 5415 -770
rect 5460 -785 5475 -770
rect 5520 -785 5535 -770
rect 5580 -785 5595 -770
rect 5640 -785 5655 -770
rect 5700 -785 5715 -770
rect 5760 -785 5775 -770
rect 5820 -785 5835 -770
rect 5880 -785 5895 -770
rect 5940 -785 5955 -770
rect 6000 -785 6015 -770
rect 6060 -785 6075 -770
rect 6120 -785 6135 -770
rect 6180 -785 6195 -770
rect 6240 -785 6255 -770
rect 6300 -785 6315 -770
rect 6360 -785 6375 -770
rect 6420 -785 6435 -770
rect 6480 -785 6495 -770
rect 6540 -785 6555 -770
rect 6600 -785 6615 -770
rect 6660 -785 6675 -770
rect 6720 -785 6735 -770
rect 6780 -785 6795 -770
rect 6840 -785 6855 -770
rect 6900 -785 6915 -770
rect 6960 -785 6975 -770
rect 7020 -785 7035 -770
rect 7080 -785 7095 -770
rect 7140 -785 7155 -770
rect 7200 -785 7215 -770
rect 7260 -785 7275 -770
rect 7320 -785 7335 -770
rect 7380 -785 7395 -770
rect 7440 -785 7455 -770
rect 7500 -785 7515 -770
rect 7560 -785 7575 -770
rect 7620 -785 7635 -770
rect 7680 -785 7695 -770
rect 7740 -785 7755 -770
rect 7800 -785 7815 -770
rect 7860 -785 7875 -770
rect 7920 -785 7935 -770
rect 7980 -785 7995 -770
rect 8040 -785 8055 -770
rect 8100 -785 8115 -770
rect 8160 -785 8175 -770
rect 8220 -785 8235 -770
rect 8280 -785 8295 -770
rect 8340 -785 8355 -770
rect 8400 -785 8415 -770
rect 8460 -785 8475 -770
rect 8520 -785 8535 -770
rect 8580 -785 8595 -770
rect 8640 -785 8655 -770
rect 8700 -785 8715 -770
rect 8760 -785 8775 -770
rect 8820 -785 8835 -770
rect 8880 -785 8895 -770
rect 8940 -785 8955 -770
rect 9000 -785 9015 -770
rect 9060 -785 9075 -770
rect 9120 -785 9135 -770
rect 9180 -785 9195 -770
rect 9240 -785 9255 -770
rect 9300 -785 9315 -770
rect 9360 -785 9375 -770
rect 9420 -785 9435 -770
rect 9480 -785 9495 -770
rect 9540 -785 9555 -770
rect 9600 -785 9615 -770
rect 9660 -785 9675 -770
rect 9720 -785 9735 -770
rect 9780 -785 9795 -770
rect 9840 -785 9855 -770
rect 9900 -785 9915 -770
rect 9960 -785 9975 -770
rect 10020 -785 10035 -770
rect 10080 -785 10095 -770
rect 10140 -785 10155 -770
rect 10200 -785 10215 -770
rect 10260 -785 10275 -770
rect 10320 -785 10335 -770
rect 10380 -785 10395 -770
rect 10440 -785 10455 -770
rect 10500 -785 10515 -770
rect 10560 -785 10575 -770
rect 10620 -785 10635 -770
rect 10680 -785 10695 -770
rect 10740 -785 10755 -770
rect 10800 -785 10815 -770
rect 10860 -785 10875 -770
rect 10920 -785 10935 -770
rect 10980 -785 10995 -770
rect 11040 -785 11055 -770
rect 11100 -785 11115 -770
rect 11160 -785 11175 -770
rect 11220 -785 11235 -770
rect 11280 -785 11295 -770
rect 11340 -785 11355 -770
rect 11400 -785 11415 -770
rect 11460 -785 11475 -770
rect 11520 -785 11535 -770
rect 11580 -785 11595 -770
rect 11640 -785 11655 -770
rect 11700 -785 11715 -770
rect 11760 -785 11775 -770
rect 11820 -785 11835 -770
rect 11880 -785 11895 -770
rect 11940 -785 11955 -770
rect 12000 -785 12015 -770
rect 12060 -785 12075 -770
rect 12120 -785 12135 -770
rect 12180 -785 12195 -770
rect 12240 -785 12255 -770
rect 12300 -785 12315 -770
rect 12360 -785 12375 -770
rect 12420 -785 12435 -770
rect 12480 -785 12495 -770
rect 12540 -785 12555 -770
rect 12600 -785 12615 -770
rect 12660 -785 12675 -770
rect 12720 -785 12735 -770
rect 12780 -785 12795 -770
rect 12840 -785 12855 -770
rect 12900 -785 12915 -770
rect 12960 -785 12975 -770
rect 13020 -785 13035 -770
rect 13080 -785 13095 -770
rect 13140 -785 13155 -770
rect 13200 -785 13215 -770
rect 13260 -785 13275 -770
rect 13320 -785 13335 -770
rect 13380 -785 13395 -770
rect 13440 -785 13455 -770
rect 13500 -785 13515 -770
rect 13560 -785 13575 -770
rect 13620 -785 13635 -770
rect 13680 -785 13695 -770
rect 13740 -785 13755 -770
rect 13800 -785 13815 -770
rect 13860 -785 13875 -770
rect 13920 -785 13935 -770
rect 13980 -785 13995 -770
rect 14040 -785 14055 -770
rect 14100 -785 14115 -770
rect 14160 -785 14175 -770
rect 14220 -785 14235 -770
rect 14280 -785 14295 -770
rect 14340 -785 14355 -770
rect 14400 -785 14415 -770
rect 14460 -785 14475 -770
rect 14520 -785 14535 -770
rect 14580 -785 14595 -770
rect 14640 -785 14655 -770
rect 14700 -785 14715 -770
rect 14760 -785 14775 -770
rect 14820 -785 14835 -770
rect 14880 -785 14895 -770
rect 14940 -785 14955 -770
rect 15000 -785 15015 -770
rect 15060 -785 15075 -770
rect 15120 -785 15135 -770
rect 15180 -785 15195 -770
rect 15240 -785 15255 -770
rect 15300 -785 15315 -770
rect 15360 -785 15375 -770
rect 15420 -785 15435 -770
rect 15480 -785 15495 -770
rect 15540 -785 15555 -770
rect 15600 -785 15615 -770
rect 15660 -785 15675 -770
rect 15720 -785 15735 -770
rect 15780 -785 15795 -770
rect 15840 -785 15855 -770
rect 15900 -785 15915 -770
rect 15960 -785 15975 -770
rect 16020 -785 16035 -770
rect 16080 -785 16095 -770
rect 16140 -785 16155 -770
rect 16200 -785 16215 -770
rect 16260 -785 16275 -770
rect 16320 -785 16335 -770
rect 16380 -785 16395 -770
rect 16440 -785 16455 -770
rect 16500 -785 16515 -770
rect 16560 -785 16575 -770
rect 16620 -785 16635 -770
rect 16680 -785 16695 -770
rect 16740 -785 16755 -770
rect 16800 -785 16815 -770
rect 16860 -785 16875 -770
rect 16920 -785 16935 -770
rect 16980 -785 16995 -770
rect 17040 -785 17055 -770
rect 17100 -785 17115 -770
rect 17160 -785 17175 -770
rect 17220 -785 17235 -770
rect 17280 -785 17295 -770
rect 17340 -785 17355 -770
rect 17400 -785 17415 -770
rect 17460 -785 17475 -770
rect 17520 -785 17535 -770
rect 17580 -785 17595 -770
rect 17640 -785 17655 -770
rect 17700 -785 17715 -770
rect 17760 -785 17775 -770
rect 17820 -785 17835 -770
rect 17880 -785 17895 -770
rect 17940 -785 17955 -770
rect 18000 -785 18015 -770
rect 18060 -785 18075 -770
rect 18120 -785 18135 -770
rect 18180 -785 18195 -770
rect 18240 -785 18255 -770
rect 18300 -785 18315 -770
rect 18360 -785 18375 -770
rect 18420 -785 18435 -770
rect 18480 -785 18495 -770
rect 18540 -785 18555 -770
rect 18600 -785 18615 -770
rect 18660 -785 18675 -770
rect 18720 -785 18735 -770
rect 18780 -785 18795 -770
rect 18840 -785 18855 -770
rect 18900 -785 18915 -770
rect 18960 -785 18975 -770
rect 19020 -785 19035 -770
rect 19080 -785 19095 -770
rect 19140 -785 19155 -770
rect 19200 -785 19215 -770
rect 19260 -785 19275 -770
rect 19320 -785 19335 -770
rect 19380 -785 19395 -770
rect 19440 -785 19455 -770
rect 19500 -785 19515 -770
rect 19560 -785 19575 -770
rect 19620 -785 19635 -770
rect 19680 -785 19695 -770
rect 19740 -785 19755 -770
rect 19800 -785 19815 -770
rect 19860 -785 19875 -770
rect 19920 -785 19935 -770
rect 19980 -785 19995 -770
rect 20040 -785 20055 -770
rect 20100 -785 20115 -770
rect 20160 -785 20175 -770
rect 20220 -785 20235 -770
rect 20280 -785 20295 -770
rect 20340 -785 20355 -770
rect 20400 -785 20415 -770
rect 20460 -785 20475 -770
rect 20520 -785 20535 -770
rect 20580 -785 20595 -770
rect 20640 -785 20655 -770
rect 20700 -785 20715 -770
rect 20760 -785 20775 -770
rect 20820 -785 20835 -770
rect 20880 -785 20895 -770
rect 20940 -785 20955 -770
rect 21000 -785 21015 -770
rect 21060 -785 21075 -770
rect 21120 -785 21135 -770
rect 21180 -785 21195 -770
rect 21240 -785 21255 -770
rect 21300 -785 21315 -770
rect 21360 -785 21375 -770
rect 21420 -785 21435 -770
rect 21480 -785 21495 -770
rect 21540 -785 21555 -770
rect 21600 -785 21615 -770
rect 21660 -785 21675 -770
rect 21720 -785 21735 -770
rect 21780 -785 21795 -770
rect 21840 -785 21855 -770
rect 21900 -785 21915 -770
rect 21960 -785 21975 -770
rect 22020 -785 22035 -770
rect 22080 -785 22095 -770
rect 22140 -785 22155 -770
rect 22200 -785 22215 -770
rect 22260 -785 22275 -770
rect 22320 -785 22335 -770
rect 22380 -785 22395 -770
rect 22440 -785 22455 -770
rect 22500 -785 22515 -770
rect 22560 -785 22575 -770
rect 22620 -785 22635 -770
rect 22680 -785 22695 -770
rect 22740 -785 22755 -770
rect 22800 -785 22815 -770
rect 22860 -785 22875 -770
rect 22920 -785 22935 -770
rect 22980 -785 22995 -770
rect 23040 -785 23055 -770
rect 23100 -785 23115 -770
rect 23160 -785 23175 -770
rect 23220 -785 23235 -770
rect 23280 -785 23295 -770
rect 23340 -785 23355 -770
rect 23400 -785 23415 -770
rect 23460 -785 23475 -770
rect 23520 -785 23535 -770
rect 23580 -785 23595 -770
rect 23640 -785 23655 -770
rect 23700 -785 23715 -770
rect 23760 -785 23775 -770
rect 23820 -785 23835 -770
rect 23880 -785 23895 -770
rect 23940 -785 23955 -770
rect 24000 -785 24015 -770
rect 24060 -785 24075 -770
rect 24120 -785 24135 -770
rect 24180 -785 24195 -770
rect 24240 -785 24255 -770
rect 24300 -785 24315 -770
rect 24360 -785 24375 -770
rect 24420 -785 24435 -770
rect 24480 -785 24495 -770
rect 24540 -785 24555 -770
rect 24600 -785 24615 -770
rect 24660 -785 24675 -770
rect 24720 -785 24735 -770
rect 24780 -785 24795 -770
rect 24840 -785 24855 -770
rect 24900 -785 24915 -770
rect 24960 -785 24975 -770
rect 25020 -785 25035 -770
rect 25080 -785 25095 -770
rect 25140 -785 25155 -770
rect 25200 -785 25215 -770
rect 25260 -785 25275 -770
rect 25320 -785 25335 -770
rect 25380 -785 25395 -770
rect 25440 -785 25455 -770
rect 25500 -785 25515 -770
rect 25560 -785 25575 -770
rect 25620 -785 25635 -770
rect 25680 -785 25695 -770
rect 25740 -785 25755 -770
rect 25800 -785 25815 -770
rect 25860 -785 25875 -770
rect 25920 -785 25935 -770
rect 25980 -785 25995 -770
rect 26040 -785 26055 -770
rect 26100 -785 26115 -770
rect 26160 -785 26175 -770
rect 26220 -785 26235 -770
rect 26280 -785 26295 -770
rect 26340 -785 26355 -770
rect 26400 -785 26415 -770
rect 26460 -785 26475 -770
rect 26520 -785 26535 -770
rect 26580 -785 26595 -770
rect 26640 -785 26655 -770
rect 26700 -785 26715 -770
rect 26760 -785 26775 -770
rect 26820 -785 26835 -770
rect 26880 -785 26895 -770
rect 26940 -785 26955 -770
rect 27000 -785 27015 -770
rect 27060 -785 27075 -770
rect 27120 -785 27135 -770
rect 27180 -785 27195 -770
rect 27240 -785 27255 -770
rect 27300 -785 27315 -770
rect 27360 -785 27375 -770
rect 27420 -785 27435 -770
rect 27480 -785 27495 -770
rect 27540 -785 27555 -770
rect 27600 -785 27615 -770
rect 27660 -785 27675 -770
rect 27720 -785 27735 -770
rect 27780 -785 27795 -770
rect 27840 -785 27855 -770
rect 27900 -785 27915 -770
rect 27960 -785 27975 -770
rect 28020 -785 28035 -770
rect 28080 -785 28095 -770
rect 28140 -785 28155 -770
rect 28200 -785 28215 -770
rect 28260 -785 28275 -770
rect 28320 -785 28335 -770
rect 28380 -785 28395 -770
rect 28440 -785 28455 -770
rect 28500 -785 28515 -770
rect 28560 -785 28575 -770
rect 28620 -785 28635 -770
rect 28680 -785 28695 -770
rect 28740 -785 28755 -770
rect 28800 -785 28815 -770
rect 28860 -785 28875 -770
rect 28920 -785 28935 -770
rect 28980 -785 28995 -770
rect 29040 -785 29055 -770
rect 29100 -785 29115 -770
rect 29160 -785 29175 -770
rect 29220 -785 29235 -770
rect 29280 -785 29295 -770
rect 29340 -785 29355 -770
rect 29400 -785 29415 -770
rect 29460 -785 29475 -770
rect 29520 -785 29535 -770
rect 29580 -785 29595 -770
rect 29640 -785 29655 -770
rect 29700 -785 29715 -770
rect 29760 -785 29775 -770
rect 29820 -785 29835 -770
rect 29880 -785 29895 -770
rect 29940 -785 29955 -770
rect 30000 -785 30015 -770
rect 30060 -785 30075 -770
rect 30120 -785 30135 -770
rect 30180 -785 30195 -770
rect 30240 -785 30255 -770
rect 30300 -785 30315 -770
rect 30360 -785 30375 -770
rect 30420 -785 30435 -770
rect 30480 -785 30495 -770
rect 30540 -785 30555 -770
rect 30600 -785 30615 -770
rect 30660 -785 30675 -770
rect 0 -800 30675 -785
<< polycont >>
rect 201 -5 221 15
rect 326 -5 346 15
rect 631 -5 651 15
rect 1666 -5 1686 15
rect 5611 -5 5631 15
rect 30685 -505 30705 -485
<< locali >>
rect -460 475 21670 495
rect -460 375 -235 475
rect -135 375 315 475
rect 415 375 865 475
rect 965 375 1415 475
rect 1515 375 1965 475
rect 2065 375 2515 475
rect 2615 375 3065 475
rect 3165 375 3615 475
rect 3715 375 4165 475
rect 4265 375 4715 475
rect 4815 375 5265 475
rect 5365 375 5815 475
rect 5915 375 6365 475
rect 6465 375 6915 475
rect 7015 375 7465 475
rect 7565 375 8015 475
rect 8115 375 8565 475
rect 8665 375 9115 475
rect 9215 375 9665 475
rect 9765 375 10215 475
rect 10315 375 10765 475
rect 10865 375 11315 475
rect 11415 375 11865 475
rect 11965 375 12415 475
rect 12515 375 12965 475
rect 13065 375 13515 475
rect 13615 375 14065 475
rect 14165 375 14615 475
rect 14715 375 15165 475
rect 15265 375 15715 475
rect 15815 375 16265 475
rect 16365 375 16815 475
rect 16915 375 17365 475
rect 17465 375 17915 475
rect 18015 375 18465 475
rect 18565 375 19015 475
rect 19115 375 19565 475
rect 19665 375 20115 475
rect 20215 375 20665 475
rect 20765 375 21215 475
rect 21315 375 21670 475
rect -460 355 21670 375
rect -460 -5 -320 355
rect 2255 305 2310 315
rect 185 275 240 285
rect 185 240 195 275
rect 230 240 240 275
rect 185 230 240 240
rect 436 265 471 275
rect 436 240 441 265
rect 466 240 471 265
rect 195 205 220 230
rect 436 225 471 240
rect 741 265 776 275
rect 741 240 746 265
rect 771 240 776 265
rect 741 225 776 240
rect 986 265 1021 275
rect 986 240 991 265
rect 1016 240 1021 265
rect 986 225 1021 240
rect 1226 265 1261 275
rect 1226 240 1231 265
rect 1256 240 1261 265
rect 1226 225 1261 240
rect 1471 265 1506 275
rect 1471 240 1476 265
rect 1501 240 1506 265
rect 1471 225 1506 240
rect 1776 265 1811 275
rect 1776 240 1781 265
rect 1806 240 1811 265
rect 1776 225 1811 240
rect 2021 265 2056 275
rect 2021 240 2026 265
rect 2051 240 2056 265
rect 2255 270 2265 305
rect 2300 270 2310 305
rect 4195 305 4250 315
rect 2255 260 2310 270
rect 2506 265 2541 275
rect 2021 225 2056 240
rect 2265 225 2290 260
rect 2506 240 2511 265
rect 2536 240 2541 265
rect 2506 225 2541 240
rect 2746 265 2781 275
rect 2746 240 2751 265
rect 2776 240 2781 265
rect 2746 225 2781 240
rect 2991 265 3026 275
rect 2991 240 2996 265
rect 3021 240 3026 265
rect 2991 225 3026 240
rect 3231 265 3266 275
rect 3231 240 3236 265
rect 3261 240 3266 265
rect 3231 225 3266 240
rect 3476 265 3511 275
rect 3476 240 3481 265
rect 3506 240 3511 265
rect 3476 225 3511 240
rect 3716 265 3751 275
rect 3716 240 3721 265
rect 3746 240 3751 265
rect 3716 225 3751 240
rect 3961 265 3996 275
rect 3961 240 3966 265
rect 3991 240 3996 265
rect 4195 270 4205 305
rect 4240 270 4250 305
rect 6445 305 6500 315
rect 4195 260 4250 270
rect 4446 265 4481 275
rect 3961 225 3996 240
rect 195 185 221 205
rect 386 185 406 200
rect 441 185 466 225
rect 506 185 526 200
rect 691 185 711 200
rect 746 185 771 225
rect 811 185 831 200
rect 936 185 956 200
rect 991 185 1016 225
rect 1056 185 1076 200
rect 1176 185 1196 200
rect 1231 185 1256 225
rect 1296 185 1316 200
rect 1421 185 1441 200
rect 1476 185 1501 225
rect 1541 185 1561 200
rect 1726 185 1746 200
rect 1781 185 1806 225
rect 1846 185 1866 200
rect 1971 185 1991 200
rect 2026 185 2051 225
rect 2091 185 2111 200
rect 2211 185 2231 200
rect 2266 185 2291 225
rect 2331 185 2351 200
rect 2456 185 2476 200
rect 2511 185 2536 225
rect 2576 185 2596 200
rect 2696 185 2716 200
rect 2751 185 2776 225
rect 2816 185 2836 200
rect 2941 185 2961 200
rect 2996 185 3021 225
rect 3061 185 3081 200
rect 3181 185 3201 200
rect 3236 185 3261 225
rect 3301 185 3321 200
rect 3426 185 3446 200
rect 3481 185 3506 225
rect 3546 185 3566 200
rect 3666 185 3686 200
rect 3721 185 3746 225
rect 3786 185 3806 200
rect 3911 185 3931 200
rect 3966 185 3991 225
rect 4205 220 4230 260
rect 4446 240 4451 265
rect 4476 240 4481 265
rect 4446 225 4481 240
rect 4686 265 4721 275
rect 4686 240 4691 265
rect 4716 240 4721 265
rect 4686 225 4721 240
rect 4931 265 4966 275
rect 4931 240 4936 265
rect 4961 240 4966 265
rect 4931 225 4966 240
rect 5171 265 5206 275
rect 5171 240 5176 265
rect 5201 240 5206 265
rect 5171 225 5206 240
rect 5416 265 5451 275
rect 5416 240 5421 265
rect 5446 240 5451 265
rect 5416 225 5451 240
rect 5721 265 5756 275
rect 5721 240 5726 265
rect 5751 240 5756 265
rect 5721 225 5756 240
rect 5966 265 6001 275
rect 5966 240 5971 265
rect 5996 240 6001 265
rect 5966 225 6001 240
rect 6206 265 6241 275
rect 6206 240 6211 265
rect 6236 240 6241 265
rect 6445 270 6455 305
rect 6490 270 6500 305
rect 9350 305 9405 315
rect 6445 260 6500 270
rect 6691 265 6726 275
rect 6206 225 6241 240
rect 6455 225 6480 260
rect 6691 240 6696 265
rect 6721 240 6726 265
rect 6691 225 6726 240
rect 6936 265 6971 275
rect 6936 240 6941 265
rect 6966 240 6971 265
rect 6936 225 6971 240
rect 7176 265 7211 275
rect 7176 240 7181 265
rect 7206 240 7211 265
rect 7176 225 7211 240
rect 7416 265 7451 275
rect 7416 240 7421 265
rect 7446 240 7451 265
rect 7416 225 7451 240
rect 7656 265 7691 275
rect 7656 240 7661 265
rect 7686 240 7691 265
rect 7656 225 7691 240
rect 7901 265 7936 275
rect 7901 240 7906 265
rect 7931 240 7936 265
rect 7901 225 7936 240
rect 8141 265 8176 275
rect 8141 240 8146 265
rect 8171 240 8176 265
rect 8141 225 8176 240
rect 8386 265 8421 275
rect 8386 240 8391 265
rect 8416 240 8421 265
rect 8386 225 8421 240
rect 8626 265 8661 275
rect 8626 240 8631 265
rect 8656 240 8661 265
rect 8626 225 8661 240
rect 8871 265 8906 275
rect 8871 240 8876 265
rect 8901 240 8906 265
rect 8871 225 8906 240
rect 9111 265 9146 275
rect 9111 240 9116 265
rect 9141 240 9146 265
rect 9350 270 9360 305
rect 9395 270 9405 305
rect 11295 305 11350 315
rect 9350 260 9405 270
rect 9601 265 9636 275
rect 9111 225 9146 240
rect 4031 185 4051 200
rect 4151 185 4171 200
rect 4206 185 4231 220
rect 4271 185 4291 200
rect 4396 185 4416 200
rect 4451 185 4476 225
rect 4516 185 4536 200
rect 4636 185 4656 200
rect 4691 185 4716 225
rect 4756 185 4776 200
rect 4881 185 4901 200
rect 4936 185 4961 225
rect 5001 185 5021 200
rect 5121 185 5141 200
rect 5176 185 5201 225
rect 5241 185 5261 200
rect 5366 185 5386 200
rect 5421 185 5446 225
rect 5486 185 5506 200
rect 5671 185 5691 200
rect 5726 185 5751 225
rect 5791 185 5811 200
rect 5916 185 5936 200
rect 5971 185 5996 225
rect 6036 185 6056 200
rect 6156 185 6176 200
rect 6211 185 6236 225
rect 6276 185 6296 200
rect 6401 185 6421 200
rect 6456 185 6481 225
rect 6521 185 6541 200
rect 6641 185 6661 200
rect 6696 185 6721 225
rect 6761 185 6781 200
rect 6886 185 6906 200
rect 6941 185 6966 225
rect 7006 185 7026 200
rect 7126 185 7146 200
rect 7181 185 7206 225
rect 7246 185 7266 200
rect 7366 185 7386 200
rect 7421 185 7446 225
rect 7486 185 7506 200
rect 7606 185 7626 200
rect 7661 185 7686 225
rect 7726 185 7746 200
rect 7851 185 7871 200
rect 7906 185 7931 225
rect 7971 185 7991 200
rect 8091 185 8111 200
rect 8146 185 8171 225
rect 8211 185 8231 200
rect 8336 185 8356 200
rect 8391 185 8416 225
rect 8456 185 8476 200
rect 8576 185 8596 200
rect 8631 185 8656 225
rect 8696 185 8716 200
rect 8821 185 8841 200
rect 8876 185 8901 225
rect 8941 185 8961 200
rect 9061 185 9081 200
rect 9116 185 9141 225
rect 9360 220 9385 260
rect 9601 240 9606 265
rect 9631 240 9636 265
rect 9601 225 9636 240
rect 9846 265 9881 275
rect 9846 240 9851 265
rect 9876 240 9881 265
rect 9846 225 9881 240
rect 10086 265 10121 275
rect 10086 240 10091 265
rect 10116 240 10121 265
rect 10086 225 10121 240
rect 10331 265 10366 275
rect 10331 240 10336 265
rect 10361 240 10366 265
rect 10331 225 10366 240
rect 10571 265 10606 275
rect 10571 240 10576 265
rect 10601 240 10606 265
rect 10571 225 10606 240
rect 10816 265 10851 275
rect 10816 240 10821 265
rect 10846 240 10851 265
rect 10816 225 10851 240
rect 11056 265 11091 275
rect 11056 240 11061 265
rect 11086 240 11091 265
rect 11295 270 11305 305
rect 11340 270 11350 305
rect 12990 305 13045 315
rect 11295 260 11350 270
rect 11541 265 11576 275
rect 11056 225 11091 240
rect 11305 225 11330 260
rect 11541 240 11546 265
rect 11571 240 11576 265
rect 11541 225 11576 240
rect 11786 265 11821 275
rect 11786 240 11791 265
rect 11816 240 11821 265
rect 11786 225 11821 240
rect 12026 265 12061 275
rect 12026 240 12031 265
rect 12056 240 12061 265
rect 12026 225 12061 240
rect 12271 265 12306 275
rect 12271 240 12276 265
rect 12301 240 12306 265
rect 12271 225 12306 240
rect 12511 265 12546 275
rect 12511 240 12516 265
rect 12541 240 12546 265
rect 12511 225 12546 240
rect 12756 265 12791 275
rect 12756 240 12761 265
rect 12786 240 12791 265
rect 12990 270 13000 305
rect 13035 270 13045 305
rect 15175 305 15230 315
rect 12990 260 13045 270
rect 13241 265 13276 275
rect 12756 225 12791 240
rect 13000 225 13025 260
rect 13241 240 13246 265
rect 13271 240 13276 265
rect 13241 225 13276 240
rect 13481 265 13516 275
rect 13481 240 13486 265
rect 13511 240 13516 265
rect 13481 225 13516 240
rect 13726 265 13761 275
rect 13726 240 13731 265
rect 13756 240 13761 265
rect 13726 225 13761 240
rect 13966 265 14001 275
rect 13966 240 13971 265
rect 13996 240 14001 265
rect 13966 225 14001 240
rect 14211 265 14246 275
rect 14211 240 14216 265
rect 14241 240 14246 265
rect 14211 225 14246 240
rect 14451 265 14486 275
rect 14451 240 14456 265
rect 14481 240 14486 265
rect 14451 225 14486 240
rect 14696 265 14731 275
rect 14696 240 14701 265
rect 14726 240 14731 265
rect 14696 225 14731 240
rect 14936 265 14971 275
rect 14936 240 14941 265
rect 14966 240 14971 265
rect 15175 270 15185 305
rect 15220 270 15230 305
rect 17355 305 17410 315
rect 15175 260 15230 270
rect 15421 265 15456 275
rect 14936 225 14971 240
rect 15185 225 15210 260
rect 15421 240 15426 265
rect 15451 240 15456 265
rect 15421 225 15456 240
rect 15666 265 15701 275
rect 15666 240 15671 265
rect 15696 240 15701 265
rect 15666 225 15701 240
rect 15906 265 15941 275
rect 15906 240 15911 265
rect 15936 240 15941 265
rect 15906 225 15941 240
rect 16151 265 16186 275
rect 16151 240 16156 265
rect 16181 240 16186 265
rect 16151 225 16186 240
rect 16391 265 16426 275
rect 16391 240 16396 265
rect 16421 240 16426 265
rect 16391 225 16426 240
rect 16636 265 16671 275
rect 16636 240 16641 265
rect 16666 240 16671 265
rect 16636 225 16671 240
rect 16876 265 16911 275
rect 16876 240 16881 265
rect 16906 240 16911 265
rect 16876 225 16911 240
rect 17121 265 17156 275
rect 17121 240 17126 265
rect 17151 240 17156 265
rect 17355 270 17365 305
rect 17400 270 17410 305
rect 19540 305 19595 315
rect 17355 260 17410 270
rect 17606 265 17641 275
rect 17121 225 17156 240
rect 17365 225 17390 260
rect 17606 240 17611 265
rect 17636 240 17641 265
rect 17606 225 17641 240
rect 17846 265 17881 275
rect 17846 240 17851 265
rect 17876 240 17881 265
rect 17846 225 17881 240
rect 18091 265 18126 275
rect 18091 240 18096 265
rect 18121 240 18126 265
rect 18091 225 18126 240
rect 18331 265 18366 275
rect 18331 240 18336 265
rect 18361 240 18366 265
rect 18331 225 18366 240
rect 18576 265 18611 275
rect 18576 240 18581 265
rect 18606 240 18611 265
rect 18576 225 18611 240
rect 18816 265 18851 275
rect 18816 240 18821 265
rect 18846 240 18851 265
rect 18816 225 18851 240
rect 19061 265 19096 275
rect 19061 240 19066 265
rect 19091 240 19096 265
rect 19061 225 19096 240
rect 19301 265 19336 275
rect 19301 240 19306 265
rect 19331 240 19336 265
rect 19540 270 19550 305
rect 19585 270 19595 305
rect 20750 305 20805 315
rect 19540 260 19595 270
rect 19786 265 19821 275
rect 19301 225 19336 240
rect 19550 225 19575 260
rect 19786 240 19791 265
rect 19816 240 19821 265
rect 19786 225 19821 240
rect 20031 265 20066 275
rect 20031 240 20036 265
rect 20061 240 20066 265
rect 20031 225 20066 240
rect 20271 265 20306 275
rect 20271 240 20276 265
rect 20301 240 20306 265
rect 20271 225 20306 240
rect 20516 265 20551 275
rect 20516 240 20521 265
rect 20546 240 20551 265
rect 20750 270 20760 305
rect 20795 270 20805 305
rect 20750 260 20805 270
rect 21001 265 21036 275
rect 20516 225 20551 240
rect 20760 225 20785 260
rect 21001 240 21006 265
rect 21031 240 21036 265
rect 21001 225 21036 240
rect 21520 265 21670 355
rect 9181 185 9201 200
rect 9306 185 9326 200
rect 9361 185 9386 220
rect 9426 185 9446 200
rect 9551 185 9571 200
rect 9606 185 9631 225
rect 9671 185 9691 200
rect 9796 185 9816 200
rect 9851 185 9876 225
rect 9916 185 9936 200
rect 10036 185 10056 200
rect 10091 185 10116 225
rect 10156 185 10176 200
rect 10281 185 10301 200
rect 10336 185 10361 225
rect 10401 185 10421 200
rect 10521 185 10541 200
rect 10576 185 10601 225
rect 10641 185 10661 200
rect 10766 185 10786 200
rect 10821 185 10846 225
rect 10886 185 10906 200
rect 11006 185 11026 200
rect 11061 185 11086 225
rect 11126 185 11146 200
rect 11251 185 11271 200
rect 11306 185 11331 225
rect 11371 185 11391 200
rect 11491 185 11511 200
rect 11546 185 11571 225
rect 11611 185 11631 200
rect 11736 185 11756 200
rect 11791 185 11816 225
rect 11856 185 11876 200
rect 11976 185 11996 200
rect 12031 185 12056 225
rect 12096 185 12116 200
rect 12221 185 12241 200
rect 12276 185 12301 225
rect 12341 185 12361 200
rect 12461 185 12481 200
rect 12516 185 12541 225
rect 12581 185 12601 200
rect 12706 185 12726 200
rect 12761 185 12786 225
rect 12826 185 12846 200
rect 12946 185 12966 200
rect 13001 185 13026 225
rect 13066 185 13086 200
rect 13191 185 13211 200
rect 13246 185 13271 225
rect 13311 185 13331 200
rect 13431 185 13451 200
rect 13486 185 13511 225
rect 13551 185 13571 200
rect 13676 185 13696 200
rect 13731 185 13756 225
rect 13796 185 13816 200
rect 13916 185 13936 200
rect 13971 185 13996 225
rect 14036 185 14056 200
rect 14161 185 14181 200
rect 14216 185 14241 225
rect 14281 185 14301 200
rect 14401 185 14421 200
rect 14456 185 14481 225
rect 14521 185 14541 200
rect 14646 185 14666 200
rect 14701 185 14726 225
rect 14766 185 14786 200
rect 14886 185 14906 200
rect 14941 185 14966 225
rect 15185 220 15211 225
rect 15006 185 15026 200
rect 15131 185 15151 200
rect 15186 185 15211 220
rect 15251 185 15271 200
rect 15371 185 15391 200
rect 15426 185 15451 225
rect 15491 185 15511 200
rect 15616 185 15636 200
rect 15671 185 15696 225
rect 15736 185 15756 200
rect 15856 185 15876 200
rect 15911 185 15936 225
rect 15976 185 15996 200
rect 16101 185 16121 200
rect 16156 185 16181 225
rect 16221 185 16241 200
rect 16341 185 16361 200
rect 16396 185 16421 225
rect 16461 185 16481 200
rect 16586 185 16606 200
rect 16641 185 16666 225
rect 16706 185 16726 200
rect 16826 185 16846 200
rect 16881 185 16906 225
rect 16946 185 16966 200
rect 17071 185 17091 200
rect 17126 185 17151 225
rect 17191 185 17211 200
rect 17311 185 17331 200
rect 17366 185 17391 225
rect 17431 185 17451 200
rect 17556 185 17576 200
rect 17611 185 17636 225
rect 17676 185 17696 200
rect 17796 185 17816 200
rect 17851 185 17876 225
rect 17916 185 17936 200
rect 18041 185 18061 200
rect 18096 185 18121 225
rect 18161 185 18181 200
rect 18281 185 18301 200
rect 18336 185 18361 225
rect 18401 185 18421 200
rect 18526 185 18546 200
rect 18581 185 18606 225
rect 18646 185 18666 200
rect 18766 185 18786 200
rect 18821 185 18846 225
rect 18886 185 18906 200
rect 19011 185 19031 200
rect 19066 185 19091 225
rect 19131 185 19151 200
rect 19251 185 19271 200
rect 19306 185 19331 225
rect 19371 185 19391 200
rect 19496 185 19516 200
rect 19551 185 19576 225
rect 19616 185 19636 200
rect 19736 185 19756 200
rect 19791 185 19816 225
rect 19856 185 19876 200
rect 19981 185 20001 200
rect 20036 185 20061 225
rect 20101 185 20121 200
rect 20221 185 20241 200
rect 20276 185 20301 225
rect 20341 185 20361 200
rect 20466 185 20486 200
rect 20521 185 20546 225
rect 20586 185 20606 200
rect 20706 185 20726 200
rect 20761 185 20786 225
rect 20826 185 20846 200
rect 20951 185 20971 200
rect 21006 185 21031 225
rect 21071 185 21091 200
rect 191 165 226 185
rect 191 140 196 165
rect 221 140 226 165
rect 191 120 226 140
rect 191 95 196 120
rect 221 95 226 120
rect 191 85 226 95
rect 251 165 286 185
rect 251 140 256 165
rect 281 140 286 165
rect 251 120 286 140
rect 251 95 256 120
rect 281 95 286 120
rect 251 85 286 95
rect 316 165 351 185
rect 316 140 321 165
rect 346 140 351 165
rect 316 120 351 140
rect 316 95 321 120
rect 346 95 351 120
rect 316 85 351 95
rect 376 165 411 185
rect 376 140 381 165
rect 406 140 411 165
rect 376 120 411 140
rect 376 95 381 120
rect 406 95 411 120
rect 376 85 411 95
rect 436 165 471 185
rect 436 140 441 165
rect 466 140 471 165
rect 436 120 471 140
rect 436 95 441 120
rect 466 95 471 120
rect 436 85 471 95
rect 496 165 531 185
rect 496 140 501 165
rect 526 140 531 165
rect 496 120 531 140
rect 496 95 501 120
rect 526 95 531 120
rect 496 85 531 95
rect 556 165 591 185
rect 556 140 561 165
rect 586 140 591 165
rect 556 120 591 140
rect 556 95 561 120
rect 586 95 591 120
rect 556 85 591 95
rect 621 165 656 185
rect 621 140 626 165
rect 651 140 656 165
rect 621 120 656 140
rect 621 95 626 120
rect 651 95 656 120
rect 621 85 656 95
rect 681 165 716 185
rect 681 140 686 165
rect 711 140 716 165
rect 681 120 716 140
rect 681 95 686 120
rect 711 95 716 120
rect 681 85 716 95
rect 741 165 776 185
rect 741 140 746 165
rect 771 140 776 165
rect 741 120 776 140
rect 741 95 746 120
rect 771 95 776 120
rect 741 85 776 95
rect 801 165 836 185
rect 801 140 806 165
rect 831 140 836 165
rect 801 120 836 140
rect 801 95 806 120
rect 831 95 836 120
rect 801 85 836 95
rect 861 165 901 185
rect 861 140 871 165
rect 896 140 901 165
rect 861 120 901 140
rect 861 95 871 120
rect 896 95 901 120
rect 861 85 901 95
rect 926 165 961 185
rect 926 140 931 165
rect 956 140 961 165
rect 926 120 961 140
rect 926 95 931 120
rect 956 95 961 120
rect 926 85 961 95
rect 986 165 1021 185
rect 986 140 991 165
rect 1016 140 1021 165
rect 986 120 1021 140
rect 986 95 991 120
rect 1016 95 1021 120
rect 986 85 1021 95
rect 1046 165 1081 185
rect 1046 140 1051 165
rect 1076 140 1081 165
rect 1046 120 1081 140
rect 1046 95 1051 120
rect 1076 95 1081 120
rect 1046 85 1081 95
rect 1106 165 1141 185
rect 1106 140 1111 165
rect 1136 140 1141 165
rect 1106 120 1141 140
rect 1106 95 1111 120
rect 1136 95 1141 120
rect 1106 85 1141 95
rect 1166 165 1201 185
rect 1166 140 1171 165
rect 1196 140 1201 165
rect 1166 120 1201 140
rect 1166 95 1171 120
rect 1196 95 1201 120
rect 1166 85 1201 95
rect 1226 165 1261 185
rect 1226 140 1231 165
rect 1256 140 1261 165
rect 1226 120 1261 140
rect 1226 95 1231 120
rect 1256 95 1261 120
rect 1226 85 1261 95
rect 1286 165 1321 185
rect 1286 140 1291 165
rect 1316 140 1321 165
rect 1286 120 1321 140
rect 1286 95 1291 120
rect 1316 95 1321 120
rect 1286 85 1321 95
rect 1346 165 1386 185
rect 1346 140 1356 165
rect 1381 140 1386 165
rect 1346 120 1386 140
rect 1346 95 1356 120
rect 1381 95 1386 120
rect 1346 85 1386 95
rect 1411 165 1446 185
rect 1411 140 1416 165
rect 1441 140 1446 165
rect 1411 120 1446 140
rect 1411 95 1416 120
rect 1441 95 1446 120
rect 1411 85 1446 95
rect 1471 165 1506 185
rect 1471 140 1476 165
rect 1501 140 1506 165
rect 1471 120 1506 140
rect 1471 95 1476 120
rect 1501 95 1506 120
rect 1471 85 1506 95
rect 1531 165 1566 185
rect 1531 140 1536 165
rect 1561 140 1566 165
rect 1531 120 1566 140
rect 1531 95 1536 120
rect 1561 95 1566 120
rect 1531 85 1566 95
rect 1591 165 1626 185
rect 1591 140 1596 165
rect 1621 140 1626 165
rect 1591 120 1626 140
rect 1591 95 1596 120
rect 1621 95 1626 120
rect 1591 85 1626 95
rect 1656 165 1691 185
rect 1656 140 1661 165
rect 1686 140 1691 165
rect 1656 120 1691 140
rect 1656 95 1661 120
rect 1686 95 1691 120
rect 1656 85 1691 95
rect 1716 165 1751 185
rect 1716 140 1721 165
rect 1746 140 1751 165
rect 1716 120 1751 140
rect 1716 95 1721 120
rect 1746 95 1751 120
rect 1716 85 1751 95
rect 1776 165 1811 185
rect 1776 140 1781 165
rect 1806 140 1811 165
rect 1776 120 1811 140
rect 1776 95 1781 120
rect 1806 95 1811 120
rect 1776 85 1811 95
rect 1836 165 1871 185
rect 1836 140 1841 165
rect 1866 140 1871 165
rect 1836 120 1871 140
rect 1836 95 1841 120
rect 1866 95 1871 120
rect 1836 85 1871 95
rect 1896 165 1936 185
rect 1896 140 1906 165
rect 1931 140 1936 165
rect 1896 120 1936 140
rect 1896 95 1906 120
rect 1931 95 1936 120
rect 1896 85 1936 95
rect 1961 165 1996 185
rect 1961 140 1966 165
rect 1991 140 1996 165
rect 1961 120 1996 140
rect 1961 95 1966 120
rect 1991 95 1996 120
rect 1961 85 1996 95
rect 2021 165 2056 185
rect 2021 140 2026 165
rect 2051 140 2056 165
rect 2021 120 2056 140
rect 2021 95 2026 120
rect 2051 95 2056 120
rect 2021 85 2056 95
rect 2081 165 2116 185
rect 2081 140 2086 165
rect 2111 140 2116 165
rect 2081 120 2116 140
rect 2081 95 2086 120
rect 2111 95 2116 120
rect 2081 85 2116 95
rect 2141 165 2176 185
rect 2141 140 2146 165
rect 2171 140 2176 165
rect 2141 120 2176 140
rect 2141 95 2146 120
rect 2171 95 2176 120
rect 2141 85 2176 95
rect 2201 165 2236 185
rect 2201 140 2206 165
rect 2231 140 2236 165
rect 2201 120 2236 140
rect 2201 95 2206 120
rect 2231 95 2236 120
rect 2201 85 2236 95
rect 2261 165 2296 185
rect 2261 140 2266 165
rect 2291 140 2296 165
rect 2261 120 2296 140
rect 2261 95 2266 120
rect 2291 95 2296 120
rect 2261 85 2296 95
rect 2321 165 2356 185
rect 2321 140 2326 165
rect 2351 140 2356 165
rect 2321 120 2356 140
rect 2321 95 2326 120
rect 2351 95 2356 120
rect 2321 85 2356 95
rect 2381 165 2421 185
rect 2381 140 2391 165
rect 2416 140 2421 165
rect 2381 120 2421 140
rect 2381 95 2391 120
rect 2416 95 2421 120
rect 2381 85 2421 95
rect 2446 165 2481 185
rect 2446 140 2451 165
rect 2476 140 2481 165
rect 2446 120 2481 140
rect 2446 95 2451 120
rect 2476 95 2481 120
rect 2446 85 2481 95
rect 2506 165 2541 185
rect 2506 140 2511 165
rect 2536 140 2541 165
rect 2506 120 2541 140
rect 2506 95 2511 120
rect 2536 95 2541 120
rect 2506 85 2541 95
rect 2566 165 2601 185
rect 2566 140 2571 165
rect 2596 140 2601 165
rect 2566 120 2601 140
rect 2566 95 2571 120
rect 2596 95 2601 120
rect 2566 85 2601 95
rect 2626 165 2661 185
rect 2626 140 2631 165
rect 2656 140 2661 165
rect 2626 120 2661 140
rect 2626 95 2631 120
rect 2656 95 2661 120
rect 2626 85 2661 95
rect 2686 165 2721 185
rect 2686 140 2691 165
rect 2716 140 2721 165
rect 2686 120 2721 140
rect 2686 95 2691 120
rect 2716 95 2721 120
rect 2686 85 2721 95
rect 2746 165 2781 185
rect 2746 140 2751 165
rect 2776 140 2781 165
rect 2746 120 2781 140
rect 2746 95 2751 120
rect 2776 95 2781 120
rect 2746 85 2781 95
rect 2806 165 2841 185
rect 2806 140 2811 165
rect 2836 140 2841 165
rect 2806 120 2841 140
rect 2806 95 2811 120
rect 2836 95 2841 120
rect 2806 85 2841 95
rect 2866 165 2906 185
rect 2866 140 2876 165
rect 2901 140 2906 165
rect 2866 120 2906 140
rect 2866 95 2876 120
rect 2901 95 2906 120
rect 2866 85 2906 95
rect 2931 165 2966 185
rect 2931 140 2936 165
rect 2961 140 2966 165
rect 2931 120 2966 140
rect 2931 95 2936 120
rect 2961 95 2966 120
rect 2931 85 2966 95
rect 2991 165 3026 185
rect 2991 140 2996 165
rect 3021 140 3026 165
rect 2991 120 3026 140
rect 2991 95 2996 120
rect 3021 95 3026 120
rect 2991 85 3026 95
rect 3051 165 3086 185
rect 3051 140 3056 165
rect 3081 140 3086 165
rect 3051 120 3086 140
rect 3051 95 3056 120
rect 3081 95 3086 120
rect 3051 85 3086 95
rect 3111 165 3146 185
rect 3111 140 3116 165
rect 3141 140 3146 165
rect 3111 120 3146 140
rect 3111 95 3116 120
rect 3141 95 3146 120
rect 3111 85 3146 95
rect 3171 165 3206 185
rect 3171 140 3176 165
rect 3201 140 3206 165
rect 3171 120 3206 140
rect 3171 95 3176 120
rect 3201 95 3206 120
rect 3171 85 3206 95
rect 3231 165 3266 185
rect 3231 140 3236 165
rect 3261 140 3266 165
rect 3231 120 3266 140
rect 3231 95 3236 120
rect 3261 95 3266 120
rect 3231 85 3266 95
rect 3291 165 3326 185
rect 3291 140 3296 165
rect 3321 140 3326 165
rect 3291 120 3326 140
rect 3291 95 3296 120
rect 3321 95 3326 120
rect 3291 85 3326 95
rect 3351 165 3391 185
rect 3351 140 3361 165
rect 3386 140 3391 165
rect 3351 120 3391 140
rect 3351 95 3361 120
rect 3386 95 3391 120
rect 3351 85 3391 95
rect 3416 165 3451 185
rect 3416 140 3421 165
rect 3446 140 3451 165
rect 3416 120 3451 140
rect 3416 95 3421 120
rect 3446 95 3451 120
rect 3416 85 3451 95
rect 3476 165 3511 185
rect 3476 140 3481 165
rect 3506 140 3511 165
rect 3476 120 3511 140
rect 3476 95 3481 120
rect 3506 95 3511 120
rect 3476 85 3511 95
rect 3536 165 3571 185
rect 3536 140 3541 165
rect 3566 140 3571 165
rect 3536 120 3571 140
rect 3536 95 3541 120
rect 3566 95 3571 120
rect 3536 85 3571 95
rect 3596 165 3631 185
rect 3596 140 3601 165
rect 3626 140 3631 165
rect 3596 120 3631 140
rect 3596 95 3601 120
rect 3626 95 3631 120
rect 3596 85 3631 95
rect 3656 165 3691 185
rect 3656 140 3661 165
rect 3686 140 3691 165
rect 3656 120 3691 140
rect 3656 95 3661 120
rect 3686 95 3691 120
rect 3656 85 3691 95
rect 3716 165 3751 185
rect 3716 140 3721 165
rect 3746 140 3751 165
rect 3716 120 3751 140
rect 3716 95 3721 120
rect 3746 95 3751 120
rect 3716 85 3751 95
rect 3776 165 3811 185
rect 3776 140 3781 165
rect 3806 140 3811 165
rect 3776 120 3811 140
rect 3776 95 3781 120
rect 3806 95 3811 120
rect 3776 85 3811 95
rect 3836 165 3876 185
rect 3836 140 3846 165
rect 3871 140 3876 165
rect 3836 120 3876 140
rect 3836 95 3846 120
rect 3871 95 3876 120
rect 3836 85 3876 95
rect 3901 165 3936 185
rect 3901 140 3906 165
rect 3931 140 3936 165
rect 3901 120 3936 140
rect 3901 95 3906 120
rect 3931 95 3936 120
rect 3901 85 3936 95
rect 3961 165 3996 185
rect 3961 140 3966 165
rect 3991 140 3996 165
rect 3961 120 3996 140
rect 3961 95 3966 120
rect 3991 95 3996 120
rect 3961 85 3996 95
rect 4021 165 4056 185
rect 4021 140 4026 165
rect 4051 140 4056 165
rect 4021 120 4056 140
rect 4021 95 4026 120
rect 4051 95 4056 120
rect 4021 85 4056 95
rect 4081 165 4116 185
rect 4081 140 4086 165
rect 4111 140 4116 165
rect 4081 120 4116 140
rect 4081 95 4086 120
rect 4111 95 4116 120
rect 4081 85 4116 95
rect 4141 165 4176 185
rect 4141 140 4146 165
rect 4171 140 4176 165
rect 4141 120 4176 140
rect 4141 95 4146 120
rect 4171 95 4176 120
rect 4141 85 4176 95
rect 4201 165 4236 185
rect 4201 140 4206 165
rect 4231 140 4236 165
rect 4201 120 4236 140
rect 4201 95 4206 120
rect 4231 95 4236 120
rect 4201 85 4236 95
rect 4261 165 4296 185
rect 4261 140 4266 165
rect 4291 140 4296 165
rect 4261 120 4296 140
rect 4261 95 4266 120
rect 4291 95 4296 120
rect 4261 85 4296 95
rect 4321 165 4361 185
rect 4321 140 4331 165
rect 4356 140 4361 165
rect 4321 120 4361 140
rect 4321 95 4331 120
rect 4356 95 4361 120
rect 4321 85 4361 95
rect 4386 165 4421 185
rect 4386 140 4391 165
rect 4416 140 4421 165
rect 4386 120 4421 140
rect 4386 95 4391 120
rect 4416 95 4421 120
rect 4386 85 4421 95
rect 4446 165 4481 185
rect 4446 140 4451 165
rect 4476 140 4481 165
rect 4446 120 4481 140
rect 4446 95 4451 120
rect 4476 95 4481 120
rect 4446 85 4481 95
rect 4506 165 4541 185
rect 4506 140 4511 165
rect 4536 140 4541 165
rect 4506 120 4541 140
rect 4506 95 4511 120
rect 4536 95 4541 120
rect 4506 85 4541 95
rect 4566 165 4601 185
rect 4566 140 4571 165
rect 4596 140 4601 165
rect 4566 120 4601 140
rect 4566 95 4571 120
rect 4596 95 4601 120
rect 4566 85 4601 95
rect 4626 165 4661 185
rect 4626 140 4631 165
rect 4656 140 4661 165
rect 4626 120 4661 140
rect 4626 95 4631 120
rect 4656 95 4661 120
rect 4626 85 4661 95
rect 4686 165 4721 185
rect 4686 140 4691 165
rect 4716 140 4721 165
rect 4686 120 4721 140
rect 4686 95 4691 120
rect 4716 95 4721 120
rect 4686 85 4721 95
rect 4746 165 4781 185
rect 4746 140 4751 165
rect 4776 140 4781 165
rect 4746 120 4781 140
rect 4746 95 4751 120
rect 4776 95 4781 120
rect 4746 85 4781 95
rect 4806 165 4846 185
rect 4806 140 4816 165
rect 4841 140 4846 165
rect 4806 120 4846 140
rect 4806 95 4816 120
rect 4841 95 4846 120
rect 4806 85 4846 95
rect 4871 165 4906 185
rect 4871 140 4876 165
rect 4901 140 4906 165
rect 4871 120 4906 140
rect 4871 95 4876 120
rect 4901 95 4906 120
rect 4871 85 4906 95
rect 4931 165 4966 185
rect 4931 140 4936 165
rect 4961 140 4966 165
rect 4931 120 4966 140
rect 4931 95 4936 120
rect 4961 95 4966 120
rect 4931 85 4966 95
rect 4991 165 5026 185
rect 4991 140 4996 165
rect 5021 140 5026 165
rect 4991 120 5026 140
rect 4991 95 4996 120
rect 5021 95 5026 120
rect 4991 85 5026 95
rect 5051 165 5086 185
rect 5051 140 5056 165
rect 5081 140 5086 165
rect 5051 120 5086 140
rect 5051 95 5056 120
rect 5081 95 5086 120
rect 5051 85 5086 95
rect 5111 165 5146 185
rect 5111 140 5116 165
rect 5141 140 5146 165
rect 5111 120 5146 140
rect 5111 95 5116 120
rect 5141 95 5146 120
rect 5111 85 5146 95
rect 5171 165 5206 185
rect 5171 140 5176 165
rect 5201 140 5206 165
rect 5171 120 5206 140
rect 5171 95 5176 120
rect 5201 95 5206 120
rect 5171 85 5206 95
rect 5231 165 5266 185
rect 5231 140 5236 165
rect 5261 140 5266 165
rect 5231 120 5266 140
rect 5231 95 5236 120
rect 5261 95 5266 120
rect 5231 85 5266 95
rect 5291 165 5331 185
rect 5291 140 5301 165
rect 5326 140 5331 165
rect 5291 120 5331 140
rect 5291 95 5301 120
rect 5326 95 5331 120
rect 5291 85 5331 95
rect 5356 165 5391 185
rect 5356 140 5361 165
rect 5386 140 5391 165
rect 5356 120 5391 140
rect 5356 95 5361 120
rect 5386 95 5391 120
rect 5356 85 5391 95
rect 5416 165 5451 185
rect 5416 140 5421 165
rect 5446 140 5451 165
rect 5416 120 5451 140
rect 5416 95 5421 120
rect 5446 95 5451 120
rect 5416 85 5451 95
rect 5476 165 5511 185
rect 5476 140 5481 165
rect 5506 140 5511 165
rect 5476 120 5511 140
rect 5476 95 5481 120
rect 5506 95 5511 120
rect 5476 85 5511 95
rect 5536 165 5571 185
rect 5536 140 5541 165
rect 5566 140 5571 165
rect 5536 120 5571 140
rect 5536 95 5541 120
rect 5566 95 5571 120
rect 5536 85 5571 95
rect 5601 165 5636 185
rect 5601 140 5606 165
rect 5631 140 5636 165
rect 5601 120 5636 140
rect 5601 95 5606 120
rect 5631 95 5636 120
rect 5601 85 5636 95
rect 5661 165 5696 185
rect 5661 140 5666 165
rect 5691 140 5696 165
rect 5661 120 5696 140
rect 5661 95 5666 120
rect 5691 95 5696 120
rect 5661 85 5696 95
rect 5721 165 5756 185
rect 5721 140 5726 165
rect 5751 140 5756 165
rect 5721 120 5756 140
rect 5721 95 5726 120
rect 5751 95 5756 120
rect 5721 85 5756 95
rect 5781 165 5816 185
rect 5781 140 5786 165
rect 5811 140 5816 165
rect 5781 120 5816 140
rect 5781 95 5786 120
rect 5811 95 5816 120
rect 5781 85 5816 95
rect 5841 165 5881 185
rect 5841 140 5851 165
rect 5876 140 5881 165
rect 5841 120 5881 140
rect 5841 95 5851 120
rect 5876 95 5881 120
rect 5841 85 5881 95
rect 5906 165 5941 185
rect 5906 140 5911 165
rect 5936 140 5941 165
rect 5906 120 5941 140
rect 5906 95 5911 120
rect 5936 95 5941 120
rect 5906 85 5941 95
rect 5966 165 6001 185
rect 5966 140 5971 165
rect 5996 140 6001 165
rect 5966 120 6001 140
rect 5966 95 5971 120
rect 5996 95 6001 120
rect 5966 85 6001 95
rect 6026 165 6061 185
rect 6026 140 6031 165
rect 6056 140 6061 165
rect 6026 120 6061 140
rect 6026 95 6031 120
rect 6056 95 6061 120
rect 6026 85 6061 95
rect 6086 165 6121 185
rect 6086 140 6091 165
rect 6116 140 6121 165
rect 6086 120 6121 140
rect 6086 95 6091 120
rect 6116 95 6121 120
rect 6086 85 6121 95
rect 6146 165 6181 185
rect 6146 140 6151 165
rect 6176 140 6181 165
rect 6146 120 6181 140
rect 6146 95 6151 120
rect 6176 95 6181 120
rect 6146 85 6181 95
rect 6206 165 6241 185
rect 6206 140 6211 165
rect 6236 140 6241 165
rect 6206 120 6241 140
rect 6206 95 6211 120
rect 6236 95 6241 120
rect 6206 85 6241 95
rect 6266 165 6301 185
rect 6266 140 6271 165
rect 6296 140 6301 165
rect 6266 120 6301 140
rect 6266 95 6271 120
rect 6296 95 6301 120
rect 6266 85 6301 95
rect 6326 165 6366 185
rect 6326 140 6336 165
rect 6361 140 6366 165
rect 6326 120 6366 140
rect 6326 95 6336 120
rect 6361 95 6366 120
rect 6326 85 6366 95
rect 6391 165 6426 185
rect 6391 140 6396 165
rect 6421 140 6426 165
rect 6391 120 6426 140
rect 6391 95 6396 120
rect 6421 95 6426 120
rect 6391 85 6426 95
rect 6451 165 6486 185
rect 6451 140 6456 165
rect 6481 140 6486 165
rect 6451 120 6486 140
rect 6451 95 6456 120
rect 6481 95 6486 120
rect 6451 85 6486 95
rect 6511 165 6546 185
rect 6511 140 6516 165
rect 6541 140 6546 165
rect 6511 120 6546 140
rect 6511 95 6516 120
rect 6541 95 6546 120
rect 6511 85 6546 95
rect 6571 165 6606 185
rect 6571 140 6576 165
rect 6601 140 6606 165
rect 6571 120 6606 140
rect 6571 95 6576 120
rect 6601 95 6606 120
rect 6571 85 6606 95
rect 6631 165 6666 185
rect 6631 140 6636 165
rect 6661 140 6666 165
rect 6631 120 6666 140
rect 6631 95 6636 120
rect 6661 95 6666 120
rect 6631 85 6666 95
rect 6691 165 6726 185
rect 6691 140 6696 165
rect 6721 140 6726 165
rect 6691 120 6726 140
rect 6691 95 6696 120
rect 6721 95 6726 120
rect 6691 85 6726 95
rect 6751 165 6786 185
rect 6751 140 6756 165
rect 6781 140 6786 165
rect 6751 120 6786 140
rect 6751 95 6756 120
rect 6781 95 6786 120
rect 6751 85 6786 95
rect 6811 165 6851 185
rect 6811 140 6821 165
rect 6846 140 6851 165
rect 6811 120 6851 140
rect 6811 95 6821 120
rect 6846 95 6851 120
rect 6811 85 6851 95
rect 6876 165 6911 185
rect 6876 140 6881 165
rect 6906 140 6911 165
rect 6876 120 6911 140
rect 6876 95 6881 120
rect 6906 95 6911 120
rect 6876 85 6911 95
rect 6936 165 6971 185
rect 6936 140 6941 165
rect 6966 140 6971 165
rect 6936 120 6971 140
rect 6936 95 6941 120
rect 6966 95 6971 120
rect 6936 85 6971 95
rect 6996 165 7031 185
rect 6996 140 7001 165
rect 7026 140 7031 165
rect 6996 120 7031 140
rect 6996 95 7001 120
rect 7026 95 7031 120
rect 6996 85 7031 95
rect 7056 165 7091 185
rect 7056 140 7061 165
rect 7086 140 7091 165
rect 7056 120 7091 140
rect 7056 95 7061 120
rect 7086 95 7091 120
rect 7056 85 7091 95
rect 7116 165 7151 185
rect 7116 140 7121 165
rect 7146 140 7151 165
rect 7116 120 7151 140
rect 7116 95 7121 120
rect 7146 95 7151 120
rect 7116 85 7151 95
rect 7176 165 7211 185
rect 7176 140 7181 165
rect 7206 140 7211 165
rect 7176 120 7211 140
rect 7176 95 7181 120
rect 7206 95 7211 120
rect 7176 85 7211 95
rect 7236 165 7271 185
rect 7236 140 7241 165
rect 7266 140 7271 165
rect 7236 120 7271 140
rect 7236 95 7241 120
rect 7266 95 7271 120
rect 7236 85 7271 95
rect 7296 165 7331 185
rect 7296 140 7301 165
rect 7326 140 7331 165
rect 7296 120 7331 140
rect 7296 95 7301 120
rect 7326 95 7331 120
rect 7296 85 7331 95
rect 7356 165 7391 185
rect 7356 140 7361 165
rect 7386 140 7391 165
rect 7356 120 7391 140
rect 7356 95 7361 120
rect 7386 95 7391 120
rect 7356 85 7391 95
rect 7416 165 7451 185
rect 7416 140 7421 165
rect 7446 140 7451 165
rect 7416 120 7451 140
rect 7416 95 7421 120
rect 7446 95 7451 120
rect 7416 85 7451 95
rect 7476 165 7511 185
rect 7476 140 7481 165
rect 7506 140 7511 165
rect 7476 120 7511 140
rect 7476 95 7481 120
rect 7506 95 7511 120
rect 7476 85 7511 95
rect 7536 165 7571 185
rect 7536 140 7541 165
rect 7566 140 7571 165
rect 7536 120 7571 140
rect 7536 95 7541 120
rect 7566 95 7571 120
rect 7536 85 7571 95
rect 7596 165 7631 185
rect 7596 140 7601 165
rect 7626 140 7631 165
rect 7596 120 7631 140
rect 7596 95 7601 120
rect 7626 95 7631 120
rect 7596 85 7631 95
rect 7656 165 7691 185
rect 7656 140 7661 165
rect 7686 140 7691 165
rect 7656 120 7691 140
rect 7656 95 7661 120
rect 7686 95 7691 120
rect 7656 85 7691 95
rect 7716 165 7751 185
rect 7716 140 7721 165
rect 7746 140 7751 165
rect 7716 120 7751 140
rect 7716 95 7721 120
rect 7746 95 7751 120
rect 7716 85 7751 95
rect 7776 165 7816 185
rect 7776 140 7786 165
rect 7811 140 7816 165
rect 7776 120 7816 140
rect 7776 95 7786 120
rect 7811 95 7816 120
rect 7776 85 7816 95
rect 7841 165 7876 185
rect 7841 140 7846 165
rect 7871 140 7876 165
rect 7841 120 7876 140
rect 7841 95 7846 120
rect 7871 95 7876 120
rect 7841 85 7876 95
rect 7901 165 7936 185
rect 7901 140 7906 165
rect 7931 140 7936 165
rect 7901 120 7936 140
rect 7901 95 7906 120
rect 7931 95 7936 120
rect 7901 85 7936 95
rect 7961 165 7996 185
rect 7961 140 7966 165
rect 7991 140 7996 165
rect 7961 120 7996 140
rect 7961 95 7966 120
rect 7991 95 7996 120
rect 7961 85 7996 95
rect 8021 165 8056 185
rect 8021 140 8026 165
rect 8051 140 8056 165
rect 8021 120 8056 140
rect 8021 95 8026 120
rect 8051 95 8056 120
rect 8021 85 8056 95
rect 8081 165 8116 185
rect 8081 140 8086 165
rect 8111 140 8116 165
rect 8081 120 8116 140
rect 8081 95 8086 120
rect 8111 95 8116 120
rect 8081 85 8116 95
rect 8141 165 8176 185
rect 8141 140 8146 165
rect 8171 140 8176 165
rect 8141 120 8176 140
rect 8141 95 8146 120
rect 8171 95 8176 120
rect 8141 85 8176 95
rect 8201 165 8236 185
rect 8201 140 8206 165
rect 8231 140 8236 165
rect 8201 120 8236 140
rect 8201 95 8206 120
rect 8231 95 8236 120
rect 8201 85 8236 95
rect 8261 165 8301 185
rect 8261 140 8271 165
rect 8296 140 8301 165
rect 8261 120 8301 140
rect 8261 95 8271 120
rect 8296 95 8301 120
rect 8261 85 8301 95
rect 8326 165 8361 185
rect 8326 140 8331 165
rect 8356 140 8361 165
rect 8326 120 8361 140
rect 8326 95 8331 120
rect 8356 95 8361 120
rect 8326 85 8361 95
rect 8386 165 8421 185
rect 8386 140 8391 165
rect 8416 140 8421 165
rect 8386 120 8421 140
rect 8386 95 8391 120
rect 8416 95 8421 120
rect 8386 85 8421 95
rect 8446 165 8481 185
rect 8446 140 8451 165
rect 8476 140 8481 165
rect 8446 120 8481 140
rect 8446 95 8451 120
rect 8476 95 8481 120
rect 8446 85 8481 95
rect 8506 165 8541 185
rect 8506 140 8511 165
rect 8536 140 8541 165
rect 8506 120 8541 140
rect 8506 95 8511 120
rect 8536 95 8541 120
rect 8506 85 8541 95
rect 8566 165 8601 185
rect 8566 140 8571 165
rect 8596 140 8601 165
rect 8566 120 8601 140
rect 8566 95 8571 120
rect 8596 95 8601 120
rect 8566 85 8601 95
rect 8626 165 8661 185
rect 8626 140 8631 165
rect 8656 140 8661 165
rect 8626 120 8661 140
rect 8626 95 8631 120
rect 8656 95 8661 120
rect 8626 85 8661 95
rect 8686 165 8721 185
rect 8686 140 8691 165
rect 8716 140 8721 165
rect 8686 120 8721 140
rect 8686 95 8691 120
rect 8716 95 8721 120
rect 8686 85 8721 95
rect 8746 165 8786 185
rect 8746 140 8756 165
rect 8781 140 8786 165
rect 8746 120 8786 140
rect 8746 95 8756 120
rect 8781 95 8786 120
rect 8746 85 8786 95
rect 8811 165 8846 185
rect 8811 140 8816 165
rect 8841 140 8846 165
rect 8811 120 8846 140
rect 8811 95 8816 120
rect 8841 95 8846 120
rect 8811 85 8846 95
rect 8871 165 8906 185
rect 8871 140 8876 165
rect 8901 140 8906 165
rect 8871 120 8906 140
rect 8871 95 8876 120
rect 8901 95 8906 120
rect 8871 85 8906 95
rect 8931 165 8966 185
rect 8931 140 8936 165
rect 8961 140 8966 165
rect 8931 120 8966 140
rect 8931 95 8936 120
rect 8961 95 8966 120
rect 8931 85 8966 95
rect 8991 165 9026 185
rect 8991 140 8996 165
rect 9021 140 9026 165
rect 8991 120 9026 140
rect 8991 95 8996 120
rect 9021 95 9026 120
rect 8991 85 9026 95
rect 9051 165 9086 185
rect 9051 140 9056 165
rect 9081 140 9086 165
rect 9051 120 9086 140
rect 9051 95 9056 120
rect 9081 95 9086 120
rect 9051 85 9086 95
rect 9111 165 9146 185
rect 9111 140 9116 165
rect 9141 140 9146 165
rect 9111 120 9146 140
rect 9111 95 9116 120
rect 9141 95 9146 120
rect 9111 85 9146 95
rect 9171 165 9206 185
rect 9171 140 9176 165
rect 9201 140 9206 165
rect 9171 120 9206 140
rect 9171 95 9176 120
rect 9201 95 9206 120
rect 9171 85 9206 95
rect 9231 165 9271 185
rect 9231 140 9241 165
rect 9266 140 9271 165
rect 9231 120 9271 140
rect 9231 95 9241 120
rect 9266 95 9271 120
rect 9231 85 9271 95
rect 9296 165 9331 185
rect 9296 140 9301 165
rect 9326 140 9331 165
rect 9296 120 9331 140
rect 9296 95 9301 120
rect 9326 95 9331 120
rect 9296 85 9331 95
rect 9356 165 9391 185
rect 9356 140 9361 165
rect 9386 140 9391 165
rect 9356 120 9391 140
rect 9356 95 9361 120
rect 9386 95 9391 120
rect 9356 85 9391 95
rect 9416 165 9451 185
rect 9416 140 9421 165
rect 9446 140 9451 165
rect 9416 120 9451 140
rect 9416 95 9421 120
rect 9446 95 9451 120
rect 9416 85 9451 95
rect 9476 165 9516 185
rect 9476 140 9486 165
rect 9511 140 9516 165
rect 9476 120 9516 140
rect 9476 95 9486 120
rect 9511 95 9516 120
rect 9476 85 9516 95
rect 9541 165 9576 185
rect 9541 140 9546 165
rect 9571 140 9576 165
rect 9541 120 9576 140
rect 9541 95 9546 120
rect 9571 95 9576 120
rect 9541 85 9576 95
rect 9601 165 9636 185
rect 9601 140 9606 165
rect 9631 140 9636 165
rect 9601 120 9636 140
rect 9601 95 9606 120
rect 9631 95 9636 120
rect 9601 85 9636 95
rect 9661 165 9696 185
rect 9661 140 9666 165
rect 9691 140 9696 165
rect 9661 120 9696 140
rect 9661 95 9666 120
rect 9691 95 9696 120
rect 9661 85 9696 95
rect 9721 165 9761 185
rect 9721 140 9731 165
rect 9756 140 9761 165
rect 9721 120 9761 140
rect 9721 95 9731 120
rect 9756 95 9761 120
rect 9721 85 9761 95
rect 9786 165 9821 185
rect 9786 140 9791 165
rect 9816 140 9821 165
rect 9786 120 9821 140
rect 9786 95 9791 120
rect 9816 95 9821 120
rect 9786 85 9821 95
rect 9846 165 9881 185
rect 9846 140 9851 165
rect 9876 140 9881 165
rect 9846 120 9881 140
rect 9846 95 9851 120
rect 9876 95 9881 120
rect 9846 85 9881 95
rect 9906 165 9941 185
rect 9906 140 9911 165
rect 9936 140 9941 165
rect 9906 120 9941 140
rect 9906 95 9911 120
rect 9936 95 9941 120
rect 9906 85 9941 95
rect 9966 165 10001 185
rect 9966 140 9971 165
rect 9996 140 10001 165
rect 9966 120 10001 140
rect 9966 95 9971 120
rect 9996 95 10001 120
rect 9966 85 10001 95
rect 10026 165 10061 185
rect 10026 140 10031 165
rect 10056 140 10061 165
rect 10026 120 10061 140
rect 10026 95 10031 120
rect 10056 95 10061 120
rect 10026 85 10061 95
rect 10086 165 10121 185
rect 10086 140 10091 165
rect 10116 140 10121 165
rect 10086 120 10121 140
rect 10086 95 10091 120
rect 10116 95 10121 120
rect 10086 85 10121 95
rect 10146 165 10181 185
rect 10146 140 10151 165
rect 10176 140 10181 165
rect 10146 120 10181 140
rect 10146 95 10151 120
rect 10176 95 10181 120
rect 10146 85 10181 95
rect 10206 165 10246 185
rect 10206 140 10216 165
rect 10241 140 10246 165
rect 10206 120 10246 140
rect 10206 95 10216 120
rect 10241 95 10246 120
rect 10206 85 10246 95
rect 10271 165 10306 185
rect 10271 140 10276 165
rect 10301 140 10306 165
rect 10271 120 10306 140
rect 10271 95 10276 120
rect 10301 95 10306 120
rect 10271 85 10306 95
rect 10331 165 10366 185
rect 10331 140 10336 165
rect 10361 140 10366 165
rect 10331 120 10366 140
rect 10331 95 10336 120
rect 10361 95 10366 120
rect 10331 85 10366 95
rect 10391 165 10426 185
rect 10391 140 10396 165
rect 10421 140 10426 165
rect 10391 120 10426 140
rect 10391 95 10396 120
rect 10421 95 10426 120
rect 10391 85 10426 95
rect 10451 165 10486 185
rect 10451 140 10456 165
rect 10481 140 10486 165
rect 10451 120 10486 140
rect 10451 95 10456 120
rect 10481 95 10486 120
rect 10451 85 10486 95
rect 10511 165 10546 185
rect 10511 140 10516 165
rect 10541 140 10546 165
rect 10511 120 10546 140
rect 10511 95 10516 120
rect 10541 95 10546 120
rect 10511 85 10546 95
rect 10571 165 10606 185
rect 10571 140 10576 165
rect 10601 140 10606 165
rect 10571 120 10606 140
rect 10571 95 10576 120
rect 10601 95 10606 120
rect 10571 85 10606 95
rect 10631 165 10666 185
rect 10631 140 10636 165
rect 10661 140 10666 165
rect 10631 120 10666 140
rect 10631 95 10636 120
rect 10661 95 10666 120
rect 10631 85 10666 95
rect 10691 165 10731 185
rect 10691 140 10701 165
rect 10726 140 10731 165
rect 10691 120 10731 140
rect 10691 95 10701 120
rect 10726 95 10731 120
rect 10691 85 10731 95
rect 10756 165 10791 185
rect 10756 140 10761 165
rect 10786 140 10791 165
rect 10756 120 10791 140
rect 10756 95 10761 120
rect 10786 95 10791 120
rect 10756 85 10791 95
rect 10816 165 10851 185
rect 10816 140 10821 165
rect 10846 140 10851 165
rect 10816 120 10851 140
rect 10816 95 10821 120
rect 10846 95 10851 120
rect 10816 85 10851 95
rect 10876 165 10911 185
rect 10876 140 10881 165
rect 10906 140 10911 165
rect 10876 120 10911 140
rect 10876 95 10881 120
rect 10906 95 10911 120
rect 10876 85 10911 95
rect 10936 165 10971 185
rect 10936 140 10941 165
rect 10966 140 10971 165
rect 10936 120 10971 140
rect 10936 95 10941 120
rect 10966 95 10971 120
rect 10936 85 10971 95
rect 10996 165 11031 185
rect 10996 140 11001 165
rect 11026 140 11031 165
rect 10996 120 11031 140
rect 10996 95 11001 120
rect 11026 95 11031 120
rect 10996 85 11031 95
rect 11056 165 11091 185
rect 11056 140 11061 165
rect 11086 140 11091 165
rect 11056 120 11091 140
rect 11056 95 11061 120
rect 11086 95 11091 120
rect 11056 85 11091 95
rect 11116 165 11151 185
rect 11116 140 11121 165
rect 11146 140 11151 165
rect 11116 120 11151 140
rect 11116 95 11121 120
rect 11146 95 11151 120
rect 11116 85 11151 95
rect 11176 165 11216 185
rect 11176 140 11186 165
rect 11211 140 11216 165
rect 11176 120 11216 140
rect 11176 95 11186 120
rect 11211 95 11216 120
rect 11176 85 11216 95
rect 11241 165 11276 185
rect 11241 140 11246 165
rect 11271 140 11276 165
rect 11241 120 11276 140
rect 11241 95 11246 120
rect 11271 95 11276 120
rect 11241 85 11276 95
rect 11301 165 11336 185
rect 11301 140 11306 165
rect 11331 140 11336 165
rect 11301 120 11336 140
rect 11301 95 11306 120
rect 11331 95 11336 120
rect 11301 85 11336 95
rect 11361 165 11396 185
rect 11361 140 11366 165
rect 11391 140 11396 165
rect 11361 120 11396 140
rect 11361 95 11366 120
rect 11391 95 11396 120
rect 11361 85 11396 95
rect 11421 165 11456 185
rect 11421 140 11426 165
rect 11451 140 11456 165
rect 11421 120 11456 140
rect 11421 95 11426 120
rect 11451 95 11456 120
rect 11421 85 11456 95
rect 11481 165 11516 185
rect 11481 140 11486 165
rect 11511 140 11516 165
rect 11481 120 11516 140
rect 11481 95 11486 120
rect 11511 95 11516 120
rect 11481 85 11516 95
rect 11541 165 11576 185
rect 11541 140 11546 165
rect 11571 140 11576 165
rect 11541 120 11576 140
rect 11541 95 11546 120
rect 11571 95 11576 120
rect 11541 85 11576 95
rect 11601 165 11636 185
rect 11601 140 11606 165
rect 11631 140 11636 165
rect 11601 120 11636 140
rect 11601 95 11606 120
rect 11631 95 11636 120
rect 11601 85 11636 95
rect 11661 165 11701 185
rect 11661 140 11671 165
rect 11696 140 11701 165
rect 11661 120 11701 140
rect 11661 95 11671 120
rect 11696 95 11701 120
rect 11661 85 11701 95
rect 11726 165 11761 185
rect 11726 140 11731 165
rect 11756 140 11761 165
rect 11726 120 11761 140
rect 11726 95 11731 120
rect 11756 95 11761 120
rect 11726 85 11761 95
rect 11786 165 11821 185
rect 11786 140 11791 165
rect 11816 140 11821 165
rect 11786 120 11821 140
rect 11786 95 11791 120
rect 11816 95 11821 120
rect 11786 85 11821 95
rect 11846 165 11881 185
rect 11846 140 11851 165
rect 11876 140 11881 165
rect 11846 120 11881 140
rect 11846 95 11851 120
rect 11876 95 11881 120
rect 11846 85 11881 95
rect 11906 165 11941 185
rect 11906 140 11911 165
rect 11936 140 11941 165
rect 11906 120 11941 140
rect 11906 95 11911 120
rect 11936 95 11941 120
rect 11906 85 11941 95
rect 11966 165 12001 185
rect 11966 140 11971 165
rect 11996 140 12001 165
rect 11966 120 12001 140
rect 11966 95 11971 120
rect 11996 95 12001 120
rect 11966 85 12001 95
rect 12026 165 12061 185
rect 12026 140 12031 165
rect 12056 140 12061 165
rect 12026 120 12061 140
rect 12026 95 12031 120
rect 12056 95 12061 120
rect 12026 85 12061 95
rect 12086 165 12121 185
rect 12086 140 12091 165
rect 12116 140 12121 165
rect 12086 120 12121 140
rect 12086 95 12091 120
rect 12116 95 12121 120
rect 12086 85 12121 95
rect 12146 165 12186 185
rect 12146 140 12156 165
rect 12181 140 12186 165
rect 12146 120 12186 140
rect 12146 95 12156 120
rect 12181 95 12186 120
rect 12146 85 12186 95
rect 12211 165 12246 185
rect 12211 140 12216 165
rect 12241 140 12246 165
rect 12211 120 12246 140
rect 12211 95 12216 120
rect 12241 95 12246 120
rect 12211 85 12246 95
rect 12271 165 12306 185
rect 12271 140 12276 165
rect 12301 140 12306 165
rect 12271 120 12306 140
rect 12271 95 12276 120
rect 12301 95 12306 120
rect 12271 85 12306 95
rect 12331 165 12366 185
rect 12331 140 12336 165
rect 12361 140 12366 165
rect 12331 120 12366 140
rect 12331 95 12336 120
rect 12361 95 12366 120
rect 12331 85 12366 95
rect 12391 165 12426 185
rect 12391 140 12396 165
rect 12421 140 12426 165
rect 12391 120 12426 140
rect 12391 95 12396 120
rect 12421 95 12426 120
rect 12391 85 12426 95
rect 12451 165 12486 185
rect 12451 140 12456 165
rect 12481 140 12486 165
rect 12451 120 12486 140
rect 12451 95 12456 120
rect 12481 95 12486 120
rect 12451 85 12486 95
rect 12511 165 12546 185
rect 12511 140 12516 165
rect 12541 140 12546 165
rect 12511 120 12546 140
rect 12511 95 12516 120
rect 12541 95 12546 120
rect 12511 85 12546 95
rect 12571 165 12606 185
rect 12571 140 12576 165
rect 12601 140 12606 165
rect 12571 120 12606 140
rect 12571 95 12576 120
rect 12601 95 12606 120
rect 12571 85 12606 95
rect 12631 165 12671 185
rect 12631 140 12641 165
rect 12666 140 12671 165
rect 12631 120 12671 140
rect 12631 95 12641 120
rect 12666 95 12671 120
rect 12631 85 12671 95
rect 12696 165 12731 185
rect 12696 140 12701 165
rect 12726 140 12731 165
rect 12696 120 12731 140
rect 12696 95 12701 120
rect 12726 95 12731 120
rect 12696 85 12731 95
rect 12756 165 12791 185
rect 12756 140 12761 165
rect 12786 140 12791 165
rect 12756 120 12791 140
rect 12756 95 12761 120
rect 12786 95 12791 120
rect 12756 85 12791 95
rect 12816 165 12851 185
rect 12816 140 12821 165
rect 12846 140 12851 165
rect 12816 120 12851 140
rect 12816 95 12821 120
rect 12846 95 12851 120
rect 12816 85 12851 95
rect 12876 165 12911 185
rect 12876 140 12881 165
rect 12906 140 12911 165
rect 12876 120 12911 140
rect 12876 95 12881 120
rect 12906 95 12911 120
rect 12876 85 12911 95
rect 12936 165 12971 185
rect 12936 140 12941 165
rect 12966 140 12971 165
rect 12936 120 12971 140
rect 12936 95 12941 120
rect 12966 95 12971 120
rect 12936 85 12971 95
rect 12996 165 13031 185
rect 12996 140 13001 165
rect 13026 140 13031 165
rect 12996 120 13031 140
rect 12996 95 13001 120
rect 13026 95 13031 120
rect 12996 85 13031 95
rect 13056 165 13091 185
rect 13056 140 13061 165
rect 13086 140 13091 165
rect 13056 120 13091 140
rect 13056 95 13061 120
rect 13086 95 13091 120
rect 13056 85 13091 95
rect 13116 165 13156 185
rect 13116 140 13126 165
rect 13151 140 13156 165
rect 13116 120 13156 140
rect 13116 95 13126 120
rect 13151 95 13156 120
rect 13116 85 13156 95
rect 13181 165 13216 185
rect 13181 140 13186 165
rect 13211 140 13216 165
rect 13181 120 13216 140
rect 13181 95 13186 120
rect 13211 95 13216 120
rect 13181 85 13216 95
rect 13241 165 13276 185
rect 13241 140 13246 165
rect 13271 140 13276 165
rect 13241 120 13276 140
rect 13241 95 13246 120
rect 13271 95 13276 120
rect 13241 85 13276 95
rect 13301 165 13336 185
rect 13301 140 13306 165
rect 13331 140 13336 165
rect 13301 120 13336 140
rect 13301 95 13306 120
rect 13331 95 13336 120
rect 13301 85 13336 95
rect 13361 165 13396 185
rect 13361 140 13366 165
rect 13391 140 13396 165
rect 13361 120 13396 140
rect 13361 95 13366 120
rect 13391 95 13396 120
rect 13361 85 13396 95
rect 13421 165 13456 185
rect 13421 140 13426 165
rect 13451 140 13456 165
rect 13421 120 13456 140
rect 13421 95 13426 120
rect 13451 95 13456 120
rect 13421 85 13456 95
rect 13481 165 13516 185
rect 13481 140 13486 165
rect 13511 140 13516 165
rect 13481 120 13516 140
rect 13481 95 13486 120
rect 13511 95 13516 120
rect 13481 85 13516 95
rect 13541 165 13576 185
rect 13541 140 13546 165
rect 13571 140 13576 165
rect 13541 120 13576 140
rect 13541 95 13546 120
rect 13571 95 13576 120
rect 13541 85 13576 95
rect 13601 165 13641 185
rect 13601 140 13611 165
rect 13636 140 13641 165
rect 13601 120 13641 140
rect 13601 95 13611 120
rect 13636 95 13641 120
rect 13601 85 13641 95
rect 13666 165 13701 185
rect 13666 140 13671 165
rect 13696 140 13701 165
rect 13666 120 13701 140
rect 13666 95 13671 120
rect 13696 95 13701 120
rect 13666 85 13701 95
rect 13726 165 13761 185
rect 13726 140 13731 165
rect 13756 140 13761 165
rect 13726 120 13761 140
rect 13726 95 13731 120
rect 13756 95 13761 120
rect 13726 85 13761 95
rect 13786 165 13821 185
rect 13786 140 13791 165
rect 13816 140 13821 165
rect 13786 120 13821 140
rect 13786 95 13791 120
rect 13816 95 13821 120
rect 13786 85 13821 95
rect 13846 165 13881 185
rect 13846 140 13851 165
rect 13876 140 13881 165
rect 13846 120 13881 140
rect 13846 95 13851 120
rect 13876 95 13881 120
rect 13846 85 13881 95
rect 13906 165 13941 185
rect 13906 140 13911 165
rect 13936 140 13941 165
rect 13906 120 13941 140
rect 13906 95 13911 120
rect 13936 95 13941 120
rect 13906 85 13941 95
rect 13966 165 14001 185
rect 13966 140 13971 165
rect 13996 140 14001 165
rect 13966 120 14001 140
rect 13966 95 13971 120
rect 13996 95 14001 120
rect 13966 85 14001 95
rect 14026 165 14061 185
rect 14026 140 14031 165
rect 14056 140 14061 165
rect 14026 120 14061 140
rect 14026 95 14031 120
rect 14056 95 14061 120
rect 14026 85 14061 95
rect 14086 165 14126 185
rect 14086 140 14096 165
rect 14121 140 14126 165
rect 14086 120 14126 140
rect 14086 95 14096 120
rect 14121 95 14126 120
rect 14086 85 14126 95
rect 14151 165 14186 185
rect 14151 140 14156 165
rect 14181 140 14186 165
rect 14151 120 14186 140
rect 14151 95 14156 120
rect 14181 95 14186 120
rect 14151 85 14186 95
rect 14211 165 14246 185
rect 14211 140 14216 165
rect 14241 140 14246 165
rect 14211 120 14246 140
rect 14211 95 14216 120
rect 14241 95 14246 120
rect 14211 85 14246 95
rect 14271 165 14306 185
rect 14271 140 14276 165
rect 14301 140 14306 165
rect 14271 120 14306 140
rect 14271 95 14276 120
rect 14301 95 14306 120
rect 14271 85 14306 95
rect 14331 165 14366 185
rect 14331 140 14336 165
rect 14361 140 14366 165
rect 14331 120 14366 140
rect 14331 95 14336 120
rect 14361 95 14366 120
rect 14331 85 14366 95
rect 14391 165 14426 185
rect 14391 140 14396 165
rect 14421 140 14426 165
rect 14391 120 14426 140
rect 14391 95 14396 120
rect 14421 95 14426 120
rect 14391 85 14426 95
rect 14451 165 14486 185
rect 14451 140 14456 165
rect 14481 140 14486 165
rect 14451 120 14486 140
rect 14451 95 14456 120
rect 14481 95 14486 120
rect 14451 85 14486 95
rect 14511 165 14546 185
rect 14511 140 14516 165
rect 14541 140 14546 165
rect 14511 120 14546 140
rect 14511 95 14516 120
rect 14541 95 14546 120
rect 14511 85 14546 95
rect 14571 165 14611 185
rect 14571 140 14581 165
rect 14606 140 14611 165
rect 14571 120 14611 140
rect 14571 95 14581 120
rect 14606 95 14611 120
rect 14571 85 14611 95
rect 14636 165 14671 185
rect 14636 140 14641 165
rect 14666 140 14671 165
rect 14636 120 14671 140
rect 14636 95 14641 120
rect 14666 95 14671 120
rect 14636 85 14671 95
rect 14696 165 14731 185
rect 14696 140 14701 165
rect 14726 140 14731 165
rect 14696 120 14731 140
rect 14696 95 14701 120
rect 14726 95 14731 120
rect 14696 85 14731 95
rect 14756 165 14791 185
rect 14756 140 14761 165
rect 14786 140 14791 165
rect 14756 120 14791 140
rect 14756 95 14761 120
rect 14786 95 14791 120
rect 14756 85 14791 95
rect 14816 165 14851 185
rect 14816 140 14821 165
rect 14846 140 14851 165
rect 14816 120 14851 140
rect 14816 95 14821 120
rect 14846 95 14851 120
rect 14816 85 14851 95
rect 14876 165 14911 185
rect 14876 140 14881 165
rect 14906 140 14911 165
rect 14876 120 14911 140
rect 14876 95 14881 120
rect 14906 95 14911 120
rect 14876 85 14911 95
rect 14936 165 14971 185
rect 14936 140 14941 165
rect 14966 140 14971 165
rect 14936 120 14971 140
rect 14936 95 14941 120
rect 14966 95 14971 120
rect 14936 85 14971 95
rect 14996 165 15031 185
rect 14996 140 15001 165
rect 15026 140 15031 165
rect 14996 120 15031 140
rect 14996 95 15001 120
rect 15026 95 15031 120
rect 14996 85 15031 95
rect 15056 165 15096 185
rect 15056 140 15066 165
rect 15091 140 15096 165
rect 15056 120 15096 140
rect 15056 95 15066 120
rect 15091 95 15096 120
rect 15056 85 15096 95
rect 15121 165 15156 185
rect 15121 140 15126 165
rect 15151 140 15156 165
rect 15121 120 15156 140
rect 15121 95 15126 120
rect 15151 95 15156 120
rect 15121 85 15156 95
rect 15181 165 15216 185
rect 15181 140 15186 165
rect 15211 140 15216 165
rect 15181 120 15216 140
rect 15181 95 15186 120
rect 15211 95 15216 120
rect 15181 85 15216 95
rect 15241 165 15276 185
rect 15241 140 15246 165
rect 15271 140 15276 165
rect 15241 120 15276 140
rect 15241 95 15246 120
rect 15271 95 15276 120
rect 15241 85 15276 95
rect 15301 165 15336 185
rect 15301 140 15306 165
rect 15331 140 15336 165
rect 15301 120 15336 140
rect 15301 95 15306 120
rect 15331 95 15336 120
rect 15301 85 15336 95
rect 15361 165 15396 185
rect 15361 140 15366 165
rect 15391 140 15396 165
rect 15361 120 15396 140
rect 15361 95 15366 120
rect 15391 95 15396 120
rect 15361 85 15396 95
rect 15421 165 15456 185
rect 15421 140 15426 165
rect 15451 140 15456 165
rect 15421 120 15456 140
rect 15421 95 15426 120
rect 15451 95 15456 120
rect 15421 85 15456 95
rect 15481 165 15516 185
rect 15481 140 15486 165
rect 15511 140 15516 165
rect 15481 120 15516 140
rect 15481 95 15486 120
rect 15511 95 15516 120
rect 15481 85 15516 95
rect 15541 165 15581 185
rect 15541 140 15551 165
rect 15576 140 15581 165
rect 15541 120 15581 140
rect 15541 95 15551 120
rect 15576 95 15581 120
rect 15541 85 15581 95
rect 15606 165 15641 185
rect 15606 140 15611 165
rect 15636 140 15641 165
rect 15606 120 15641 140
rect 15606 95 15611 120
rect 15636 95 15641 120
rect 15606 85 15641 95
rect 15666 165 15701 185
rect 15666 140 15671 165
rect 15696 140 15701 165
rect 15666 120 15701 140
rect 15666 95 15671 120
rect 15696 95 15701 120
rect 15666 85 15701 95
rect 15726 165 15761 185
rect 15726 140 15731 165
rect 15756 140 15761 165
rect 15726 120 15761 140
rect 15726 95 15731 120
rect 15756 95 15761 120
rect 15726 85 15761 95
rect 15786 165 15821 185
rect 15786 140 15791 165
rect 15816 140 15821 165
rect 15786 120 15821 140
rect 15786 95 15791 120
rect 15816 95 15821 120
rect 15786 85 15821 95
rect 15846 165 15881 185
rect 15846 140 15851 165
rect 15876 140 15881 165
rect 15846 120 15881 140
rect 15846 95 15851 120
rect 15876 95 15881 120
rect 15846 85 15881 95
rect 15906 165 15941 185
rect 15906 140 15911 165
rect 15936 140 15941 165
rect 15906 120 15941 140
rect 15906 95 15911 120
rect 15936 95 15941 120
rect 15906 85 15941 95
rect 15966 165 16001 185
rect 15966 140 15971 165
rect 15996 140 16001 165
rect 15966 120 16001 140
rect 15966 95 15971 120
rect 15996 95 16001 120
rect 15966 85 16001 95
rect 16026 165 16066 185
rect 16026 140 16036 165
rect 16061 140 16066 165
rect 16026 120 16066 140
rect 16026 95 16036 120
rect 16061 95 16066 120
rect 16026 85 16066 95
rect 16091 165 16126 185
rect 16091 140 16096 165
rect 16121 140 16126 165
rect 16091 120 16126 140
rect 16091 95 16096 120
rect 16121 95 16126 120
rect 16091 85 16126 95
rect 16151 165 16186 185
rect 16151 140 16156 165
rect 16181 140 16186 165
rect 16151 120 16186 140
rect 16151 95 16156 120
rect 16181 95 16186 120
rect 16151 85 16186 95
rect 16211 165 16246 185
rect 16211 140 16216 165
rect 16241 140 16246 165
rect 16211 120 16246 140
rect 16211 95 16216 120
rect 16241 95 16246 120
rect 16211 85 16246 95
rect 16271 165 16306 185
rect 16271 140 16276 165
rect 16301 140 16306 165
rect 16271 120 16306 140
rect 16271 95 16276 120
rect 16301 95 16306 120
rect 16271 85 16306 95
rect 16331 165 16366 185
rect 16331 140 16336 165
rect 16361 140 16366 165
rect 16331 120 16366 140
rect 16331 95 16336 120
rect 16361 95 16366 120
rect 16331 85 16366 95
rect 16391 165 16426 185
rect 16391 140 16396 165
rect 16421 140 16426 165
rect 16391 120 16426 140
rect 16391 95 16396 120
rect 16421 95 16426 120
rect 16391 85 16426 95
rect 16451 165 16486 185
rect 16451 140 16456 165
rect 16481 140 16486 165
rect 16451 120 16486 140
rect 16451 95 16456 120
rect 16481 95 16486 120
rect 16451 85 16486 95
rect 16511 165 16551 185
rect 16511 140 16521 165
rect 16546 140 16551 165
rect 16511 120 16551 140
rect 16511 95 16521 120
rect 16546 95 16551 120
rect 16511 85 16551 95
rect 16576 165 16611 185
rect 16576 140 16581 165
rect 16606 140 16611 165
rect 16576 120 16611 140
rect 16576 95 16581 120
rect 16606 95 16611 120
rect 16576 85 16611 95
rect 16636 165 16671 185
rect 16636 140 16641 165
rect 16666 140 16671 165
rect 16636 120 16671 140
rect 16636 95 16641 120
rect 16666 95 16671 120
rect 16636 85 16671 95
rect 16696 165 16731 185
rect 16696 140 16701 165
rect 16726 140 16731 165
rect 16696 120 16731 140
rect 16696 95 16701 120
rect 16726 95 16731 120
rect 16696 85 16731 95
rect 16756 165 16791 185
rect 16756 140 16761 165
rect 16786 140 16791 165
rect 16756 120 16791 140
rect 16756 95 16761 120
rect 16786 95 16791 120
rect 16756 85 16791 95
rect 16816 165 16851 185
rect 16816 140 16821 165
rect 16846 140 16851 165
rect 16816 120 16851 140
rect 16816 95 16821 120
rect 16846 95 16851 120
rect 16816 85 16851 95
rect 16876 165 16911 185
rect 16876 140 16881 165
rect 16906 140 16911 165
rect 16876 120 16911 140
rect 16876 95 16881 120
rect 16906 95 16911 120
rect 16876 85 16911 95
rect 16936 165 16971 185
rect 16936 140 16941 165
rect 16966 140 16971 165
rect 16936 120 16971 140
rect 16936 95 16941 120
rect 16966 95 16971 120
rect 16936 85 16971 95
rect 16996 165 17036 185
rect 16996 140 17006 165
rect 17031 140 17036 165
rect 16996 120 17036 140
rect 16996 95 17006 120
rect 17031 95 17036 120
rect 16996 85 17036 95
rect 17061 165 17096 185
rect 17061 140 17066 165
rect 17091 140 17096 165
rect 17061 120 17096 140
rect 17061 95 17066 120
rect 17091 95 17096 120
rect 17061 85 17096 95
rect 17121 165 17156 185
rect 17121 140 17126 165
rect 17151 140 17156 165
rect 17121 120 17156 140
rect 17121 95 17126 120
rect 17151 95 17156 120
rect 17121 85 17156 95
rect 17181 165 17216 185
rect 17181 140 17186 165
rect 17211 140 17216 165
rect 17181 120 17216 140
rect 17181 95 17186 120
rect 17211 95 17216 120
rect 17181 85 17216 95
rect 17241 165 17276 185
rect 17241 140 17246 165
rect 17271 140 17276 165
rect 17241 120 17276 140
rect 17241 95 17246 120
rect 17271 95 17276 120
rect 17241 85 17276 95
rect 17301 165 17336 185
rect 17301 140 17306 165
rect 17331 140 17336 165
rect 17301 120 17336 140
rect 17301 95 17306 120
rect 17331 95 17336 120
rect 17301 85 17336 95
rect 17361 165 17396 185
rect 17361 140 17366 165
rect 17391 140 17396 165
rect 17361 120 17396 140
rect 17361 95 17366 120
rect 17391 95 17396 120
rect 17361 85 17396 95
rect 17421 165 17456 185
rect 17421 140 17426 165
rect 17451 140 17456 165
rect 17421 120 17456 140
rect 17421 95 17426 120
rect 17451 95 17456 120
rect 17421 85 17456 95
rect 17481 165 17521 185
rect 17481 140 17491 165
rect 17516 140 17521 165
rect 17481 120 17521 140
rect 17481 95 17491 120
rect 17516 95 17521 120
rect 17481 85 17521 95
rect 17546 165 17581 185
rect 17546 140 17551 165
rect 17576 140 17581 165
rect 17546 120 17581 140
rect 17546 95 17551 120
rect 17576 95 17581 120
rect 17546 85 17581 95
rect 17606 165 17641 185
rect 17606 140 17611 165
rect 17636 140 17641 165
rect 17606 120 17641 140
rect 17606 95 17611 120
rect 17636 95 17641 120
rect 17606 85 17641 95
rect 17666 165 17701 185
rect 17666 140 17671 165
rect 17696 140 17701 165
rect 17666 120 17701 140
rect 17666 95 17671 120
rect 17696 95 17701 120
rect 17666 85 17701 95
rect 17726 165 17761 185
rect 17726 140 17731 165
rect 17756 140 17761 165
rect 17726 120 17761 140
rect 17726 95 17731 120
rect 17756 95 17761 120
rect 17726 85 17761 95
rect 17786 165 17821 185
rect 17786 140 17791 165
rect 17816 140 17821 165
rect 17786 120 17821 140
rect 17786 95 17791 120
rect 17816 95 17821 120
rect 17786 85 17821 95
rect 17846 165 17881 185
rect 17846 140 17851 165
rect 17876 140 17881 165
rect 17846 120 17881 140
rect 17846 95 17851 120
rect 17876 95 17881 120
rect 17846 85 17881 95
rect 17906 165 17941 185
rect 17906 140 17911 165
rect 17936 140 17941 165
rect 17906 120 17941 140
rect 17906 95 17911 120
rect 17936 95 17941 120
rect 17906 85 17941 95
rect 17966 165 18006 185
rect 17966 140 17976 165
rect 18001 140 18006 165
rect 17966 120 18006 140
rect 17966 95 17976 120
rect 18001 95 18006 120
rect 17966 85 18006 95
rect 18031 165 18066 185
rect 18031 140 18036 165
rect 18061 140 18066 165
rect 18031 120 18066 140
rect 18031 95 18036 120
rect 18061 95 18066 120
rect 18031 85 18066 95
rect 18091 165 18126 185
rect 18091 140 18096 165
rect 18121 140 18126 165
rect 18091 120 18126 140
rect 18091 95 18096 120
rect 18121 95 18126 120
rect 18091 85 18126 95
rect 18151 165 18186 185
rect 18151 140 18156 165
rect 18181 140 18186 165
rect 18151 120 18186 140
rect 18151 95 18156 120
rect 18181 95 18186 120
rect 18151 85 18186 95
rect 18211 165 18246 185
rect 18211 140 18216 165
rect 18241 140 18246 165
rect 18211 120 18246 140
rect 18211 95 18216 120
rect 18241 95 18246 120
rect 18211 85 18246 95
rect 18271 165 18306 185
rect 18271 140 18276 165
rect 18301 140 18306 165
rect 18271 120 18306 140
rect 18271 95 18276 120
rect 18301 95 18306 120
rect 18271 85 18306 95
rect 18331 165 18366 185
rect 18331 140 18336 165
rect 18361 140 18366 165
rect 18331 120 18366 140
rect 18331 95 18336 120
rect 18361 95 18366 120
rect 18331 85 18366 95
rect 18391 165 18426 185
rect 18391 140 18396 165
rect 18421 140 18426 165
rect 18391 120 18426 140
rect 18391 95 18396 120
rect 18421 95 18426 120
rect 18391 85 18426 95
rect 18451 165 18491 185
rect 18451 140 18461 165
rect 18486 140 18491 165
rect 18451 120 18491 140
rect 18451 95 18461 120
rect 18486 95 18491 120
rect 18451 85 18491 95
rect 18516 165 18551 185
rect 18516 140 18521 165
rect 18546 140 18551 165
rect 18516 120 18551 140
rect 18516 95 18521 120
rect 18546 95 18551 120
rect 18516 85 18551 95
rect 18576 165 18611 185
rect 18576 140 18581 165
rect 18606 140 18611 165
rect 18576 120 18611 140
rect 18576 95 18581 120
rect 18606 95 18611 120
rect 18576 85 18611 95
rect 18636 165 18671 185
rect 18636 140 18641 165
rect 18666 140 18671 165
rect 18636 120 18671 140
rect 18636 95 18641 120
rect 18666 95 18671 120
rect 18636 85 18671 95
rect 18696 165 18731 185
rect 18696 140 18701 165
rect 18726 140 18731 165
rect 18696 120 18731 140
rect 18696 95 18701 120
rect 18726 95 18731 120
rect 18696 85 18731 95
rect 18756 165 18791 185
rect 18756 140 18761 165
rect 18786 140 18791 165
rect 18756 120 18791 140
rect 18756 95 18761 120
rect 18786 95 18791 120
rect 18756 85 18791 95
rect 18816 165 18851 185
rect 18816 140 18821 165
rect 18846 140 18851 165
rect 18816 120 18851 140
rect 18816 95 18821 120
rect 18846 95 18851 120
rect 18816 85 18851 95
rect 18876 165 18911 185
rect 18876 140 18881 165
rect 18906 140 18911 165
rect 18876 120 18911 140
rect 18876 95 18881 120
rect 18906 95 18911 120
rect 18876 85 18911 95
rect 18936 165 18976 185
rect 18936 140 18946 165
rect 18971 140 18976 165
rect 18936 120 18976 140
rect 18936 95 18946 120
rect 18971 95 18976 120
rect 18936 85 18976 95
rect 19001 165 19036 185
rect 19001 140 19006 165
rect 19031 140 19036 165
rect 19001 120 19036 140
rect 19001 95 19006 120
rect 19031 95 19036 120
rect 19001 85 19036 95
rect 19061 165 19096 185
rect 19061 140 19066 165
rect 19091 140 19096 165
rect 19061 120 19096 140
rect 19061 95 19066 120
rect 19091 95 19096 120
rect 19061 85 19096 95
rect 19121 165 19156 185
rect 19121 140 19126 165
rect 19151 140 19156 165
rect 19121 120 19156 140
rect 19121 95 19126 120
rect 19151 95 19156 120
rect 19121 85 19156 95
rect 19181 165 19216 185
rect 19181 140 19186 165
rect 19211 140 19216 165
rect 19181 120 19216 140
rect 19181 95 19186 120
rect 19211 95 19216 120
rect 19181 85 19216 95
rect 19241 165 19276 185
rect 19241 140 19246 165
rect 19271 140 19276 165
rect 19241 120 19276 140
rect 19241 95 19246 120
rect 19271 95 19276 120
rect 19241 85 19276 95
rect 19301 165 19336 185
rect 19301 140 19306 165
rect 19331 140 19336 165
rect 19301 120 19336 140
rect 19301 95 19306 120
rect 19331 95 19336 120
rect 19301 85 19336 95
rect 19361 165 19396 185
rect 19361 140 19366 165
rect 19391 140 19396 165
rect 19361 120 19396 140
rect 19361 95 19366 120
rect 19391 95 19396 120
rect 19361 85 19396 95
rect 19421 165 19461 185
rect 19421 140 19431 165
rect 19456 140 19461 165
rect 19421 120 19461 140
rect 19421 95 19431 120
rect 19456 95 19461 120
rect 19421 85 19461 95
rect 19486 165 19521 185
rect 19486 140 19491 165
rect 19516 140 19521 165
rect 19486 120 19521 140
rect 19486 95 19491 120
rect 19516 95 19521 120
rect 19486 85 19521 95
rect 19546 165 19581 185
rect 19546 140 19551 165
rect 19576 140 19581 165
rect 19546 120 19581 140
rect 19546 95 19551 120
rect 19576 95 19581 120
rect 19546 85 19581 95
rect 19606 165 19641 185
rect 19606 140 19611 165
rect 19636 140 19641 165
rect 19606 120 19641 140
rect 19606 95 19611 120
rect 19636 95 19641 120
rect 19606 85 19641 95
rect 19666 165 19701 185
rect 19666 140 19671 165
rect 19696 140 19701 165
rect 19666 120 19701 140
rect 19666 95 19671 120
rect 19696 95 19701 120
rect 19666 85 19701 95
rect 19726 165 19761 185
rect 19726 140 19731 165
rect 19756 140 19761 165
rect 19726 120 19761 140
rect 19726 95 19731 120
rect 19756 95 19761 120
rect 19726 85 19761 95
rect 19786 165 19821 185
rect 19786 140 19791 165
rect 19816 140 19821 165
rect 19786 120 19821 140
rect 19786 95 19791 120
rect 19816 95 19821 120
rect 19786 85 19821 95
rect 19846 165 19881 185
rect 19846 140 19851 165
rect 19876 140 19881 165
rect 19846 120 19881 140
rect 19846 95 19851 120
rect 19876 95 19881 120
rect 19846 85 19881 95
rect 19906 165 19946 185
rect 19906 140 19916 165
rect 19941 140 19946 165
rect 19906 120 19946 140
rect 19906 95 19916 120
rect 19941 95 19946 120
rect 19906 85 19946 95
rect 19971 165 20006 185
rect 19971 140 19976 165
rect 20001 140 20006 165
rect 19971 120 20006 140
rect 19971 95 19976 120
rect 20001 95 20006 120
rect 19971 85 20006 95
rect 20031 165 20066 185
rect 20031 140 20036 165
rect 20061 140 20066 165
rect 20031 120 20066 140
rect 20031 95 20036 120
rect 20061 95 20066 120
rect 20031 85 20066 95
rect 20091 165 20126 185
rect 20091 140 20096 165
rect 20121 140 20126 165
rect 20091 120 20126 140
rect 20091 95 20096 120
rect 20121 95 20126 120
rect 20091 85 20126 95
rect 20151 165 20186 185
rect 20151 140 20156 165
rect 20181 140 20186 165
rect 20151 120 20186 140
rect 20151 95 20156 120
rect 20181 95 20186 120
rect 20151 85 20186 95
rect 20211 165 20246 185
rect 20211 140 20216 165
rect 20241 140 20246 165
rect 20211 120 20246 140
rect 20211 95 20216 120
rect 20241 95 20246 120
rect 20211 85 20246 95
rect 20271 165 20306 185
rect 20271 140 20276 165
rect 20301 140 20306 165
rect 20271 120 20306 140
rect 20271 95 20276 120
rect 20301 95 20306 120
rect 20271 85 20306 95
rect 20331 165 20366 185
rect 20331 140 20336 165
rect 20361 140 20366 165
rect 20331 120 20366 140
rect 20331 95 20336 120
rect 20361 95 20366 120
rect 20331 85 20366 95
rect 20391 165 20431 185
rect 20391 140 20401 165
rect 20426 140 20431 165
rect 20391 120 20431 140
rect 20391 95 20401 120
rect 20426 95 20431 120
rect 20391 85 20431 95
rect 20456 165 20491 185
rect 20456 140 20461 165
rect 20486 140 20491 165
rect 20456 120 20491 140
rect 20456 95 20461 120
rect 20486 95 20491 120
rect 20456 85 20491 95
rect 20516 165 20551 185
rect 20516 140 20521 165
rect 20546 140 20551 165
rect 20516 120 20551 140
rect 20516 95 20521 120
rect 20546 95 20551 120
rect 20516 85 20551 95
rect 20576 165 20611 185
rect 20576 140 20581 165
rect 20606 140 20611 165
rect 20576 120 20611 140
rect 20576 95 20581 120
rect 20606 95 20611 120
rect 20576 85 20611 95
rect 20636 165 20671 185
rect 20636 140 20641 165
rect 20666 140 20671 165
rect 20636 120 20671 140
rect 20636 95 20641 120
rect 20666 95 20671 120
rect 20636 85 20671 95
rect 20696 165 20731 185
rect 20696 140 20701 165
rect 20726 140 20731 165
rect 20696 120 20731 140
rect 20696 95 20701 120
rect 20726 95 20731 120
rect 20696 85 20731 95
rect 20756 165 20791 185
rect 20756 140 20761 165
rect 20786 140 20791 165
rect 20756 120 20791 140
rect 20756 95 20761 120
rect 20786 95 20791 120
rect 20756 85 20791 95
rect 20816 165 20851 185
rect 20816 140 20821 165
rect 20846 140 20851 165
rect 20816 120 20851 140
rect 20816 95 20821 120
rect 20846 95 20851 120
rect 20816 85 20851 95
rect 20876 165 20916 185
rect 20876 140 20886 165
rect 20911 140 20916 165
rect 20876 120 20916 140
rect 20876 95 20886 120
rect 20911 95 20916 120
rect 20876 85 20916 95
rect 20941 165 20976 185
rect 20941 140 20946 165
rect 20971 140 20976 165
rect 20941 120 20976 140
rect 20941 95 20946 120
rect 20971 95 20976 120
rect 20941 85 20976 95
rect 21001 165 21036 185
rect 21001 140 21006 165
rect 21031 140 21036 165
rect 21001 120 21036 140
rect 21001 95 21006 120
rect 21031 95 21036 120
rect 21001 85 21036 95
rect 21061 165 21096 185
rect 21061 140 21066 165
rect 21091 140 21096 165
rect 21061 120 21096 140
rect 21061 95 21066 120
rect 21091 95 21096 120
rect 21061 85 21096 95
rect 21121 165 21156 185
rect 21121 140 21126 165
rect 21151 140 21156 165
rect 21121 120 21156 140
rect 21121 95 21126 120
rect 21151 95 21156 120
rect 21121 85 21156 95
rect 21520 165 21545 265
rect 21645 165 21670 265
rect 191 15 231 25
rect -190 -5 201 15
rect 221 -5 231 15
rect -460 -105 -440 -5
rect -340 -105 -320 -5
rect 191 -15 231 -5
rect 256 15 281 85
rect 326 75 346 85
rect 441 75 461 85
rect 316 15 356 25
rect 256 -5 326 15
rect 346 -5 356 15
rect 256 -70 281 -5
rect 316 -15 356 -5
rect 501 15 526 85
rect 561 75 581 85
rect 631 75 651 85
rect 746 75 766 85
rect 866 75 896 85
rect 866 55 876 75
rect 991 75 1011 85
rect 1111 75 1136 85
rect 1111 55 1116 75
rect 1231 75 1251 85
rect 1351 75 1381 85
rect 1351 55 1361 75
rect 1476 75 1496 85
rect 621 15 661 25
rect 501 -5 631 15
rect 651 -5 661 15
rect 326 -70 346 -65
rect 446 -50 466 -45
rect 501 -70 526 -5
rect 621 -15 661 -5
rect 1536 15 1561 85
rect 1596 75 1616 85
rect 1666 75 1686 85
rect 1781 75 1801 85
rect 1901 75 1931 85
rect 1901 55 1911 75
rect 2026 75 2046 85
rect 2146 75 2171 85
rect 2146 55 2151 75
rect 2266 75 2286 85
rect 2386 75 2416 85
rect 2386 55 2396 75
rect 2511 75 2531 85
rect 2631 75 2656 85
rect 2631 55 2636 75
rect 2751 75 2771 85
rect 2871 75 2901 85
rect 2871 55 2881 75
rect 2996 75 3016 85
rect 3116 75 3141 85
rect 3116 55 3121 75
rect 3236 75 3256 85
rect 3356 75 3386 85
rect 3356 55 3366 75
rect 3481 75 3501 85
rect 3596 75 3626 85
rect 3596 55 3606 75
rect 3721 75 3741 85
rect 3841 75 3871 85
rect 3841 55 3851 75
rect 3966 75 3986 85
rect 4086 75 4111 85
rect 4086 55 4091 75
rect 4206 75 4226 85
rect 4326 75 4356 85
rect 4326 55 4336 75
rect 4451 75 4471 85
rect 4571 75 4596 85
rect 4571 55 4576 75
rect 4691 75 4711 85
rect 4811 75 4841 85
rect 4811 55 4821 75
rect 4936 75 4956 85
rect 5056 75 5081 85
rect 5056 55 5061 75
rect 5176 75 5196 85
rect 5296 75 5326 85
rect 5296 55 5306 75
rect 5421 75 5441 85
rect 1656 15 1696 25
rect 1536 -5 1666 15
rect 1686 -5 1696 15
rect 631 -70 651 -65
rect 751 -50 771 -45
rect 866 -65 876 -50
rect 866 -70 896 -65
rect 996 -50 1016 -45
rect 1111 -65 1116 -50
rect 1111 -70 1136 -65
rect 1236 -50 1256 -45
rect 1351 -65 1361 -50
rect 1351 -70 1381 -65
rect 1481 -50 1501 -45
rect 1536 -70 1561 -5
rect 1656 -15 1696 -5
rect 5481 15 5506 85
rect 5541 75 5561 85
rect 5611 75 5631 85
rect 5726 75 5746 85
rect 5846 75 5876 85
rect 5846 55 5856 75
rect 5971 75 5991 85
rect 6091 75 6116 85
rect 6091 55 6096 75
rect 6211 75 6231 85
rect 6331 75 6361 85
rect 6331 55 6341 75
rect 6456 75 6476 85
rect 6576 75 6601 85
rect 6576 55 6581 75
rect 6696 75 6716 85
rect 6816 75 6846 85
rect 6816 55 6826 75
rect 6941 75 6961 85
rect 7061 75 7086 85
rect 7061 55 7066 75
rect 7181 75 7201 85
rect 7301 75 7326 85
rect 7301 55 7306 75
rect 7421 75 7441 85
rect 7536 75 7566 85
rect 7536 55 7546 75
rect 7661 75 7681 85
rect 7781 75 7811 85
rect 7781 55 7791 75
rect 7906 75 7926 85
rect 8026 75 8051 85
rect 8026 55 8031 75
rect 8146 75 8166 85
rect 8266 75 8296 85
rect 8266 55 8276 75
rect 8391 75 8411 85
rect 8511 75 8536 85
rect 8511 55 8516 75
rect 8631 75 8651 85
rect 8751 75 8781 85
rect 8751 55 8761 75
rect 8876 75 8896 85
rect 8996 75 9021 85
rect 8996 55 9001 75
rect 9116 75 9136 85
rect 9236 75 9266 85
rect 9236 55 9246 75
rect 9361 75 9381 85
rect 9481 75 9511 85
rect 9481 55 9491 75
rect 9606 75 9626 85
rect 9726 75 9756 85
rect 9726 55 9736 75
rect 9851 75 9871 85
rect 9971 75 9996 85
rect 9971 55 9976 75
rect 10091 75 10111 85
rect 10211 75 10241 85
rect 10211 55 10221 75
rect 10336 75 10356 85
rect 10456 75 10481 85
rect 10456 55 10461 75
rect 10576 75 10596 85
rect 10696 75 10726 85
rect 10696 55 10706 75
rect 10821 75 10841 85
rect 10941 75 10966 85
rect 10941 55 10946 75
rect 11061 75 11081 85
rect 11181 75 11211 85
rect 11181 55 11191 75
rect 11306 75 11326 85
rect 11421 75 11451 85
rect 11421 55 11431 75
rect 11546 75 11566 85
rect 11666 75 11696 85
rect 11666 55 11676 75
rect 11791 75 11811 85
rect 11911 75 11936 85
rect 11911 55 11916 75
rect 12031 75 12051 85
rect 12151 75 12181 85
rect 12151 55 12161 75
rect 12276 75 12296 85
rect 12396 75 12421 85
rect 12396 55 12401 75
rect 12516 75 12536 85
rect 12636 75 12666 85
rect 12636 55 12646 75
rect 12761 75 12781 85
rect 12881 75 12906 85
rect 12881 55 12886 75
rect 13001 75 13021 85
rect 13121 75 13151 85
rect 13121 55 13131 75
rect 13246 75 13266 85
rect 13366 75 13391 85
rect 13366 55 13371 75
rect 13486 75 13506 85
rect 13606 75 13636 85
rect 13606 55 13616 75
rect 13731 75 13751 85
rect 13851 75 13876 85
rect 13851 55 13856 75
rect 13971 75 13991 85
rect 14091 75 14121 85
rect 14091 55 14101 75
rect 14216 75 14236 85
rect 14336 75 14361 85
rect 14336 55 14341 75
rect 14456 75 14476 85
rect 14576 75 14606 85
rect 14576 55 14586 75
rect 14701 75 14721 85
rect 14821 75 14846 85
rect 14821 55 14826 75
rect 14941 75 14961 85
rect 15061 75 15091 85
rect 15061 55 15071 75
rect 15186 75 15206 85
rect 15301 75 15331 85
rect 15301 55 15311 75
rect 15426 75 15446 85
rect 15546 75 15576 85
rect 15546 55 15556 75
rect 15671 75 15691 85
rect 15791 75 15816 85
rect 15791 55 15796 75
rect 15911 75 15931 85
rect 16031 75 16061 85
rect 16031 55 16041 75
rect 16156 75 16176 85
rect 16276 75 16301 85
rect 16276 55 16281 75
rect 16396 75 16416 85
rect 16516 75 16546 85
rect 16516 55 16526 75
rect 16641 75 16661 85
rect 16761 75 16786 85
rect 16761 55 16766 75
rect 16881 75 16901 85
rect 17001 75 17031 85
rect 17001 55 17011 75
rect 17126 75 17146 85
rect 17246 75 17271 85
rect 17246 55 17251 75
rect 17366 75 17386 85
rect 17486 75 17516 85
rect 17486 55 17496 75
rect 17611 75 17631 85
rect 17731 75 17756 85
rect 17731 55 17736 75
rect 17851 75 17871 85
rect 17971 75 18001 85
rect 17971 55 17981 75
rect 18096 75 18116 85
rect 18216 75 18241 85
rect 18216 55 18221 75
rect 18336 75 18356 85
rect 18456 75 18486 85
rect 18456 55 18466 75
rect 18581 75 18601 85
rect 18701 75 18726 85
rect 18701 55 18706 75
rect 18821 75 18841 85
rect 18941 75 18971 85
rect 18941 55 18951 75
rect 19066 75 19086 85
rect 19181 75 19211 85
rect 19181 55 19191 75
rect 19306 75 19326 85
rect 19426 75 19456 85
rect 19426 55 19436 75
rect 19551 75 19571 85
rect 19671 75 19696 85
rect 19671 55 19676 75
rect 19791 75 19811 85
rect 19911 75 19941 85
rect 19911 55 19921 75
rect 20036 75 20056 85
rect 20156 75 20181 85
rect 20156 55 20161 75
rect 20276 75 20296 85
rect 20396 75 20426 85
rect 20396 55 20406 75
rect 20521 75 20541 85
rect 20641 75 20666 85
rect 20641 55 20646 75
rect 20761 75 20781 85
rect 20881 75 20911 85
rect 20881 55 20891 75
rect 21006 75 21026 85
rect 5601 15 5641 25
rect 5481 -5 5611 15
rect 5631 -5 5641 15
rect 21066 10 21091 85
rect 21126 75 21146 85
rect 21520 15 21670 165
rect 1666 -70 1686 -65
rect 1786 -50 1806 -45
rect 1901 -65 1911 -50
rect 1901 -70 1931 -65
rect 2031 -50 2051 -45
rect 2146 -65 2151 -50
rect 2146 -70 2171 -65
rect 2271 -50 2291 -45
rect 2386 -65 2396 -50
rect 2386 -70 2416 -65
rect 2516 -50 2536 -45
rect 2631 -65 2636 -50
rect 2631 -70 2656 -65
rect 2756 -50 2776 -45
rect 2871 -65 2881 -50
rect 2871 -70 2901 -65
rect 3001 -50 3021 -45
rect 3116 -65 3121 -50
rect 3116 -70 3141 -65
rect 3241 -50 3261 -45
rect 3356 -65 3366 -50
rect 3356 -70 3386 -65
rect 3486 -50 3506 -45
rect 3596 -65 3606 -50
rect 3596 -70 3626 -65
rect 3726 -50 3746 -45
rect 3841 -65 3851 -50
rect 3841 -70 3871 -65
rect 3971 -50 3991 -45
rect 4086 -65 4091 -50
rect 4086 -70 4111 -65
rect 4211 -50 4231 -45
rect 4326 -65 4336 -50
rect 4326 -70 4356 -65
rect 4456 -50 4476 -45
rect 4571 -65 4576 -50
rect 4571 -70 4596 -65
rect 4696 -50 4716 -45
rect 4811 -65 4821 -50
rect 4811 -70 4841 -65
rect 4941 -50 4961 -45
rect 5056 -65 5061 -50
rect 5056 -70 5081 -65
rect 5181 -50 5201 -45
rect 5296 -65 5306 -50
rect 5296 -70 5326 -65
rect 5426 -50 5446 -45
rect 5481 -70 5506 -5
rect 5601 -15 5641 -5
rect 21065 -10 21160 10
rect 21520 -5 31200 15
rect 5611 -70 5631 -65
rect 5731 -50 5751 -45
rect 5846 -65 5856 -50
rect 5846 -70 5876 -65
rect 5976 -50 5996 -45
rect 6091 -65 6096 -50
rect 6091 -70 6116 -65
rect 6216 -50 6236 -45
rect 6331 -65 6341 -50
rect 6331 -70 6361 -65
rect 6461 -50 6481 -45
rect 6576 -65 6581 -50
rect 6576 -70 6601 -65
rect 6701 -50 6721 -45
rect 6816 -65 6826 -50
rect 6816 -70 6846 -65
rect 6946 -50 6966 -45
rect 7061 -65 7066 -50
rect 7061 -70 7086 -65
rect 7186 -50 7206 -45
rect 7301 -65 7306 -50
rect 7301 -70 7326 -65
rect 7426 -50 7446 -45
rect 7536 -65 7546 -50
rect 7536 -70 7566 -65
rect 7666 -50 7686 -45
rect 7781 -65 7791 -50
rect 7781 -70 7811 -65
rect 7911 -50 7931 -45
rect 8026 -65 8031 -50
rect 8026 -70 8051 -65
rect 8151 -50 8171 -45
rect 8266 -65 8276 -50
rect 8266 -70 8296 -65
rect 8396 -50 8416 -45
rect 8511 -65 8516 -50
rect 8511 -70 8536 -65
rect 8636 -50 8656 -45
rect 8751 -65 8761 -50
rect 8751 -70 8781 -65
rect 8881 -50 8901 -45
rect 8996 -65 9001 -50
rect 8996 -70 9021 -65
rect 9121 -50 9141 -45
rect 9236 -65 9246 -50
rect 9236 -70 9266 -65
rect 9366 -50 9386 -45
rect 9481 -65 9491 -50
rect 9481 -70 9511 -65
rect 9611 -50 9631 -45
rect 9726 -65 9736 -50
rect 9726 -70 9756 -65
rect 9856 -50 9876 -45
rect 9971 -65 9976 -50
rect 9971 -70 9996 -65
rect 10096 -50 10116 -45
rect 10211 -65 10221 -50
rect 10211 -70 10241 -65
rect 10341 -50 10361 -45
rect 10456 -65 10461 -50
rect 10456 -70 10481 -65
rect 10581 -50 10601 -45
rect 10696 -65 10706 -50
rect 10696 -70 10726 -65
rect 10826 -50 10846 -45
rect 10941 -65 10946 -50
rect 10941 -70 10966 -65
rect 11066 -50 11086 -45
rect 11181 -65 11191 -50
rect 11181 -70 11211 -65
rect 11311 -50 11331 -45
rect 11421 -65 11431 -50
rect 11421 -70 11451 -65
rect 11551 -50 11571 -45
rect 11666 -65 11676 -50
rect 11666 -70 11696 -65
rect 11796 -50 11816 -45
rect 11911 -65 11916 -50
rect 11911 -70 11936 -65
rect 12036 -50 12056 -45
rect 12151 -65 12161 -50
rect 12151 -70 12181 -65
rect 12281 -50 12301 -45
rect 12396 -65 12401 -50
rect 12396 -70 12421 -65
rect 12521 -50 12541 -45
rect 12636 -65 12646 -50
rect 12636 -70 12666 -65
rect 12766 -50 12786 -45
rect 12881 -65 12886 -50
rect 12881 -70 12906 -65
rect 13006 -50 13026 -45
rect 13121 -65 13131 -50
rect 13121 -70 13151 -65
rect 13251 -50 13271 -45
rect 13366 -65 13371 -50
rect 13366 -70 13391 -65
rect 13491 -50 13511 -45
rect 13606 -65 13616 -50
rect 13606 -70 13636 -65
rect 13736 -50 13756 -45
rect 13851 -65 13856 -50
rect 13851 -70 13876 -65
rect 13976 -50 13996 -45
rect 14091 -65 14101 -50
rect 14091 -70 14121 -65
rect 14221 -50 14241 -45
rect 14336 -65 14341 -50
rect 14336 -70 14361 -65
rect 14461 -50 14481 -45
rect 14576 -65 14586 -50
rect 14576 -70 14606 -65
rect 14706 -50 14726 -45
rect 14821 -65 14826 -50
rect 14821 -70 14846 -65
rect 14946 -50 14966 -45
rect 15061 -65 15071 -50
rect 15061 -70 15091 -65
rect 15191 -50 15211 -45
rect 15301 -65 15311 -50
rect 15301 -70 15331 -65
rect 15431 -50 15451 -45
rect 15546 -65 15556 -50
rect 15546 -70 15576 -65
rect 15676 -50 15696 -45
rect 15791 -65 15796 -50
rect 15791 -70 15816 -65
rect 15916 -50 15936 -45
rect 16031 -65 16041 -50
rect 16031 -70 16061 -65
rect 16161 -50 16181 -45
rect 16276 -65 16281 -50
rect 16276 -70 16301 -65
rect 16401 -50 16421 -45
rect 16516 -65 16526 -50
rect 16516 -70 16546 -65
rect 16646 -50 16666 -45
rect 16761 -65 16766 -50
rect 16761 -70 16786 -65
rect 16886 -50 16906 -45
rect 17001 -65 17011 -50
rect 17001 -70 17031 -65
rect 17131 -50 17151 -45
rect 17246 -65 17251 -50
rect 17246 -70 17271 -65
rect 17371 -50 17391 -45
rect 17486 -65 17496 -50
rect 17486 -70 17516 -65
rect 17616 -50 17636 -45
rect 17731 -65 17736 -50
rect 17731 -70 17756 -65
rect 17856 -50 17876 -45
rect 17971 -65 17981 -50
rect 17971 -70 18001 -65
rect 18101 -50 18121 -45
rect 18216 -65 18221 -50
rect 18216 -70 18241 -65
rect 18341 -50 18361 -45
rect 18456 -65 18466 -50
rect 18456 -70 18486 -65
rect 18586 -50 18606 -45
rect 18701 -65 18706 -50
rect 18701 -70 18726 -65
rect 18826 -50 18846 -45
rect 18941 -65 18951 -50
rect 18941 -70 18971 -65
rect 19071 -50 19091 -45
rect 19181 -65 19191 -50
rect 19181 -70 19211 -65
rect 19311 -50 19331 -45
rect 19426 -65 19436 -50
rect 19426 -70 19456 -65
rect 19556 -50 19576 -45
rect 19671 -65 19676 -50
rect 19671 -70 19696 -65
rect 19796 -50 19816 -45
rect 19911 -65 19921 -50
rect 19911 -70 19941 -65
rect 20041 -50 20061 -45
rect 20156 -65 20161 -50
rect 20156 -70 20181 -65
rect 20281 -50 20301 -45
rect 20396 -65 20406 -50
rect 20396 -70 20426 -65
rect 20526 -50 20546 -45
rect 20641 -65 20646 -50
rect 20641 -70 20666 -65
rect 20766 -50 20786 -45
rect 20881 -65 20891 -50
rect 20881 -70 20911 -65
rect 21011 -50 21031 -45
rect 21066 -70 21091 -10
rect -460 -190 -320 -105
rect 191 -85 226 -70
rect 191 -110 196 -85
rect 221 -110 226 -85
rect 191 -120 226 -110
rect 251 -85 286 -70
rect 251 -110 256 -85
rect 281 -110 286 -85
rect 251 -120 286 -110
rect 316 -85 351 -70
rect 316 -110 321 -85
rect 346 -110 351 -85
rect 316 -120 351 -110
rect 376 -85 411 -70
rect 376 -110 381 -85
rect 406 -110 411 -85
rect 376 -120 411 -110
rect 436 -85 471 -70
rect 436 -110 441 -85
rect 466 -110 471 -85
rect 436 -120 471 -110
rect 496 -85 531 -70
rect 496 -110 501 -85
rect 526 -110 531 -85
rect 496 -120 531 -110
rect 556 -85 591 -70
rect 556 -110 561 -85
rect 586 -110 591 -85
rect 556 -120 591 -110
rect 621 -85 656 -70
rect 621 -110 626 -85
rect 651 -110 656 -85
rect 621 -120 656 -110
rect 681 -85 716 -70
rect 681 -110 686 -85
rect 711 -110 716 -85
rect 681 -120 716 -110
rect 741 -85 776 -70
rect 741 -110 746 -85
rect 771 -110 776 -85
rect 741 -120 776 -110
rect 801 -85 836 -70
rect 801 -110 806 -85
rect 831 -110 836 -85
rect 801 -120 836 -110
rect 861 -85 901 -70
rect 861 -110 871 -85
rect 896 -110 901 -85
rect 861 -120 901 -110
rect 926 -85 961 -70
rect 926 -110 931 -85
rect 956 -110 961 -85
rect 926 -120 961 -110
rect 986 -85 1021 -70
rect 986 -110 991 -85
rect 1016 -110 1021 -85
rect 986 -120 1021 -110
rect 1046 -85 1081 -70
rect 1046 -110 1051 -85
rect 1076 -110 1081 -85
rect 1046 -120 1081 -110
rect 1106 -85 1141 -70
rect 1106 -110 1111 -85
rect 1136 -110 1141 -85
rect 1106 -120 1141 -110
rect 1166 -85 1201 -70
rect 1166 -110 1171 -85
rect 1196 -110 1201 -85
rect 1166 -120 1201 -110
rect 1226 -85 1261 -70
rect 1226 -110 1231 -85
rect 1256 -110 1261 -85
rect 1226 -120 1261 -110
rect 1286 -85 1321 -70
rect 1286 -110 1291 -85
rect 1316 -110 1321 -85
rect 1286 -120 1321 -110
rect 1346 -85 1386 -70
rect 1346 -110 1356 -85
rect 1381 -110 1386 -85
rect 1346 -120 1386 -110
rect 1411 -85 1446 -70
rect 1411 -110 1416 -85
rect 1441 -110 1446 -85
rect 1411 -120 1446 -110
rect 1471 -85 1506 -70
rect 1471 -110 1476 -85
rect 1501 -110 1506 -85
rect 1471 -120 1506 -110
rect 1531 -85 1566 -70
rect 1531 -110 1536 -85
rect 1561 -110 1566 -85
rect 1531 -120 1566 -110
rect 1591 -85 1626 -70
rect 1591 -110 1596 -85
rect 1621 -110 1626 -85
rect 1591 -120 1626 -110
rect 1656 -85 1691 -70
rect 1656 -110 1661 -85
rect 1686 -110 1691 -85
rect 1656 -120 1691 -110
rect 1716 -85 1751 -70
rect 1716 -110 1721 -85
rect 1746 -110 1751 -85
rect 1716 -120 1751 -110
rect 1776 -85 1811 -70
rect 1776 -110 1781 -85
rect 1806 -110 1811 -85
rect 1776 -120 1811 -110
rect 1836 -85 1871 -70
rect 1836 -110 1841 -85
rect 1866 -110 1871 -85
rect 1836 -120 1871 -110
rect 1896 -85 1936 -70
rect 1896 -110 1906 -85
rect 1931 -110 1936 -85
rect 1896 -120 1936 -110
rect 1961 -85 1996 -70
rect 1961 -110 1966 -85
rect 1991 -110 1996 -85
rect 1961 -120 1996 -110
rect 2021 -85 2056 -70
rect 2021 -110 2026 -85
rect 2051 -110 2056 -85
rect 2021 -120 2056 -110
rect 2081 -85 2116 -70
rect 2081 -110 2086 -85
rect 2111 -110 2116 -85
rect 2081 -120 2116 -110
rect 2141 -85 2176 -70
rect 2141 -110 2146 -85
rect 2171 -110 2176 -85
rect 2141 -120 2176 -110
rect 2201 -85 2236 -70
rect 2201 -110 2206 -85
rect 2231 -110 2236 -85
rect 2201 -120 2236 -110
rect 2261 -85 2296 -70
rect 2261 -110 2266 -85
rect 2291 -110 2296 -85
rect 2261 -120 2296 -110
rect 2321 -85 2356 -70
rect 2321 -110 2326 -85
rect 2351 -110 2356 -85
rect 2321 -120 2356 -110
rect 2381 -85 2421 -70
rect 2381 -110 2391 -85
rect 2416 -110 2421 -85
rect 2381 -120 2421 -110
rect 2446 -85 2481 -70
rect 2446 -110 2451 -85
rect 2476 -110 2481 -85
rect 2446 -120 2481 -110
rect 2506 -85 2541 -70
rect 2506 -110 2511 -85
rect 2536 -110 2541 -85
rect 2506 -120 2541 -110
rect 2566 -85 2601 -70
rect 2566 -110 2571 -85
rect 2596 -110 2601 -85
rect 2566 -120 2601 -110
rect 2626 -85 2661 -70
rect 2626 -110 2631 -85
rect 2656 -110 2661 -85
rect 2626 -120 2661 -110
rect 2686 -85 2721 -70
rect 2686 -110 2691 -85
rect 2716 -110 2721 -85
rect 2686 -120 2721 -110
rect 2746 -85 2781 -70
rect 2746 -110 2751 -85
rect 2776 -110 2781 -85
rect 2746 -120 2781 -110
rect 2806 -85 2841 -70
rect 2806 -110 2811 -85
rect 2836 -110 2841 -85
rect 2806 -120 2841 -110
rect 2866 -85 2906 -70
rect 2866 -110 2876 -85
rect 2901 -110 2906 -85
rect 2866 -120 2906 -110
rect 2931 -85 2966 -70
rect 2931 -110 2936 -85
rect 2961 -110 2966 -85
rect 2931 -120 2966 -110
rect 2991 -85 3026 -70
rect 2991 -110 2996 -85
rect 3021 -110 3026 -85
rect 2991 -120 3026 -110
rect 3051 -85 3086 -70
rect 3051 -110 3056 -85
rect 3081 -110 3086 -85
rect 3051 -120 3086 -110
rect 3111 -85 3146 -70
rect 3111 -110 3116 -85
rect 3141 -110 3146 -85
rect 3111 -120 3146 -110
rect 3171 -85 3206 -70
rect 3171 -110 3176 -85
rect 3201 -110 3206 -85
rect 3171 -120 3206 -110
rect 3231 -85 3266 -70
rect 3231 -110 3236 -85
rect 3261 -110 3266 -85
rect 3231 -120 3266 -110
rect 3291 -85 3326 -70
rect 3291 -110 3296 -85
rect 3321 -110 3326 -85
rect 3291 -120 3326 -110
rect 3351 -85 3391 -70
rect 3351 -110 3361 -85
rect 3386 -110 3391 -85
rect 3351 -120 3391 -110
rect 3416 -85 3451 -70
rect 3416 -110 3421 -85
rect 3446 -110 3451 -85
rect 3416 -120 3451 -110
rect 3476 -85 3511 -70
rect 3476 -110 3481 -85
rect 3506 -110 3511 -85
rect 3476 -120 3511 -110
rect 3536 -85 3571 -70
rect 3536 -110 3541 -85
rect 3566 -110 3571 -85
rect 3536 -120 3571 -110
rect 3596 -85 3631 -70
rect 3596 -110 3601 -85
rect 3626 -110 3631 -85
rect 3596 -120 3631 -110
rect 3656 -85 3691 -70
rect 3656 -110 3661 -85
rect 3686 -110 3691 -85
rect 3656 -120 3691 -110
rect 3716 -85 3751 -70
rect 3716 -110 3721 -85
rect 3746 -110 3751 -85
rect 3716 -120 3751 -110
rect 3776 -85 3811 -70
rect 3776 -110 3781 -85
rect 3806 -110 3811 -85
rect 3776 -120 3811 -110
rect 3836 -85 3876 -70
rect 3836 -110 3846 -85
rect 3871 -110 3876 -85
rect 3836 -120 3876 -110
rect 3901 -85 3936 -70
rect 3901 -110 3906 -85
rect 3931 -110 3936 -85
rect 3901 -120 3936 -110
rect 3961 -85 3996 -70
rect 3961 -110 3966 -85
rect 3991 -110 3996 -85
rect 3961 -120 3996 -110
rect 4021 -85 4056 -70
rect 4021 -110 4026 -85
rect 4051 -110 4056 -85
rect 4021 -120 4056 -110
rect 4081 -85 4116 -70
rect 4081 -110 4086 -85
rect 4111 -110 4116 -85
rect 4081 -120 4116 -110
rect 4141 -85 4176 -70
rect 4141 -110 4146 -85
rect 4171 -110 4176 -85
rect 4141 -120 4176 -110
rect 4201 -85 4236 -70
rect 4201 -110 4206 -85
rect 4231 -110 4236 -85
rect 4201 -120 4236 -110
rect 4261 -85 4296 -70
rect 4261 -110 4266 -85
rect 4291 -110 4296 -85
rect 4261 -120 4296 -110
rect 4321 -85 4361 -70
rect 4321 -110 4331 -85
rect 4356 -110 4361 -85
rect 4321 -120 4361 -110
rect 4386 -85 4421 -70
rect 4386 -110 4391 -85
rect 4416 -110 4421 -85
rect 4386 -120 4421 -110
rect 4446 -85 4481 -70
rect 4446 -110 4451 -85
rect 4476 -110 4481 -85
rect 4446 -120 4481 -110
rect 4506 -85 4541 -70
rect 4506 -110 4511 -85
rect 4536 -110 4541 -85
rect 4506 -120 4541 -110
rect 4566 -85 4601 -70
rect 4566 -110 4571 -85
rect 4596 -110 4601 -85
rect 4566 -120 4601 -110
rect 4626 -85 4661 -70
rect 4626 -110 4631 -85
rect 4656 -110 4661 -85
rect 4626 -120 4661 -110
rect 4686 -85 4721 -70
rect 4686 -110 4691 -85
rect 4716 -110 4721 -85
rect 4686 -120 4721 -110
rect 4746 -85 4781 -70
rect 4746 -110 4751 -85
rect 4776 -110 4781 -85
rect 4746 -120 4781 -110
rect 4806 -85 4846 -70
rect 4806 -110 4816 -85
rect 4841 -110 4846 -85
rect 4806 -120 4846 -110
rect 4871 -85 4906 -70
rect 4871 -110 4876 -85
rect 4901 -110 4906 -85
rect 4871 -120 4906 -110
rect 4931 -85 4966 -70
rect 4931 -110 4936 -85
rect 4961 -110 4966 -85
rect 4931 -120 4966 -110
rect 4991 -85 5026 -70
rect 4991 -110 4996 -85
rect 5021 -110 5026 -85
rect 4991 -120 5026 -110
rect 5051 -85 5086 -70
rect 5051 -110 5056 -85
rect 5081 -110 5086 -85
rect 5051 -120 5086 -110
rect 5111 -85 5146 -70
rect 5111 -110 5116 -85
rect 5141 -110 5146 -85
rect 5111 -120 5146 -110
rect 5171 -85 5206 -70
rect 5171 -110 5176 -85
rect 5201 -110 5206 -85
rect 5171 -120 5206 -110
rect 5231 -85 5266 -70
rect 5231 -110 5236 -85
rect 5261 -110 5266 -85
rect 5231 -120 5266 -110
rect 5291 -85 5331 -70
rect 5291 -110 5301 -85
rect 5326 -110 5331 -85
rect 5291 -120 5331 -110
rect 5356 -85 5391 -70
rect 5356 -110 5361 -85
rect 5386 -110 5391 -85
rect 5356 -120 5391 -110
rect 5416 -85 5451 -70
rect 5416 -110 5421 -85
rect 5446 -110 5451 -85
rect 5416 -120 5451 -110
rect 5476 -85 5511 -70
rect 5476 -110 5481 -85
rect 5506 -110 5511 -85
rect 5476 -120 5511 -110
rect 5536 -85 5571 -70
rect 5536 -110 5541 -85
rect 5566 -110 5571 -85
rect 5536 -120 5571 -110
rect 5601 -85 5636 -70
rect 5601 -110 5606 -85
rect 5631 -110 5636 -85
rect 5601 -120 5636 -110
rect 5661 -85 5696 -70
rect 5661 -110 5666 -85
rect 5691 -110 5696 -85
rect 5661 -120 5696 -110
rect 5721 -85 5756 -70
rect 5721 -110 5726 -85
rect 5751 -110 5756 -85
rect 5721 -120 5756 -110
rect 5781 -85 5816 -70
rect 5781 -110 5786 -85
rect 5811 -110 5816 -85
rect 5781 -120 5816 -110
rect 5841 -85 5881 -70
rect 5841 -110 5851 -85
rect 5876 -110 5881 -85
rect 5841 -120 5881 -110
rect 5906 -85 5941 -70
rect 5906 -110 5911 -85
rect 5936 -110 5941 -85
rect 5906 -120 5941 -110
rect 5966 -85 6001 -70
rect 5966 -110 5971 -85
rect 5996 -110 6001 -85
rect 5966 -120 6001 -110
rect 6026 -85 6061 -70
rect 6026 -110 6031 -85
rect 6056 -110 6061 -85
rect 6026 -120 6061 -110
rect 6086 -85 6121 -70
rect 6086 -110 6091 -85
rect 6116 -110 6121 -85
rect 6086 -120 6121 -110
rect 6146 -85 6181 -70
rect 6146 -110 6151 -85
rect 6176 -110 6181 -85
rect 6146 -120 6181 -110
rect 6206 -85 6241 -70
rect 6206 -110 6211 -85
rect 6236 -110 6241 -85
rect 6206 -120 6241 -110
rect 6266 -85 6301 -70
rect 6266 -110 6271 -85
rect 6296 -110 6301 -85
rect 6266 -120 6301 -110
rect 6326 -85 6366 -70
rect 6326 -110 6336 -85
rect 6361 -110 6366 -85
rect 6326 -120 6366 -110
rect 6391 -85 6426 -70
rect 6391 -110 6396 -85
rect 6421 -110 6426 -85
rect 6391 -120 6426 -110
rect 6451 -85 6486 -70
rect 6451 -110 6456 -85
rect 6481 -110 6486 -85
rect 6451 -120 6486 -110
rect 6511 -85 6546 -70
rect 6511 -110 6516 -85
rect 6541 -110 6546 -85
rect 6511 -120 6546 -110
rect 6571 -85 6606 -70
rect 6571 -110 6576 -85
rect 6601 -110 6606 -85
rect 6571 -120 6606 -110
rect 6631 -85 6666 -70
rect 6631 -110 6636 -85
rect 6661 -110 6666 -85
rect 6631 -120 6666 -110
rect 6691 -85 6726 -70
rect 6691 -110 6696 -85
rect 6721 -110 6726 -85
rect 6691 -120 6726 -110
rect 6751 -85 6786 -70
rect 6751 -110 6756 -85
rect 6781 -110 6786 -85
rect 6751 -120 6786 -110
rect 6811 -85 6851 -70
rect 6811 -110 6821 -85
rect 6846 -110 6851 -85
rect 6811 -120 6851 -110
rect 6876 -85 6911 -70
rect 6876 -110 6881 -85
rect 6906 -110 6911 -85
rect 6876 -120 6911 -110
rect 6936 -85 6971 -70
rect 6936 -110 6941 -85
rect 6966 -110 6971 -85
rect 6936 -120 6971 -110
rect 6996 -85 7031 -70
rect 6996 -110 7001 -85
rect 7026 -110 7031 -85
rect 6996 -120 7031 -110
rect 7056 -85 7091 -70
rect 7056 -110 7061 -85
rect 7086 -110 7091 -85
rect 7056 -120 7091 -110
rect 7116 -85 7151 -70
rect 7116 -110 7121 -85
rect 7146 -110 7151 -85
rect 7116 -120 7151 -110
rect 7176 -85 7211 -70
rect 7176 -110 7181 -85
rect 7206 -110 7211 -85
rect 7176 -120 7211 -110
rect 7236 -85 7271 -70
rect 7236 -110 7241 -85
rect 7266 -110 7271 -85
rect 7236 -120 7271 -110
rect 7296 -85 7331 -70
rect 7296 -110 7301 -85
rect 7326 -110 7331 -85
rect 7296 -120 7331 -110
rect 7356 -85 7391 -70
rect 7356 -110 7361 -85
rect 7386 -110 7391 -85
rect 7356 -120 7391 -110
rect 7416 -85 7451 -70
rect 7416 -110 7421 -85
rect 7446 -110 7451 -85
rect 7416 -120 7451 -110
rect 7476 -85 7511 -70
rect 7476 -110 7481 -85
rect 7506 -110 7511 -85
rect 7476 -120 7511 -110
rect 7536 -85 7571 -70
rect 7536 -110 7541 -85
rect 7566 -110 7571 -85
rect 7536 -120 7571 -110
rect 7596 -85 7631 -70
rect 7596 -110 7601 -85
rect 7626 -110 7631 -85
rect 7596 -120 7631 -110
rect 7656 -85 7691 -70
rect 7656 -110 7661 -85
rect 7686 -110 7691 -85
rect 7656 -120 7691 -110
rect 7716 -85 7751 -70
rect 7716 -110 7721 -85
rect 7746 -110 7751 -85
rect 7716 -120 7751 -110
rect 7776 -85 7816 -70
rect 7776 -110 7786 -85
rect 7811 -110 7816 -85
rect 7776 -120 7816 -110
rect 7841 -85 7876 -70
rect 7841 -110 7846 -85
rect 7871 -110 7876 -85
rect 7841 -120 7876 -110
rect 7901 -85 7936 -70
rect 7901 -110 7906 -85
rect 7931 -110 7936 -85
rect 7901 -120 7936 -110
rect 7961 -85 7996 -70
rect 7961 -110 7966 -85
rect 7991 -110 7996 -85
rect 7961 -120 7996 -110
rect 8021 -85 8056 -70
rect 8021 -110 8026 -85
rect 8051 -110 8056 -85
rect 8021 -120 8056 -110
rect 8081 -85 8116 -70
rect 8081 -110 8086 -85
rect 8111 -110 8116 -85
rect 8081 -120 8116 -110
rect 8141 -85 8176 -70
rect 8141 -110 8146 -85
rect 8171 -110 8176 -85
rect 8141 -120 8176 -110
rect 8201 -85 8236 -70
rect 8201 -110 8206 -85
rect 8231 -110 8236 -85
rect 8201 -120 8236 -110
rect 8261 -85 8301 -70
rect 8261 -110 8271 -85
rect 8296 -110 8301 -85
rect 8261 -120 8301 -110
rect 8326 -85 8361 -70
rect 8326 -110 8331 -85
rect 8356 -110 8361 -85
rect 8326 -120 8361 -110
rect 8386 -85 8421 -70
rect 8386 -110 8391 -85
rect 8416 -110 8421 -85
rect 8386 -120 8421 -110
rect 8446 -85 8481 -70
rect 8446 -110 8451 -85
rect 8476 -110 8481 -85
rect 8446 -120 8481 -110
rect 8506 -85 8541 -70
rect 8506 -110 8511 -85
rect 8536 -110 8541 -85
rect 8506 -120 8541 -110
rect 8566 -85 8601 -70
rect 8566 -110 8571 -85
rect 8596 -110 8601 -85
rect 8566 -120 8601 -110
rect 8626 -85 8661 -70
rect 8626 -110 8631 -85
rect 8656 -110 8661 -85
rect 8626 -120 8661 -110
rect 8686 -85 8721 -70
rect 8686 -110 8691 -85
rect 8716 -110 8721 -85
rect 8686 -120 8721 -110
rect 8746 -85 8786 -70
rect 8746 -110 8756 -85
rect 8781 -110 8786 -85
rect 8746 -120 8786 -110
rect 8811 -85 8846 -70
rect 8811 -110 8816 -85
rect 8841 -110 8846 -85
rect 8811 -120 8846 -110
rect 8871 -85 8906 -70
rect 8871 -110 8876 -85
rect 8901 -110 8906 -85
rect 8871 -120 8906 -110
rect 8931 -85 8966 -70
rect 8931 -110 8936 -85
rect 8961 -110 8966 -85
rect 8931 -120 8966 -110
rect 8991 -85 9026 -70
rect 8991 -110 8996 -85
rect 9021 -110 9026 -85
rect 8991 -120 9026 -110
rect 9051 -85 9086 -70
rect 9051 -110 9056 -85
rect 9081 -110 9086 -85
rect 9051 -120 9086 -110
rect 9111 -85 9146 -70
rect 9111 -110 9116 -85
rect 9141 -110 9146 -85
rect 9111 -120 9146 -110
rect 9171 -85 9206 -70
rect 9171 -110 9176 -85
rect 9201 -110 9206 -85
rect 9171 -120 9206 -110
rect 9231 -85 9271 -70
rect 9231 -110 9241 -85
rect 9266 -110 9271 -85
rect 9231 -120 9271 -110
rect 9296 -85 9331 -70
rect 9296 -110 9301 -85
rect 9326 -110 9331 -85
rect 9296 -120 9331 -110
rect 9356 -85 9391 -70
rect 9356 -110 9361 -85
rect 9386 -110 9391 -85
rect 9356 -120 9391 -110
rect 9416 -85 9451 -70
rect 9416 -110 9421 -85
rect 9446 -110 9451 -85
rect 9416 -120 9451 -110
rect 9476 -85 9516 -70
rect 9476 -110 9486 -85
rect 9511 -110 9516 -85
rect 9476 -120 9516 -110
rect 9541 -85 9576 -70
rect 9541 -110 9546 -85
rect 9571 -110 9576 -85
rect 9541 -120 9576 -110
rect 9601 -85 9636 -70
rect 9601 -110 9606 -85
rect 9631 -110 9636 -85
rect 9601 -120 9636 -110
rect 9661 -85 9696 -70
rect 9661 -110 9666 -85
rect 9691 -110 9696 -85
rect 9661 -120 9696 -110
rect 9721 -85 9761 -70
rect 9721 -110 9731 -85
rect 9756 -110 9761 -85
rect 9721 -120 9761 -110
rect 9786 -85 9821 -70
rect 9786 -110 9791 -85
rect 9816 -110 9821 -85
rect 9786 -120 9821 -110
rect 9846 -85 9881 -70
rect 9846 -110 9851 -85
rect 9876 -110 9881 -85
rect 9846 -120 9881 -110
rect 9906 -85 9941 -70
rect 9906 -110 9911 -85
rect 9936 -110 9941 -85
rect 9906 -120 9941 -110
rect 9966 -85 10001 -70
rect 9966 -110 9971 -85
rect 9996 -110 10001 -85
rect 9966 -120 10001 -110
rect 10026 -85 10061 -70
rect 10026 -110 10031 -85
rect 10056 -110 10061 -85
rect 10026 -120 10061 -110
rect 10086 -85 10121 -70
rect 10086 -110 10091 -85
rect 10116 -110 10121 -85
rect 10086 -120 10121 -110
rect 10146 -85 10181 -70
rect 10146 -110 10151 -85
rect 10176 -110 10181 -85
rect 10146 -120 10181 -110
rect 10206 -85 10246 -70
rect 10206 -110 10216 -85
rect 10241 -110 10246 -85
rect 10206 -120 10246 -110
rect 10271 -85 10306 -70
rect 10271 -110 10276 -85
rect 10301 -110 10306 -85
rect 10271 -120 10306 -110
rect 10331 -85 10366 -70
rect 10331 -110 10336 -85
rect 10361 -110 10366 -85
rect 10331 -120 10366 -110
rect 10391 -85 10426 -70
rect 10391 -110 10396 -85
rect 10421 -110 10426 -85
rect 10391 -120 10426 -110
rect 10451 -85 10486 -70
rect 10451 -110 10456 -85
rect 10481 -110 10486 -85
rect 10451 -120 10486 -110
rect 10511 -85 10546 -70
rect 10511 -110 10516 -85
rect 10541 -110 10546 -85
rect 10511 -120 10546 -110
rect 10571 -85 10606 -70
rect 10571 -110 10576 -85
rect 10601 -110 10606 -85
rect 10571 -120 10606 -110
rect 10631 -85 10666 -70
rect 10631 -110 10636 -85
rect 10661 -110 10666 -85
rect 10631 -120 10666 -110
rect 10691 -85 10731 -70
rect 10691 -110 10701 -85
rect 10726 -110 10731 -85
rect 10691 -120 10731 -110
rect 10756 -85 10791 -70
rect 10756 -110 10761 -85
rect 10786 -110 10791 -85
rect 10756 -120 10791 -110
rect 10816 -85 10851 -70
rect 10816 -110 10821 -85
rect 10846 -110 10851 -85
rect 10816 -120 10851 -110
rect 10876 -85 10911 -70
rect 10876 -110 10881 -85
rect 10906 -110 10911 -85
rect 10876 -120 10911 -110
rect 10936 -85 10971 -70
rect 10936 -110 10941 -85
rect 10966 -110 10971 -85
rect 10936 -120 10971 -110
rect 10996 -85 11031 -70
rect 10996 -110 11001 -85
rect 11026 -110 11031 -85
rect 10996 -120 11031 -110
rect 11056 -85 11091 -70
rect 11056 -110 11061 -85
rect 11086 -110 11091 -85
rect 11056 -120 11091 -110
rect 11116 -85 11151 -70
rect 11116 -110 11121 -85
rect 11146 -110 11151 -85
rect 11116 -120 11151 -110
rect 11176 -85 11216 -70
rect 11176 -110 11186 -85
rect 11211 -110 11216 -85
rect 11176 -120 11216 -110
rect 11241 -85 11276 -70
rect 11241 -110 11246 -85
rect 11271 -110 11276 -85
rect 11241 -120 11276 -110
rect 11301 -85 11336 -70
rect 11301 -110 11306 -85
rect 11331 -110 11336 -85
rect 11301 -120 11336 -110
rect 11361 -85 11396 -70
rect 11361 -110 11366 -85
rect 11391 -110 11396 -85
rect 11361 -120 11396 -110
rect 11421 -85 11456 -70
rect 11421 -110 11426 -85
rect 11451 -110 11456 -85
rect 11421 -120 11456 -110
rect 11481 -85 11516 -70
rect 11481 -110 11486 -85
rect 11511 -110 11516 -85
rect 11481 -120 11516 -110
rect 11541 -85 11576 -70
rect 11541 -110 11546 -85
rect 11571 -110 11576 -85
rect 11541 -120 11576 -110
rect 11601 -85 11636 -70
rect 11601 -110 11606 -85
rect 11631 -110 11636 -85
rect 11601 -120 11636 -110
rect 11661 -85 11701 -70
rect 11661 -110 11671 -85
rect 11696 -110 11701 -85
rect 11661 -120 11701 -110
rect 11726 -85 11761 -70
rect 11726 -110 11731 -85
rect 11756 -110 11761 -85
rect 11726 -120 11761 -110
rect 11786 -85 11821 -70
rect 11786 -110 11791 -85
rect 11816 -110 11821 -85
rect 11786 -120 11821 -110
rect 11846 -85 11881 -70
rect 11846 -110 11851 -85
rect 11876 -110 11881 -85
rect 11846 -120 11881 -110
rect 11906 -85 11941 -70
rect 11906 -110 11911 -85
rect 11936 -110 11941 -85
rect 11906 -120 11941 -110
rect 11966 -85 12001 -70
rect 11966 -110 11971 -85
rect 11996 -110 12001 -85
rect 11966 -120 12001 -110
rect 12026 -85 12061 -70
rect 12026 -110 12031 -85
rect 12056 -110 12061 -85
rect 12026 -120 12061 -110
rect 12086 -85 12121 -70
rect 12086 -110 12091 -85
rect 12116 -110 12121 -85
rect 12086 -120 12121 -110
rect 12146 -85 12186 -70
rect 12146 -110 12156 -85
rect 12181 -110 12186 -85
rect 12146 -120 12186 -110
rect 12211 -85 12246 -70
rect 12211 -110 12216 -85
rect 12241 -110 12246 -85
rect 12211 -120 12246 -110
rect 12271 -85 12306 -70
rect 12271 -110 12276 -85
rect 12301 -110 12306 -85
rect 12271 -120 12306 -110
rect 12331 -85 12366 -70
rect 12331 -110 12336 -85
rect 12361 -110 12366 -85
rect 12331 -120 12366 -110
rect 12391 -85 12426 -70
rect 12391 -110 12396 -85
rect 12421 -110 12426 -85
rect 12391 -120 12426 -110
rect 12451 -85 12486 -70
rect 12451 -110 12456 -85
rect 12481 -110 12486 -85
rect 12451 -120 12486 -110
rect 12511 -85 12546 -70
rect 12511 -110 12516 -85
rect 12541 -110 12546 -85
rect 12511 -120 12546 -110
rect 12571 -85 12606 -70
rect 12571 -110 12576 -85
rect 12601 -110 12606 -85
rect 12571 -120 12606 -110
rect 12631 -85 12671 -70
rect 12631 -110 12641 -85
rect 12666 -110 12671 -85
rect 12631 -120 12671 -110
rect 12696 -85 12731 -70
rect 12696 -110 12701 -85
rect 12726 -110 12731 -85
rect 12696 -120 12731 -110
rect 12756 -85 12791 -70
rect 12756 -110 12761 -85
rect 12786 -110 12791 -85
rect 12756 -120 12791 -110
rect 12816 -85 12851 -70
rect 12816 -110 12821 -85
rect 12846 -110 12851 -85
rect 12816 -120 12851 -110
rect 12876 -85 12911 -70
rect 12876 -110 12881 -85
rect 12906 -110 12911 -85
rect 12876 -120 12911 -110
rect 12936 -85 12971 -70
rect 12936 -110 12941 -85
rect 12966 -110 12971 -85
rect 12936 -120 12971 -110
rect 12996 -85 13031 -70
rect 12996 -110 13001 -85
rect 13026 -110 13031 -85
rect 12996 -120 13031 -110
rect 13056 -85 13091 -70
rect 13056 -110 13061 -85
rect 13086 -110 13091 -85
rect 13056 -120 13091 -110
rect 13116 -85 13156 -70
rect 13116 -110 13126 -85
rect 13151 -110 13156 -85
rect 13116 -120 13156 -110
rect 13181 -85 13216 -70
rect 13181 -110 13186 -85
rect 13211 -110 13216 -85
rect 13181 -120 13216 -110
rect 13241 -85 13276 -70
rect 13241 -110 13246 -85
rect 13271 -110 13276 -85
rect 13241 -120 13276 -110
rect 13301 -85 13336 -70
rect 13301 -110 13306 -85
rect 13331 -110 13336 -85
rect 13301 -120 13336 -110
rect 13361 -85 13396 -70
rect 13361 -110 13366 -85
rect 13391 -110 13396 -85
rect 13361 -120 13396 -110
rect 13421 -85 13456 -70
rect 13421 -110 13426 -85
rect 13451 -110 13456 -85
rect 13421 -120 13456 -110
rect 13481 -85 13516 -70
rect 13481 -110 13486 -85
rect 13511 -110 13516 -85
rect 13481 -120 13516 -110
rect 13541 -85 13576 -70
rect 13541 -110 13546 -85
rect 13571 -110 13576 -85
rect 13541 -120 13576 -110
rect 13601 -85 13641 -70
rect 13601 -110 13611 -85
rect 13636 -110 13641 -85
rect 13601 -120 13641 -110
rect 13666 -85 13701 -70
rect 13666 -110 13671 -85
rect 13696 -110 13701 -85
rect 13666 -120 13701 -110
rect 13726 -85 13761 -70
rect 13726 -110 13731 -85
rect 13756 -110 13761 -85
rect 13726 -120 13761 -110
rect 13786 -85 13821 -70
rect 13786 -110 13791 -85
rect 13816 -110 13821 -85
rect 13786 -120 13821 -110
rect 13846 -85 13881 -70
rect 13846 -110 13851 -85
rect 13876 -110 13881 -85
rect 13846 -120 13881 -110
rect 13906 -85 13941 -70
rect 13906 -110 13911 -85
rect 13936 -110 13941 -85
rect 13906 -120 13941 -110
rect 13966 -85 14001 -70
rect 13966 -110 13971 -85
rect 13996 -110 14001 -85
rect 13966 -120 14001 -110
rect 14026 -85 14061 -70
rect 14026 -110 14031 -85
rect 14056 -110 14061 -85
rect 14026 -120 14061 -110
rect 14086 -85 14126 -70
rect 14086 -110 14096 -85
rect 14121 -110 14126 -85
rect 14086 -120 14126 -110
rect 14151 -85 14186 -70
rect 14151 -110 14156 -85
rect 14181 -110 14186 -85
rect 14151 -120 14186 -110
rect 14211 -85 14246 -70
rect 14211 -110 14216 -85
rect 14241 -110 14246 -85
rect 14211 -120 14246 -110
rect 14271 -85 14306 -70
rect 14271 -110 14276 -85
rect 14301 -110 14306 -85
rect 14271 -120 14306 -110
rect 14331 -85 14366 -70
rect 14331 -110 14336 -85
rect 14361 -110 14366 -85
rect 14331 -120 14366 -110
rect 14391 -85 14426 -70
rect 14391 -110 14396 -85
rect 14421 -110 14426 -85
rect 14391 -120 14426 -110
rect 14451 -85 14486 -70
rect 14451 -110 14456 -85
rect 14481 -110 14486 -85
rect 14451 -120 14486 -110
rect 14511 -85 14546 -70
rect 14511 -110 14516 -85
rect 14541 -110 14546 -85
rect 14511 -120 14546 -110
rect 14571 -85 14611 -70
rect 14571 -110 14581 -85
rect 14606 -110 14611 -85
rect 14571 -120 14611 -110
rect 14636 -85 14671 -70
rect 14636 -110 14641 -85
rect 14666 -110 14671 -85
rect 14636 -120 14671 -110
rect 14696 -85 14731 -70
rect 14696 -110 14701 -85
rect 14726 -110 14731 -85
rect 14696 -120 14731 -110
rect 14756 -85 14791 -70
rect 14756 -110 14761 -85
rect 14786 -110 14791 -85
rect 14756 -120 14791 -110
rect 14816 -85 14851 -70
rect 14816 -110 14821 -85
rect 14846 -110 14851 -85
rect 14816 -120 14851 -110
rect 14876 -85 14911 -70
rect 14876 -110 14881 -85
rect 14906 -110 14911 -85
rect 14876 -120 14911 -110
rect 14936 -85 14971 -70
rect 14936 -110 14941 -85
rect 14966 -110 14971 -85
rect 14936 -120 14971 -110
rect 14996 -85 15031 -70
rect 14996 -110 15001 -85
rect 15026 -110 15031 -85
rect 14996 -120 15031 -110
rect 15056 -85 15096 -70
rect 15056 -110 15066 -85
rect 15091 -110 15096 -85
rect 15056 -120 15096 -110
rect 15121 -85 15156 -70
rect 15121 -110 15126 -85
rect 15151 -110 15156 -85
rect 15121 -120 15156 -110
rect 15181 -85 15216 -70
rect 15181 -110 15186 -85
rect 15211 -110 15216 -85
rect 15181 -120 15216 -110
rect 15241 -85 15276 -70
rect 15241 -110 15246 -85
rect 15271 -110 15276 -85
rect 15241 -120 15276 -110
rect 15301 -85 15336 -70
rect 15301 -110 15306 -85
rect 15331 -110 15336 -85
rect 15301 -120 15336 -110
rect 15361 -85 15396 -70
rect 15361 -110 15366 -85
rect 15391 -110 15396 -85
rect 15361 -120 15396 -110
rect 15421 -85 15456 -70
rect 15421 -110 15426 -85
rect 15451 -110 15456 -85
rect 15421 -120 15456 -110
rect 15481 -85 15516 -70
rect 15481 -110 15486 -85
rect 15511 -110 15516 -85
rect 15481 -120 15516 -110
rect 15541 -85 15581 -70
rect 15541 -110 15551 -85
rect 15576 -110 15581 -85
rect 15541 -120 15581 -110
rect 15606 -85 15641 -70
rect 15606 -110 15611 -85
rect 15636 -110 15641 -85
rect 15606 -120 15641 -110
rect 15666 -85 15701 -70
rect 15666 -110 15671 -85
rect 15696 -110 15701 -85
rect 15666 -120 15701 -110
rect 15726 -85 15761 -70
rect 15726 -110 15731 -85
rect 15756 -110 15761 -85
rect 15726 -120 15761 -110
rect 15786 -85 15821 -70
rect 15786 -110 15791 -85
rect 15816 -110 15821 -85
rect 15786 -120 15821 -110
rect 15846 -85 15881 -70
rect 15846 -110 15851 -85
rect 15876 -110 15881 -85
rect 15846 -120 15881 -110
rect 15906 -85 15941 -70
rect 15906 -110 15911 -85
rect 15936 -110 15941 -85
rect 15906 -120 15941 -110
rect 15966 -85 16001 -70
rect 15966 -110 15971 -85
rect 15996 -110 16001 -85
rect 15966 -120 16001 -110
rect 16026 -85 16066 -70
rect 16026 -110 16036 -85
rect 16061 -110 16066 -85
rect 16026 -120 16066 -110
rect 16091 -85 16126 -70
rect 16091 -110 16096 -85
rect 16121 -110 16126 -85
rect 16091 -120 16126 -110
rect 16151 -85 16186 -70
rect 16151 -110 16156 -85
rect 16181 -110 16186 -85
rect 16151 -120 16186 -110
rect 16211 -85 16246 -70
rect 16211 -110 16216 -85
rect 16241 -110 16246 -85
rect 16211 -120 16246 -110
rect 16271 -85 16306 -70
rect 16271 -110 16276 -85
rect 16301 -110 16306 -85
rect 16271 -120 16306 -110
rect 16331 -85 16366 -70
rect 16331 -110 16336 -85
rect 16361 -110 16366 -85
rect 16331 -120 16366 -110
rect 16391 -85 16426 -70
rect 16391 -110 16396 -85
rect 16421 -110 16426 -85
rect 16391 -120 16426 -110
rect 16451 -85 16486 -70
rect 16451 -110 16456 -85
rect 16481 -110 16486 -85
rect 16451 -120 16486 -110
rect 16511 -85 16551 -70
rect 16511 -110 16521 -85
rect 16546 -110 16551 -85
rect 16511 -120 16551 -110
rect 16576 -85 16611 -70
rect 16576 -110 16581 -85
rect 16606 -110 16611 -85
rect 16576 -120 16611 -110
rect 16636 -85 16671 -70
rect 16636 -110 16641 -85
rect 16666 -110 16671 -85
rect 16636 -120 16671 -110
rect 16696 -85 16731 -70
rect 16696 -110 16701 -85
rect 16726 -110 16731 -85
rect 16696 -120 16731 -110
rect 16756 -85 16791 -70
rect 16756 -110 16761 -85
rect 16786 -110 16791 -85
rect 16756 -120 16791 -110
rect 16816 -85 16851 -70
rect 16816 -110 16821 -85
rect 16846 -110 16851 -85
rect 16816 -120 16851 -110
rect 16876 -85 16911 -70
rect 16876 -110 16881 -85
rect 16906 -110 16911 -85
rect 16876 -120 16911 -110
rect 16936 -85 16971 -70
rect 16936 -110 16941 -85
rect 16966 -110 16971 -85
rect 16936 -120 16971 -110
rect 16996 -85 17036 -70
rect 16996 -110 17006 -85
rect 17031 -110 17036 -85
rect 16996 -120 17036 -110
rect 17061 -85 17096 -70
rect 17061 -110 17066 -85
rect 17091 -110 17096 -85
rect 17061 -120 17096 -110
rect 17121 -85 17156 -70
rect 17121 -110 17126 -85
rect 17151 -110 17156 -85
rect 17121 -120 17156 -110
rect 17181 -85 17216 -70
rect 17181 -110 17186 -85
rect 17211 -110 17216 -85
rect 17181 -120 17216 -110
rect 17241 -85 17276 -70
rect 17241 -110 17246 -85
rect 17271 -110 17276 -85
rect 17241 -120 17276 -110
rect 17301 -85 17336 -70
rect 17301 -110 17306 -85
rect 17331 -110 17336 -85
rect 17301 -120 17336 -110
rect 17361 -85 17396 -70
rect 17361 -110 17366 -85
rect 17391 -110 17396 -85
rect 17361 -120 17396 -110
rect 17421 -85 17456 -70
rect 17421 -110 17426 -85
rect 17451 -110 17456 -85
rect 17421 -120 17456 -110
rect 17481 -85 17521 -70
rect 17481 -110 17491 -85
rect 17516 -110 17521 -85
rect 17481 -120 17521 -110
rect 17546 -85 17581 -70
rect 17546 -110 17551 -85
rect 17576 -110 17581 -85
rect 17546 -120 17581 -110
rect 17606 -85 17641 -70
rect 17606 -110 17611 -85
rect 17636 -110 17641 -85
rect 17606 -120 17641 -110
rect 17666 -85 17701 -70
rect 17666 -110 17671 -85
rect 17696 -110 17701 -85
rect 17666 -120 17701 -110
rect 17726 -85 17761 -70
rect 17726 -110 17731 -85
rect 17756 -110 17761 -85
rect 17726 -120 17761 -110
rect 17786 -85 17821 -70
rect 17786 -110 17791 -85
rect 17816 -110 17821 -85
rect 17786 -120 17821 -110
rect 17846 -85 17881 -70
rect 17846 -110 17851 -85
rect 17876 -110 17881 -85
rect 17846 -120 17881 -110
rect 17906 -85 17941 -70
rect 17906 -110 17911 -85
rect 17936 -110 17941 -85
rect 17906 -120 17941 -110
rect 17966 -85 18006 -70
rect 17966 -110 17976 -85
rect 18001 -110 18006 -85
rect 17966 -120 18006 -110
rect 18031 -85 18066 -70
rect 18031 -110 18036 -85
rect 18061 -110 18066 -85
rect 18031 -120 18066 -110
rect 18091 -85 18126 -70
rect 18091 -110 18096 -85
rect 18121 -110 18126 -85
rect 18091 -120 18126 -110
rect 18151 -85 18186 -70
rect 18151 -110 18156 -85
rect 18181 -110 18186 -85
rect 18151 -120 18186 -110
rect 18211 -85 18246 -70
rect 18211 -110 18216 -85
rect 18241 -110 18246 -85
rect 18211 -120 18246 -110
rect 18271 -85 18306 -70
rect 18271 -110 18276 -85
rect 18301 -110 18306 -85
rect 18271 -120 18306 -110
rect 18331 -85 18366 -70
rect 18331 -110 18336 -85
rect 18361 -110 18366 -85
rect 18331 -120 18366 -110
rect 18391 -85 18426 -70
rect 18391 -110 18396 -85
rect 18421 -110 18426 -85
rect 18391 -120 18426 -110
rect 18451 -85 18491 -70
rect 18451 -110 18461 -85
rect 18486 -110 18491 -85
rect 18451 -120 18491 -110
rect 18516 -85 18551 -70
rect 18516 -110 18521 -85
rect 18546 -110 18551 -85
rect 18516 -120 18551 -110
rect 18576 -85 18611 -70
rect 18576 -110 18581 -85
rect 18606 -110 18611 -85
rect 18576 -120 18611 -110
rect 18636 -85 18671 -70
rect 18636 -110 18641 -85
rect 18666 -110 18671 -85
rect 18636 -120 18671 -110
rect 18696 -85 18731 -70
rect 18696 -110 18701 -85
rect 18726 -110 18731 -85
rect 18696 -120 18731 -110
rect 18756 -85 18791 -70
rect 18756 -110 18761 -85
rect 18786 -110 18791 -85
rect 18756 -120 18791 -110
rect 18816 -85 18851 -70
rect 18816 -110 18821 -85
rect 18846 -110 18851 -85
rect 18816 -120 18851 -110
rect 18876 -85 18911 -70
rect 18876 -110 18881 -85
rect 18906 -110 18911 -85
rect 18876 -120 18911 -110
rect 18936 -85 18976 -70
rect 18936 -110 18946 -85
rect 18971 -110 18976 -85
rect 18936 -120 18976 -110
rect 19001 -85 19036 -70
rect 19001 -110 19006 -85
rect 19031 -110 19036 -85
rect 19001 -120 19036 -110
rect 19061 -85 19096 -70
rect 19061 -110 19066 -85
rect 19091 -110 19096 -85
rect 19061 -120 19096 -110
rect 19121 -85 19156 -70
rect 19121 -110 19126 -85
rect 19151 -110 19156 -85
rect 19121 -120 19156 -110
rect 19181 -85 19216 -70
rect 19181 -110 19186 -85
rect 19211 -110 19216 -85
rect 19181 -120 19216 -110
rect 19241 -85 19276 -70
rect 19241 -110 19246 -85
rect 19271 -110 19276 -85
rect 19241 -120 19276 -110
rect 19301 -85 19336 -70
rect 19301 -110 19306 -85
rect 19331 -110 19336 -85
rect 19301 -120 19336 -110
rect 19361 -85 19396 -70
rect 19361 -110 19366 -85
rect 19391 -110 19396 -85
rect 19361 -120 19396 -110
rect 19421 -85 19461 -70
rect 19421 -110 19431 -85
rect 19456 -110 19461 -85
rect 19421 -120 19461 -110
rect 19486 -85 19521 -70
rect 19486 -110 19491 -85
rect 19516 -110 19521 -85
rect 19486 -120 19521 -110
rect 19546 -85 19581 -70
rect 19546 -110 19551 -85
rect 19576 -110 19581 -85
rect 19546 -120 19581 -110
rect 19606 -85 19641 -70
rect 19606 -110 19611 -85
rect 19636 -110 19641 -85
rect 19606 -120 19641 -110
rect 19666 -85 19701 -70
rect 19666 -110 19671 -85
rect 19696 -110 19701 -85
rect 19666 -120 19701 -110
rect 19726 -85 19761 -70
rect 19726 -110 19731 -85
rect 19756 -110 19761 -85
rect 19726 -120 19761 -110
rect 19786 -85 19821 -70
rect 19786 -110 19791 -85
rect 19816 -110 19821 -85
rect 19786 -120 19821 -110
rect 19846 -85 19881 -70
rect 19846 -110 19851 -85
rect 19876 -110 19881 -85
rect 19846 -120 19881 -110
rect 19906 -85 19946 -70
rect 19906 -110 19916 -85
rect 19941 -110 19946 -85
rect 19906 -120 19946 -110
rect 19971 -85 20006 -70
rect 19971 -110 19976 -85
rect 20001 -110 20006 -85
rect 19971 -120 20006 -110
rect 20031 -85 20066 -70
rect 20031 -110 20036 -85
rect 20061 -110 20066 -85
rect 20031 -120 20066 -110
rect 20091 -85 20126 -70
rect 20091 -110 20096 -85
rect 20121 -110 20126 -85
rect 20091 -120 20126 -110
rect 20151 -85 20186 -70
rect 20151 -110 20156 -85
rect 20181 -110 20186 -85
rect 20151 -120 20186 -110
rect 20211 -85 20246 -70
rect 20211 -110 20216 -85
rect 20241 -110 20246 -85
rect 20211 -120 20246 -110
rect 20271 -85 20306 -70
rect 20271 -110 20276 -85
rect 20301 -110 20306 -85
rect 20271 -120 20306 -110
rect 20331 -85 20366 -70
rect 20331 -110 20336 -85
rect 20361 -110 20366 -85
rect 20331 -120 20366 -110
rect 20391 -85 20431 -70
rect 20391 -110 20401 -85
rect 20426 -110 20431 -85
rect 20391 -120 20431 -110
rect 20456 -85 20491 -70
rect 20456 -110 20461 -85
rect 20486 -110 20491 -85
rect 20456 -120 20491 -110
rect 20516 -85 20551 -70
rect 20516 -110 20521 -85
rect 20546 -110 20551 -85
rect 20516 -120 20551 -110
rect 20576 -85 20611 -70
rect 20576 -110 20581 -85
rect 20606 -110 20611 -85
rect 20576 -120 20611 -110
rect 20636 -85 20671 -70
rect 20636 -110 20641 -85
rect 20666 -110 20671 -85
rect 20636 -120 20671 -110
rect 20696 -85 20731 -70
rect 20696 -110 20701 -85
rect 20726 -110 20731 -85
rect 20696 -120 20731 -110
rect 20756 -85 20791 -70
rect 20756 -110 20761 -85
rect 20786 -110 20791 -85
rect 20756 -120 20791 -110
rect 20816 -85 20851 -70
rect 20816 -110 20821 -85
rect 20846 -110 20851 -85
rect 20816 -120 20851 -110
rect 20876 -85 20916 -70
rect 20876 -110 20886 -85
rect 20911 -110 20916 -85
rect 20876 -120 20916 -110
rect 20941 -85 20976 -70
rect 20941 -110 20946 -85
rect 20971 -110 20976 -85
rect 20941 -120 20976 -110
rect 21001 -85 21036 -70
rect 21001 -110 21006 -85
rect 21031 -110 21036 -85
rect 21001 -120 21036 -110
rect 21061 -85 21096 -70
rect 21061 -110 21066 -85
rect 21091 -110 21096 -85
rect 21061 -120 21096 -110
rect 21121 -85 21156 -70
rect 21121 -110 21126 -85
rect 21151 -110 21156 -85
rect 21121 -120 21156 -110
rect 21520 -105 21765 -5
rect 21865 -105 22315 -5
rect 22415 -105 22865 -5
rect 22965 -105 23415 -5
rect 23515 -105 23965 -5
rect 24065 -105 24515 -5
rect 24615 -105 25065 -5
rect 25165 -105 25615 -5
rect 25715 -105 26165 -5
rect 26265 -105 26715 -5
rect 26815 -105 27265 -5
rect 27365 -105 27815 -5
rect 27915 -105 28365 -5
rect 28465 -105 28915 -5
rect 29015 -105 29465 -5
rect 29565 -105 30015 -5
rect 30115 -105 30565 -5
rect 30665 -105 31200 -5
rect 191 -170 211 -120
rect 386 -125 406 -120
rect 436 -170 456 -120
rect 506 -125 526 -120
rect 691 -125 711 -120
rect 741 -170 761 -120
rect 811 -125 831 -120
rect 936 -125 956 -120
rect 986 -170 1006 -120
rect 1056 -125 1076 -120
rect 1176 -125 1196 -120
rect 1226 -170 1246 -120
rect 1296 -125 1316 -120
rect 1421 -125 1441 -120
rect 1471 -170 1491 -120
rect 1541 -125 1561 -120
rect 1726 -125 1746 -120
rect 1776 -170 1796 -120
rect 1846 -125 1866 -120
rect 1971 -125 1991 -120
rect 2021 -170 2041 -120
rect 2091 -125 2111 -120
rect 2211 -125 2231 -120
rect 2261 -170 2281 -120
rect 2331 -125 2351 -120
rect 2456 -125 2476 -120
rect 2506 -170 2526 -120
rect 2576 -125 2596 -120
rect 2696 -125 2716 -120
rect 2746 -170 2766 -120
rect 2816 -125 2836 -120
rect 2941 -125 2961 -120
rect 2991 -170 3011 -120
rect 3061 -125 3081 -120
rect 3181 -125 3201 -120
rect 3231 -170 3251 -120
rect 3301 -125 3321 -120
rect 3426 -125 3446 -120
rect 3476 -170 3496 -120
rect 3546 -125 3566 -120
rect 3666 -125 3686 -120
rect 3716 -170 3736 -120
rect 3786 -125 3806 -120
rect 3911 -125 3931 -120
rect 3961 -170 3981 -120
rect 4031 -125 4051 -120
rect 4151 -125 4171 -120
rect 4201 -170 4221 -120
rect 4271 -125 4291 -120
rect 4396 -125 4416 -120
rect -460 -240 -415 -190
rect -365 -240 -320 -190
rect -460 -555 -320 -240
rect 1625 -200 1685 -190
rect 1625 -240 1635 -200
rect 1675 -240 1685 -200
rect 1625 -250 1685 -240
rect 4050 -195 4110 -185
rect 4446 -170 4466 -120
rect 4516 -125 4536 -120
rect 4636 -125 4656 -120
rect 4686 -170 4706 -120
rect 4756 -125 4776 -120
rect 4881 -125 4901 -120
rect 4931 -170 4951 -120
rect 5001 -125 5021 -120
rect 5121 -125 5141 -120
rect 5171 -170 5191 -120
rect 5241 -125 5261 -120
rect 5366 -125 5386 -120
rect 5416 -170 5436 -120
rect 5486 -125 5506 -120
rect 5671 -125 5691 -120
rect 5721 -170 5741 -120
rect 5791 -125 5811 -120
rect 5916 -125 5936 -120
rect 5966 -170 5986 -120
rect 6036 -125 6056 -120
rect 6156 -125 6176 -120
rect 6206 -170 6226 -120
rect 6276 -125 6296 -120
rect 6451 -155 6471 -120
rect 6521 -125 6541 -120
rect 6641 -125 6661 -120
rect 6450 -160 6470 -155
rect 6335 -180 6470 -160
rect 6691 -170 6711 -120
rect 6761 -125 6781 -120
rect 6886 -125 6906 -120
rect 4050 -235 4060 -195
rect 4100 -235 4110 -195
rect 4050 -245 4110 -235
rect 6335 -250 6355 -180
rect 6936 -170 6956 -120
rect 7006 -125 7026 -120
rect 7126 -125 7146 -120
rect 7176 -170 7196 -120
rect 7246 -125 7266 -120
rect 7366 -125 7386 -120
rect 7416 -170 7436 -120
rect 7486 -125 7506 -120
rect 7606 -125 7626 -120
rect 7656 -170 7676 -120
rect 7726 -125 7746 -120
rect 7851 -125 7871 -120
rect 7901 -140 7921 -120
rect 7900 -150 7921 -140
rect 7971 -125 7991 -120
rect 8091 -125 8111 -120
rect 7900 -165 7920 -150
rect 7775 -185 7920 -165
rect 8141 -170 8161 -120
rect 8211 -125 8231 -120
rect 8336 -125 8356 -120
rect 25 -320 45 -315
rect 95 -320 115 -270
rect 145 -320 165 -315
rect 265 -320 285 -315
rect 335 -320 355 -270
rect 385 -320 405 -315
rect 505 -320 525 -315
rect 575 -320 595 -270
rect 625 -320 645 -315
rect 745 -320 765 -315
rect 815 -320 835 -270
rect 865 -320 885 -315
rect 985 -320 1005 -315
rect 1055 -320 1075 -270
rect 1105 -320 1125 -315
rect 1225 -320 1245 -315
rect 1295 -320 1315 -270
rect 1345 -320 1365 -315
rect 1465 -320 1485 -315
rect 1535 -320 1555 -270
rect 1585 -320 1605 -315
rect 1705 -320 1725 -315
rect 1775 -320 1795 -270
rect 1825 -320 1845 -315
rect 1945 -320 1965 -315
rect 2015 -320 2035 -270
rect 2065 -320 2085 -315
rect 2185 -320 2205 -315
rect 2255 -320 2275 -270
rect 2305 -320 2325 -315
rect 2425 -320 2445 -315
rect 2495 -320 2515 -270
rect 2545 -320 2565 -315
rect 2665 -320 2685 -315
rect 2735 -320 2755 -270
rect 2785 -320 2805 -315
rect 2905 -320 2925 -315
rect 2975 -320 2995 -270
rect 3025 -320 3045 -315
rect 3145 -320 3165 -315
rect 3215 -320 3235 -270
rect 3265 -320 3285 -315
rect 3385 -320 3405 -315
rect 3455 -320 3475 -270
rect 3505 -320 3525 -315
rect 3625 -320 3645 -315
rect 3695 -320 3715 -270
rect 3745 -320 3765 -315
rect 3865 -320 3885 -315
rect 3935 -320 3955 -270
rect 3985 -320 4005 -315
rect 4105 -320 4125 -315
rect 4175 -320 4195 -270
rect 4225 -320 4245 -315
rect 4345 -320 4365 -315
rect 4415 -320 4435 -270
rect 4465 -320 4485 -315
rect 4585 -320 4605 -315
rect 4655 -320 4675 -270
rect 4705 -320 4725 -315
rect 4825 -320 4845 -315
rect 4895 -320 4915 -270
rect 4945 -320 4965 -315
rect 5065 -320 5085 -315
rect 5135 -320 5155 -270
rect 5185 -320 5205 -315
rect 5305 -320 5325 -315
rect 5375 -320 5395 -270
rect 5425 -320 5445 -315
rect 5545 -320 5565 -315
rect 5615 -320 5635 -270
rect 5665 -320 5685 -315
rect 5785 -320 5805 -315
rect 5855 -320 5875 -270
rect 5905 -320 5925 -315
rect 6025 -320 6045 -315
rect 6095 -320 6115 -270
rect 6445 -220 6505 -210
rect 6445 -260 6455 -220
rect 6495 -260 6505 -220
rect 7775 -250 7795 -185
rect 8386 -170 8406 -120
rect 8456 -125 8476 -120
rect 8576 -125 8596 -120
rect 8626 -170 8646 -120
rect 8696 -125 8716 -120
rect 8821 -125 8841 -120
rect 8871 -170 8891 -120
rect 8941 -125 8961 -120
rect 9061 -125 9081 -120
rect 9111 -170 9131 -120
rect 9181 -125 9201 -120
rect 9306 -125 9326 -120
rect 9356 -170 9376 -120
rect 9426 -125 9446 -120
rect 9601 -145 9621 -120
rect 9671 -125 9691 -120
rect 9796 -125 9816 -120
rect 9600 -150 9621 -145
rect 9600 -160 9620 -150
rect 9455 -180 9620 -160
rect 9846 -170 9866 -120
rect 9916 -125 9936 -120
rect 10036 -125 10056 -120
rect 6445 -270 6505 -260
rect 6145 -320 6165 -315
rect 6265 -320 6285 -315
rect 6335 -320 6355 -270
rect 6385 -320 6405 -315
rect 6505 -320 6525 -315
rect 6575 -320 6595 -270
rect 6625 -320 6645 -315
rect 6745 -320 6765 -315
rect 6815 -320 6835 -270
rect 6865 -320 6885 -315
rect 6985 -320 7005 -315
rect 7055 -320 7075 -270
rect 7105 -320 7125 -315
rect 7225 -320 7245 -315
rect 7295 -320 7315 -270
rect 7345 -320 7365 -315
rect 7465 -320 7485 -315
rect 7535 -320 7555 -270
rect 7870 -220 7930 -210
rect 7870 -260 7880 -220
rect 7920 -260 7930 -220
rect 9455 -250 9475 -180
rect 10086 -170 10106 -120
rect 10156 -125 10176 -120
rect 10281 -125 10301 -120
rect 10331 -170 10351 -120
rect 10401 -125 10421 -120
rect 10521 -125 10541 -120
rect 10571 -170 10591 -120
rect 10641 -125 10661 -120
rect 10766 -125 10786 -120
rect 10816 -170 10836 -120
rect 10886 -125 10906 -120
rect 11006 -125 11026 -120
rect 11056 -170 11076 -120
rect 11126 -125 11146 -120
rect 11251 -125 11271 -120
rect 11301 -170 11321 -120
rect 11371 -125 11391 -120
rect 11491 -125 11511 -120
rect 11541 -170 11561 -120
rect 11611 -125 11631 -120
rect 11736 -125 11756 -120
rect 11786 -170 11806 -120
rect 11856 -125 11876 -120
rect 11976 -125 11996 -120
rect 12026 -150 12046 -120
rect 12096 -125 12116 -120
rect 12221 -125 12241 -120
rect 12025 -170 12045 -150
rect 11855 -190 12045 -170
rect 12271 -170 12291 -120
rect 12341 -125 12361 -120
rect 12461 -125 12481 -120
rect 12511 -170 12531 -120
rect 12581 -125 12601 -120
rect 12706 -125 12726 -120
rect 12756 -170 12776 -120
rect 12826 -125 12846 -120
rect 12946 -125 12966 -120
rect 12996 -170 13016 -120
rect 13066 -125 13086 -120
rect 13191 -125 13211 -120
rect 13241 -170 13261 -120
rect 13311 -125 13331 -120
rect 13431 -125 13451 -120
rect 13481 -170 13501 -120
rect 13551 -125 13571 -120
rect 13676 -125 13696 -120
rect 13726 -170 13746 -120
rect 13796 -125 13816 -120
rect 13916 -125 13936 -120
rect 13966 -145 13986 -120
rect 14036 -125 14056 -120
rect 14161 -125 14181 -120
rect 13965 -150 13986 -145
rect 13965 -165 13985 -150
rect 13780 -190 13985 -165
rect 14211 -170 14231 -120
rect 14281 -125 14301 -120
rect 14401 -125 14421 -120
rect 14451 -170 14471 -120
rect 14521 -125 14541 -120
rect 14646 -125 14666 -120
rect 14696 -170 14716 -120
rect 14766 -125 14786 -120
rect 14886 -125 14906 -120
rect 14936 -170 14956 -120
rect 15006 -125 15026 -120
rect 15131 -125 15151 -120
rect 15181 -170 15201 -120
rect 15251 -125 15271 -120
rect 15371 -125 15391 -120
rect 15421 -170 15441 -120
rect 15491 -125 15511 -120
rect 15616 -125 15636 -120
rect 15666 -170 15686 -120
rect 15736 -125 15756 -120
rect 15856 -125 15876 -120
rect 15906 -140 15926 -120
rect 15905 -145 15926 -140
rect 15976 -125 15996 -120
rect 16101 -125 16121 -120
rect 15905 -165 15925 -145
rect 15750 -185 15925 -165
rect 16151 -170 16171 -120
rect 16221 -125 16241 -120
rect 16341 -125 16361 -120
rect 7870 -270 7930 -260
rect 7585 -320 7605 -315
rect 7705 -320 7725 -315
rect 7775 -320 7795 -270
rect 7825 -320 7845 -315
rect 7945 -320 7965 -315
rect 8015 -320 8035 -270
rect 8065 -320 8085 -315
rect 8185 -320 8205 -315
rect 8255 -320 8275 -270
rect 8305 -320 8325 -315
rect 8425 -320 8445 -315
rect 8495 -320 8515 -270
rect 8545 -320 8565 -315
rect 8665 -320 8685 -315
rect 8735 -320 8755 -270
rect 8785 -320 8805 -315
rect 8905 -320 8925 -315
rect 8975 -320 8995 -270
rect 9025 -320 9045 -315
rect 9145 -320 9165 -315
rect 9215 -320 9235 -270
rect 9560 -210 9620 -200
rect 9560 -250 9570 -210
rect 9610 -250 9620 -210
rect 11855 -250 11880 -190
rect 11940 -220 12000 -210
rect 9560 -260 9620 -250
rect 9265 -320 9285 -315
rect 9385 -320 9405 -315
rect 9455 -320 9475 -270
rect 9505 -320 9525 -315
rect 9625 -320 9645 -315
rect 9695 -320 9715 -270
rect 9745 -320 9765 -315
rect 9865 -320 9885 -315
rect 9935 -320 9955 -270
rect 9985 -320 10005 -315
rect 10105 -320 10125 -315
rect 10175 -320 10195 -270
rect 10225 -320 10245 -315
rect 10345 -320 10365 -315
rect 10415 -320 10435 -270
rect 10465 -320 10485 -315
rect 10585 -320 10605 -315
rect 10655 -320 10675 -270
rect 10705 -320 10725 -315
rect 10825 -320 10845 -315
rect 10895 -320 10915 -270
rect 10945 -320 10965 -315
rect 11065 -320 11085 -315
rect 11135 -320 11155 -270
rect 11185 -320 11205 -315
rect 11305 -320 11325 -315
rect 11375 -320 11395 -270
rect 11425 -320 11445 -315
rect 11545 -320 11565 -315
rect 11615 -320 11635 -270
rect 11940 -260 11950 -220
rect 11990 -260 12000 -220
rect 13780 -230 13800 -190
rect 13775 -250 13800 -230
rect 13860 -220 13920 -210
rect 11940 -270 12000 -260
rect 11665 -320 11685 -315
rect 11785 -320 11805 -315
rect 11855 -320 11875 -270
rect 11905 -320 11925 -315
rect 12025 -320 12045 -315
rect 12095 -320 12115 -270
rect 12145 -320 12165 -315
rect 12265 -320 12285 -315
rect 12335 -320 12355 -270
rect 12385 -320 12405 -315
rect 12505 -320 12525 -315
rect 12575 -320 12595 -270
rect 12625 -320 12645 -315
rect 12745 -320 12765 -315
rect 12815 -320 12835 -270
rect 12865 -320 12885 -315
rect 12985 -320 13005 -315
rect 13055 -320 13075 -270
rect 13105 -320 13125 -315
rect 13225 -320 13245 -315
rect 13295 -320 13315 -270
rect 13345 -320 13365 -315
rect 13465 -320 13485 -315
rect 13535 -320 13555 -270
rect 13860 -260 13870 -220
rect 13910 -260 13920 -220
rect 15750 -250 15770 -185
rect 16391 -170 16411 -120
rect 16461 -125 16481 -120
rect 16586 -125 16606 -120
rect 16636 -170 16656 -120
rect 16706 -125 16726 -120
rect 16826 -125 16846 -120
rect 16876 -170 16896 -120
rect 16946 -125 16966 -120
rect 17071 -125 17091 -120
rect 17121 -170 17141 -120
rect 17191 -125 17211 -120
rect 17311 -125 17331 -120
rect 17361 -170 17381 -120
rect 17431 -125 17451 -120
rect 17556 -125 17576 -120
rect 17606 -170 17626 -120
rect 17676 -125 17696 -120
rect 17796 -125 17816 -120
rect 17846 -170 17866 -120
rect 17916 -125 17936 -120
rect 18041 -125 18061 -120
rect 18091 -170 18111 -120
rect 18161 -125 18181 -120
rect 18281 -125 18301 -120
rect 18331 -170 18351 -120
rect 18401 -125 18421 -120
rect 18526 -125 18546 -120
rect 18576 -170 18596 -120
rect 18646 -125 18666 -120
rect 18766 -125 18786 -120
rect 18816 -170 18836 -120
rect 18886 -125 18906 -120
rect 19011 -125 19031 -120
rect 19061 -170 19081 -120
rect 19131 -125 19151 -120
rect 19251 -125 19271 -120
rect 19301 -170 19321 -120
rect 19371 -125 19391 -120
rect 19496 -125 19516 -120
rect 19546 -170 19566 -120
rect 19616 -125 19636 -120
rect 19736 -125 19756 -120
rect 19786 -170 19806 -120
rect 19856 -125 19876 -120
rect 19981 -125 20001 -120
rect 20031 -170 20051 -120
rect 20101 -125 20121 -120
rect 20221 -125 20241 -120
rect 20271 -170 20291 -120
rect 20341 -125 20361 -120
rect 20466 -125 20486 -120
rect 20516 -170 20536 -120
rect 20586 -125 20606 -120
rect 20706 -125 20726 -120
rect 20756 -170 20776 -120
rect 20826 -125 20846 -120
rect 20951 -125 20971 -120
rect 21001 -170 21021 -120
rect 21071 -125 21091 -120
rect 21520 -125 31200 -105
rect 17695 -210 17755 -200
rect 13860 -270 13920 -260
rect 13585 -320 13605 -315
rect 13705 -320 13725 -315
rect 13775 -320 13795 -270
rect 13825 -320 13845 -315
rect 13945 -320 13965 -315
rect 14015 -320 14035 -270
rect 14065 -320 14085 -315
rect 14185 -320 14205 -315
rect 14255 -320 14275 -270
rect 14305 -320 14325 -315
rect 14425 -320 14445 -315
rect 14495 -320 14515 -270
rect 14545 -320 14565 -315
rect 14665 -320 14685 -315
rect 14735 -320 14755 -270
rect 14785 -320 14805 -315
rect 14905 -320 14925 -315
rect 14975 -320 14995 -270
rect 15025 -320 15045 -315
rect 15145 -320 15165 -315
rect 15215 -320 15235 -270
rect 15265 -320 15285 -315
rect 15385 -320 15405 -315
rect 15455 -320 15475 -270
rect 15715 -270 15770 -250
rect 15805 -220 15865 -210
rect 15805 -260 15815 -220
rect 15855 -260 15865 -220
rect 17695 -250 17705 -210
rect 17745 -250 17755 -210
rect 19635 -210 19695 -200
rect 19635 -250 19645 -210
rect 19685 -250 19695 -210
rect 31060 -220 31200 -125
rect 15805 -270 15865 -260
rect 15505 -320 15525 -315
rect 15625 -320 15645 -315
rect 15695 -320 15715 -270
rect 15745 -320 15765 -315
rect 15865 -320 15885 -315
rect 15935 -320 15955 -270
rect 15985 -320 16005 -315
rect 16105 -320 16125 -315
rect 16175 -320 16195 -270
rect 16225 -320 16245 -315
rect 16345 -320 16365 -315
rect 16415 -320 16435 -270
rect 16465 -320 16485 -315
rect 16585 -320 16605 -315
rect 16655 -320 16675 -270
rect 16705 -320 16725 -315
rect 16825 -320 16845 -315
rect 16895 -320 16915 -270
rect 16945 -320 16965 -315
rect 17065 -320 17085 -315
rect 17135 -320 17155 -270
rect 17185 -320 17205 -315
rect 17305 -320 17325 -315
rect 17375 -320 17395 -270
rect 17695 -260 17755 -250
rect 17425 -320 17445 -315
rect 17545 -320 17565 -315
rect 17615 -320 17635 -270
rect 17665 -320 17685 -315
rect 17785 -320 17805 -315
rect 17855 -320 17875 -270
rect 17905 -320 17925 -315
rect 18025 -320 18045 -315
rect 18095 -320 18115 -270
rect 18145 -320 18165 -315
rect 18265 -320 18285 -315
rect 18335 -320 18355 -270
rect 18385 -320 18405 -315
rect 18505 -320 18525 -315
rect 18575 -320 18595 -270
rect 18625 -320 18645 -315
rect 18745 -320 18765 -315
rect 18815 -320 18835 -270
rect 18865 -320 18885 -315
rect 18985 -320 19005 -315
rect 19055 -320 19075 -270
rect 19105 -320 19125 -315
rect 19225 -320 19245 -315
rect 19295 -320 19315 -270
rect 19635 -260 19695 -250
rect 19345 -320 19365 -315
rect 19465 -320 19485 -315
rect 19535 -320 19555 -270
rect 19585 -320 19605 -315
rect 19705 -320 19725 -315
rect 19775 -320 19795 -270
rect 19825 -320 19845 -315
rect 19945 -320 19965 -315
rect 20015 -320 20035 -270
rect 20065 -320 20085 -315
rect 20185 -320 20205 -315
rect 20255 -320 20275 -270
rect 20305 -320 20325 -315
rect 20425 -320 20445 -315
rect 20495 -320 20515 -270
rect 20545 -320 20565 -315
rect 20665 -320 20685 -315
rect 20735 -320 20755 -270
rect 20785 -320 20805 -315
rect 20905 -320 20925 -315
rect 20975 -320 20995 -270
rect 21025 -320 21045 -315
rect 21145 -320 21165 -315
rect 21215 -320 21235 -270
rect 21265 -320 21285 -315
rect 21385 -320 21405 -315
rect 21455 -320 21475 -270
rect 21505 -320 21525 -315
rect 21625 -320 21645 -315
rect 21695 -320 21715 -270
rect 21745 -320 21765 -315
rect 21865 -320 21885 -315
rect 21935 -320 21955 -270
rect 21985 -320 22005 -315
rect 22105 -320 22125 -315
rect 22175 -320 22195 -270
rect 22225 -320 22245 -315
rect 22345 -320 22365 -315
rect 22415 -320 22435 -270
rect 22465 -320 22485 -315
rect 22585 -320 22605 -315
rect 22655 -320 22675 -270
rect 22705 -320 22725 -315
rect 22825 -320 22845 -315
rect 22895 -320 22915 -270
rect 22945 -320 22965 -315
rect 23065 -320 23085 -315
rect 23135 -320 23155 -270
rect 23185 -320 23205 -315
rect 23305 -320 23325 -315
rect 23375 -320 23395 -270
rect 23425 -320 23445 -315
rect 23545 -320 23565 -315
rect 23615 -320 23635 -270
rect 23665 -320 23685 -315
rect 23785 -320 23805 -315
rect 23855 -320 23875 -270
rect 23905 -320 23925 -315
rect 24025 -320 24045 -315
rect 24095 -320 24115 -270
rect 24145 -320 24165 -315
rect 24265 -320 24285 -315
rect 24335 -320 24355 -270
rect 24385 -320 24405 -315
rect 24505 -320 24525 -315
rect 24575 -320 24595 -270
rect 24625 -320 24645 -315
rect 24745 -320 24765 -315
rect 24815 -320 24835 -270
rect 24865 -320 24885 -315
rect 24985 -320 25005 -315
rect 25055 -320 25075 -270
rect 25105 -320 25125 -315
rect 25225 -320 25245 -315
rect 25295 -320 25315 -270
rect 25345 -320 25365 -315
rect 25465 -320 25485 -315
rect 25535 -320 25555 -270
rect 25585 -320 25605 -315
rect 25705 -320 25725 -315
rect 25775 -320 25795 -270
rect 25825 -320 25845 -315
rect 25945 -320 25965 -315
rect 26015 -320 26035 -270
rect 26065 -320 26085 -315
rect 26185 -320 26205 -315
rect 26255 -320 26275 -270
rect 26305 -320 26325 -315
rect 26425 -320 26445 -315
rect 26495 -320 26515 -270
rect 26545 -320 26565 -315
rect 26665 -320 26685 -315
rect 26735 -320 26755 -270
rect 26785 -320 26805 -315
rect 26905 -320 26925 -315
rect 26975 -320 26995 -270
rect 27025 -320 27045 -315
rect 27145 -320 27165 -315
rect 27215 -320 27235 -270
rect 27265 -320 27285 -315
rect 27385 -320 27405 -315
rect 27455 -320 27475 -270
rect 27505 -320 27525 -315
rect 27625 -320 27645 -315
rect 27695 -320 27715 -270
rect 27745 -320 27765 -315
rect 27865 -320 27885 -315
rect 27935 -320 27955 -270
rect 27985 -320 28005 -315
rect 28105 -320 28125 -315
rect 28175 -320 28195 -270
rect 28225 -320 28245 -315
rect 28345 -320 28365 -315
rect 28415 -320 28435 -270
rect 28465 -320 28485 -315
rect 28585 -320 28605 -315
rect 28655 -320 28675 -270
rect 28705 -320 28725 -315
rect 28825 -320 28845 -315
rect 28895 -320 28915 -270
rect 28945 -320 28965 -315
rect 29065 -320 29085 -315
rect 29135 -320 29155 -270
rect 29185 -320 29205 -315
rect 29305 -320 29325 -315
rect 29375 -320 29395 -270
rect 29425 -320 29445 -315
rect 29545 -320 29565 -315
rect 29615 -320 29635 -270
rect 29665 -320 29685 -315
rect 29785 -320 29805 -315
rect 29855 -320 29875 -270
rect 29905 -320 29925 -315
rect 30025 -320 30045 -315
rect 30095 -320 30115 -270
rect 30145 -320 30165 -315
rect 30265 -320 30285 -315
rect 30335 -320 30355 -270
rect 30385 -320 30405 -315
rect 30505 -320 30525 -315
rect 30575 -320 30595 -270
rect 30625 -320 30645 -315
rect 31060 -320 31080 -220
rect 31180 -320 31200 -220
rect -40 -335 -5 -320
rect -40 -360 -35 -335
rect -10 -360 -5 -335
rect -40 -380 -5 -360
rect -40 -405 -35 -380
rect -10 -405 -5 -380
rect -40 -420 -5 -405
rect 20 -335 55 -320
rect 20 -360 25 -335
rect 50 -360 55 -335
rect 20 -380 55 -360
rect 20 -405 25 -380
rect 50 -405 55 -380
rect 20 -420 55 -405
rect 80 -335 115 -320
rect 80 -360 85 -335
rect 110 -360 115 -335
rect 80 -380 115 -360
rect 80 -405 85 -380
rect 110 -405 115 -380
rect 80 -420 115 -405
rect 140 -335 175 -320
rect 140 -360 145 -335
rect 170 -360 175 -335
rect 140 -380 175 -360
rect 140 -405 145 -380
rect 170 -405 175 -380
rect 140 -420 175 -405
rect 200 -335 235 -320
rect 200 -360 205 -335
rect 230 -360 235 -335
rect 200 -380 235 -360
rect 200 -405 205 -380
rect 230 -405 235 -380
rect 200 -420 235 -405
rect 260 -335 295 -320
rect 260 -360 265 -335
rect 290 -360 295 -335
rect 260 -380 295 -360
rect 260 -405 265 -380
rect 290 -405 295 -380
rect 260 -420 295 -405
rect 320 -335 355 -320
rect 320 -360 325 -335
rect 350 -360 355 -335
rect 320 -380 355 -360
rect 320 -405 325 -380
rect 350 -405 355 -380
rect 320 -420 355 -405
rect 380 -335 415 -320
rect 380 -360 385 -335
rect 410 -360 415 -335
rect 380 -380 415 -360
rect 380 -405 385 -380
rect 410 -405 415 -380
rect 380 -420 415 -405
rect 440 -335 475 -320
rect 440 -360 445 -335
rect 470 -360 475 -335
rect 440 -380 475 -360
rect 440 -405 445 -380
rect 470 -405 475 -380
rect 440 -420 475 -405
rect 500 -335 535 -320
rect 500 -360 505 -335
rect 530 -360 535 -335
rect 500 -380 535 -360
rect 500 -405 505 -380
rect 530 -405 535 -380
rect 500 -420 535 -405
rect 560 -335 595 -320
rect 560 -360 565 -335
rect 590 -360 595 -335
rect 560 -380 595 -360
rect 560 -405 565 -380
rect 590 -405 595 -380
rect 560 -420 595 -405
rect 620 -335 655 -320
rect 620 -360 625 -335
rect 650 -360 655 -335
rect 620 -380 655 -360
rect 620 -405 625 -380
rect 650 -405 655 -380
rect 620 -420 655 -405
rect 680 -335 715 -320
rect 680 -360 685 -335
rect 710 -360 715 -335
rect 680 -380 715 -360
rect 680 -405 685 -380
rect 710 -405 715 -380
rect 680 -420 715 -405
rect 740 -335 775 -320
rect 740 -360 745 -335
rect 770 -360 775 -335
rect 740 -380 775 -360
rect 740 -405 745 -380
rect 770 -405 775 -380
rect 740 -420 775 -405
rect 800 -335 835 -320
rect 800 -360 805 -335
rect 830 -360 835 -335
rect 800 -380 835 -360
rect 800 -405 805 -380
rect 830 -405 835 -380
rect 800 -420 835 -405
rect 860 -335 895 -320
rect 860 -360 865 -335
rect 890 -360 895 -335
rect 860 -380 895 -360
rect 860 -405 865 -380
rect 890 -405 895 -380
rect 860 -420 895 -405
rect 920 -335 955 -320
rect 920 -360 925 -335
rect 950 -360 955 -335
rect 920 -380 955 -360
rect 920 -405 925 -380
rect 950 -405 955 -380
rect 920 -420 955 -405
rect 980 -335 1015 -320
rect 980 -360 985 -335
rect 1010 -360 1015 -335
rect 980 -380 1015 -360
rect 980 -405 985 -380
rect 1010 -405 1015 -380
rect 980 -420 1015 -405
rect 1040 -335 1075 -320
rect 1040 -360 1045 -335
rect 1070 -360 1075 -335
rect 1040 -380 1075 -360
rect 1040 -405 1045 -380
rect 1070 -405 1075 -380
rect 1040 -420 1075 -405
rect 1100 -335 1135 -320
rect 1100 -360 1105 -335
rect 1130 -360 1135 -335
rect 1100 -380 1135 -360
rect 1100 -405 1105 -380
rect 1130 -405 1135 -380
rect 1100 -420 1135 -405
rect 1160 -335 1195 -320
rect 1160 -360 1165 -335
rect 1190 -360 1195 -335
rect 1160 -380 1195 -360
rect 1160 -405 1165 -380
rect 1190 -405 1195 -380
rect 1160 -420 1195 -405
rect 1220 -335 1255 -320
rect 1220 -360 1225 -335
rect 1250 -360 1255 -335
rect 1220 -380 1255 -360
rect 1220 -405 1225 -380
rect 1250 -405 1255 -380
rect 1220 -420 1255 -405
rect 1280 -335 1315 -320
rect 1280 -360 1285 -335
rect 1310 -360 1315 -335
rect 1280 -380 1315 -360
rect 1280 -405 1285 -380
rect 1310 -405 1315 -380
rect 1280 -420 1315 -405
rect 1340 -335 1375 -320
rect 1340 -360 1345 -335
rect 1370 -360 1375 -335
rect 1340 -380 1375 -360
rect 1340 -405 1345 -380
rect 1370 -405 1375 -380
rect 1340 -420 1375 -405
rect 1400 -335 1435 -320
rect 1400 -360 1405 -335
rect 1430 -360 1435 -335
rect 1400 -380 1435 -360
rect 1400 -405 1405 -380
rect 1430 -405 1435 -380
rect 1400 -420 1435 -405
rect 1460 -335 1495 -320
rect 1460 -360 1465 -335
rect 1490 -360 1495 -335
rect 1460 -380 1495 -360
rect 1460 -405 1465 -380
rect 1490 -405 1495 -380
rect 1460 -420 1495 -405
rect 1520 -335 1555 -320
rect 1520 -360 1525 -335
rect 1550 -360 1555 -335
rect 1520 -380 1555 -360
rect 1520 -405 1525 -380
rect 1550 -405 1555 -380
rect 1520 -420 1555 -405
rect 1580 -335 1615 -320
rect 1580 -360 1585 -335
rect 1610 -360 1615 -335
rect 1580 -380 1615 -360
rect 1580 -405 1585 -380
rect 1610 -405 1615 -380
rect 1580 -420 1615 -405
rect 1640 -335 1675 -320
rect 1640 -360 1645 -335
rect 1670 -360 1675 -335
rect 1640 -380 1675 -360
rect 1640 -405 1645 -380
rect 1670 -405 1675 -380
rect 1640 -420 1675 -405
rect 1700 -335 1735 -320
rect 1700 -360 1705 -335
rect 1730 -360 1735 -335
rect 1700 -380 1735 -360
rect 1700 -405 1705 -380
rect 1730 -405 1735 -380
rect 1700 -420 1735 -405
rect 1760 -335 1795 -320
rect 1760 -360 1765 -335
rect 1790 -360 1795 -335
rect 1760 -380 1795 -360
rect 1760 -405 1765 -380
rect 1790 -405 1795 -380
rect 1760 -420 1795 -405
rect 1820 -335 1855 -320
rect 1820 -360 1825 -335
rect 1850 -360 1855 -335
rect 1820 -380 1855 -360
rect 1820 -405 1825 -380
rect 1850 -405 1855 -380
rect 1820 -420 1855 -405
rect 1880 -335 1915 -320
rect 1880 -360 1885 -335
rect 1910 -360 1915 -335
rect 1880 -380 1915 -360
rect 1880 -405 1885 -380
rect 1910 -405 1915 -380
rect 1880 -420 1915 -405
rect 1940 -335 1975 -320
rect 1940 -360 1945 -335
rect 1970 -360 1975 -335
rect 1940 -380 1975 -360
rect 1940 -405 1945 -380
rect 1970 -405 1975 -380
rect 1940 -420 1975 -405
rect 2000 -335 2035 -320
rect 2000 -360 2005 -335
rect 2030 -360 2035 -335
rect 2000 -380 2035 -360
rect 2000 -405 2005 -380
rect 2030 -405 2035 -380
rect 2000 -420 2035 -405
rect 2060 -335 2095 -320
rect 2060 -360 2065 -335
rect 2090 -360 2095 -335
rect 2060 -380 2095 -360
rect 2060 -405 2065 -380
rect 2090 -405 2095 -380
rect 2060 -420 2095 -405
rect 2120 -335 2155 -320
rect 2120 -360 2125 -335
rect 2150 -360 2155 -335
rect 2120 -380 2155 -360
rect 2120 -405 2125 -380
rect 2150 -405 2155 -380
rect 2120 -420 2155 -405
rect 2180 -335 2215 -320
rect 2180 -360 2185 -335
rect 2210 -360 2215 -335
rect 2180 -380 2215 -360
rect 2180 -405 2185 -380
rect 2210 -405 2215 -380
rect 2180 -420 2215 -405
rect 2240 -335 2275 -320
rect 2240 -360 2245 -335
rect 2270 -360 2275 -335
rect 2240 -380 2275 -360
rect 2240 -405 2245 -380
rect 2270 -405 2275 -380
rect 2240 -420 2275 -405
rect 2300 -335 2335 -320
rect 2300 -360 2305 -335
rect 2330 -360 2335 -335
rect 2300 -380 2335 -360
rect 2300 -405 2305 -380
rect 2330 -405 2335 -380
rect 2300 -420 2335 -405
rect 2360 -335 2395 -320
rect 2360 -360 2365 -335
rect 2390 -360 2395 -335
rect 2360 -380 2395 -360
rect 2360 -405 2365 -380
rect 2390 -405 2395 -380
rect 2360 -420 2395 -405
rect 2420 -335 2455 -320
rect 2420 -360 2425 -335
rect 2450 -360 2455 -335
rect 2420 -380 2455 -360
rect 2420 -405 2425 -380
rect 2450 -405 2455 -380
rect 2420 -420 2455 -405
rect 2480 -335 2515 -320
rect 2480 -360 2485 -335
rect 2510 -360 2515 -335
rect 2480 -380 2515 -360
rect 2480 -405 2485 -380
rect 2510 -405 2515 -380
rect 2480 -420 2515 -405
rect 2540 -335 2575 -320
rect 2540 -360 2545 -335
rect 2570 -360 2575 -335
rect 2540 -380 2575 -360
rect 2540 -405 2545 -380
rect 2570 -405 2575 -380
rect 2540 -420 2575 -405
rect 2600 -335 2635 -320
rect 2600 -360 2605 -335
rect 2630 -360 2635 -335
rect 2600 -380 2635 -360
rect 2600 -405 2605 -380
rect 2630 -405 2635 -380
rect 2600 -420 2635 -405
rect 2660 -335 2695 -320
rect 2660 -360 2665 -335
rect 2690 -360 2695 -335
rect 2660 -380 2695 -360
rect 2660 -405 2665 -380
rect 2690 -405 2695 -380
rect 2660 -420 2695 -405
rect 2720 -335 2755 -320
rect 2720 -360 2725 -335
rect 2750 -360 2755 -335
rect 2720 -380 2755 -360
rect 2720 -405 2725 -380
rect 2750 -405 2755 -380
rect 2720 -420 2755 -405
rect 2780 -335 2815 -320
rect 2780 -360 2785 -335
rect 2810 -360 2815 -335
rect 2780 -380 2815 -360
rect 2780 -405 2785 -380
rect 2810 -405 2815 -380
rect 2780 -420 2815 -405
rect 2840 -335 2875 -320
rect 2840 -360 2845 -335
rect 2870 -360 2875 -335
rect 2840 -380 2875 -360
rect 2840 -405 2845 -380
rect 2870 -405 2875 -380
rect 2840 -420 2875 -405
rect 2900 -335 2935 -320
rect 2900 -360 2905 -335
rect 2930 -360 2935 -335
rect 2900 -380 2935 -360
rect 2900 -405 2905 -380
rect 2930 -405 2935 -380
rect 2900 -420 2935 -405
rect 2960 -335 2995 -320
rect 2960 -360 2965 -335
rect 2990 -360 2995 -335
rect 2960 -380 2995 -360
rect 2960 -405 2965 -380
rect 2990 -405 2995 -380
rect 2960 -420 2995 -405
rect 3020 -335 3055 -320
rect 3020 -360 3025 -335
rect 3050 -360 3055 -335
rect 3020 -380 3055 -360
rect 3020 -405 3025 -380
rect 3050 -405 3055 -380
rect 3020 -420 3055 -405
rect 3080 -335 3115 -320
rect 3080 -360 3085 -335
rect 3110 -360 3115 -335
rect 3080 -380 3115 -360
rect 3080 -405 3085 -380
rect 3110 -405 3115 -380
rect 3080 -420 3115 -405
rect 3140 -335 3175 -320
rect 3140 -360 3145 -335
rect 3170 -360 3175 -335
rect 3140 -380 3175 -360
rect 3140 -405 3145 -380
rect 3170 -405 3175 -380
rect 3140 -420 3175 -405
rect 3200 -335 3235 -320
rect 3200 -360 3205 -335
rect 3230 -360 3235 -335
rect 3200 -380 3235 -360
rect 3200 -405 3205 -380
rect 3230 -405 3235 -380
rect 3200 -420 3235 -405
rect 3260 -335 3295 -320
rect 3260 -360 3265 -335
rect 3290 -360 3295 -335
rect 3260 -380 3295 -360
rect 3260 -405 3265 -380
rect 3290 -405 3295 -380
rect 3260 -420 3295 -405
rect 3320 -335 3355 -320
rect 3320 -360 3325 -335
rect 3350 -360 3355 -335
rect 3320 -380 3355 -360
rect 3320 -405 3325 -380
rect 3350 -405 3355 -380
rect 3320 -420 3355 -405
rect 3380 -335 3415 -320
rect 3380 -360 3385 -335
rect 3410 -360 3415 -335
rect 3380 -380 3415 -360
rect 3380 -405 3385 -380
rect 3410 -405 3415 -380
rect 3380 -420 3415 -405
rect 3440 -335 3475 -320
rect 3440 -360 3445 -335
rect 3470 -360 3475 -335
rect 3440 -380 3475 -360
rect 3440 -405 3445 -380
rect 3470 -405 3475 -380
rect 3440 -420 3475 -405
rect 3500 -335 3535 -320
rect 3500 -360 3505 -335
rect 3530 -360 3535 -335
rect 3500 -380 3535 -360
rect 3500 -405 3505 -380
rect 3530 -405 3535 -380
rect 3500 -420 3535 -405
rect 3560 -335 3595 -320
rect 3560 -360 3565 -335
rect 3590 -360 3595 -335
rect 3560 -380 3595 -360
rect 3560 -405 3565 -380
rect 3590 -405 3595 -380
rect 3560 -420 3595 -405
rect 3620 -335 3655 -320
rect 3620 -360 3625 -335
rect 3650 -360 3655 -335
rect 3620 -380 3655 -360
rect 3620 -405 3625 -380
rect 3650 -405 3655 -380
rect 3620 -420 3655 -405
rect 3680 -335 3715 -320
rect 3680 -360 3685 -335
rect 3710 -360 3715 -335
rect 3680 -380 3715 -360
rect 3680 -405 3685 -380
rect 3710 -405 3715 -380
rect 3680 -420 3715 -405
rect 3740 -335 3775 -320
rect 3740 -360 3745 -335
rect 3770 -360 3775 -335
rect 3740 -380 3775 -360
rect 3740 -405 3745 -380
rect 3770 -405 3775 -380
rect 3740 -420 3775 -405
rect 3800 -335 3835 -320
rect 3800 -360 3805 -335
rect 3830 -360 3835 -335
rect 3800 -380 3835 -360
rect 3800 -405 3805 -380
rect 3830 -405 3835 -380
rect 3800 -420 3835 -405
rect 3860 -335 3895 -320
rect 3860 -360 3865 -335
rect 3890 -360 3895 -335
rect 3860 -380 3895 -360
rect 3860 -405 3865 -380
rect 3890 -405 3895 -380
rect 3860 -420 3895 -405
rect 3920 -335 3955 -320
rect 3920 -360 3925 -335
rect 3950 -360 3955 -335
rect 3920 -380 3955 -360
rect 3920 -405 3925 -380
rect 3950 -405 3955 -380
rect 3920 -420 3955 -405
rect 3980 -335 4015 -320
rect 3980 -360 3985 -335
rect 4010 -360 4015 -335
rect 3980 -380 4015 -360
rect 3980 -405 3985 -380
rect 4010 -405 4015 -380
rect 3980 -420 4015 -405
rect 4040 -335 4075 -320
rect 4040 -360 4045 -335
rect 4070 -360 4075 -335
rect 4040 -380 4075 -360
rect 4040 -405 4045 -380
rect 4070 -405 4075 -380
rect 4040 -420 4075 -405
rect 4100 -335 4135 -320
rect 4100 -360 4105 -335
rect 4130 -360 4135 -335
rect 4100 -380 4135 -360
rect 4100 -405 4105 -380
rect 4130 -405 4135 -380
rect 4100 -420 4135 -405
rect 4160 -335 4195 -320
rect 4160 -360 4165 -335
rect 4190 -360 4195 -335
rect 4160 -380 4195 -360
rect 4160 -405 4165 -380
rect 4190 -405 4195 -380
rect 4160 -420 4195 -405
rect 4220 -335 4255 -320
rect 4220 -360 4225 -335
rect 4250 -360 4255 -335
rect 4220 -380 4255 -360
rect 4220 -405 4225 -380
rect 4250 -405 4255 -380
rect 4220 -420 4255 -405
rect 4280 -335 4315 -320
rect 4280 -360 4285 -335
rect 4310 -360 4315 -335
rect 4280 -380 4315 -360
rect 4280 -405 4285 -380
rect 4310 -405 4315 -380
rect 4280 -420 4315 -405
rect 4340 -335 4375 -320
rect 4340 -360 4345 -335
rect 4370 -360 4375 -335
rect 4340 -380 4375 -360
rect 4340 -405 4345 -380
rect 4370 -405 4375 -380
rect 4340 -420 4375 -405
rect 4400 -335 4435 -320
rect 4400 -360 4405 -335
rect 4430 -360 4435 -335
rect 4400 -380 4435 -360
rect 4400 -405 4405 -380
rect 4430 -405 4435 -380
rect 4400 -420 4435 -405
rect 4460 -335 4495 -320
rect 4460 -360 4465 -335
rect 4490 -360 4495 -335
rect 4460 -380 4495 -360
rect 4460 -405 4465 -380
rect 4490 -405 4495 -380
rect 4460 -420 4495 -405
rect 4520 -335 4555 -320
rect 4520 -360 4525 -335
rect 4550 -360 4555 -335
rect 4520 -380 4555 -360
rect 4520 -405 4525 -380
rect 4550 -405 4555 -380
rect 4520 -420 4555 -405
rect 4580 -335 4615 -320
rect 4580 -360 4585 -335
rect 4610 -360 4615 -335
rect 4580 -380 4615 -360
rect 4580 -405 4585 -380
rect 4610 -405 4615 -380
rect 4580 -420 4615 -405
rect 4640 -335 4675 -320
rect 4640 -360 4645 -335
rect 4670 -360 4675 -335
rect 4640 -380 4675 -360
rect 4640 -405 4645 -380
rect 4670 -405 4675 -380
rect 4640 -420 4675 -405
rect 4700 -335 4735 -320
rect 4700 -360 4705 -335
rect 4730 -360 4735 -335
rect 4700 -380 4735 -360
rect 4700 -405 4705 -380
rect 4730 -405 4735 -380
rect 4700 -420 4735 -405
rect 4760 -335 4795 -320
rect 4760 -360 4765 -335
rect 4790 -360 4795 -335
rect 4760 -380 4795 -360
rect 4760 -405 4765 -380
rect 4790 -405 4795 -380
rect 4760 -420 4795 -405
rect 4820 -335 4855 -320
rect 4820 -360 4825 -335
rect 4850 -360 4855 -335
rect 4820 -380 4855 -360
rect 4820 -405 4825 -380
rect 4850 -405 4855 -380
rect 4820 -420 4855 -405
rect 4880 -335 4915 -320
rect 4880 -360 4885 -335
rect 4910 -360 4915 -335
rect 4880 -380 4915 -360
rect 4880 -405 4885 -380
rect 4910 -405 4915 -380
rect 4880 -420 4915 -405
rect 4940 -335 4975 -320
rect 4940 -360 4945 -335
rect 4970 -360 4975 -335
rect 4940 -380 4975 -360
rect 4940 -405 4945 -380
rect 4970 -405 4975 -380
rect 4940 -420 4975 -405
rect 5000 -335 5035 -320
rect 5000 -360 5005 -335
rect 5030 -360 5035 -335
rect 5000 -380 5035 -360
rect 5000 -405 5005 -380
rect 5030 -405 5035 -380
rect 5000 -420 5035 -405
rect 5060 -335 5095 -320
rect 5060 -360 5065 -335
rect 5090 -360 5095 -335
rect 5060 -380 5095 -360
rect 5060 -405 5065 -380
rect 5090 -405 5095 -380
rect 5060 -420 5095 -405
rect 5120 -335 5155 -320
rect 5120 -360 5125 -335
rect 5150 -360 5155 -335
rect 5120 -380 5155 -360
rect 5120 -405 5125 -380
rect 5150 -405 5155 -380
rect 5120 -420 5155 -405
rect 5180 -335 5215 -320
rect 5180 -360 5185 -335
rect 5210 -360 5215 -335
rect 5180 -380 5215 -360
rect 5180 -405 5185 -380
rect 5210 -405 5215 -380
rect 5180 -420 5215 -405
rect 5240 -335 5275 -320
rect 5240 -360 5245 -335
rect 5270 -360 5275 -335
rect 5240 -380 5275 -360
rect 5240 -405 5245 -380
rect 5270 -405 5275 -380
rect 5240 -420 5275 -405
rect 5300 -335 5335 -320
rect 5300 -360 5305 -335
rect 5330 -360 5335 -335
rect 5300 -380 5335 -360
rect 5300 -405 5305 -380
rect 5330 -405 5335 -380
rect 5300 -420 5335 -405
rect 5360 -335 5395 -320
rect 5360 -360 5365 -335
rect 5390 -360 5395 -335
rect 5360 -380 5395 -360
rect 5360 -405 5365 -380
rect 5390 -405 5395 -380
rect 5360 -420 5395 -405
rect 5420 -335 5455 -320
rect 5420 -360 5425 -335
rect 5450 -360 5455 -335
rect 5420 -380 5455 -360
rect 5420 -405 5425 -380
rect 5450 -405 5455 -380
rect 5420 -420 5455 -405
rect 5480 -335 5515 -320
rect 5480 -360 5485 -335
rect 5510 -360 5515 -335
rect 5480 -380 5515 -360
rect 5480 -405 5485 -380
rect 5510 -405 5515 -380
rect 5480 -420 5515 -405
rect 5540 -335 5575 -320
rect 5540 -360 5545 -335
rect 5570 -360 5575 -335
rect 5540 -380 5575 -360
rect 5540 -405 5545 -380
rect 5570 -405 5575 -380
rect 5540 -420 5575 -405
rect 5600 -335 5635 -320
rect 5600 -360 5605 -335
rect 5630 -360 5635 -335
rect 5600 -380 5635 -360
rect 5600 -405 5605 -380
rect 5630 -405 5635 -380
rect 5600 -420 5635 -405
rect 5660 -335 5695 -320
rect 5660 -360 5665 -335
rect 5690 -360 5695 -335
rect 5660 -380 5695 -360
rect 5660 -405 5665 -380
rect 5690 -405 5695 -380
rect 5660 -420 5695 -405
rect 5720 -335 5755 -320
rect 5720 -360 5725 -335
rect 5750 -360 5755 -335
rect 5720 -380 5755 -360
rect 5720 -405 5725 -380
rect 5750 -405 5755 -380
rect 5720 -420 5755 -405
rect 5780 -335 5815 -320
rect 5780 -360 5785 -335
rect 5810 -360 5815 -335
rect 5780 -380 5815 -360
rect 5780 -405 5785 -380
rect 5810 -405 5815 -380
rect 5780 -420 5815 -405
rect 5840 -335 5875 -320
rect 5840 -360 5845 -335
rect 5870 -360 5875 -335
rect 5840 -380 5875 -360
rect 5840 -405 5845 -380
rect 5870 -405 5875 -380
rect 5840 -420 5875 -405
rect 5900 -335 5935 -320
rect 5900 -360 5905 -335
rect 5930 -360 5935 -335
rect 5900 -380 5935 -360
rect 5900 -405 5905 -380
rect 5930 -405 5935 -380
rect 5900 -420 5935 -405
rect 5960 -335 5995 -320
rect 5960 -360 5965 -335
rect 5990 -360 5995 -335
rect 5960 -380 5995 -360
rect 5960 -405 5965 -380
rect 5990 -405 5995 -380
rect 5960 -420 5995 -405
rect 6020 -335 6055 -320
rect 6020 -360 6025 -335
rect 6050 -360 6055 -335
rect 6020 -380 6055 -360
rect 6020 -405 6025 -380
rect 6050 -405 6055 -380
rect 6020 -420 6055 -405
rect 6080 -335 6115 -320
rect 6080 -360 6085 -335
rect 6110 -360 6115 -335
rect 6080 -380 6115 -360
rect 6080 -405 6085 -380
rect 6110 -405 6115 -380
rect 6080 -420 6115 -405
rect 6140 -335 6175 -320
rect 6140 -360 6145 -335
rect 6170 -360 6175 -335
rect 6140 -380 6175 -360
rect 6140 -405 6145 -380
rect 6170 -405 6175 -380
rect 6140 -420 6175 -405
rect 6200 -335 6235 -320
rect 6200 -360 6205 -335
rect 6230 -360 6235 -335
rect 6200 -380 6235 -360
rect 6200 -405 6205 -380
rect 6230 -405 6235 -380
rect 6200 -420 6235 -405
rect 6260 -335 6295 -320
rect 6260 -360 6265 -335
rect 6290 -360 6295 -335
rect 6260 -380 6295 -360
rect 6260 -405 6265 -380
rect 6290 -405 6295 -380
rect 6260 -420 6295 -405
rect 6320 -335 6355 -320
rect 6320 -360 6325 -335
rect 6350 -360 6355 -335
rect 6320 -380 6355 -360
rect 6320 -405 6325 -380
rect 6350 -405 6355 -380
rect 6320 -420 6355 -405
rect 6380 -335 6415 -320
rect 6380 -360 6385 -335
rect 6410 -360 6415 -335
rect 6380 -380 6415 -360
rect 6380 -405 6385 -380
rect 6410 -405 6415 -380
rect 6380 -420 6415 -405
rect 6440 -335 6475 -320
rect 6440 -360 6445 -335
rect 6470 -360 6475 -335
rect 6440 -380 6475 -360
rect 6440 -405 6445 -380
rect 6470 -405 6475 -380
rect 6440 -420 6475 -405
rect 6500 -335 6535 -320
rect 6500 -360 6505 -335
rect 6530 -360 6535 -335
rect 6500 -380 6535 -360
rect 6500 -405 6505 -380
rect 6530 -405 6535 -380
rect 6500 -420 6535 -405
rect 6560 -335 6595 -320
rect 6560 -360 6565 -335
rect 6590 -360 6595 -335
rect 6560 -380 6595 -360
rect 6560 -405 6565 -380
rect 6590 -405 6595 -380
rect 6560 -420 6595 -405
rect 6620 -335 6655 -320
rect 6620 -360 6625 -335
rect 6650 -360 6655 -335
rect 6620 -380 6655 -360
rect 6620 -405 6625 -380
rect 6650 -405 6655 -380
rect 6620 -420 6655 -405
rect 6680 -335 6715 -320
rect 6680 -360 6685 -335
rect 6710 -360 6715 -335
rect 6680 -380 6715 -360
rect 6680 -405 6685 -380
rect 6710 -405 6715 -380
rect 6680 -420 6715 -405
rect 6740 -335 6775 -320
rect 6740 -360 6745 -335
rect 6770 -360 6775 -335
rect 6740 -380 6775 -360
rect 6740 -405 6745 -380
rect 6770 -405 6775 -380
rect 6740 -420 6775 -405
rect 6800 -335 6835 -320
rect 6800 -360 6805 -335
rect 6830 -360 6835 -335
rect 6800 -380 6835 -360
rect 6800 -405 6805 -380
rect 6830 -405 6835 -380
rect 6800 -420 6835 -405
rect 6860 -335 6895 -320
rect 6860 -360 6865 -335
rect 6890 -360 6895 -335
rect 6860 -380 6895 -360
rect 6860 -405 6865 -380
rect 6890 -405 6895 -380
rect 6860 -420 6895 -405
rect 6920 -335 6955 -320
rect 6920 -360 6925 -335
rect 6950 -360 6955 -335
rect 6920 -380 6955 -360
rect 6920 -405 6925 -380
rect 6950 -405 6955 -380
rect 6920 -420 6955 -405
rect 6980 -335 7015 -320
rect 6980 -360 6985 -335
rect 7010 -360 7015 -335
rect 6980 -380 7015 -360
rect 6980 -405 6985 -380
rect 7010 -405 7015 -380
rect 6980 -420 7015 -405
rect 7040 -335 7075 -320
rect 7040 -360 7045 -335
rect 7070 -360 7075 -335
rect 7040 -380 7075 -360
rect 7040 -405 7045 -380
rect 7070 -405 7075 -380
rect 7040 -420 7075 -405
rect 7100 -335 7135 -320
rect 7100 -360 7105 -335
rect 7130 -360 7135 -335
rect 7100 -380 7135 -360
rect 7100 -405 7105 -380
rect 7130 -405 7135 -380
rect 7100 -420 7135 -405
rect 7160 -335 7195 -320
rect 7160 -360 7165 -335
rect 7190 -360 7195 -335
rect 7160 -380 7195 -360
rect 7160 -405 7165 -380
rect 7190 -405 7195 -380
rect 7160 -420 7195 -405
rect 7220 -335 7255 -320
rect 7220 -360 7225 -335
rect 7250 -360 7255 -335
rect 7220 -380 7255 -360
rect 7220 -405 7225 -380
rect 7250 -405 7255 -380
rect 7220 -420 7255 -405
rect 7280 -335 7315 -320
rect 7280 -360 7285 -335
rect 7310 -360 7315 -335
rect 7280 -380 7315 -360
rect 7280 -405 7285 -380
rect 7310 -405 7315 -380
rect 7280 -420 7315 -405
rect 7340 -335 7375 -320
rect 7340 -360 7345 -335
rect 7370 -360 7375 -335
rect 7340 -380 7375 -360
rect 7340 -405 7345 -380
rect 7370 -405 7375 -380
rect 7340 -420 7375 -405
rect 7400 -335 7435 -320
rect 7400 -360 7405 -335
rect 7430 -360 7435 -335
rect 7400 -380 7435 -360
rect 7400 -405 7405 -380
rect 7430 -405 7435 -380
rect 7400 -420 7435 -405
rect 7460 -335 7495 -320
rect 7460 -360 7465 -335
rect 7490 -360 7495 -335
rect 7460 -380 7495 -360
rect 7460 -405 7465 -380
rect 7490 -405 7495 -380
rect 7460 -420 7495 -405
rect 7520 -335 7555 -320
rect 7520 -360 7525 -335
rect 7550 -360 7555 -335
rect 7520 -380 7555 -360
rect 7520 -405 7525 -380
rect 7550 -405 7555 -380
rect 7520 -420 7555 -405
rect 7580 -335 7615 -320
rect 7580 -360 7585 -335
rect 7610 -360 7615 -335
rect 7580 -380 7615 -360
rect 7580 -405 7585 -380
rect 7610 -405 7615 -380
rect 7580 -420 7615 -405
rect 7640 -335 7675 -320
rect 7640 -360 7645 -335
rect 7670 -360 7675 -335
rect 7640 -380 7675 -360
rect 7640 -405 7645 -380
rect 7670 -405 7675 -380
rect 7640 -420 7675 -405
rect 7700 -335 7735 -320
rect 7700 -360 7705 -335
rect 7730 -360 7735 -335
rect 7700 -380 7735 -360
rect 7700 -405 7705 -380
rect 7730 -405 7735 -380
rect 7700 -420 7735 -405
rect 7760 -335 7795 -320
rect 7760 -360 7765 -335
rect 7790 -360 7795 -335
rect 7760 -380 7795 -360
rect 7760 -405 7765 -380
rect 7790 -405 7795 -380
rect 7760 -420 7795 -405
rect 7820 -335 7855 -320
rect 7820 -360 7825 -335
rect 7850 -360 7855 -335
rect 7820 -380 7855 -360
rect 7820 -405 7825 -380
rect 7850 -405 7855 -380
rect 7820 -420 7855 -405
rect 7880 -335 7915 -320
rect 7880 -360 7885 -335
rect 7910 -360 7915 -335
rect 7880 -380 7915 -360
rect 7880 -405 7885 -380
rect 7910 -405 7915 -380
rect 7880 -420 7915 -405
rect 7940 -335 7975 -320
rect 7940 -360 7945 -335
rect 7970 -360 7975 -335
rect 7940 -380 7975 -360
rect 7940 -405 7945 -380
rect 7970 -405 7975 -380
rect 7940 -420 7975 -405
rect 8000 -335 8035 -320
rect 8000 -360 8005 -335
rect 8030 -360 8035 -335
rect 8000 -380 8035 -360
rect 8000 -405 8005 -380
rect 8030 -405 8035 -380
rect 8000 -420 8035 -405
rect 8060 -335 8095 -320
rect 8060 -360 8065 -335
rect 8090 -360 8095 -335
rect 8060 -380 8095 -360
rect 8060 -405 8065 -380
rect 8090 -405 8095 -380
rect 8060 -420 8095 -405
rect 8120 -335 8155 -320
rect 8120 -360 8125 -335
rect 8150 -360 8155 -335
rect 8120 -380 8155 -360
rect 8120 -405 8125 -380
rect 8150 -405 8155 -380
rect 8120 -420 8155 -405
rect 8180 -335 8215 -320
rect 8180 -360 8185 -335
rect 8210 -360 8215 -335
rect 8180 -380 8215 -360
rect 8180 -405 8185 -380
rect 8210 -405 8215 -380
rect 8180 -420 8215 -405
rect 8240 -335 8275 -320
rect 8240 -360 8245 -335
rect 8270 -360 8275 -335
rect 8240 -380 8275 -360
rect 8240 -405 8245 -380
rect 8270 -405 8275 -380
rect 8240 -420 8275 -405
rect 8300 -335 8335 -320
rect 8300 -360 8305 -335
rect 8330 -360 8335 -335
rect 8300 -380 8335 -360
rect 8300 -405 8305 -380
rect 8330 -405 8335 -380
rect 8300 -420 8335 -405
rect 8360 -335 8395 -320
rect 8360 -360 8365 -335
rect 8390 -360 8395 -335
rect 8360 -380 8395 -360
rect 8360 -405 8365 -380
rect 8390 -405 8395 -380
rect 8360 -420 8395 -405
rect 8420 -335 8455 -320
rect 8420 -360 8425 -335
rect 8450 -360 8455 -335
rect 8420 -380 8455 -360
rect 8420 -405 8425 -380
rect 8450 -405 8455 -380
rect 8420 -420 8455 -405
rect 8480 -335 8515 -320
rect 8480 -360 8485 -335
rect 8510 -360 8515 -335
rect 8480 -380 8515 -360
rect 8480 -405 8485 -380
rect 8510 -405 8515 -380
rect 8480 -420 8515 -405
rect 8540 -335 8575 -320
rect 8540 -360 8545 -335
rect 8570 -360 8575 -335
rect 8540 -380 8575 -360
rect 8540 -405 8545 -380
rect 8570 -405 8575 -380
rect 8540 -420 8575 -405
rect 8600 -335 8635 -320
rect 8600 -360 8605 -335
rect 8630 -360 8635 -335
rect 8600 -380 8635 -360
rect 8600 -405 8605 -380
rect 8630 -405 8635 -380
rect 8600 -420 8635 -405
rect 8660 -335 8695 -320
rect 8660 -360 8665 -335
rect 8690 -360 8695 -335
rect 8660 -380 8695 -360
rect 8660 -405 8665 -380
rect 8690 -405 8695 -380
rect 8660 -420 8695 -405
rect 8720 -335 8755 -320
rect 8720 -360 8725 -335
rect 8750 -360 8755 -335
rect 8720 -380 8755 -360
rect 8720 -405 8725 -380
rect 8750 -405 8755 -380
rect 8720 -420 8755 -405
rect 8780 -335 8815 -320
rect 8780 -360 8785 -335
rect 8810 -360 8815 -335
rect 8780 -380 8815 -360
rect 8780 -405 8785 -380
rect 8810 -405 8815 -380
rect 8780 -420 8815 -405
rect 8840 -335 8875 -320
rect 8840 -360 8845 -335
rect 8870 -360 8875 -335
rect 8840 -380 8875 -360
rect 8840 -405 8845 -380
rect 8870 -405 8875 -380
rect 8840 -420 8875 -405
rect 8900 -335 8935 -320
rect 8900 -360 8905 -335
rect 8930 -360 8935 -335
rect 8900 -380 8935 -360
rect 8900 -405 8905 -380
rect 8930 -405 8935 -380
rect 8900 -420 8935 -405
rect 8960 -335 8995 -320
rect 8960 -360 8965 -335
rect 8990 -360 8995 -335
rect 8960 -380 8995 -360
rect 8960 -405 8965 -380
rect 8990 -405 8995 -380
rect 8960 -420 8995 -405
rect 9020 -335 9055 -320
rect 9020 -360 9025 -335
rect 9050 -360 9055 -335
rect 9020 -380 9055 -360
rect 9020 -405 9025 -380
rect 9050 -405 9055 -380
rect 9020 -420 9055 -405
rect 9080 -335 9115 -320
rect 9080 -360 9085 -335
rect 9110 -360 9115 -335
rect 9080 -380 9115 -360
rect 9080 -405 9085 -380
rect 9110 -405 9115 -380
rect 9080 -420 9115 -405
rect 9140 -335 9175 -320
rect 9140 -360 9145 -335
rect 9170 -360 9175 -335
rect 9140 -380 9175 -360
rect 9140 -405 9145 -380
rect 9170 -405 9175 -380
rect 9140 -420 9175 -405
rect 9200 -335 9235 -320
rect 9200 -360 9205 -335
rect 9230 -360 9235 -335
rect 9200 -380 9235 -360
rect 9200 -405 9205 -380
rect 9230 -405 9235 -380
rect 9200 -420 9235 -405
rect 9260 -335 9295 -320
rect 9260 -360 9265 -335
rect 9290 -360 9295 -335
rect 9260 -380 9295 -360
rect 9260 -405 9265 -380
rect 9290 -405 9295 -380
rect 9260 -420 9295 -405
rect 9320 -335 9355 -320
rect 9320 -360 9325 -335
rect 9350 -360 9355 -335
rect 9320 -380 9355 -360
rect 9320 -405 9325 -380
rect 9350 -405 9355 -380
rect 9320 -420 9355 -405
rect 9380 -335 9415 -320
rect 9380 -360 9385 -335
rect 9410 -360 9415 -335
rect 9380 -380 9415 -360
rect 9380 -405 9385 -380
rect 9410 -405 9415 -380
rect 9380 -420 9415 -405
rect 9440 -335 9475 -320
rect 9440 -360 9445 -335
rect 9470 -360 9475 -335
rect 9440 -380 9475 -360
rect 9440 -405 9445 -380
rect 9470 -405 9475 -380
rect 9440 -420 9475 -405
rect 9500 -335 9535 -320
rect 9500 -360 9505 -335
rect 9530 -360 9535 -335
rect 9500 -380 9535 -360
rect 9500 -405 9505 -380
rect 9530 -405 9535 -380
rect 9500 -420 9535 -405
rect 9560 -335 9595 -320
rect 9560 -360 9565 -335
rect 9590 -360 9595 -335
rect 9560 -380 9595 -360
rect 9560 -405 9565 -380
rect 9590 -405 9595 -380
rect 9560 -420 9595 -405
rect 9620 -335 9655 -320
rect 9620 -360 9625 -335
rect 9650 -360 9655 -335
rect 9620 -380 9655 -360
rect 9620 -405 9625 -380
rect 9650 -405 9655 -380
rect 9620 -420 9655 -405
rect 9680 -335 9715 -320
rect 9680 -360 9685 -335
rect 9710 -360 9715 -335
rect 9680 -380 9715 -360
rect 9680 -405 9685 -380
rect 9710 -405 9715 -380
rect 9680 -420 9715 -405
rect 9740 -335 9775 -320
rect 9740 -360 9745 -335
rect 9770 -360 9775 -335
rect 9740 -380 9775 -360
rect 9740 -405 9745 -380
rect 9770 -405 9775 -380
rect 9740 -420 9775 -405
rect 9800 -335 9835 -320
rect 9800 -360 9805 -335
rect 9830 -360 9835 -335
rect 9800 -380 9835 -360
rect 9800 -405 9805 -380
rect 9830 -405 9835 -380
rect 9800 -420 9835 -405
rect 9860 -335 9895 -320
rect 9860 -360 9865 -335
rect 9890 -360 9895 -335
rect 9860 -380 9895 -360
rect 9860 -405 9865 -380
rect 9890 -405 9895 -380
rect 9860 -420 9895 -405
rect 9920 -335 9955 -320
rect 9920 -360 9925 -335
rect 9950 -360 9955 -335
rect 9920 -380 9955 -360
rect 9920 -405 9925 -380
rect 9950 -405 9955 -380
rect 9920 -420 9955 -405
rect 9980 -335 10015 -320
rect 9980 -360 9985 -335
rect 10010 -360 10015 -335
rect 9980 -380 10015 -360
rect 9980 -405 9985 -380
rect 10010 -405 10015 -380
rect 9980 -420 10015 -405
rect 10040 -335 10075 -320
rect 10040 -360 10045 -335
rect 10070 -360 10075 -335
rect 10040 -380 10075 -360
rect 10040 -405 10045 -380
rect 10070 -405 10075 -380
rect 10040 -420 10075 -405
rect 10100 -335 10135 -320
rect 10100 -360 10105 -335
rect 10130 -360 10135 -335
rect 10100 -380 10135 -360
rect 10100 -405 10105 -380
rect 10130 -405 10135 -380
rect 10100 -420 10135 -405
rect 10160 -335 10195 -320
rect 10160 -360 10165 -335
rect 10190 -360 10195 -335
rect 10160 -380 10195 -360
rect 10160 -405 10165 -380
rect 10190 -405 10195 -380
rect 10160 -420 10195 -405
rect 10220 -335 10255 -320
rect 10220 -360 10225 -335
rect 10250 -360 10255 -335
rect 10220 -380 10255 -360
rect 10220 -405 10225 -380
rect 10250 -405 10255 -380
rect 10220 -420 10255 -405
rect 10280 -335 10315 -320
rect 10280 -360 10285 -335
rect 10310 -360 10315 -335
rect 10280 -380 10315 -360
rect 10280 -405 10285 -380
rect 10310 -405 10315 -380
rect 10280 -420 10315 -405
rect 10340 -335 10375 -320
rect 10340 -360 10345 -335
rect 10370 -360 10375 -335
rect 10340 -380 10375 -360
rect 10340 -405 10345 -380
rect 10370 -405 10375 -380
rect 10340 -420 10375 -405
rect 10400 -335 10435 -320
rect 10400 -360 10405 -335
rect 10430 -360 10435 -335
rect 10400 -380 10435 -360
rect 10400 -405 10405 -380
rect 10430 -405 10435 -380
rect 10400 -420 10435 -405
rect 10460 -335 10495 -320
rect 10460 -360 10465 -335
rect 10490 -360 10495 -335
rect 10460 -380 10495 -360
rect 10460 -405 10465 -380
rect 10490 -405 10495 -380
rect 10460 -420 10495 -405
rect 10520 -335 10555 -320
rect 10520 -360 10525 -335
rect 10550 -360 10555 -335
rect 10520 -380 10555 -360
rect 10520 -405 10525 -380
rect 10550 -405 10555 -380
rect 10520 -420 10555 -405
rect 10580 -335 10615 -320
rect 10580 -360 10585 -335
rect 10610 -360 10615 -335
rect 10580 -380 10615 -360
rect 10580 -405 10585 -380
rect 10610 -405 10615 -380
rect 10580 -420 10615 -405
rect 10640 -335 10675 -320
rect 10640 -360 10645 -335
rect 10670 -360 10675 -335
rect 10640 -380 10675 -360
rect 10640 -405 10645 -380
rect 10670 -405 10675 -380
rect 10640 -420 10675 -405
rect 10700 -335 10735 -320
rect 10700 -360 10705 -335
rect 10730 -360 10735 -335
rect 10700 -380 10735 -360
rect 10700 -405 10705 -380
rect 10730 -405 10735 -380
rect 10700 -420 10735 -405
rect 10760 -335 10795 -320
rect 10760 -360 10765 -335
rect 10790 -360 10795 -335
rect 10760 -380 10795 -360
rect 10760 -405 10765 -380
rect 10790 -405 10795 -380
rect 10760 -420 10795 -405
rect 10820 -335 10855 -320
rect 10820 -360 10825 -335
rect 10850 -360 10855 -335
rect 10820 -380 10855 -360
rect 10820 -405 10825 -380
rect 10850 -405 10855 -380
rect 10820 -420 10855 -405
rect 10880 -335 10915 -320
rect 10880 -360 10885 -335
rect 10910 -360 10915 -335
rect 10880 -380 10915 -360
rect 10880 -405 10885 -380
rect 10910 -405 10915 -380
rect 10880 -420 10915 -405
rect 10940 -335 10975 -320
rect 10940 -360 10945 -335
rect 10970 -360 10975 -335
rect 10940 -380 10975 -360
rect 10940 -405 10945 -380
rect 10970 -405 10975 -380
rect 10940 -420 10975 -405
rect 11000 -335 11035 -320
rect 11000 -360 11005 -335
rect 11030 -360 11035 -335
rect 11000 -380 11035 -360
rect 11000 -405 11005 -380
rect 11030 -405 11035 -380
rect 11000 -420 11035 -405
rect 11060 -335 11095 -320
rect 11060 -360 11065 -335
rect 11090 -360 11095 -335
rect 11060 -380 11095 -360
rect 11060 -405 11065 -380
rect 11090 -405 11095 -380
rect 11060 -420 11095 -405
rect 11120 -335 11155 -320
rect 11120 -360 11125 -335
rect 11150 -360 11155 -335
rect 11120 -380 11155 -360
rect 11120 -405 11125 -380
rect 11150 -405 11155 -380
rect 11120 -420 11155 -405
rect 11180 -335 11215 -320
rect 11180 -360 11185 -335
rect 11210 -360 11215 -335
rect 11180 -380 11215 -360
rect 11180 -405 11185 -380
rect 11210 -405 11215 -380
rect 11180 -420 11215 -405
rect 11240 -335 11275 -320
rect 11240 -360 11245 -335
rect 11270 -360 11275 -335
rect 11240 -380 11275 -360
rect 11240 -405 11245 -380
rect 11270 -405 11275 -380
rect 11240 -420 11275 -405
rect 11300 -335 11335 -320
rect 11300 -360 11305 -335
rect 11330 -360 11335 -335
rect 11300 -380 11335 -360
rect 11300 -405 11305 -380
rect 11330 -405 11335 -380
rect 11300 -420 11335 -405
rect 11360 -335 11395 -320
rect 11360 -360 11365 -335
rect 11390 -360 11395 -335
rect 11360 -380 11395 -360
rect 11360 -405 11365 -380
rect 11390 -405 11395 -380
rect 11360 -420 11395 -405
rect 11420 -335 11455 -320
rect 11420 -360 11425 -335
rect 11450 -360 11455 -335
rect 11420 -380 11455 -360
rect 11420 -405 11425 -380
rect 11450 -405 11455 -380
rect 11420 -420 11455 -405
rect 11480 -335 11515 -320
rect 11480 -360 11485 -335
rect 11510 -360 11515 -335
rect 11480 -380 11515 -360
rect 11480 -405 11485 -380
rect 11510 -405 11515 -380
rect 11480 -420 11515 -405
rect 11540 -335 11575 -320
rect 11540 -360 11545 -335
rect 11570 -360 11575 -335
rect 11540 -380 11575 -360
rect 11540 -405 11545 -380
rect 11570 -405 11575 -380
rect 11540 -420 11575 -405
rect 11600 -335 11635 -320
rect 11600 -360 11605 -335
rect 11630 -360 11635 -335
rect 11600 -380 11635 -360
rect 11600 -405 11605 -380
rect 11630 -405 11635 -380
rect 11600 -420 11635 -405
rect 11660 -335 11695 -320
rect 11660 -360 11665 -335
rect 11690 -360 11695 -335
rect 11660 -380 11695 -360
rect 11660 -405 11665 -380
rect 11690 -405 11695 -380
rect 11660 -420 11695 -405
rect 11720 -335 11755 -320
rect 11720 -360 11725 -335
rect 11750 -360 11755 -335
rect 11720 -380 11755 -360
rect 11720 -405 11725 -380
rect 11750 -405 11755 -380
rect 11720 -420 11755 -405
rect 11780 -335 11815 -320
rect 11780 -360 11785 -335
rect 11810 -360 11815 -335
rect 11780 -380 11815 -360
rect 11780 -405 11785 -380
rect 11810 -405 11815 -380
rect 11780 -420 11815 -405
rect 11840 -335 11875 -320
rect 11840 -360 11845 -335
rect 11870 -360 11875 -335
rect 11840 -380 11875 -360
rect 11840 -405 11845 -380
rect 11870 -405 11875 -380
rect 11840 -420 11875 -405
rect 11900 -335 11935 -320
rect 11900 -360 11905 -335
rect 11930 -360 11935 -335
rect 11900 -380 11935 -360
rect 11900 -405 11905 -380
rect 11930 -405 11935 -380
rect 11900 -420 11935 -405
rect 11960 -335 11995 -320
rect 11960 -360 11965 -335
rect 11990 -360 11995 -335
rect 11960 -380 11995 -360
rect 11960 -405 11965 -380
rect 11990 -405 11995 -380
rect 11960 -420 11995 -405
rect 12020 -335 12055 -320
rect 12020 -360 12025 -335
rect 12050 -360 12055 -335
rect 12020 -380 12055 -360
rect 12020 -405 12025 -380
rect 12050 -405 12055 -380
rect 12020 -420 12055 -405
rect 12080 -335 12115 -320
rect 12080 -360 12085 -335
rect 12110 -360 12115 -335
rect 12080 -380 12115 -360
rect 12080 -405 12085 -380
rect 12110 -405 12115 -380
rect 12080 -420 12115 -405
rect 12140 -335 12175 -320
rect 12140 -360 12145 -335
rect 12170 -360 12175 -335
rect 12140 -380 12175 -360
rect 12140 -405 12145 -380
rect 12170 -405 12175 -380
rect 12140 -420 12175 -405
rect 12200 -335 12235 -320
rect 12200 -360 12205 -335
rect 12230 -360 12235 -335
rect 12200 -380 12235 -360
rect 12200 -405 12205 -380
rect 12230 -405 12235 -380
rect 12200 -420 12235 -405
rect 12260 -335 12295 -320
rect 12260 -360 12265 -335
rect 12290 -360 12295 -335
rect 12260 -380 12295 -360
rect 12260 -405 12265 -380
rect 12290 -405 12295 -380
rect 12260 -420 12295 -405
rect 12320 -335 12355 -320
rect 12320 -360 12325 -335
rect 12350 -360 12355 -335
rect 12320 -380 12355 -360
rect 12320 -405 12325 -380
rect 12350 -405 12355 -380
rect 12320 -420 12355 -405
rect 12380 -335 12415 -320
rect 12380 -360 12385 -335
rect 12410 -360 12415 -335
rect 12380 -380 12415 -360
rect 12380 -405 12385 -380
rect 12410 -405 12415 -380
rect 12380 -420 12415 -405
rect 12440 -335 12475 -320
rect 12440 -360 12445 -335
rect 12470 -360 12475 -335
rect 12440 -380 12475 -360
rect 12440 -405 12445 -380
rect 12470 -405 12475 -380
rect 12440 -420 12475 -405
rect 12500 -335 12535 -320
rect 12500 -360 12505 -335
rect 12530 -360 12535 -335
rect 12500 -380 12535 -360
rect 12500 -405 12505 -380
rect 12530 -405 12535 -380
rect 12500 -420 12535 -405
rect 12560 -335 12595 -320
rect 12560 -360 12565 -335
rect 12590 -360 12595 -335
rect 12560 -380 12595 -360
rect 12560 -405 12565 -380
rect 12590 -405 12595 -380
rect 12560 -420 12595 -405
rect 12620 -335 12655 -320
rect 12620 -360 12625 -335
rect 12650 -360 12655 -335
rect 12620 -380 12655 -360
rect 12620 -405 12625 -380
rect 12650 -405 12655 -380
rect 12620 -420 12655 -405
rect 12680 -335 12715 -320
rect 12680 -360 12685 -335
rect 12710 -360 12715 -335
rect 12680 -380 12715 -360
rect 12680 -405 12685 -380
rect 12710 -405 12715 -380
rect 12680 -420 12715 -405
rect 12740 -335 12775 -320
rect 12740 -360 12745 -335
rect 12770 -360 12775 -335
rect 12740 -380 12775 -360
rect 12740 -405 12745 -380
rect 12770 -405 12775 -380
rect 12740 -420 12775 -405
rect 12800 -335 12835 -320
rect 12800 -360 12805 -335
rect 12830 -360 12835 -335
rect 12800 -380 12835 -360
rect 12800 -405 12805 -380
rect 12830 -405 12835 -380
rect 12800 -420 12835 -405
rect 12860 -335 12895 -320
rect 12860 -360 12865 -335
rect 12890 -360 12895 -335
rect 12860 -380 12895 -360
rect 12860 -405 12865 -380
rect 12890 -405 12895 -380
rect 12860 -420 12895 -405
rect 12920 -335 12955 -320
rect 12920 -360 12925 -335
rect 12950 -360 12955 -335
rect 12920 -380 12955 -360
rect 12920 -405 12925 -380
rect 12950 -405 12955 -380
rect 12920 -420 12955 -405
rect 12980 -335 13015 -320
rect 12980 -360 12985 -335
rect 13010 -360 13015 -335
rect 12980 -380 13015 -360
rect 12980 -405 12985 -380
rect 13010 -405 13015 -380
rect 12980 -420 13015 -405
rect 13040 -335 13075 -320
rect 13040 -360 13045 -335
rect 13070 -360 13075 -335
rect 13040 -380 13075 -360
rect 13040 -405 13045 -380
rect 13070 -405 13075 -380
rect 13040 -420 13075 -405
rect 13100 -335 13135 -320
rect 13100 -360 13105 -335
rect 13130 -360 13135 -335
rect 13100 -380 13135 -360
rect 13100 -405 13105 -380
rect 13130 -405 13135 -380
rect 13100 -420 13135 -405
rect 13160 -335 13195 -320
rect 13160 -360 13165 -335
rect 13190 -360 13195 -335
rect 13160 -380 13195 -360
rect 13160 -405 13165 -380
rect 13190 -405 13195 -380
rect 13160 -420 13195 -405
rect 13220 -335 13255 -320
rect 13220 -360 13225 -335
rect 13250 -360 13255 -335
rect 13220 -380 13255 -360
rect 13220 -405 13225 -380
rect 13250 -405 13255 -380
rect 13220 -420 13255 -405
rect 13280 -335 13315 -320
rect 13280 -360 13285 -335
rect 13310 -360 13315 -335
rect 13280 -380 13315 -360
rect 13280 -405 13285 -380
rect 13310 -405 13315 -380
rect 13280 -420 13315 -405
rect 13340 -335 13375 -320
rect 13340 -360 13345 -335
rect 13370 -360 13375 -335
rect 13340 -380 13375 -360
rect 13340 -405 13345 -380
rect 13370 -405 13375 -380
rect 13340 -420 13375 -405
rect 13400 -335 13435 -320
rect 13400 -360 13405 -335
rect 13430 -360 13435 -335
rect 13400 -380 13435 -360
rect 13400 -405 13405 -380
rect 13430 -405 13435 -380
rect 13400 -420 13435 -405
rect 13460 -335 13495 -320
rect 13460 -360 13465 -335
rect 13490 -360 13495 -335
rect 13460 -380 13495 -360
rect 13460 -405 13465 -380
rect 13490 -405 13495 -380
rect 13460 -420 13495 -405
rect 13520 -335 13555 -320
rect 13520 -360 13525 -335
rect 13550 -360 13555 -335
rect 13520 -380 13555 -360
rect 13520 -405 13525 -380
rect 13550 -405 13555 -380
rect 13520 -420 13555 -405
rect 13580 -335 13615 -320
rect 13580 -360 13585 -335
rect 13610 -360 13615 -335
rect 13580 -380 13615 -360
rect 13580 -405 13585 -380
rect 13610 -405 13615 -380
rect 13580 -420 13615 -405
rect 13640 -335 13675 -320
rect 13640 -360 13645 -335
rect 13670 -360 13675 -335
rect 13640 -380 13675 -360
rect 13640 -405 13645 -380
rect 13670 -405 13675 -380
rect 13640 -420 13675 -405
rect 13700 -335 13735 -320
rect 13700 -360 13705 -335
rect 13730 -360 13735 -335
rect 13700 -380 13735 -360
rect 13700 -405 13705 -380
rect 13730 -405 13735 -380
rect 13700 -420 13735 -405
rect 13760 -335 13795 -320
rect 13760 -360 13765 -335
rect 13790 -360 13795 -335
rect 13760 -380 13795 -360
rect 13760 -405 13765 -380
rect 13790 -405 13795 -380
rect 13760 -420 13795 -405
rect 13820 -335 13855 -320
rect 13820 -360 13825 -335
rect 13850 -360 13855 -335
rect 13820 -380 13855 -360
rect 13820 -405 13825 -380
rect 13850 -405 13855 -380
rect 13820 -420 13855 -405
rect 13880 -335 13915 -320
rect 13880 -360 13885 -335
rect 13910 -360 13915 -335
rect 13880 -380 13915 -360
rect 13880 -405 13885 -380
rect 13910 -405 13915 -380
rect 13880 -420 13915 -405
rect 13940 -335 13975 -320
rect 13940 -360 13945 -335
rect 13970 -360 13975 -335
rect 13940 -380 13975 -360
rect 13940 -405 13945 -380
rect 13970 -405 13975 -380
rect 13940 -420 13975 -405
rect 14000 -335 14035 -320
rect 14000 -360 14005 -335
rect 14030 -360 14035 -335
rect 14000 -380 14035 -360
rect 14000 -405 14005 -380
rect 14030 -405 14035 -380
rect 14000 -420 14035 -405
rect 14060 -335 14095 -320
rect 14060 -360 14065 -335
rect 14090 -360 14095 -335
rect 14060 -380 14095 -360
rect 14060 -405 14065 -380
rect 14090 -405 14095 -380
rect 14060 -420 14095 -405
rect 14120 -335 14155 -320
rect 14120 -360 14125 -335
rect 14150 -360 14155 -335
rect 14120 -380 14155 -360
rect 14120 -405 14125 -380
rect 14150 -405 14155 -380
rect 14120 -420 14155 -405
rect 14180 -335 14215 -320
rect 14180 -360 14185 -335
rect 14210 -360 14215 -335
rect 14180 -380 14215 -360
rect 14180 -405 14185 -380
rect 14210 -405 14215 -380
rect 14180 -420 14215 -405
rect 14240 -335 14275 -320
rect 14240 -360 14245 -335
rect 14270 -360 14275 -335
rect 14240 -380 14275 -360
rect 14240 -405 14245 -380
rect 14270 -405 14275 -380
rect 14240 -420 14275 -405
rect 14300 -335 14335 -320
rect 14300 -360 14305 -335
rect 14330 -360 14335 -335
rect 14300 -380 14335 -360
rect 14300 -405 14305 -380
rect 14330 -405 14335 -380
rect 14300 -420 14335 -405
rect 14360 -335 14395 -320
rect 14360 -360 14365 -335
rect 14390 -360 14395 -335
rect 14360 -380 14395 -360
rect 14360 -405 14365 -380
rect 14390 -405 14395 -380
rect 14360 -420 14395 -405
rect 14420 -335 14455 -320
rect 14420 -360 14425 -335
rect 14450 -360 14455 -335
rect 14420 -380 14455 -360
rect 14420 -405 14425 -380
rect 14450 -405 14455 -380
rect 14420 -420 14455 -405
rect 14480 -335 14515 -320
rect 14480 -360 14485 -335
rect 14510 -360 14515 -335
rect 14480 -380 14515 -360
rect 14480 -405 14485 -380
rect 14510 -405 14515 -380
rect 14480 -420 14515 -405
rect 14540 -335 14575 -320
rect 14540 -360 14545 -335
rect 14570 -360 14575 -335
rect 14540 -380 14575 -360
rect 14540 -405 14545 -380
rect 14570 -405 14575 -380
rect 14540 -420 14575 -405
rect 14600 -335 14635 -320
rect 14600 -360 14605 -335
rect 14630 -360 14635 -335
rect 14600 -380 14635 -360
rect 14600 -405 14605 -380
rect 14630 -405 14635 -380
rect 14600 -420 14635 -405
rect 14660 -335 14695 -320
rect 14660 -360 14665 -335
rect 14690 -360 14695 -335
rect 14660 -380 14695 -360
rect 14660 -405 14665 -380
rect 14690 -405 14695 -380
rect 14660 -420 14695 -405
rect 14720 -335 14755 -320
rect 14720 -360 14725 -335
rect 14750 -360 14755 -335
rect 14720 -380 14755 -360
rect 14720 -405 14725 -380
rect 14750 -405 14755 -380
rect 14720 -420 14755 -405
rect 14780 -335 14815 -320
rect 14780 -360 14785 -335
rect 14810 -360 14815 -335
rect 14780 -380 14815 -360
rect 14780 -405 14785 -380
rect 14810 -405 14815 -380
rect 14780 -420 14815 -405
rect 14840 -335 14875 -320
rect 14840 -360 14845 -335
rect 14870 -360 14875 -335
rect 14840 -380 14875 -360
rect 14840 -405 14845 -380
rect 14870 -405 14875 -380
rect 14840 -420 14875 -405
rect 14900 -335 14935 -320
rect 14900 -360 14905 -335
rect 14930 -360 14935 -335
rect 14900 -380 14935 -360
rect 14900 -405 14905 -380
rect 14930 -405 14935 -380
rect 14900 -420 14935 -405
rect 14960 -335 14995 -320
rect 14960 -360 14965 -335
rect 14990 -360 14995 -335
rect 14960 -380 14995 -360
rect 14960 -405 14965 -380
rect 14990 -405 14995 -380
rect 14960 -420 14995 -405
rect 15020 -335 15055 -320
rect 15020 -360 15025 -335
rect 15050 -360 15055 -335
rect 15020 -380 15055 -360
rect 15020 -405 15025 -380
rect 15050 -405 15055 -380
rect 15020 -420 15055 -405
rect 15080 -335 15115 -320
rect 15080 -360 15085 -335
rect 15110 -360 15115 -335
rect 15080 -380 15115 -360
rect 15080 -405 15085 -380
rect 15110 -405 15115 -380
rect 15080 -420 15115 -405
rect 15140 -335 15175 -320
rect 15140 -360 15145 -335
rect 15170 -360 15175 -335
rect 15140 -380 15175 -360
rect 15140 -405 15145 -380
rect 15170 -405 15175 -380
rect 15140 -420 15175 -405
rect 15200 -335 15235 -320
rect 15200 -360 15205 -335
rect 15230 -360 15235 -335
rect 15200 -380 15235 -360
rect 15200 -405 15205 -380
rect 15230 -405 15235 -380
rect 15200 -420 15235 -405
rect 15260 -335 15295 -320
rect 15260 -360 15265 -335
rect 15290 -360 15295 -335
rect 15260 -380 15295 -360
rect 15260 -405 15265 -380
rect 15290 -405 15295 -380
rect 15260 -420 15295 -405
rect 15320 -335 15355 -320
rect 15320 -360 15325 -335
rect 15350 -360 15355 -335
rect 15320 -380 15355 -360
rect 15320 -405 15325 -380
rect 15350 -405 15355 -380
rect 15320 -420 15355 -405
rect 15380 -335 15415 -320
rect 15380 -360 15385 -335
rect 15410 -360 15415 -335
rect 15380 -380 15415 -360
rect 15380 -405 15385 -380
rect 15410 -405 15415 -380
rect 15380 -420 15415 -405
rect 15440 -335 15475 -320
rect 15440 -360 15445 -335
rect 15470 -360 15475 -335
rect 15440 -380 15475 -360
rect 15440 -405 15445 -380
rect 15470 -405 15475 -380
rect 15440 -420 15475 -405
rect 15500 -335 15535 -320
rect 15500 -360 15505 -335
rect 15530 -360 15535 -335
rect 15500 -380 15535 -360
rect 15500 -405 15505 -380
rect 15530 -405 15535 -380
rect 15500 -420 15535 -405
rect 15560 -335 15595 -320
rect 15560 -360 15565 -335
rect 15590 -360 15595 -335
rect 15560 -380 15595 -360
rect 15560 -405 15565 -380
rect 15590 -405 15595 -380
rect 15560 -420 15595 -405
rect 15620 -335 15655 -320
rect 15620 -360 15625 -335
rect 15650 -360 15655 -335
rect 15620 -380 15655 -360
rect 15620 -405 15625 -380
rect 15650 -405 15655 -380
rect 15620 -420 15655 -405
rect 15680 -335 15715 -320
rect 15680 -360 15685 -335
rect 15710 -360 15715 -335
rect 15680 -380 15715 -360
rect 15680 -405 15685 -380
rect 15710 -405 15715 -380
rect 15680 -420 15715 -405
rect 15740 -335 15775 -320
rect 15740 -360 15745 -335
rect 15770 -360 15775 -335
rect 15740 -380 15775 -360
rect 15740 -405 15745 -380
rect 15770 -405 15775 -380
rect 15740 -420 15775 -405
rect 15800 -335 15835 -320
rect 15800 -360 15805 -335
rect 15830 -360 15835 -335
rect 15800 -380 15835 -360
rect 15800 -405 15805 -380
rect 15830 -405 15835 -380
rect 15800 -420 15835 -405
rect 15860 -335 15895 -320
rect 15860 -360 15865 -335
rect 15890 -360 15895 -335
rect 15860 -380 15895 -360
rect 15860 -405 15865 -380
rect 15890 -405 15895 -380
rect 15860 -420 15895 -405
rect 15920 -335 15955 -320
rect 15920 -360 15925 -335
rect 15950 -360 15955 -335
rect 15920 -380 15955 -360
rect 15920 -405 15925 -380
rect 15950 -405 15955 -380
rect 15920 -420 15955 -405
rect 15980 -335 16015 -320
rect 15980 -360 15985 -335
rect 16010 -360 16015 -335
rect 15980 -380 16015 -360
rect 15980 -405 15985 -380
rect 16010 -405 16015 -380
rect 15980 -420 16015 -405
rect 16040 -335 16075 -320
rect 16040 -360 16045 -335
rect 16070 -360 16075 -335
rect 16040 -380 16075 -360
rect 16040 -405 16045 -380
rect 16070 -405 16075 -380
rect 16040 -420 16075 -405
rect 16100 -335 16135 -320
rect 16100 -360 16105 -335
rect 16130 -360 16135 -335
rect 16100 -380 16135 -360
rect 16100 -405 16105 -380
rect 16130 -405 16135 -380
rect 16100 -420 16135 -405
rect 16160 -335 16195 -320
rect 16160 -360 16165 -335
rect 16190 -360 16195 -335
rect 16160 -380 16195 -360
rect 16160 -405 16165 -380
rect 16190 -405 16195 -380
rect 16160 -420 16195 -405
rect 16220 -335 16255 -320
rect 16220 -360 16225 -335
rect 16250 -360 16255 -335
rect 16220 -380 16255 -360
rect 16220 -405 16225 -380
rect 16250 -405 16255 -380
rect 16220 -420 16255 -405
rect 16280 -335 16315 -320
rect 16280 -360 16285 -335
rect 16310 -360 16315 -335
rect 16280 -380 16315 -360
rect 16280 -405 16285 -380
rect 16310 -405 16315 -380
rect 16280 -420 16315 -405
rect 16340 -335 16375 -320
rect 16340 -360 16345 -335
rect 16370 -360 16375 -335
rect 16340 -380 16375 -360
rect 16340 -405 16345 -380
rect 16370 -405 16375 -380
rect 16340 -420 16375 -405
rect 16400 -335 16435 -320
rect 16400 -360 16405 -335
rect 16430 -360 16435 -335
rect 16400 -380 16435 -360
rect 16400 -405 16405 -380
rect 16430 -405 16435 -380
rect 16400 -420 16435 -405
rect 16460 -335 16495 -320
rect 16460 -360 16465 -335
rect 16490 -360 16495 -335
rect 16460 -380 16495 -360
rect 16460 -405 16465 -380
rect 16490 -405 16495 -380
rect 16460 -420 16495 -405
rect 16520 -335 16555 -320
rect 16520 -360 16525 -335
rect 16550 -360 16555 -335
rect 16520 -380 16555 -360
rect 16520 -405 16525 -380
rect 16550 -405 16555 -380
rect 16520 -420 16555 -405
rect 16580 -335 16615 -320
rect 16580 -360 16585 -335
rect 16610 -360 16615 -335
rect 16580 -380 16615 -360
rect 16580 -405 16585 -380
rect 16610 -405 16615 -380
rect 16580 -420 16615 -405
rect 16640 -335 16675 -320
rect 16640 -360 16645 -335
rect 16670 -360 16675 -335
rect 16640 -380 16675 -360
rect 16640 -405 16645 -380
rect 16670 -405 16675 -380
rect 16640 -420 16675 -405
rect 16700 -335 16735 -320
rect 16700 -360 16705 -335
rect 16730 -360 16735 -335
rect 16700 -380 16735 -360
rect 16700 -405 16705 -380
rect 16730 -405 16735 -380
rect 16700 -420 16735 -405
rect 16760 -335 16795 -320
rect 16760 -360 16765 -335
rect 16790 -360 16795 -335
rect 16760 -380 16795 -360
rect 16760 -405 16765 -380
rect 16790 -405 16795 -380
rect 16760 -420 16795 -405
rect 16820 -335 16855 -320
rect 16820 -360 16825 -335
rect 16850 -360 16855 -335
rect 16820 -380 16855 -360
rect 16820 -405 16825 -380
rect 16850 -405 16855 -380
rect 16820 -420 16855 -405
rect 16880 -335 16915 -320
rect 16880 -360 16885 -335
rect 16910 -360 16915 -335
rect 16880 -380 16915 -360
rect 16880 -405 16885 -380
rect 16910 -405 16915 -380
rect 16880 -420 16915 -405
rect 16940 -335 16975 -320
rect 16940 -360 16945 -335
rect 16970 -360 16975 -335
rect 16940 -380 16975 -360
rect 16940 -405 16945 -380
rect 16970 -405 16975 -380
rect 16940 -420 16975 -405
rect 17000 -335 17035 -320
rect 17000 -360 17005 -335
rect 17030 -360 17035 -335
rect 17000 -380 17035 -360
rect 17000 -405 17005 -380
rect 17030 -405 17035 -380
rect 17000 -420 17035 -405
rect 17060 -335 17095 -320
rect 17060 -360 17065 -335
rect 17090 -360 17095 -335
rect 17060 -380 17095 -360
rect 17060 -405 17065 -380
rect 17090 -405 17095 -380
rect 17060 -420 17095 -405
rect 17120 -335 17155 -320
rect 17120 -360 17125 -335
rect 17150 -360 17155 -335
rect 17120 -380 17155 -360
rect 17120 -405 17125 -380
rect 17150 -405 17155 -380
rect 17120 -420 17155 -405
rect 17180 -335 17215 -320
rect 17180 -360 17185 -335
rect 17210 -360 17215 -335
rect 17180 -380 17215 -360
rect 17180 -405 17185 -380
rect 17210 -405 17215 -380
rect 17180 -420 17215 -405
rect 17240 -335 17275 -320
rect 17240 -360 17245 -335
rect 17270 -360 17275 -335
rect 17240 -380 17275 -360
rect 17240 -405 17245 -380
rect 17270 -405 17275 -380
rect 17240 -420 17275 -405
rect 17300 -335 17335 -320
rect 17300 -360 17305 -335
rect 17330 -360 17335 -335
rect 17300 -380 17335 -360
rect 17300 -405 17305 -380
rect 17330 -405 17335 -380
rect 17300 -420 17335 -405
rect 17360 -335 17395 -320
rect 17360 -360 17365 -335
rect 17390 -360 17395 -335
rect 17360 -380 17395 -360
rect 17360 -405 17365 -380
rect 17390 -405 17395 -380
rect 17360 -420 17395 -405
rect 17420 -335 17455 -320
rect 17420 -360 17425 -335
rect 17450 -360 17455 -335
rect 17420 -380 17455 -360
rect 17420 -405 17425 -380
rect 17450 -405 17455 -380
rect 17420 -420 17455 -405
rect 17480 -335 17515 -320
rect 17480 -360 17485 -335
rect 17510 -360 17515 -335
rect 17480 -380 17515 -360
rect 17480 -405 17485 -380
rect 17510 -405 17515 -380
rect 17480 -420 17515 -405
rect 17540 -335 17575 -320
rect 17540 -360 17545 -335
rect 17570 -360 17575 -335
rect 17540 -380 17575 -360
rect 17540 -405 17545 -380
rect 17570 -405 17575 -380
rect 17540 -420 17575 -405
rect 17600 -335 17635 -320
rect 17600 -360 17605 -335
rect 17630 -360 17635 -335
rect 17600 -380 17635 -360
rect 17600 -405 17605 -380
rect 17630 -405 17635 -380
rect 17600 -420 17635 -405
rect 17660 -335 17695 -320
rect 17660 -360 17665 -335
rect 17690 -360 17695 -335
rect 17660 -380 17695 -360
rect 17660 -405 17665 -380
rect 17690 -405 17695 -380
rect 17660 -420 17695 -405
rect 17720 -335 17755 -320
rect 17720 -360 17725 -335
rect 17750 -360 17755 -335
rect 17720 -380 17755 -360
rect 17720 -405 17725 -380
rect 17750 -405 17755 -380
rect 17720 -420 17755 -405
rect 17780 -335 17815 -320
rect 17780 -360 17785 -335
rect 17810 -360 17815 -335
rect 17780 -380 17815 -360
rect 17780 -405 17785 -380
rect 17810 -405 17815 -380
rect 17780 -420 17815 -405
rect 17840 -335 17875 -320
rect 17840 -360 17845 -335
rect 17870 -360 17875 -335
rect 17840 -380 17875 -360
rect 17840 -405 17845 -380
rect 17870 -405 17875 -380
rect 17840 -420 17875 -405
rect 17900 -335 17935 -320
rect 17900 -360 17905 -335
rect 17930 -360 17935 -335
rect 17900 -380 17935 -360
rect 17900 -405 17905 -380
rect 17930 -405 17935 -380
rect 17900 -420 17935 -405
rect 17960 -335 17995 -320
rect 17960 -360 17965 -335
rect 17990 -360 17995 -335
rect 17960 -380 17995 -360
rect 17960 -405 17965 -380
rect 17990 -405 17995 -380
rect 17960 -420 17995 -405
rect 18020 -335 18055 -320
rect 18020 -360 18025 -335
rect 18050 -360 18055 -335
rect 18020 -380 18055 -360
rect 18020 -405 18025 -380
rect 18050 -405 18055 -380
rect 18020 -420 18055 -405
rect 18080 -335 18115 -320
rect 18080 -360 18085 -335
rect 18110 -360 18115 -335
rect 18080 -380 18115 -360
rect 18080 -405 18085 -380
rect 18110 -405 18115 -380
rect 18080 -420 18115 -405
rect 18140 -335 18175 -320
rect 18140 -360 18145 -335
rect 18170 -360 18175 -335
rect 18140 -380 18175 -360
rect 18140 -405 18145 -380
rect 18170 -405 18175 -380
rect 18140 -420 18175 -405
rect 18200 -335 18235 -320
rect 18200 -360 18205 -335
rect 18230 -360 18235 -335
rect 18200 -380 18235 -360
rect 18200 -405 18205 -380
rect 18230 -405 18235 -380
rect 18200 -420 18235 -405
rect 18260 -335 18295 -320
rect 18260 -360 18265 -335
rect 18290 -360 18295 -335
rect 18260 -380 18295 -360
rect 18260 -405 18265 -380
rect 18290 -405 18295 -380
rect 18260 -420 18295 -405
rect 18320 -335 18355 -320
rect 18320 -360 18325 -335
rect 18350 -360 18355 -335
rect 18320 -380 18355 -360
rect 18320 -405 18325 -380
rect 18350 -405 18355 -380
rect 18320 -420 18355 -405
rect 18380 -335 18415 -320
rect 18380 -360 18385 -335
rect 18410 -360 18415 -335
rect 18380 -380 18415 -360
rect 18380 -405 18385 -380
rect 18410 -405 18415 -380
rect 18380 -420 18415 -405
rect 18440 -335 18475 -320
rect 18440 -360 18445 -335
rect 18470 -360 18475 -335
rect 18440 -380 18475 -360
rect 18440 -405 18445 -380
rect 18470 -405 18475 -380
rect 18440 -420 18475 -405
rect 18500 -335 18535 -320
rect 18500 -360 18505 -335
rect 18530 -360 18535 -335
rect 18500 -380 18535 -360
rect 18500 -405 18505 -380
rect 18530 -405 18535 -380
rect 18500 -420 18535 -405
rect 18560 -335 18595 -320
rect 18560 -360 18565 -335
rect 18590 -360 18595 -335
rect 18560 -380 18595 -360
rect 18560 -405 18565 -380
rect 18590 -405 18595 -380
rect 18560 -420 18595 -405
rect 18620 -335 18655 -320
rect 18620 -360 18625 -335
rect 18650 -360 18655 -335
rect 18620 -380 18655 -360
rect 18620 -405 18625 -380
rect 18650 -405 18655 -380
rect 18620 -420 18655 -405
rect 18680 -335 18715 -320
rect 18680 -360 18685 -335
rect 18710 -360 18715 -335
rect 18680 -380 18715 -360
rect 18680 -405 18685 -380
rect 18710 -405 18715 -380
rect 18680 -420 18715 -405
rect 18740 -335 18775 -320
rect 18740 -360 18745 -335
rect 18770 -360 18775 -335
rect 18740 -380 18775 -360
rect 18740 -405 18745 -380
rect 18770 -405 18775 -380
rect 18740 -420 18775 -405
rect 18800 -335 18835 -320
rect 18800 -360 18805 -335
rect 18830 -360 18835 -335
rect 18800 -380 18835 -360
rect 18800 -405 18805 -380
rect 18830 -405 18835 -380
rect 18800 -420 18835 -405
rect 18860 -335 18895 -320
rect 18860 -360 18865 -335
rect 18890 -360 18895 -335
rect 18860 -380 18895 -360
rect 18860 -405 18865 -380
rect 18890 -405 18895 -380
rect 18860 -420 18895 -405
rect 18920 -335 18955 -320
rect 18920 -360 18925 -335
rect 18950 -360 18955 -335
rect 18920 -380 18955 -360
rect 18920 -405 18925 -380
rect 18950 -405 18955 -380
rect 18920 -420 18955 -405
rect 18980 -335 19015 -320
rect 18980 -360 18985 -335
rect 19010 -360 19015 -335
rect 18980 -380 19015 -360
rect 18980 -405 18985 -380
rect 19010 -405 19015 -380
rect 18980 -420 19015 -405
rect 19040 -335 19075 -320
rect 19040 -360 19045 -335
rect 19070 -360 19075 -335
rect 19040 -380 19075 -360
rect 19040 -405 19045 -380
rect 19070 -405 19075 -380
rect 19040 -420 19075 -405
rect 19100 -335 19135 -320
rect 19100 -360 19105 -335
rect 19130 -360 19135 -335
rect 19100 -380 19135 -360
rect 19100 -405 19105 -380
rect 19130 -405 19135 -380
rect 19100 -420 19135 -405
rect 19160 -335 19195 -320
rect 19160 -360 19165 -335
rect 19190 -360 19195 -335
rect 19160 -380 19195 -360
rect 19160 -405 19165 -380
rect 19190 -405 19195 -380
rect 19160 -420 19195 -405
rect 19220 -335 19255 -320
rect 19220 -360 19225 -335
rect 19250 -360 19255 -335
rect 19220 -380 19255 -360
rect 19220 -405 19225 -380
rect 19250 -405 19255 -380
rect 19220 -420 19255 -405
rect 19280 -335 19315 -320
rect 19280 -360 19285 -335
rect 19310 -360 19315 -335
rect 19280 -380 19315 -360
rect 19280 -405 19285 -380
rect 19310 -405 19315 -380
rect 19280 -420 19315 -405
rect 19340 -335 19375 -320
rect 19340 -360 19345 -335
rect 19370 -360 19375 -335
rect 19340 -380 19375 -360
rect 19340 -405 19345 -380
rect 19370 -405 19375 -380
rect 19340 -420 19375 -405
rect 19400 -335 19435 -320
rect 19400 -360 19405 -335
rect 19430 -360 19435 -335
rect 19400 -380 19435 -360
rect 19400 -405 19405 -380
rect 19430 -405 19435 -380
rect 19400 -420 19435 -405
rect 19460 -335 19495 -320
rect 19460 -360 19465 -335
rect 19490 -360 19495 -335
rect 19460 -380 19495 -360
rect 19460 -405 19465 -380
rect 19490 -405 19495 -380
rect 19460 -420 19495 -405
rect 19520 -335 19555 -320
rect 19520 -360 19525 -335
rect 19550 -360 19555 -335
rect 19520 -380 19555 -360
rect 19520 -405 19525 -380
rect 19550 -405 19555 -380
rect 19520 -420 19555 -405
rect 19580 -335 19615 -320
rect 19580 -360 19585 -335
rect 19610 -360 19615 -335
rect 19580 -380 19615 -360
rect 19580 -405 19585 -380
rect 19610 -405 19615 -380
rect 19580 -420 19615 -405
rect 19640 -335 19675 -320
rect 19640 -360 19645 -335
rect 19670 -360 19675 -335
rect 19640 -380 19675 -360
rect 19640 -405 19645 -380
rect 19670 -405 19675 -380
rect 19640 -420 19675 -405
rect 19700 -335 19735 -320
rect 19700 -360 19705 -335
rect 19730 -360 19735 -335
rect 19700 -380 19735 -360
rect 19700 -405 19705 -380
rect 19730 -405 19735 -380
rect 19700 -420 19735 -405
rect 19760 -335 19795 -320
rect 19760 -360 19765 -335
rect 19790 -360 19795 -335
rect 19760 -380 19795 -360
rect 19760 -405 19765 -380
rect 19790 -405 19795 -380
rect 19760 -420 19795 -405
rect 19820 -335 19855 -320
rect 19820 -360 19825 -335
rect 19850 -360 19855 -335
rect 19820 -380 19855 -360
rect 19820 -405 19825 -380
rect 19850 -405 19855 -380
rect 19820 -420 19855 -405
rect 19880 -335 19915 -320
rect 19880 -360 19885 -335
rect 19910 -360 19915 -335
rect 19880 -380 19915 -360
rect 19880 -405 19885 -380
rect 19910 -405 19915 -380
rect 19880 -420 19915 -405
rect 19940 -335 19975 -320
rect 19940 -360 19945 -335
rect 19970 -360 19975 -335
rect 19940 -380 19975 -360
rect 19940 -405 19945 -380
rect 19970 -405 19975 -380
rect 19940 -420 19975 -405
rect 20000 -335 20035 -320
rect 20000 -360 20005 -335
rect 20030 -360 20035 -335
rect 20000 -380 20035 -360
rect 20000 -405 20005 -380
rect 20030 -405 20035 -380
rect 20000 -420 20035 -405
rect 20060 -335 20095 -320
rect 20060 -360 20065 -335
rect 20090 -360 20095 -335
rect 20060 -380 20095 -360
rect 20060 -405 20065 -380
rect 20090 -405 20095 -380
rect 20060 -420 20095 -405
rect 20120 -335 20155 -320
rect 20120 -360 20125 -335
rect 20150 -360 20155 -335
rect 20120 -380 20155 -360
rect 20120 -405 20125 -380
rect 20150 -405 20155 -380
rect 20120 -420 20155 -405
rect 20180 -335 20215 -320
rect 20180 -360 20185 -335
rect 20210 -360 20215 -335
rect 20180 -380 20215 -360
rect 20180 -405 20185 -380
rect 20210 -405 20215 -380
rect 20180 -420 20215 -405
rect 20240 -335 20275 -320
rect 20240 -360 20245 -335
rect 20270 -360 20275 -335
rect 20240 -380 20275 -360
rect 20240 -405 20245 -380
rect 20270 -405 20275 -380
rect 20240 -420 20275 -405
rect 20300 -335 20335 -320
rect 20300 -360 20305 -335
rect 20330 -360 20335 -335
rect 20300 -380 20335 -360
rect 20300 -405 20305 -380
rect 20330 -405 20335 -380
rect 20300 -420 20335 -405
rect 20360 -335 20395 -320
rect 20360 -360 20365 -335
rect 20390 -360 20395 -335
rect 20360 -380 20395 -360
rect 20360 -405 20365 -380
rect 20390 -405 20395 -380
rect 20360 -420 20395 -405
rect 20420 -335 20455 -320
rect 20420 -360 20425 -335
rect 20450 -360 20455 -335
rect 20420 -380 20455 -360
rect 20420 -405 20425 -380
rect 20450 -405 20455 -380
rect 20420 -420 20455 -405
rect 20480 -335 20515 -320
rect 20480 -360 20485 -335
rect 20510 -360 20515 -335
rect 20480 -380 20515 -360
rect 20480 -405 20485 -380
rect 20510 -405 20515 -380
rect 20480 -420 20515 -405
rect 20540 -335 20575 -320
rect 20540 -360 20545 -335
rect 20570 -360 20575 -335
rect 20540 -380 20575 -360
rect 20540 -405 20545 -380
rect 20570 -405 20575 -380
rect 20540 -420 20575 -405
rect 20600 -335 20635 -320
rect 20600 -360 20605 -335
rect 20630 -360 20635 -335
rect 20600 -380 20635 -360
rect 20600 -405 20605 -380
rect 20630 -405 20635 -380
rect 20600 -420 20635 -405
rect 20660 -335 20695 -320
rect 20660 -360 20665 -335
rect 20690 -360 20695 -335
rect 20660 -380 20695 -360
rect 20660 -405 20665 -380
rect 20690 -405 20695 -380
rect 20660 -420 20695 -405
rect 20720 -335 20755 -320
rect 20720 -360 20725 -335
rect 20750 -360 20755 -335
rect 20720 -380 20755 -360
rect 20720 -405 20725 -380
rect 20750 -405 20755 -380
rect 20720 -420 20755 -405
rect 20780 -335 20815 -320
rect 20780 -360 20785 -335
rect 20810 -360 20815 -335
rect 20780 -380 20815 -360
rect 20780 -405 20785 -380
rect 20810 -405 20815 -380
rect 20780 -420 20815 -405
rect 20840 -335 20875 -320
rect 20840 -360 20845 -335
rect 20870 -360 20875 -335
rect 20840 -380 20875 -360
rect 20840 -405 20845 -380
rect 20870 -405 20875 -380
rect 20840 -420 20875 -405
rect 20900 -335 20935 -320
rect 20900 -360 20905 -335
rect 20930 -360 20935 -335
rect 20900 -380 20935 -360
rect 20900 -405 20905 -380
rect 20930 -405 20935 -380
rect 20900 -420 20935 -405
rect 20960 -335 20995 -320
rect 20960 -360 20965 -335
rect 20990 -360 20995 -335
rect 20960 -380 20995 -360
rect 20960 -405 20965 -380
rect 20990 -405 20995 -380
rect 20960 -420 20995 -405
rect 21020 -335 21055 -320
rect 21020 -360 21025 -335
rect 21050 -360 21055 -335
rect 21020 -380 21055 -360
rect 21020 -405 21025 -380
rect 21050 -405 21055 -380
rect 21020 -420 21055 -405
rect 21080 -335 21115 -320
rect 21080 -360 21085 -335
rect 21110 -360 21115 -335
rect 21080 -380 21115 -360
rect 21080 -405 21085 -380
rect 21110 -405 21115 -380
rect 21080 -420 21115 -405
rect 21140 -335 21175 -320
rect 21140 -360 21145 -335
rect 21170 -360 21175 -335
rect 21140 -380 21175 -360
rect 21140 -405 21145 -380
rect 21170 -405 21175 -380
rect 21140 -420 21175 -405
rect 21200 -335 21235 -320
rect 21200 -360 21205 -335
rect 21230 -360 21235 -335
rect 21200 -380 21235 -360
rect 21200 -405 21205 -380
rect 21230 -405 21235 -380
rect 21200 -420 21235 -405
rect 21260 -335 21295 -320
rect 21260 -360 21265 -335
rect 21290 -360 21295 -335
rect 21260 -380 21295 -360
rect 21260 -405 21265 -380
rect 21290 -405 21295 -380
rect 21260 -420 21295 -405
rect 21320 -335 21355 -320
rect 21320 -360 21325 -335
rect 21350 -360 21355 -335
rect 21320 -380 21355 -360
rect 21320 -405 21325 -380
rect 21350 -405 21355 -380
rect 21320 -420 21355 -405
rect 21380 -335 21415 -320
rect 21380 -360 21385 -335
rect 21410 -360 21415 -335
rect 21380 -380 21415 -360
rect 21380 -405 21385 -380
rect 21410 -405 21415 -380
rect 21380 -420 21415 -405
rect 21440 -335 21475 -320
rect 21440 -360 21445 -335
rect 21470 -360 21475 -335
rect 21440 -380 21475 -360
rect 21440 -405 21445 -380
rect 21470 -405 21475 -380
rect 21440 -420 21475 -405
rect 21500 -335 21535 -320
rect 21500 -360 21505 -335
rect 21530 -360 21535 -335
rect 21500 -380 21535 -360
rect 21500 -405 21505 -380
rect 21530 -405 21535 -380
rect 21500 -420 21535 -405
rect 21560 -335 21595 -320
rect 21560 -360 21565 -335
rect 21590 -360 21595 -335
rect 21560 -380 21595 -360
rect 21560 -405 21565 -380
rect 21590 -405 21595 -380
rect 21560 -420 21595 -405
rect 21620 -335 21655 -320
rect 21620 -360 21625 -335
rect 21650 -360 21655 -335
rect 21620 -380 21655 -360
rect 21620 -405 21625 -380
rect 21650 -405 21655 -380
rect 21620 -420 21655 -405
rect 21680 -335 21715 -320
rect 21680 -360 21685 -335
rect 21710 -360 21715 -335
rect 21680 -380 21715 -360
rect 21680 -405 21685 -380
rect 21710 -405 21715 -380
rect 21680 -420 21715 -405
rect 21740 -335 21775 -320
rect 21740 -360 21745 -335
rect 21770 -360 21775 -335
rect 21740 -380 21775 -360
rect 21740 -405 21745 -380
rect 21770 -405 21775 -380
rect 21740 -420 21775 -405
rect 21800 -335 21835 -320
rect 21800 -360 21805 -335
rect 21830 -360 21835 -335
rect 21800 -380 21835 -360
rect 21800 -405 21805 -380
rect 21830 -405 21835 -380
rect 21800 -420 21835 -405
rect 21860 -335 21895 -320
rect 21860 -360 21865 -335
rect 21890 -360 21895 -335
rect 21860 -380 21895 -360
rect 21860 -405 21865 -380
rect 21890 -405 21895 -380
rect 21860 -420 21895 -405
rect 21920 -335 21955 -320
rect 21920 -360 21925 -335
rect 21950 -360 21955 -335
rect 21920 -380 21955 -360
rect 21920 -405 21925 -380
rect 21950 -405 21955 -380
rect 21920 -420 21955 -405
rect 21980 -335 22015 -320
rect 21980 -360 21985 -335
rect 22010 -360 22015 -335
rect 21980 -380 22015 -360
rect 21980 -405 21985 -380
rect 22010 -405 22015 -380
rect 21980 -420 22015 -405
rect 22040 -335 22075 -320
rect 22040 -360 22045 -335
rect 22070 -360 22075 -335
rect 22040 -380 22075 -360
rect 22040 -405 22045 -380
rect 22070 -405 22075 -380
rect 22040 -420 22075 -405
rect 22100 -335 22135 -320
rect 22100 -360 22105 -335
rect 22130 -360 22135 -335
rect 22100 -380 22135 -360
rect 22100 -405 22105 -380
rect 22130 -405 22135 -380
rect 22100 -420 22135 -405
rect 22160 -335 22195 -320
rect 22160 -360 22165 -335
rect 22190 -360 22195 -335
rect 22160 -380 22195 -360
rect 22160 -405 22165 -380
rect 22190 -405 22195 -380
rect 22160 -420 22195 -405
rect 22220 -335 22255 -320
rect 22220 -360 22225 -335
rect 22250 -360 22255 -335
rect 22220 -380 22255 -360
rect 22220 -405 22225 -380
rect 22250 -405 22255 -380
rect 22220 -420 22255 -405
rect 22280 -335 22315 -320
rect 22280 -360 22285 -335
rect 22310 -360 22315 -335
rect 22280 -380 22315 -360
rect 22280 -405 22285 -380
rect 22310 -405 22315 -380
rect 22280 -420 22315 -405
rect 22340 -335 22375 -320
rect 22340 -360 22345 -335
rect 22370 -360 22375 -335
rect 22340 -380 22375 -360
rect 22340 -405 22345 -380
rect 22370 -405 22375 -380
rect 22340 -420 22375 -405
rect 22400 -335 22435 -320
rect 22400 -360 22405 -335
rect 22430 -360 22435 -335
rect 22400 -380 22435 -360
rect 22400 -405 22405 -380
rect 22430 -405 22435 -380
rect 22400 -420 22435 -405
rect 22460 -335 22495 -320
rect 22460 -360 22465 -335
rect 22490 -360 22495 -335
rect 22460 -380 22495 -360
rect 22460 -405 22465 -380
rect 22490 -405 22495 -380
rect 22460 -420 22495 -405
rect 22520 -335 22555 -320
rect 22520 -360 22525 -335
rect 22550 -360 22555 -335
rect 22520 -380 22555 -360
rect 22520 -405 22525 -380
rect 22550 -405 22555 -380
rect 22520 -420 22555 -405
rect 22580 -335 22615 -320
rect 22580 -360 22585 -335
rect 22610 -360 22615 -335
rect 22580 -380 22615 -360
rect 22580 -405 22585 -380
rect 22610 -405 22615 -380
rect 22580 -420 22615 -405
rect 22640 -335 22675 -320
rect 22640 -360 22645 -335
rect 22670 -360 22675 -335
rect 22640 -380 22675 -360
rect 22640 -405 22645 -380
rect 22670 -405 22675 -380
rect 22640 -420 22675 -405
rect 22700 -335 22735 -320
rect 22700 -360 22705 -335
rect 22730 -360 22735 -335
rect 22700 -380 22735 -360
rect 22700 -405 22705 -380
rect 22730 -405 22735 -380
rect 22700 -420 22735 -405
rect 22760 -335 22795 -320
rect 22760 -360 22765 -335
rect 22790 -360 22795 -335
rect 22760 -380 22795 -360
rect 22760 -405 22765 -380
rect 22790 -405 22795 -380
rect 22760 -420 22795 -405
rect 22820 -335 22855 -320
rect 22820 -360 22825 -335
rect 22850 -360 22855 -335
rect 22820 -380 22855 -360
rect 22820 -405 22825 -380
rect 22850 -405 22855 -380
rect 22820 -420 22855 -405
rect 22880 -335 22915 -320
rect 22880 -360 22885 -335
rect 22910 -360 22915 -335
rect 22880 -380 22915 -360
rect 22880 -405 22885 -380
rect 22910 -405 22915 -380
rect 22880 -420 22915 -405
rect 22940 -335 22975 -320
rect 22940 -360 22945 -335
rect 22970 -360 22975 -335
rect 22940 -380 22975 -360
rect 22940 -405 22945 -380
rect 22970 -405 22975 -380
rect 22940 -420 22975 -405
rect 23000 -335 23035 -320
rect 23000 -360 23005 -335
rect 23030 -360 23035 -335
rect 23000 -380 23035 -360
rect 23000 -405 23005 -380
rect 23030 -405 23035 -380
rect 23000 -420 23035 -405
rect 23060 -335 23095 -320
rect 23060 -360 23065 -335
rect 23090 -360 23095 -335
rect 23060 -380 23095 -360
rect 23060 -405 23065 -380
rect 23090 -405 23095 -380
rect 23060 -420 23095 -405
rect 23120 -335 23155 -320
rect 23120 -360 23125 -335
rect 23150 -360 23155 -335
rect 23120 -380 23155 -360
rect 23120 -405 23125 -380
rect 23150 -405 23155 -380
rect 23120 -420 23155 -405
rect 23180 -335 23215 -320
rect 23180 -360 23185 -335
rect 23210 -360 23215 -335
rect 23180 -380 23215 -360
rect 23180 -405 23185 -380
rect 23210 -405 23215 -380
rect 23180 -420 23215 -405
rect 23240 -335 23275 -320
rect 23240 -360 23245 -335
rect 23270 -360 23275 -335
rect 23240 -380 23275 -360
rect 23240 -405 23245 -380
rect 23270 -405 23275 -380
rect 23240 -420 23275 -405
rect 23300 -335 23335 -320
rect 23300 -360 23305 -335
rect 23330 -360 23335 -335
rect 23300 -380 23335 -360
rect 23300 -405 23305 -380
rect 23330 -405 23335 -380
rect 23300 -420 23335 -405
rect 23360 -335 23395 -320
rect 23360 -360 23365 -335
rect 23390 -360 23395 -335
rect 23360 -380 23395 -360
rect 23360 -405 23365 -380
rect 23390 -405 23395 -380
rect 23360 -420 23395 -405
rect 23420 -335 23455 -320
rect 23420 -360 23425 -335
rect 23450 -360 23455 -335
rect 23420 -380 23455 -360
rect 23420 -405 23425 -380
rect 23450 -405 23455 -380
rect 23420 -420 23455 -405
rect 23480 -335 23515 -320
rect 23480 -360 23485 -335
rect 23510 -360 23515 -335
rect 23480 -380 23515 -360
rect 23480 -405 23485 -380
rect 23510 -405 23515 -380
rect 23480 -420 23515 -405
rect 23540 -335 23575 -320
rect 23540 -360 23545 -335
rect 23570 -360 23575 -335
rect 23540 -380 23575 -360
rect 23540 -405 23545 -380
rect 23570 -405 23575 -380
rect 23540 -420 23575 -405
rect 23600 -335 23635 -320
rect 23600 -360 23605 -335
rect 23630 -360 23635 -335
rect 23600 -380 23635 -360
rect 23600 -405 23605 -380
rect 23630 -405 23635 -380
rect 23600 -420 23635 -405
rect 23660 -335 23695 -320
rect 23660 -360 23665 -335
rect 23690 -360 23695 -335
rect 23660 -380 23695 -360
rect 23660 -405 23665 -380
rect 23690 -405 23695 -380
rect 23660 -420 23695 -405
rect 23720 -335 23755 -320
rect 23720 -360 23725 -335
rect 23750 -360 23755 -335
rect 23720 -380 23755 -360
rect 23720 -405 23725 -380
rect 23750 -405 23755 -380
rect 23720 -420 23755 -405
rect 23780 -335 23815 -320
rect 23780 -360 23785 -335
rect 23810 -360 23815 -335
rect 23780 -380 23815 -360
rect 23780 -405 23785 -380
rect 23810 -405 23815 -380
rect 23780 -420 23815 -405
rect 23840 -335 23875 -320
rect 23840 -360 23845 -335
rect 23870 -360 23875 -335
rect 23840 -380 23875 -360
rect 23840 -405 23845 -380
rect 23870 -405 23875 -380
rect 23840 -420 23875 -405
rect 23900 -335 23935 -320
rect 23900 -360 23905 -335
rect 23930 -360 23935 -335
rect 23900 -380 23935 -360
rect 23900 -405 23905 -380
rect 23930 -405 23935 -380
rect 23900 -420 23935 -405
rect 23960 -335 23995 -320
rect 23960 -360 23965 -335
rect 23990 -360 23995 -335
rect 23960 -380 23995 -360
rect 23960 -405 23965 -380
rect 23990 -405 23995 -380
rect 23960 -420 23995 -405
rect 24020 -335 24055 -320
rect 24020 -360 24025 -335
rect 24050 -360 24055 -335
rect 24020 -380 24055 -360
rect 24020 -405 24025 -380
rect 24050 -405 24055 -380
rect 24020 -420 24055 -405
rect 24080 -335 24115 -320
rect 24080 -360 24085 -335
rect 24110 -360 24115 -335
rect 24080 -380 24115 -360
rect 24080 -405 24085 -380
rect 24110 -405 24115 -380
rect 24080 -420 24115 -405
rect 24140 -335 24175 -320
rect 24140 -360 24145 -335
rect 24170 -360 24175 -335
rect 24140 -380 24175 -360
rect 24140 -405 24145 -380
rect 24170 -405 24175 -380
rect 24140 -420 24175 -405
rect 24200 -335 24235 -320
rect 24200 -360 24205 -335
rect 24230 -360 24235 -335
rect 24200 -380 24235 -360
rect 24200 -405 24205 -380
rect 24230 -405 24235 -380
rect 24200 -420 24235 -405
rect 24260 -335 24295 -320
rect 24260 -360 24265 -335
rect 24290 -360 24295 -335
rect 24260 -380 24295 -360
rect 24260 -405 24265 -380
rect 24290 -405 24295 -380
rect 24260 -420 24295 -405
rect 24320 -335 24355 -320
rect 24320 -360 24325 -335
rect 24350 -360 24355 -335
rect 24320 -380 24355 -360
rect 24320 -405 24325 -380
rect 24350 -405 24355 -380
rect 24320 -420 24355 -405
rect 24380 -335 24415 -320
rect 24380 -360 24385 -335
rect 24410 -360 24415 -335
rect 24380 -380 24415 -360
rect 24380 -405 24385 -380
rect 24410 -405 24415 -380
rect 24380 -420 24415 -405
rect 24440 -335 24475 -320
rect 24440 -360 24445 -335
rect 24470 -360 24475 -335
rect 24440 -380 24475 -360
rect 24440 -405 24445 -380
rect 24470 -405 24475 -380
rect 24440 -420 24475 -405
rect 24500 -335 24535 -320
rect 24500 -360 24505 -335
rect 24530 -360 24535 -335
rect 24500 -380 24535 -360
rect 24500 -405 24505 -380
rect 24530 -405 24535 -380
rect 24500 -420 24535 -405
rect 24560 -335 24595 -320
rect 24560 -360 24565 -335
rect 24590 -360 24595 -335
rect 24560 -380 24595 -360
rect 24560 -405 24565 -380
rect 24590 -405 24595 -380
rect 24560 -420 24595 -405
rect 24620 -335 24655 -320
rect 24620 -360 24625 -335
rect 24650 -360 24655 -335
rect 24620 -380 24655 -360
rect 24620 -405 24625 -380
rect 24650 -405 24655 -380
rect 24620 -420 24655 -405
rect 24680 -335 24715 -320
rect 24680 -360 24685 -335
rect 24710 -360 24715 -335
rect 24680 -380 24715 -360
rect 24680 -405 24685 -380
rect 24710 -405 24715 -380
rect 24680 -420 24715 -405
rect 24740 -335 24775 -320
rect 24740 -360 24745 -335
rect 24770 -360 24775 -335
rect 24740 -380 24775 -360
rect 24740 -405 24745 -380
rect 24770 -405 24775 -380
rect 24740 -420 24775 -405
rect 24800 -335 24835 -320
rect 24800 -360 24805 -335
rect 24830 -360 24835 -335
rect 24800 -380 24835 -360
rect 24800 -405 24805 -380
rect 24830 -405 24835 -380
rect 24800 -420 24835 -405
rect 24860 -335 24895 -320
rect 24860 -360 24865 -335
rect 24890 -360 24895 -335
rect 24860 -380 24895 -360
rect 24860 -405 24865 -380
rect 24890 -405 24895 -380
rect 24860 -420 24895 -405
rect 24920 -335 24955 -320
rect 24920 -360 24925 -335
rect 24950 -360 24955 -335
rect 24920 -380 24955 -360
rect 24920 -405 24925 -380
rect 24950 -405 24955 -380
rect 24920 -420 24955 -405
rect 24980 -335 25015 -320
rect 24980 -360 24985 -335
rect 25010 -360 25015 -335
rect 24980 -380 25015 -360
rect 24980 -405 24985 -380
rect 25010 -405 25015 -380
rect 24980 -420 25015 -405
rect 25040 -335 25075 -320
rect 25040 -360 25045 -335
rect 25070 -360 25075 -335
rect 25040 -380 25075 -360
rect 25040 -405 25045 -380
rect 25070 -405 25075 -380
rect 25040 -420 25075 -405
rect 25100 -335 25135 -320
rect 25100 -360 25105 -335
rect 25130 -360 25135 -335
rect 25100 -380 25135 -360
rect 25100 -405 25105 -380
rect 25130 -405 25135 -380
rect 25100 -420 25135 -405
rect 25160 -335 25195 -320
rect 25160 -360 25165 -335
rect 25190 -360 25195 -335
rect 25160 -380 25195 -360
rect 25160 -405 25165 -380
rect 25190 -405 25195 -380
rect 25160 -420 25195 -405
rect 25220 -335 25255 -320
rect 25220 -360 25225 -335
rect 25250 -360 25255 -335
rect 25220 -380 25255 -360
rect 25220 -405 25225 -380
rect 25250 -405 25255 -380
rect 25220 -420 25255 -405
rect 25280 -335 25315 -320
rect 25280 -360 25285 -335
rect 25310 -360 25315 -335
rect 25280 -380 25315 -360
rect 25280 -405 25285 -380
rect 25310 -405 25315 -380
rect 25280 -420 25315 -405
rect 25340 -335 25375 -320
rect 25340 -360 25345 -335
rect 25370 -360 25375 -335
rect 25340 -380 25375 -360
rect 25340 -405 25345 -380
rect 25370 -405 25375 -380
rect 25340 -420 25375 -405
rect 25400 -335 25435 -320
rect 25400 -360 25405 -335
rect 25430 -360 25435 -335
rect 25400 -380 25435 -360
rect 25400 -405 25405 -380
rect 25430 -405 25435 -380
rect 25400 -420 25435 -405
rect 25460 -335 25495 -320
rect 25460 -360 25465 -335
rect 25490 -360 25495 -335
rect 25460 -380 25495 -360
rect 25460 -405 25465 -380
rect 25490 -405 25495 -380
rect 25460 -420 25495 -405
rect 25520 -335 25555 -320
rect 25520 -360 25525 -335
rect 25550 -360 25555 -335
rect 25520 -380 25555 -360
rect 25520 -405 25525 -380
rect 25550 -405 25555 -380
rect 25520 -420 25555 -405
rect 25580 -335 25615 -320
rect 25580 -360 25585 -335
rect 25610 -360 25615 -335
rect 25580 -380 25615 -360
rect 25580 -405 25585 -380
rect 25610 -405 25615 -380
rect 25580 -420 25615 -405
rect 25640 -335 25675 -320
rect 25640 -360 25645 -335
rect 25670 -360 25675 -335
rect 25640 -380 25675 -360
rect 25640 -405 25645 -380
rect 25670 -405 25675 -380
rect 25640 -420 25675 -405
rect 25700 -335 25735 -320
rect 25700 -360 25705 -335
rect 25730 -360 25735 -335
rect 25700 -380 25735 -360
rect 25700 -405 25705 -380
rect 25730 -405 25735 -380
rect 25700 -420 25735 -405
rect 25760 -335 25795 -320
rect 25760 -360 25765 -335
rect 25790 -360 25795 -335
rect 25760 -380 25795 -360
rect 25760 -405 25765 -380
rect 25790 -405 25795 -380
rect 25760 -420 25795 -405
rect 25820 -335 25855 -320
rect 25820 -360 25825 -335
rect 25850 -360 25855 -335
rect 25820 -380 25855 -360
rect 25820 -405 25825 -380
rect 25850 -405 25855 -380
rect 25820 -420 25855 -405
rect 25880 -335 25915 -320
rect 25880 -360 25885 -335
rect 25910 -360 25915 -335
rect 25880 -380 25915 -360
rect 25880 -405 25885 -380
rect 25910 -405 25915 -380
rect 25880 -420 25915 -405
rect 25940 -335 25975 -320
rect 25940 -360 25945 -335
rect 25970 -360 25975 -335
rect 25940 -380 25975 -360
rect 25940 -405 25945 -380
rect 25970 -405 25975 -380
rect 25940 -420 25975 -405
rect 26000 -335 26035 -320
rect 26000 -360 26005 -335
rect 26030 -360 26035 -335
rect 26000 -380 26035 -360
rect 26000 -405 26005 -380
rect 26030 -405 26035 -380
rect 26000 -420 26035 -405
rect 26060 -335 26095 -320
rect 26060 -360 26065 -335
rect 26090 -360 26095 -335
rect 26060 -380 26095 -360
rect 26060 -405 26065 -380
rect 26090 -405 26095 -380
rect 26060 -420 26095 -405
rect 26120 -335 26155 -320
rect 26120 -360 26125 -335
rect 26150 -360 26155 -335
rect 26120 -380 26155 -360
rect 26120 -405 26125 -380
rect 26150 -405 26155 -380
rect 26120 -420 26155 -405
rect 26180 -335 26215 -320
rect 26180 -360 26185 -335
rect 26210 -360 26215 -335
rect 26180 -380 26215 -360
rect 26180 -405 26185 -380
rect 26210 -405 26215 -380
rect 26180 -420 26215 -405
rect 26240 -335 26275 -320
rect 26240 -360 26245 -335
rect 26270 -360 26275 -335
rect 26240 -380 26275 -360
rect 26240 -405 26245 -380
rect 26270 -405 26275 -380
rect 26240 -420 26275 -405
rect 26300 -335 26335 -320
rect 26300 -360 26305 -335
rect 26330 -360 26335 -335
rect 26300 -380 26335 -360
rect 26300 -405 26305 -380
rect 26330 -405 26335 -380
rect 26300 -420 26335 -405
rect 26360 -335 26395 -320
rect 26360 -360 26365 -335
rect 26390 -360 26395 -335
rect 26360 -380 26395 -360
rect 26360 -405 26365 -380
rect 26390 -405 26395 -380
rect 26360 -420 26395 -405
rect 26420 -335 26455 -320
rect 26420 -360 26425 -335
rect 26450 -360 26455 -335
rect 26420 -380 26455 -360
rect 26420 -405 26425 -380
rect 26450 -405 26455 -380
rect 26420 -420 26455 -405
rect 26480 -335 26515 -320
rect 26480 -360 26485 -335
rect 26510 -360 26515 -335
rect 26480 -380 26515 -360
rect 26480 -405 26485 -380
rect 26510 -405 26515 -380
rect 26480 -420 26515 -405
rect 26540 -335 26575 -320
rect 26540 -360 26545 -335
rect 26570 -360 26575 -335
rect 26540 -380 26575 -360
rect 26540 -405 26545 -380
rect 26570 -405 26575 -380
rect 26540 -420 26575 -405
rect 26600 -335 26635 -320
rect 26600 -360 26605 -335
rect 26630 -360 26635 -335
rect 26600 -380 26635 -360
rect 26600 -405 26605 -380
rect 26630 -405 26635 -380
rect 26600 -420 26635 -405
rect 26660 -335 26695 -320
rect 26660 -360 26665 -335
rect 26690 -360 26695 -335
rect 26660 -380 26695 -360
rect 26660 -405 26665 -380
rect 26690 -405 26695 -380
rect 26660 -420 26695 -405
rect 26720 -335 26755 -320
rect 26720 -360 26725 -335
rect 26750 -360 26755 -335
rect 26720 -380 26755 -360
rect 26720 -405 26725 -380
rect 26750 -405 26755 -380
rect 26720 -420 26755 -405
rect 26780 -335 26815 -320
rect 26780 -360 26785 -335
rect 26810 -360 26815 -335
rect 26780 -380 26815 -360
rect 26780 -405 26785 -380
rect 26810 -405 26815 -380
rect 26780 -420 26815 -405
rect 26840 -335 26875 -320
rect 26840 -360 26845 -335
rect 26870 -360 26875 -335
rect 26840 -380 26875 -360
rect 26840 -405 26845 -380
rect 26870 -405 26875 -380
rect 26840 -420 26875 -405
rect 26900 -335 26935 -320
rect 26900 -360 26905 -335
rect 26930 -360 26935 -335
rect 26900 -380 26935 -360
rect 26900 -405 26905 -380
rect 26930 -405 26935 -380
rect 26900 -420 26935 -405
rect 26960 -335 26995 -320
rect 26960 -360 26965 -335
rect 26990 -360 26995 -335
rect 26960 -380 26995 -360
rect 26960 -405 26965 -380
rect 26990 -405 26995 -380
rect 26960 -420 26995 -405
rect 27020 -335 27055 -320
rect 27020 -360 27025 -335
rect 27050 -360 27055 -335
rect 27020 -380 27055 -360
rect 27020 -405 27025 -380
rect 27050 -405 27055 -380
rect 27020 -420 27055 -405
rect 27080 -335 27115 -320
rect 27080 -360 27085 -335
rect 27110 -360 27115 -335
rect 27080 -380 27115 -360
rect 27080 -405 27085 -380
rect 27110 -405 27115 -380
rect 27080 -420 27115 -405
rect 27140 -335 27175 -320
rect 27140 -360 27145 -335
rect 27170 -360 27175 -335
rect 27140 -380 27175 -360
rect 27140 -405 27145 -380
rect 27170 -405 27175 -380
rect 27140 -420 27175 -405
rect 27200 -335 27235 -320
rect 27200 -360 27205 -335
rect 27230 -360 27235 -335
rect 27200 -380 27235 -360
rect 27200 -405 27205 -380
rect 27230 -405 27235 -380
rect 27200 -420 27235 -405
rect 27260 -335 27295 -320
rect 27260 -360 27265 -335
rect 27290 -360 27295 -335
rect 27260 -380 27295 -360
rect 27260 -405 27265 -380
rect 27290 -405 27295 -380
rect 27260 -420 27295 -405
rect 27320 -335 27355 -320
rect 27320 -360 27325 -335
rect 27350 -360 27355 -335
rect 27320 -380 27355 -360
rect 27320 -405 27325 -380
rect 27350 -405 27355 -380
rect 27320 -420 27355 -405
rect 27380 -335 27415 -320
rect 27380 -360 27385 -335
rect 27410 -360 27415 -335
rect 27380 -380 27415 -360
rect 27380 -405 27385 -380
rect 27410 -405 27415 -380
rect 27380 -420 27415 -405
rect 27440 -335 27475 -320
rect 27440 -360 27445 -335
rect 27470 -360 27475 -335
rect 27440 -380 27475 -360
rect 27440 -405 27445 -380
rect 27470 -405 27475 -380
rect 27440 -420 27475 -405
rect 27500 -335 27535 -320
rect 27500 -360 27505 -335
rect 27530 -360 27535 -335
rect 27500 -380 27535 -360
rect 27500 -405 27505 -380
rect 27530 -405 27535 -380
rect 27500 -420 27535 -405
rect 27560 -335 27595 -320
rect 27560 -360 27565 -335
rect 27590 -360 27595 -335
rect 27560 -380 27595 -360
rect 27560 -405 27565 -380
rect 27590 -405 27595 -380
rect 27560 -420 27595 -405
rect 27620 -335 27655 -320
rect 27620 -360 27625 -335
rect 27650 -360 27655 -335
rect 27620 -380 27655 -360
rect 27620 -405 27625 -380
rect 27650 -405 27655 -380
rect 27620 -420 27655 -405
rect 27680 -335 27715 -320
rect 27680 -360 27685 -335
rect 27710 -360 27715 -335
rect 27680 -380 27715 -360
rect 27680 -405 27685 -380
rect 27710 -405 27715 -380
rect 27680 -420 27715 -405
rect 27740 -335 27775 -320
rect 27740 -360 27745 -335
rect 27770 -360 27775 -335
rect 27740 -380 27775 -360
rect 27740 -405 27745 -380
rect 27770 -405 27775 -380
rect 27740 -420 27775 -405
rect 27800 -335 27835 -320
rect 27800 -360 27805 -335
rect 27830 -360 27835 -335
rect 27800 -380 27835 -360
rect 27800 -405 27805 -380
rect 27830 -405 27835 -380
rect 27800 -420 27835 -405
rect 27860 -335 27895 -320
rect 27860 -360 27865 -335
rect 27890 -360 27895 -335
rect 27860 -380 27895 -360
rect 27860 -405 27865 -380
rect 27890 -405 27895 -380
rect 27860 -420 27895 -405
rect 27920 -335 27955 -320
rect 27920 -360 27925 -335
rect 27950 -360 27955 -335
rect 27920 -380 27955 -360
rect 27920 -405 27925 -380
rect 27950 -405 27955 -380
rect 27920 -420 27955 -405
rect 27980 -335 28015 -320
rect 27980 -360 27985 -335
rect 28010 -360 28015 -335
rect 27980 -380 28015 -360
rect 27980 -405 27985 -380
rect 28010 -405 28015 -380
rect 27980 -420 28015 -405
rect 28040 -335 28075 -320
rect 28040 -360 28045 -335
rect 28070 -360 28075 -335
rect 28040 -380 28075 -360
rect 28040 -405 28045 -380
rect 28070 -405 28075 -380
rect 28040 -420 28075 -405
rect 28100 -335 28135 -320
rect 28100 -360 28105 -335
rect 28130 -360 28135 -335
rect 28100 -380 28135 -360
rect 28100 -405 28105 -380
rect 28130 -405 28135 -380
rect 28100 -420 28135 -405
rect 28160 -335 28195 -320
rect 28160 -360 28165 -335
rect 28190 -360 28195 -335
rect 28160 -380 28195 -360
rect 28160 -405 28165 -380
rect 28190 -405 28195 -380
rect 28160 -420 28195 -405
rect 28220 -335 28255 -320
rect 28220 -360 28225 -335
rect 28250 -360 28255 -335
rect 28220 -380 28255 -360
rect 28220 -405 28225 -380
rect 28250 -405 28255 -380
rect 28220 -420 28255 -405
rect 28280 -335 28315 -320
rect 28280 -360 28285 -335
rect 28310 -360 28315 -335
rect 28280 -380 28315 -360
rect 28280 -405 28285 -380
rect 28310 -405 28315 -380
rect 28280 -420 28315 -405
rect 28340 -335 28375 -320
rect 28340 -360 28345 -335
rect 28370 -360 28375 -335
rect 28340 -380 28375 -360
rect 28340 -405 28345 -380
rect 28370 -405 28375 -380
rect 28340 -420 28375 -405
rect 28400 -335 28435 -320
rect 28400 -360 28405 -335
rect 28430 -360 28435 -335
rect 28400 -380 28435 -360
rect 28400 -405 28405 -380
rect 28430 -405 28435 -380
rect 28400 -420 28435 -405
rect 28460 -335 28495 -320
rect 28460 -360 28465 -335
rect 28490 -360 28495 -335
rect 28460 -380 28495 -360
rect 28460 -405 28465 -380
rect 28490 -405 28495 -380
rect 28460 -420 28495 -405
rect 28520 -335 28555 -320
rect 28520 -360 28525 -335
rect 28550 -360 28555 -335
rect 28520 -380 28555 -360
rect 28520 -405 28525 -380
rect 28550 -405 28555 -380
rect 28520 -420 28555 -405
rect 28580 -335 28615 -320
rect 28580 -360 28585 -335
rect 28610 -360 28615 -335
rect 28580 -380 28615 -360
rect 28580 -405 28585 -380
rect 28610 -405 28615 -380
rect 28580 -420 28615 -405
rect 28640 -335 28675 -320
rect 28640 -360 28645 -335
rect 28670 -360 28675 -335
rect 28640 -380 28675 -360
rect 28640 -405 28645 -380
rect 28670 -405 28675 -380
rect 28640 -420 28675 -405
rect 28700 -335 28735 -320
rect 28700 -360 28705 -335
rect 28730 -360 28735 -335
rect 28700 -380 28735 -360
rect 28700 -405 28705 -380
rect 28730 -405 28735 -380
rect 28700 -420 28735 -405
rect 28760 -335 28795 -320
rect 28760 -360 28765 -335
rect 28790 -360 28795 -335
rect 28760 -380 28795 -360
rect 28760 -405 28765 -380
rect 28790 -405 28795 -380
rect 28760 -420 28795 -405
rect 28820 -335 28855 -320
rect 28820 -360 28825 -335
rect 28850 -360 28855 -335
rect 28820 -380 28855 -360
rect 28820 -405 28825 -380
rect 28850 -405 28855 -380
rect 28820 -420 28855 -405
rect 28880 -335 28915 -320
rect 28880 -360 28885 -335
rect 28910 -360 28915 -335
rect 28880 -380 28915 -360
rect 28880 -405 28885 -380
rect 28910 -405 28915 -380
rect 28880 -420 28915 -405
rect 28940 -335 28975 -320
rect 28940 -360 28945 -335
rect 28970 -360 28975 -335
rect 28940 -380 28975 -360
rect 28940 -405 28945 -380
rect 28970 -405 28975 -380
rect 28940 -420 28975 -405
rect 29000 -335 29035 -320
rect 29000 -360 29005 -335
rect 29030 -360 29035 -335
rect 29000 -380 29035 -360
rect 29000 -405 29005 -380
rect 29030 -405 29035 -380
rect 29000 -420 29035 -405
rect 29060 -335 29095 -320
rect 29060 -360 29065 -335
rect 29090 -360 29095 -335
rect 29060 -380 29095 -360
rect 29060 -405 29065 -380
rect 29090 -405 29095 -380
rect 29060 -420 29095 -405
rect 29120 -335 29155 -320
rect 29120 -360 29125 -335
rect 29150 -360 29155 -335
rect 29120 -380 29155 -360
rect 29120 -405 29125 -380
rect 29150 -405 29155 -380
rect 29120 -420 29155 -405
rect 29180 -335 29215 -320
rect 29180 -360 29185 -335
rect 29210 -360 29215 -335
rect 29180 -380 29215 -360
rect 29180 -405 29185 -380
rect 29210 -405 29215 -380
rect 29180 -420 29215 -405
rect 29240 -335 29275 -320
rect 29240 -360 29245 -335
rect 29270 -360 29275 -335
rect 29240 -380 29275 -360
rect 29240 -405 29245 -380
rect 29270 -405 29275 -380
rect 29240 -420 29275 -405
rect 29300 -335 29335 -320
rect 29300 -360 29305 -335
rect 29330 -360 29335 -335
rect 29300 -380 29335 -360
rect 29300 -405 29305 -380
rect 29330 -405 29335 -380
rect 29300 -420 29335 -405
rect 29360 -335 29395 -320
rect 29360 -360 29365 -335
rect 29390 -360 29395 -335
rect 29360 -380 29395 -360
rect 29360 -405 29365 -380
rect 29390 -405 29395 -380
rect 29360 -420 29395 -405
rect 29420 -335 29455 -320
rect 29420 -360 29425 -335
rect 29450 -360 29455 -335
rect 29420 -380 29455 -360
rect 29420 -405 29425 -380
rect 29450 -405 29455 -380
rect 29420 -420 29455 -405
rect 29480 -335 29515 -320
rect 29480 -360 29485 -335
rect 29510 -360 29515 -335
rect 29480 -380 29515 -360
rect 29480 -405 29485 -380
rect 29510 -405 29515 -380
rect 29480 -420 29515 -405
rect 29540 -335 29575 -320
rect 29540 -360 29545 -335
rect 29570 -360 29575 -335
rect 29540 -380 29575 -360
rect 29540 -405 29545 -380
rect 29570 -405 29575 -380
rect 29540 -420 29575 -405
rect 29600 -335 29635 -320
rect 29600 -360 29605 -335
rect 29630 -360 29635 -335
rect 29600 -380 29635 -360
rect 29600 -405 29605 -380
rect 29630 -405 29635 -380
rect 29600 -420 29635 -405
rect 29660 -335 29695 -320
rect 29660 -360 29665 -335
rect 29690 -360 29695 -335
rect 29660 -380 29695 -360
rect 29660 -405 29665 -380
rect 29690 -405 29695 -380
rect 29660 -420 29695 -405
rect 29720 -335 29755 -320
rect 29720 -360 29725 -335
rect 29750 -360 29755 -335
rect 29720 -380 29755 -360
rect 29720 -405 29725 -380
rect 29750 -405 29755 -380
rect 29720 -420 29755 -405
rect 29780 -335 29815 -320
rect 29780 -360 29785 -335
rect 29810 -360 29815 -335
rect 29780 -380 29815 -360
rect 29780 -405 29785 -380
rect 29810 -405 29815 -380
rect 29780 -420 29815 -405
rect 29840 -335 29875 -320
rect 29840 -360 29845 -335
rect 29870 -360 29875 -335
rect 29840 -380 29875 -360
rect 29840 -405 29845 -380
rect 29870 -405 29875 -380
rect 29840 -420 29875 -405
rect 29900 -335 29935 -320
rect 29900 -360 29905 -335
rect 29930 -360 29935 -335
rect 29900 -380 29935 -360
rect 29900 -405 29905 -380
rect 29930 -405 29935 -380
rect 29900 -420 29935 -405
rect 29960 -335 29995 -320
rect 29960 -360 29965 -335
rect 29990 -360 29995 -335
rect 29960 -380 29995 -360
rect 29960 -405 29965 -380
rect 29990 -405 29995 -380
rect 29960 -420 29995 -405
rect 30020 -335 30055 -320
rect 30020 -360 30025 -335
rect 30050 -360 30055 -335
rect 30020 -380 30055 -360
rect 30020 -405 30025 -380
rect 30050 -405 30055 -380
rect 30020 -420 30055 -405
rect 30080 -335 30115 -320
rect 30080 -360 30085 -335
rect 30110 -360 30115 -335
rect 30080 -380 30115 -360
rect 30080 -405 30085 -380
rect 30110 -405 30115 -380
rect 30080 -420 30115 -405
rect 30140 -335 30175 -320
rect 30140 -360 30145 -335
rect 30170 -360 30175 -335
rect 30140 -380 30175 -360
rect 30140 -405 30145 -380
rect 30170 -405 30175 -380
rect 30140 -420 30175 -405
rect 30200 -335 30235 -320
rect 30200 -360 30205 -335
rect 30230 -360 30235 -335
rect 30200 -380 30235 -360
rect 30200 -405 30205 -380
rect 30230 -405 30235 -380
rect 30200 -420 30235 -405
rect 30260 -335 30295 -320
rect 30260 -360 30265 -335
rect 30290 -360 30295 -335
rect 30260 -380 30295 -360
rect 30260 -405 30265 -380
rect 30290 -405 30295 -380
rect 30260 -420 30295 -405
rect 30320 -335 30355 -320
rect 30320 -360 30325 -335
rect 30350 -360 30355 -335
rect 30320 -380 30355 -360
rect 30320 -405 30325 -380
rect 30350 -405 30355 -380
rect 30320 -420 30355 -405
rect 30380 -335 30415 -320
rect 30380 -360 30385 -335
rect 30410 -360 30415 -335
rect 30380 -380 30415 -360
rect 30380 -405 30385 -380
rect 30410 -405 30415 -380
rect 30380 -420 30415 -405
rect 30440 -335 30475 -320
rect 30440 -360 30445 -335
rect 30470 -360 30475 -335
rect 30440 -380 30475 -360
rect 30440 -405 30445 -380
rect 30470 -405 30475 -380
rect 30440 -420 30475 -405
rect 30500 -335 30535 -320
rect 30500 -360 30505 -335
rect 30530 -360 30535 -335
rect 30500 -380 30535 -360
rect 30500 -405 30505 -380
rect 30530 -405 30535 -380
rect 30500 -420 30535 -405
rect 30560 -335 30595 -320
rect 30560 -360 30565 -335
rect 30590 -360 30595 -335
rect 30560 -380 30595 -360
rect 30560 -405 30565 -380
rect 30590 -405 30595 -380
rect 30560 -420 30595 -405
rect 30620 -335 30655 -320
rect 30620 -360 30625 -335
rect 30650 -360 30655 -335
rect 30620 -380 30655 -360
rect 30620 -405 30625 -380
rect 30650 -405 30655 -380
rect 30620 -420 30655 -405
rect 30680 -335 30715 -320
rect 30680 -360 30685 -335
rect 30710 -360 30715 -335
rect 30680 -380 30715 -360
rect 30680 -405 30685 -380
rect 30710 -405 30715 -380
rect 30680 -420 30715 -405
rect 25 -495 50 -420
rect 85 -445 105 -440
rect 205 -440 210 -420
rect 205 -445 225 -440
rect 325 -445 345 -440
rect 445 -440 450 -420
rect 445 -445 465 -440
rect 565 -445 585 -440
rect 685 -440 690 -420
rect 685 -445 705 -440
rect 805 -445 825 -440
rect 925 -440 930 -420
rect 925 -445 945 -440
rect 1045 -445 1065 -440
rect 1165 -440 1170 -420
rect 1165 -445 1185 -440
rect 1285 -445 1305 -440
rect 1405 -440 1410 -420
rect 1405 -445 1425 -440
rect 1525 -445 1545 -440
rect 1645 -440 1650 -420
rect 1645 -445 1665 -440
rect 1765 -445 1785 -440
rect 1885 -440 1890 -420
rect 1885 -445 1905 -440
rect 2005 -445 2025 -440
rect 2125 -440 2130 -420
rect 2125 -445 2145 -440
rect 2245 -445 2265 -440
rect 2365 -440 2370 -420
rect 2365 -445 2385 -440
rect 2485 -445 2505 -440
rect 2605 -440 2610 -420
rect 2605 -445 2625 -440
rect 2725 -445 2745 -440
rect 2845 -440 2850 -420
rect 2845 -445 2865 -440
rect 2965 -445 2985 -440
rect 3085 -440 3090 -420
rect 3085 -445 3105 -440
rect 3205 -445 3225 -440
rect 3325 -440 3330 -420
rect 3325 -445 3345 -440
rect 3445 -445 3465 -440
rect 3565 -440 3570 -420
rect 3565 -445 3585 -440
rect 3685 -445 3705 -440
rect 3805 -440 3810 -420
rect 3805 -445 3825 -440
rect 3925 -445 3945 -440
rect 4045 -440 4050 -420
rect 4045 -445 4065 -440
rect 4165 -445 4185 -440
rect 4285 -440 4290 -420
rect 4285 -445 4305 -440
rect 4405 -445 4425 -440
rect 4525 -440 4530 -420
rect 4525 -445 4545 -440
rect 4645 -445 4665 -440
rect 4765 -440 4770 -420
rect 4765 -445 4785 -440
rect 4885 -445 4905 -440
rect 5005 -440 5010 -420
rect 5005 -445 5025 -440
rect 5125 -445 5145 -440
rect 5245 -440 5250 -420
rect 5245 -445 5265 -440
rect 5365 -445 5385 -440
rect 5485 -440 5490 -420
rect 5485 -445 5505 -440
rect 5605 -445 5625 -440
rect 5725 -440 5730 -420
rect 5725 -445 5745 -440
rect 5845 -445 5865 -440
rect 5965 -440 5970 -420
rect 5965 -445 5985 -440
rect 6085 -445 6105 -440
rect 6205 -440 6210 -420
rect 6205 -445 6225 -440
rect 6325 -445 6345 -440
rect 6445 -440 6450 -420
rect 6445 -445 6465 -440
rect 6565 -445 6585 -440
rect 6685 -440 6690 -420
rect 6685 -445 6705 -440
rect 6805 -445 6825 -440
rect 6925 -440 6930 -420
rect 6925 -445 6945 -440
rect 7045 -445 7065 -440
rect 7165 -440 7170 -420
rect 7165 -445 7185 -440
rect 7285 -445 7305 -440
rect 7405 -440 7410 -420
rect 7405 -445 7425 -440
rect 7525 -445 7545 -440
rect 7645 -440 7650 -420
rect 7645 -445 7665 -440
rect 7765 -445 7785 -440
rect 7885 -440 7890 -420
rect 7885 -445 7905 -440
rect 8005 -445 8025 -440
rect 8125 -440 8130 -420
rect 8125 -445 8145 -440
rect 8245 -445 8265 -440
rect 8365 -440 8370 -420
rect 8365 -445 8385 -440
rect 8485 -445 8505 -440
rect 8605 -440 8610 -420
rect 8605 -445 8625 -440
rect 8725 -445 8745 -440
rect 8845 -440 8850 -420
rect 8845 -445 8865 -440
rect 8965 -445 8985 -440
rect 9085 -440 9090 -420
rect 9085 -445 9105 -440
rect 9205 -445 9225 -440
rect 9325 -440 9330 -420
rect 9325 -445 9345 -440
rect 9445 -445 9465 -440
rect 9565 -440 9570 -420
rect 9565 -445 9585 -440
rect 9685 -445 9705 -440
rect 9805 -440 9810 -420
rect 9805 -445 9825 -440
rect 9925 -445 9945 -440
rect 10045 -440 10050 -420
rect 10045 -445 10065 -440
rect 10165 -445 10185 -440
rect 10285 -440 10290 -420
rect 10285 -445 10305 -440
rect 10405 -445 10425 -440
rect 10525 -440 10530 -420
rect 10525 -445 10545 -440
rect 10645 -445 10665 -440
rect 10765 -440 10770 -420
rect 10765 -445 10785 -440
rect 10885 -445 10905 -440
rect 11005 -440 11010 -420
rect 11005 -445 11025 -440
rect 11125 -445 11145 -440
rect 11245 -440 11250 -420
rect 11245 -445 11265 -440
rect 11365 -445 11385 -440
rect 11485 -440 11490 -420
rect 11485 -445 11505 -440
rect 11605 -445 11625 -440
rect 11725 -440 11730 -420
rect 11725 -445 11745 -440
rect 11845 -445 11865 -440
rect 11965 -440 11970 -420
rect 11965 -445 11985 -440
rect 12085 -445 12105 -440
rect 12205 -440 12210 -420
rect 12205 -445 12225 -440
rect 12325 -445 12345 -440
rect 12445 -440 12450 -420
rect 12445 -445 12465 -440
rect 12565 -445 12585 -440
rect 12685 -440 12690 -420
rect 12685 -445 12705 -440
rect 12805 -445 12825 -440
rect 12925 -440 12930 -420
rect 12925 -445 12945 -440
rect 13045 -445 13065 -440
rect 13165 -440 13170 -420
rect 13165 -445 13185 -440
rect 13285 -445 13305 -440
rect 13405 -440 13410 -420
rect 13405 -445 13425 -440
rect 13525 -445 13545 -440
rect 13645 -440 13650 -420
rect 13645 -445 13665 -440
rect 13765 -445 13785 -440
rect 13885 -440 13890 -420
rect 13885 -445 13905 -440
rect 14005 -445 14025 -440
rect 14125 -440 14130 -420
rect 14125 -445 14145 -440
rect 14245 -445 14265 -440
rect 14365 -440 14370 -420
rect 14365 -445 14385 -440
rect 14485 -445 14505 -440
rect 14605 -440 14610 -420
rect 14605 -445 14625 -440
rect 14725 -445 14745 -440
rect 14845 -440 14850 -420
rect 14845 -445 14865 -440
rect 14965 -445 14985 -440
rect 15085 -440 15090 -420
rect 15085 -445 15105 -440
rect 15205 -445 15225 -440
rect 15325 -440 15330 -420
rect 15325 -445 15345 -440
rect 15445 -445 15465 -440
rect 15565 -440 15570 -420
rect 15565 -445 15585 -440
rect 15685 -445 15705 -440
rect 15805 -440 15810 -420
rect 15805 -445 15825 -440
rect 15925 -445 15945 -440
rect 16045 -440 16050 -420
rect 16045 -445 16065 -440
rect 16165 -445 16185 -440
rect 16285 -440 16290 -420
rect 16285 -445 16305 -440
rect 16405 -445 16425 -440
rect 16525 -440 16530 -420
rect 16525 -445 16545 -440
rect 16645 -445 16665 -440
rect 16765 -440 16770 -420
rect 16765 -445 16785 -440
rect 16885 -445 16905 -440
rect 17005 -440 17010 -420
rect 17005 -445 17025 -440
rect 17125 -445 17145 -440
rect 17245 -440 17250 -420
rect 17245 -445 17265 -440
rect 17365 -445 17385 -440
rect 17485 -440 17490 -420
rect 17485 -445 17505 -440
rect 17605 -445 17625 -440
rect 17725 -440 17730 -420
rect 17725 -445 17745 -440
rect 17845 -445 17865 -440
rect 17965 -440 17970 -420
rect 17965 -445 17985 -440
rect 18085 -445 18105 -440
rect 18205 -440 18210 -420
rect 18205 -445 18225 -440
rect 18325 -445 18345 -440
rect 18445 -440 18450 -420
rect 18445 -445 18465 -440
rect 18565 -445 18585 -440
rect 18685 -440 18690 -420
rect 18685 -445 18705 -440
rect 18805 -445 18825 -440
rect 18925 -440 18930 -420
rect 18925 -445 18945 -440
rect 19045 -445 19065 -440
rect 19165 -440 19170 -420
rect 19165 -445 19185 -440
rect 19285 -445 19305 -440
rect 19405 -440 19410 -420
rect 19405 -445 19425 -440
rect 19525 -445 19545 -440
rect 19645 -440 19650 -420
rect 19645 -445 19665 -440
rect 19765 -445 19785 -440
rect 19885 -440 19890 -420
rect 19885 -445 19905 -440
rect 20005 -445 20025 -440
rect 20125 -440 20130 -420
rect 20125 -445 20145 -440
rect 20245 -445 20265 -440
rect 20365 -440 20370 -420
rect 20365 -445 20385 -440
rect 20485 -445 20505 -440
rect 20605 -440 20610 -420
rect 20605 -445 20625 -440
rect 20725 -445 20745 -440
rect 20845 -440 20850 -420
rect 20845 -445 20865 -440
rect 20965 -445 20985 -440
rect 21085 -440 21090 -420
rect 21085 -445 21105 -440
rect 21205 -445 21225 -440
rect 21325 -440 21330 -420
rect 21325 -445 21345 -440
rect 21445 -445 21465 -440
rect 21565 -440 21570 -420
rect 21565 -445 21585 -440
rect 21685 -445 21705 -440
rect 21805 -440 21810 -420
rect 21805 -445 21825 -440
rect 21925 -445 21945 -440
rect 22045 -440 22050 -420
rect 22045 -445 22065 -440
rect 22165 -445 22185 -440
rect 22285 -440 22290 -420
rect 22285 -445 22305 -440
rect 22405 -445 22425 -440
rect 22525 -440 22530 -420
rect 22525 -445 22545 -440
rect 22645 -445 22665 -440
rect 22765 -440 22770 -420
rect 22765 -445 22785 -440
rect 22885 -445 22905 -440
rect 23005 -440 23010 -420
rect 23005 -445 23025 -440
rect 23125 -445 23145 -440
rect 23245 -440 23250 -420
rect 23245 -445 23265 -440
rect 23365 -445 23385 -440
rect 23485 -440 23490 -420
rect 23485 -445 23505 -440
rect 23605 -445 23625 -440
rect 23725 -440 23730 -420
rect 23725 -445 23745 -440
rect 23845 -445 23865 -440
rect 23965 -440 23970 -420
rect 23965 -445 23985 -440
rect 24085 -445 24105 -440
rect 24205 -440 24210 -420
rect 24205 -445 24225 -440
rect 24325 -445 24345 -440
rect 24445 -440 24450 -420
rect 24445 -445 24465 -440
rect 24565 -445 24585 -440
rect 24685 -440 24690 -420
rect 24685 -445 24705 -440
rect 24805 -445 24825 -440
rect 24925 -440 24930 -420
rect 24925 -445 24945 -440
rect 25045 -445 25065 -440
rect 25165 -440 25170 -420
rect 25165 -445 25185 -440
rect 25285 -445 25305 -440
rect 25405 -440 25410 -420
rect 25405 -445 25425 -440
rect 25525 -445 25545 -440
rect 25645 -440 25650 -420
rect 25645 -445 25665 -440
rect 25765 -445 25785 -440
rect 25885 -440 25890 -420
rect 25885 -445 25905 -440
rect 26005 -445 26025 -440
rect 26125 -440 26130 -420
rect 26125 -445 26145 -440
rect 26245 -445 26265 -440
rect 26365 -440 26370 -420
rect 26365 -445 26385 -440
rect 26485 -445 26505 -440
rect 26605 -440 26610 -420
rect 26605 -445 26625 -440
rect 26725 -445 26745 -440
rect 26845 -440 26850 -420
rect 26845 -445 26865 -440
rect 26965 -445 26985 -440
rect 27085 -440 27090 -420
rect 27085 -445 27105 -440
rect 27205 -445 27225 -440
rect 27325 -440 27330 -420
rect 27325 -445 27345 -440
rect 27445 -445 27465 -440
rect 27565 -440 27570 -420
rect 27565 -445 27585 -440
rect 27685 -445 27705 -440
rect 27805 -440 27810 -420
rect 27805 -445 27825 -440
rect 27925 -445 27945 -440
rect 28045 -440 28050 -420
rect 28045 -445 28065 -440
rect 28165 -445 28185 -440
rect 28285 -440 28290 -420
rect 28285 -445 28305 -440
rect 28405 -445 28425 -440
rect 28525 -440 28530 -420
rect 28525 -445 28545 -440
rect 28645 -445 28665 -440
rect 28765 -440 28770 -420
rect 28765 -445 28785 -440
rect 28885 -445 28905 -440
rect 29005 -440 29010 -420
rect 29005 -445 29025 -440
rect 29125 -445 29145 -440
rect 29245 -440 29250 -420
rect 29245 -445 29265 -440
rect 29365 -445 29385 -440
rect 29485 -440 29490 -420
rect 29485 -445 29505 -440
rect 29605 -445 29625 -440
rect 29725 -440 29730 -420
rect 29725 -445 29745 -440
rect 29845 -445 29865 -440
rect 29965 -440 29970 -420
rect 29965 -445 29985 -440
rect 30085 -445 30105 -440
rect 30205 -440 30210 -420
rect 30205 -445 30225 -440
rect 30325 -445 30345 -440
rect 30445 -440 30450 -420
rect 30445 -445 30465 -440
rect 30565 -445 30585 -440
rect 30685 -425 30705 -420
rect -190 -515 50 -495
rect 30675 -485 30715 -475
rect 30675 -505 30685 -485
rect 30705 -505 30740 -485
rect 30675 -515 30715 -505
rect -460 -655 -440 -555
rect -340 -655 -320 -555
rect -30 -575 -10 -565
rect 25 -575 50 -515
rect 90 -575 110 -565
rect 205 -565 210 -545
rect 205 -575 230 -565
rect 330 -575 350 -565
rect 445 -565 450 -545
rect 445 -575 470 -565
rect 570 -575 590 -565
rect 685 -565 690 -545
rect 685 -575 710 -565
rect 810 -575 830 -565
rect 925 -565 930 -545
rect 925 -575 950 -565
rect 1050 -575 1070 -565
rect 1165 -565 1170 -545
rect 1165 -575 1190 -565
rect 1290 -575 1310 -565
rect 1405 -565 1410 -545
rect 1405 -575 1430 -565
rect 1530 -575 1550 -565
rect 1645 -565 1650 -545
rect 1645 -575 1670 -565
rect 1770 -575 1790 -565
rect 1885 -565 1890 -545
rect 1885 -575 1910 -565
rect 2010 -575 2030 -565
rect 2125 -565 2130 -545
rect 2125 -575 2150 -565
rect 2250 -575 2270 -565
rect 2365 -565 2370 -545
rect 2365 -575 2390 -565
rect 2490 -575 2510 -565
rect 2605 -565 2610 -545
rect 2605 -575 2630 -565
rect 2730 -575 2750 -565
rect 2845 -565 2850 -545
rect 2845 -575 2870 -565
rect 2970 -575 2990 -565
rect 3085 -565 3090 -545
rect 3085 -575 3110 -565
rect 3210 -575 3230 -565
rect 3325 -565 3330 -545
rect 3325 -575 3350 -565
rect 3450 -575 3470 -565
rect 3565 -565 3570 -545
rect 3565 -575 3590 -565
rect 3690 -575 3710 -565
rect 3805 -565 3810 -545
rect 3805 -575 3830 -565
rect 3930 -575 3950 -565
rect 4045 -565 4050 -545
rect 4045 -575 4070 -565
rect 4170 -575 4190 -565
rect 4285 -565 4290 -545
rect 4285 -575 4310 -565
rect 4410 -575 4430 -565
rect 4525 -565 4530 -545
rect 4525 -575 4550 -565
rect 4650 -575 4670 -565
rect 4765 -565 4770 -545
rect 4765 -575 4790 -565
rect 4890 -575 4910 -565
rect 5005 -565 5010 -545
rect 5005 -575 5030 -565
rect 5130 -575 5150 -565
rect 5245 -565 5250 -545
rect 5245 -575 5270 -565
rect 5370 -575 5390 -565
rect 5485 -565 5490 -545
rect 5485 -575 5510 -565
rect 5610 -575 5630 -565
rect 5725 -565 5730 -545
rect 5725 -575 5750 -565
rect 5850 -575 5870 -565
rect 5965 -565 5970 -545
rect 5965 -575 5990 -565
rect 6090 -575 6110 -565
rect 6205 -565 6210 -545
rect 6205 -575 6230 -565
rect 6330 -575 6350 -565
rect 6445 -565 6450 -545
rect 6445 -575 6470 -565
rect 6570 -575 6590 -565
rect 6685 -565 6690 -545
rect 6685 -575 6710 -565
rect 6810 -575 6830 -565
rect 6925 -565 6930 -545
rect 6925 -575 6950 -565
rect 7050 -575 7070 -565
rect 7165 -565 7170 -545
rect 7165 -575 7190 -565
rect 7290 -575 7310 -565
rect 7405 -565 7410 -545
rect 7405 -575 7430 -565
rect 7530 -575 7550 -565
rect 7645 -565 7650 -545
rect 7645 -575 7670 -565
rect 7770 -575 7790 -565
rect 7885 -565 7890 -545
rect 7885 -575 7910 -565
rect 8010 -575 8030 -565
rect 8125 -565 8130 -545
rect 8125 -575 8150 -565
rect 8250 -575 8270 -565
rect 8365 -565 8370 -545
rect 8365 -575 8390 -565
rect 8490 -575 8510 -565
rect 8605 -565 8610 -545
rect 8605 -575 8630 -565
rect 8730 -575 8750 -565
rect 8845 -565 8850 -545
rect 8845 -575 8870 -565
rect 8970 -575 8990 -565
rect 9085 -565 9090 -545
rect 9085 -575 9110 -565
rect 9210 -575 9230 -565
rect 9325 -565 9330 -545
rect 9325 -575 9350 -565
rect 9450 -575 9470 -565
rect 9565 -565 9570 -545
rect 9565 -575 9590 -565
rect 9690 -575 9710 -565
rect 9805 -565 9810 -545
rect 9805 -575 9830 -565
rect 9930 -575 9950 -565
rect 10045 -565 10050 -545
rect 10045 -575 10070 -565
rect 10170 -575 10190 -565
rect 10285 -565 10290 -545
rect 10285 -575 10310 -565
rect 10410 -575 10430 -565
rect 10525 -565 10530 -545
rect 10525 -575 10550 -565
rect 10650 -575 10670 -565
rect 10765 -565 10770 -545
rect 10765 -575 10790 -565
rect 10890 -575 10910 -565
rect 11005 -565 11010 -545
rect 11005 -575 11030 -565
rect 11130 -575 11150 -565
rect 11245 -565 11250 -545
rect 11245 -575 11270 -565
rect 11370 -575 11390 -565
rect 11485 -565 11490 -545
rect 11485 -575 11510 -565
rect 11610 -575 11630 -565
rect 11725 -565 11730 -545
rect 11725 -575 11750 -565
rect 11850 -575 11870 -565
rect 11965 -565 11970 -545
rect 11965 -575 11990 -565
rect 12090 -575 12110 -565
rect 12205 -565 12210 -545
rect 12205 -575 12230 -565
rect 12330 -575 12350 -565
rect 12445 -565 12450 -545
rect 12445 -575 12470 -565
rect 12570 -575 12590 -565
rect 12685 -565 12690 -545
rect 12685 -575 12710 -565
rect 12810 -575 12830 -565
rect 12925 -565 12930 -545
rect 12925 -575 12950 -565
rect 13050 -575 13070 -565
rect 13165 -565 13170 -545
rect 13165 -575 13190 -565
rect 13290 -575 13310 -565
rect 13405 -565 13410 -545
rect 13405 -575 13430 -565
rect 13530 -575 13550 -565
rect 13645 -565 13650 -545
rect 13645 -575 13670 -565
rect 13770 -575 13790 -565
rect 13885 -565 13890 -545
rect 13885 -575 13910 -565
rect 14010 -575 14030 -565
rect 14125 -565 14130 -545
rect 14125 -575 14150 -565
rect 14250 -575 14270 -565
rect 14365 -565 14370 -545
rect 14365 -575 14390 -565
rect 14490 -575 14510 -565
rect 14605 -565 14610 -545
rect 14605 -575 14630 -565
rect 14730 -575 14750 -565
rect 14845 -565 14850 -545
rect 14845 -575 14870 -565
rect 14970 -575 14990 -565
rect 15085 -565 15090 -545
rect 15085 -575 15110 -565
rect 15210 -575 15230 -565
rect 15325 -565 15330 -545
rect 15325 -575 15350 -565
rect 15450 -575 15470 -565
rect 15565 -565 15570 -545
rect 15565 -575 15590 -565
rect 15690 -575 15710 -565
rect 15805 -565 15810 -545
rect 15805 -575 15830 -565
rect 15930 -575 15950 -565
rect 16045 -565 16050 -545
rect 16045 -575 16070 -565
rect 16170 -575 16190 -565
rect 16285 -565 16290 -545
rect 16285 -575 16310 -565
rect 16410 -575 16430 -565
rect 16525 -565 16530 -545
rect 16525 -575 16550 -565
rect 16650 -575 16670 -565
rect 16765 -565 16770 -545
rect 16765 -575 16790 -565
rect 16890 -575 16910 -565
rect 17005 -565 17010 -545
rect 17005 -575 17030 -565
rect 17130 -575 17150 -565
rect 17245 -565 17250 -545
rect 17245 -575 17270 -565
rect 17370 -575 17390 -565
rect 17485 -565 17490 -545
rect 17485 -575 17510 -565
rect 17610 -575 17630 -565
rect 17725 -565 17730 -545
rect 17725 -575 17750 -565
rect 17850 -575 17870 -565
rect 17965 -565 17970 -545
rect 17965 -575 17990 -565
rect 18090 -575 18110 -565
rect 18205 -565 18210 -545
rect 18205 -575 18230 -565
rect 18330 -575 18350 -565
rect 18445 -565 18450 -545
rect 18445 -575 18470 -565
rect 18570 -575 18590 -565
rect 18685 -565 18690 -545
rect 18685 -575 18710 -565
rect 18810 -575 18830 -565
rect 18925 -565 18930 -545
rect 18925 -575 18950 -565
rect 19050 -575 19070 -565
rect 19165 -565 19170 -545
rect 19165 -575 19190 -565
rect 19290 -575 19310 -565
rect 19405 -565 19410 -545
rect 19405 -575 19430 -565
rect 19530 -575 19550 -565
rect 19645 -565 19650 -545
rect 19645 -575 19670 -565
rect 19770 -575 19790 -565
rect 19885 -565 19890 -545
rect 19885 -575 19910 -565
rect 20010 -575 20030 -565
rect 20125 -565 20130 -545
rect 20125 -575 20150 -565
rect 20250 -575 20270 -565
rect 20365 -565 20370 -545
rect 20365 -575 20390 -565
rect 20490 -575 20510 -565
rect 20605 -565 20610 -545
rect 20605 -575 20630 -565
rect 20730 -575 20750 -565
rect 20845 -565 20850 -545
rect 20845 -575 20870 -565
rect 20970 -575 20990 -565
rect 21085 -565 21090 -545
rect 21085 -575 21110 -565
rect 21210 -575 21230 -565
rect 21325 -565 21330 -545
rect 21325 -575 21350 -565
rect 21450 -575 21470 -565
rect 21565 -565 21570 -545
rect 21565 -575 21590 -565
rect 21690 -575 21710 -565
rect 21805 -565 21810 -545
rect 21805 -575 21830 -565
rect 21930 -575 21950 -565
rect 22045 -565 22050 -545
rect 22045 -575 22070 -565
rect 22170 -575 22190 -565
rect 22285 -565 22290 -545
rect 22285 -575 22310 -565
rect 22410 -575 22430 -565
rect 22525 -565 22530 -545
rect 22525 -575 22550 -565
rect 22650 -575 22670 -565
rect 22765 -565 22770 -545
rect 22765 -575 22790 -565
rect 22890 -575 22910 -565
rect 23005 -565 23010 -545
rect 23005 -575 23030 -565
rect 23130 -575 23150 -565
rect 23245 -565 23250 -545
rect 23245 -575 23270 -565
rect 23370 -575 23390 -565
rect 23485 -565 23490 -545
rect 23485 -575 23510 -565
rect 23610 -575 23630 -565
rect 23725 -565 23730 -545
rect 23725 -575 23750 -565
rect 23850 -575 23870 -565
rect 23965 -565 23970 -545
rect 23965 -575 23990 -565
rect 24090 -575 24110 -565
rect 24205 -565 24210 -545
rect 24205 -575 24230 -565
rect 24330 -575 24350 -565
rect 24445 -565 24450 -545
rect 24445 -575 24470 -565
rect 24570 -575 24590 -565
rect 24685 -565 24690 -545
rect 24685 -575 24710 -565
rect 24810 -575 24830 -565
rect 24925 -565 24930 -545
rect 24925 -575 24950 -565
rect 25050 -575 25070 -565
rect 25165 -565 25170 -545
rect 25165 -575 25190 -565
rect 25290 -575 25310 -565
rect 25405 -565 25410 -545
rect 25405 -575 25430 -565
rect 25530 -575 25550 -565
rect 25645 -565 25650 -545
rect 25645 -575 25670 -565
rect 25770 -575 25790 -565
rect 25885 -565 25890 -545
rect 25885 -575 25910 -565
rect 26010 -575 26030 -565
rect 26125 -565 26130 -545
rect 26125 -575 26150 -565
rect 26250 -575 26270 -565
rect 26365 -565 26370 -545
rect 26365 -575 26390 -565
rect 26490 -575 26510 -565
rect 26605 -565 26610 -545
rect 26605 -575 26630 -565
rect 26730 -575 26750 -565
rect 26845 -565 26850 -545
rect 26845 -575 26870 -565
rect 26970 -575 26990 -565
rect 27085 -565 27090 -545
rect 27085 -575 27110 -565
rect 27210 -575 27230 -565
rect 27325 -565 27330 -545
rect 27325 -575 27350 -565
rect 27450 -575 27470 -565
rect 27565 -565 27570 -545
rect 27565 -575 27590 -565
rect 27690 -575 27710 -565
rect 27805 -565 27810 -545
rect 27805 -575 27830 -565
rect 27930 -575 27950 -565
rect 28045 -565 28050 -545
rect 28045 -575 28070 -565
rect 28170 -575 28190 -565
rect 28285 -565 28290 -545
rect 28285 -575 28310 -565
rect 28410 -575 28430 -565
rect 28525 -565 28530 -545
rect 28525 -575 28550 -565
rect 28650 -575 28670 -565
rect 28765 -565 28770 -545
rect 28765 -575 28790 -565
rect 28890 -575 28910 -565
rect 29005 -565 29010 -545
rect 29005 -575 29030 -565
rect 29130 -575 29150 -565
rect 29245 -565 29250 -545
rect 29245 -575 29270 -565
rect 29370 -575 29390 -565
rect 29485 -565 29490 -545
rect 29485 -575 29510 -565
rect 29610 -575 29630 -565
rect 29725 -565 29730 -545
rect 29725 -575 29750 -565
rect 29850 -575 29870 -565
rect 29965 -565 29970 -545
rect 29965 -575 29990 -565
rect 30090 -575 30110 -565
rect 30205 -565 30210 -545
rect 30205 -575 30230 -565
rect 30330 -575 30350 -565
rect 30445 -565 30450 -545
rect 30445 -575 30470 -565
rect 30570 -575 30590 -565
rect 30685 -575 30705 -565
rect -460 -945 -320 -655
rect -40 -585 -5 -575
rect -40 -610 -35 -585
rect -10 -610 -5 -585
rect -40 -630 -5 -610
rect -40 -655 -35 -630
rect -10 -655 -5 -630
rect -40 -675 -5 -655
rect -40 -700 -35 -675
rect -10 -700 -5 -675
rect -40 -725 -5 -700
rect -40 -750 -35 -725
rect -10 -750 -5 -725
rect -40 -770 -5 -750
rect 20 -585 55 -575
rect 20 -610 25 -585
rect 50 -610 55 -585
rect 20 -630 55 -610
rect 20 -655 25 -630
rect 50 -655 55 -630
rect 20 -675 55 -655
rect 20 -700 25 -675
rect 50 -700 55 -675
rect 20 -725 55 -700
rect 20 -750 25 -725
rect 50 -750 55 -725
rect 20 -770 55 -750
rect 80 -585 115 -575
rect 80 -610 85 -585
rect 110 -610 115 -585
rect 80 -630 115 -610
rect 80 -655 85 -630
rect 110 -655 115 -630
rect 80 -675 115 -655
rect 80 -700 85 -675
rect 110 -700 115 -675
rect 80 -725 115 -700
rect 80 -750 85 -725
rect 110 -750 115 -725
rect 80 -770 115 -750
rect 140 -585 175 -575
rect 140 -610 145 -585
rect 170 -610 175 -585
rect 140 -630 175 -610
rect 140 -655 145 -630
rect 170 -655 175 -630
rect 140 -675 175 -655
rect 140 -700 145 -675
rect 170 -700 175 -675
rect 140 -725 175 -700
rect 140 -750 145 -725
rect 170 -750 175 -725
rect 140 -770 175 -750
rect 200 -585 235 -575
rect 200 -610 205 -585
rect 230 -610 235 -585
rect 200 -630 235 -610
rect 200 -655 205 -630
rect 230 -655 235 -630
rect 200 -675 235 -655
rect 200 -700 205 -675
rect 230 -700 235 -675
rect 200 -725 235 -700
rect 200 -750 205 -725
rect 230 -750 235 -725
rect 200 -770 235 -750
rect 260 -585 295 -575
rect 260 -610 265 -585
rect 290 -610 295 -585
rect 260 -630 295 -610
rect 260 -655 265 -630
rect 290 -655 295 -630
rect 260 -675 295 -655
rect 260 -700 265 -675
rect 290 -700 295 -675
rect 260 -725 295 -700
rect 260 -750 265 -725
rect 290 -750 295 -725
rect 260 -770 295 -750
rect 320 -585 355 -575
rect 320 -610 325 -585
rect 350 -610 355 -585
rect 320 -630 355 -610
rect 320 -655 325 -630
rect 350 -655 355 -630
rect 320 -675 355 -655
rect 320 -700 325 -675
rect 350 -700 355 -675
rect 320 -725 355 -700
rect 320 -750 325 -725
rect 350 -750 355 -725
rect 320 -770 355 -750
rect 380 -585 415 -575
rect 380 -610 385 -585
rect 410 -610 415 -585
rect 380 -630 415 -610
rect 380 -655 385 -630
rect 410 -655 415 -630
rect 380 -675 415 -655
rect 380 -700 385 -675
rect 410 -700 415 -675
rect 380 -725 415 -700
rect 380 -750 385 -725
rect 410 -750 415 -725
rect 380 -770 415 -750
rect 440 -585 475 -575
rect 440 -610 445 -585
rect 470 -610 475 -585
rect 440 -630 475 -610
rect 440 -655 445 -630
rect 470 -655 475 -630
rect 440 -675 475 -655
rect 440 -700 445 -675
rect 470 -700 475 -675
rect 440 -725 475 -700
rect 440 -750 445 -725
rect 470 -750 475 -725
rect 440 -770 475 -750
rect 500 -585 535 -575
rect 500 -610 505 -585
rect 530 -610 535 -585
rect 500 -630 535 -610
rect 500 -655 505 -630
rect 530 -655 535 -630
rect 500 -675 535 -655
rect 500 -700 505 -675
rect 530 -700 535 -675
rect 500 -725 535 -700
rect 500 -750 505 -725
rect 530 -750 535 -725
rect 500 -770 535 -750
rect 560 -585 595 -575
rect 560 -610 565 -585
rect 590 -610 595 -585
rect 560 -630 595 -610
rect 560 -655 565 -630
rect 590 -655 595 -630
rect 560 -675 595 -655
rect 560 -700 565 -675
rect 590 -700 595 -675
rect 560 -725 595 -700
rect 560 -750 565 -725
rect 590 -750 595 -725
rect 560 -770 595 -750
rect 620 -585 655 -575
rect 620 -610 625 -585
rect 650 -610 655 -585
rect 620 -630 655 -610
rect 620 -655 625 -630
rect 650 -655 655 -630
rect 620 -675 655 -655
rect 620 -700 625 -675
rect 650 -700 655 -675
rect 620 -725 655 -700
rect 620 -750 625 -725
rect 650 -750 655 -725
rect 620 -770 655 -750
rect 680 -585 715 -575
rect 680 -610 685 -585
rect 710 -610 715 -585
rect 680 -630 715 -610
rect 680 -655 685 -630
rect 710 -655 715 -630
rect 680 -675 715 -655
rect 680 -700 685 -675
rect 710 -700 715 -675
rect 680 -725 715 -700
rect 680 -750 685 -725
rect 710 -750 715 -725
rect 680 -770 715 -750
rect 740 -585 775 -575
rect 740 -610 745 -585
rect 770 -610 775 -585
rect 740 -630 775 -610
rect 740 -655 745 -630
rect 770 -655 775 -630
rect 740 -675 775 -655
rect 740 -700 745 -675
rect 770 -700 775 -675
rect 740 -725 775 -700
rect 740 -750 745 -725
rect 770 -750 775 -725
rect 740 -770 775 -750
rect 800 -585 835 -575
rect 800 -610 805 -585
rect 830 -610 835 -585
rect 800 -630 835 -610
rect 800 -655 805 -630
rect 830 -655 835 -630
rect 800 -675 835 -655
rect 800 -700 805 -675
rect 830 -700 835 -675
rect 800 -725 835 -700
rect 800 -750 805 -725
rect 830 -750 835 -725
rect 800 -770 835 -750
rect 860 -585 895 -575
rect 860 -610 865 -585
rect 890 -610 895 -585
rect 860 -630 895 -610
rect 860 -655 865 -630
rect 890 -655 895 -630
rect 860 -675 895 -655
rect 860 -700 865 -675
rect 890 -700 895 -675
rect 860 -725 895 -700
rect 860 -750 865 -725
rect 890 -750 895 -725
rect 860 -770 895 -750
rect 920 -585 955 -575
rect 920 -610 925 -585
rect 950 -610 955 -585
rect 920 -630 955 -610
rect 920 -655 925 -630
rect 950 -655 955 -630
rect 920 -675 955 -655
rect 920 -700 925 -675
rect 950 -700 955 -675
rect 920 -725 955 -700
rect 920 -750 925 -725
rect 950 -750 955 -725
rect 920 -770 955 -750
rect 980 -585 1015 -575
rect 980 -610 985 -585
rect 1010 -610 1015 -585
rect 980 -630 1015 -610
rect 980 -655 985 -630
rect 1010 -655 1015 -630
rect 980 -675 1015 -655
rect 980 -700 985 -675
rect 1010 -700 1015 -675
rect 980 -725 1015 -700
rect 980 -750 985 -725
rect 1010 -750 1015 -725
rect 980 -770 1015 -750
rect 1040 -585 1075 -575
rect 1040 -610 1045 -585
rect 1070 -610 1075 -585
rect 1040 -630 1075 -610
rect 1040 -655 1045 -630
rect 1070 -655 1075 -630
rect 1040 -675 1075 -655
rect 1040 -700 1045 -675
rect 1070 -700 1075 -675
rect 1040 -725 1075 -700
rect 1040 -750 1045 -725
rect 1070 -750 1075 -725
rect 1040 -770 1075 -750
rect 1100 -585 1135 -575
rect 1100 -610 1105 -585
rect 1130 -610 1135 -585
rect 1100 -630 1135 -610
rect 1100 -655 1105 -630
rect 1130 -655 1135 -630
rect 1100 -675 1135 -655
rect 1100 -700 1105 -675
rect 1130 -700 1135 -675
rect 1100 -725 1135 -700
rect 1100 -750 1105 -725
rect 1130 -750 1135 -725
rect 1100 -770 1135 -750
rect 1160 -585 1195 -575
rect 1160 -610 1165 -585
rect 1190 -610 1195 -585
rect 1160 -630 1195 -610
rect 1160 -655 1165 -630
rect 1190 -655 1195 -630
rect 1160 -675 1195 -655
rect 1160 -700 1165 -675
rect 1190 -700 1195 -675
rect 1160 -725 1195 -700
rect 1160 -750 1165 -725
rect 1190 -750 1195 -725
rect 1160 -770 1195 -750
rect 1220 -585 1255 -575
rect 1220 -610 1225 -585
rect 1250 -610 1255 -585
rect 1220 -630 1255 -610
rect 1220 -655 1225 -630
rect 1250 -655 1255 -630
rect 1220 -675 1255 -655
rect 1220 -700 1225 -675
rect 1250 -700 1255 -675
rect 1220 -725 1255 -700
rect 1220 -750 1225 -725
rect 1250 -750 1255 -725
rect 1220 -770 1255 -750
rect 1280 -585 1315 -575
rect 1280 -610 1285 -585
rect 1310 -610 1315 -585
rect 1280 -630 1315 -610
rect 1280 -655 1285 -630
rect 1310 -655 1315 -630
rect 1280 -675 1315 -655
rect 1280 -700 1285 -675
rect 1310 -700 1315 -675
rect 1280 -725 1315 -700
rect 1280 -750 1285 -725
rect 1310 -750 1315 -725
rect 1280 -770 1315 -750
rect 1340 -585 1375 -575
rect 1340 -610 1345 -585
rect 1370 -610 1375 -585
rect 1340 -630 1375 -610
rect 1340 -655 1345 -630
rect 1370 -655 1375 -630
rect 1340 -675 1375 -655
rect 1340 -700 1345 -675
rect 1370 -700 1375 -675
rect 1340 -725 1375 -700
rect 1340 -750 1345 -725
rect 1370 -750 1375 -725
rect 1340 -770 1375 -750
rect 1400 -585 1435 -575
rect 1400 -610 1405 -585
rect 1430 -610 1435 -585
rect 1400 -630 1435 -610
rect 1400 -655 1405 -630
rect 1430 -655 1435 -630
rect 1400 -675 1435 -655
rect 1400 -700 1405 -675
rect 1430 -700 1435 -675
rect 1400 -725 1435 -700
rect 1400 -750 1405 -725
rect 1430 -750 1435 -725
rect 1400 -770 1435 -750
rect 1460 -585 1495 -575
rect 1460 -610 1465 -585
rect 1490 -610 1495 -585
rect 1460 -630 1495 -610
rect 1460 -655 1465 -630
rect 1490 -655 1495 -630
rect 1460 -675 1495 -655
rect 1460 -700 1465 -675
rect 1490 -700 1495 -675
rect 1460 -725 1495 -700
rect 1460 -750 1465 -725
rect 1490 -750 1495 -725
rect 1460 -770 1495 -750
rect 1520 -585 1555 -575
rect 1520 -610 1525 -585
rect 1550 -610 1555 -585
rect 1520 -630 1555 -610
rect 1520 -655 1525 -630
rect 1550 -655 1555 -630
rect 1520 -675 1555 -655
rect 1520 -700 1525 -675
rect 1550 -700 1555 -675
rect 1520 -725 1555 -700
rect 1520 -750 1525 -725
rect 1550 -750 1555 -725
rect 1520 -770 1555 -750
rect 1580 -585 1615 -575
rect 1580 -610 1585 -585
rect 1610 -610 1615 -585
rect 1580 -630 1615 -610
rect 1580 -655 1585 -630
rect 1610 -655 1615 -630
rect 1580 -675 1615 -655
rect 1580 -700 1585 -675
rect 1610 -700 1615 -675
rect 1580 -725 1615 -700
rect 1580 -750 1585 -725
rect 1610 -750 1615 -725
rect 1580 -770 1615 -750
rect 1640 -585 1675 -575
rect 1640 -610 1645 -585
rect 1670 -610 1675 -585
rect 1640 -630 1675 -610
rect 1640 -655 1645 -630
rect 1670 -655 1675 -630
rect 1640 -675 1675 -655
rect 1640 -700 1645 -675
rect 1670 -700 1675 -675
rect 1640 -725 1675 -700
rect 1640 -750 1645 -725
rect 1670 -750 1675 -725
rect 1640 -770 1675 -750
rect 1700 -585 1735 -575
rect 1700 -610 1705 -585
rect 1730 -610 1735 -585
rect 1700 -630 1735 -610
rect 1700 -655 1705 -630
rect 1730 -655 1735 -630
rect 1700 -675 1735 -655
rect 1700 -700 1705 -675
rect 1730 -700 1735 -675
rect 1700 -725 1735 -700
rect 1700 -750 1705 -725
rect 1730 -750 1735 -725
rect 1700 -770 1735 -750
rect 1760 -585 1795 -575
rect 1760 -610 1765 -585
rect 1790 -610 1795 -585
rect 1760 -630 1795 -610
rect 1760 -655 1765 -630
rect 1790 -655 1795 -630
rect 1760 -675 1795 -655
rect 1760 -700 1765 -675
rect 1790 -700 1795 -675
rect 1760 -725 1795 -700
rect 1760 -750 1765 -725
rect 1790 -750 1795 -725
rect 1760 -770 1795 -750
rect 1820 -585 1855 -575
rect 1820 -610 1825 -585
rect 1850 -610 1855 -585
rect 1820 -630 1855 -610
rect 1820 -655 1825 -630
rect 1850 -655 1855 -630
rect 1820 -675 1855 -655
rect 1820 -700 1825 -675
rect 1850 -700 1855 -675
rect 1820 -725 1855 -700
rect 1820 -750 1825 -725
rect 1850 -750 1855 -725
rect 1820 -770 1855 -750
rect 1880 -585 1915 -575
rect 1880 -610 1885 -585
rect 1910 -610 1915 -585
rect 1880 -630 1915 -610
rect 1880 -655 1885 -630
rect 1910 -655 1915 -630
rect 1880 -675 1915 -655
rect 1880 -700 1885 -675
rect 1910 -700 1915 -675
rect 1880 -725 1915 -700
rect 1880 -750 1885 -725
rect 1910 -750 1915 -725
rect 1880 -770 1915 -750
rect 1940 -585 1975 -575
rect 1940 -610 1945 -585
rect 1970 -610 1975 -585
rect 1940 -630 1975 -610
rect 1940 -655 1945 -630
rect 1970 -655 1975 -630
rect 1940 -675 1975 -655
rect 1940 -700 1945 -675
rect 1970 -700 1975 -675
rect 1940 -725 1975 -700
rect 1940 -750 1945 -725
rect 1970 -750 1975 -725
rect 1940 -770 1975 -750
rect 2000 -585 2035 -575
rect 2000 -610 2005 -585
rect 2030 -610 2035 -585
rect 2000 -630 2035 -610
rect 2000 -655 2005 -630
rect 2030 -655 2035 -630
rect 2000 -675 2035 -655
rect 2000 -700 2005 -675
rect 2030 -700 2035 -675
rect 2000 -725 2035 -700
rect 2000 -750 2005 -725
rect 2030 -750 2035 -725
rect 2000 -770 2035 -750
rect 2060 -585 2095 -575
rect 2060 -610 2065 -585
rect 2090 -610 2095 -585
rect 2060 -630 2095 -610
rect 2060 -655 2065 -630
rect 2090 -655 2095 -630
rect 2060 -675 2095 -655
rect 2060 -700 2065 -675
rect 2090 -700 2095 -675
rect 2060 -725 2095 -700
rect 2060 -750 2065 -725
rect 2090 -750 2095 -725
rect 2060 -770 2095 -750
rect 2120 -585 2155 -575
rect 2120 -610 2125 -585
rect 2150 -610 2155 -585
rect 2120 -630 2155 -610
rect 2120 -655 2125 -630
rect 2150 -655 2155 -630
rect 2120 -675 2155 -655
rect 2120 -700 2125 -675
rect 2150 -700 2155 -675
rect 2120 -725 2155 -700
rect 2120 -750 2125 -725
rect 2150 -750 2155 -725
rect 2120 -770 2155 -750
rect 2180 -585 2215 -575
rect 2180 -610 2185 -585
rect 2210 -610 2215 -585
rect 2180 -630 2215 -610
rect 2180 -655 2185 -630
rect 2210 -655 2215 -630
rect 2180 -675 2215 -655
rect 2180 -700 2185 -675
rect 2210 -700 2215 -675
rect 2180 -725 2215 -700
rect 2180 -750 2185 -725
rect 2210 -750 2215 -725
rect 2180 -770 2215 -750
rect 2240 -585 2275 -575
rect 2240 -610 2245 -585
rect 2270 -610 2275 -585
rect 2240 -630 2275 -610
rect 2240 -655 2245 -630
rect 2270 -655 2275 -630
rect 2240 -675 2275 -655
rect 2240 -700 2245 -675
rect 2270 -700 2275 -675
rect 2240 -725 2275 -700
rect 2240 -750 2245 -725
rect 2270 -750 2275 -725
rect 2240 -770 2275 -750
rect 2300 -585 2335 -575
rect 2300 -610 2305 -585
rect 2330 -610 2335 -585
rect 2300 -630 2335 -610
rect 2300 -655 2305 -630
rect 2330 -655 2335 -630
rect 2300 -675 2335 -655
rect 2300 -700 2305 -675
rect 2330 -700 2335 -675
rect 2300 -725 2335 -700
rect 2300 -750 2305 -725
rect 2330 -750 2335 -725
rect 2300 -770 2335 -750
rect 2360 -585 2395 -575
rect 2360 -610 2365 -585
rect 2390 -610 2395 -585
rect 2360 -630 2395 -610
rect 2360 -655 2365 -630
rect 2390 -655 2395 -630
rect 2360 -675 2395 -655
rect 2360 -700 2365 -675
rect 2390 -700 2395 -675
rect 2360 -725 2395 -700
rect 2360 -750 2365 -725
rect 2390 -750 2395 -725
rect 2360 -770 2395 -750
rect 2420 -585 2455 -575
rect 2420 -610 2425 -585
rect 2450 -610 2455 -585
rect 2420 -630 2455 -610
rect 2420 -655 2425 -630
rect 2450 -655 2455 -630
rect 2420 -675 2455 -655
rect 2420 -700 2425 -675
rect 2450 -700 2455 -675
rect 2420 -725 2455 -700
rect 2420 -750 2425 -725
rect 2450 -750 2455 -725
rect 2420 -770 2455 -750
rect 2480 -585 2515 -575
rect 2480 -610 2485 -585
rect 2510 -610 2515 -585
rect 2480 -630 2515 -610
rect 2480 -655 2485 -630
rect 2510 -655 2515 -630
rect 2480 -675 2515 -655
rect 2480 -700 2485 -675
rect 2510 -700 2515 -675
rect 2480 -725 2515 -700
rect 2480 -750 2485 -725
rect 2510 -750 2515 -725
rect 2480 -770 2515 -750
rect 2540 -585 2575 -575
rect 2540 -610 2545 -585
rect 2570 -610 2575 -585
rect 2540 -630 2575 -610
rect 2540 -655 2545 -630
rect 2570 -655 2575 -630
rect 2540 -675 2575 -655
rect 2540 -700 2545 -675
rect 2570 -700 2575 -675
rect 2540 -725 2575 -700
rect 2540 -750 2545 -725
rect 2570 -750 2575 -725
rect 2540 -770 2575 -750
rect 2600 -585 2635 -575
rect 2600 -610 2605 -585
rect 2630 -610 2635 -585
rect 2600 -630 2635 -610
rect 2600 -655 2605 -630
rect 2630 -655 2635 -630
rect 2600 -675 2635 -655
rect 2600 -700 2605 -675
rect 2630 -700 2635 -675
rect 2600 -725 2635 -700
rect 2600 -750 2605 -725
rect 2630 -750 2635 -725
rect 2600 -770 2635 -750
rect 2660 -585 2695 -575
rect 2660 -610 2665 -585
rect 2690 -610 2695 -585
rect 2660 -630 2695 -610
rect 2660 -655 2665 -630
rect 2690 -655 2695 -630
rect 2660 -675 2695 -655
rect 2660 -700 2665 -675
rect 2690 -700 2695 -675
rect 2660 -725 2695 -700
rect 2660 -750 2665 -725
rect 2690 -750 2695 -725
rect 2660 -770 2695 -750
rect 2720 -585 2755 -575
rect 2720 -610 2725 -585
rect 2750 -610 2755 -585
rect 2720 -630 2755 -610
rect 2720 -655 2725 -630
rect 2750 -655 2755 -630
rect 2720 -675 2755 -655
rect 2720 -700 2725 -675
rect 2750 -700 2755 -675
rect 2720 -725 2755 -700
rect 2720 -750 2725 -725
rect 2750 -750 2755 -725
rect 2720 -770 2755 -750
rect 2780 -585 2815 -575
rect 2780 -610 2785 -585
rect 2810 -610 2815 -585
rect 2780 -630 2815 -610
rect 2780 -655 2785 -630
rect 2810 -655 2815 -630
rect 2780 -675 2815 -655
rect 2780 -700 2785 -675
rect 2810 -700 2815 -675
rect 2780 -725 2815 -700
rect 2780 -750 2785 -725
rect 2810 -750 2815 -725
rect 2780 -770 2815 -750
rect 2840 -585 2875 -575
rect 2840 -610 2845 -585
rect 2870 -610 2875 -585
rect 2840 -630 2875 -610
rect 2840 -655 2845 -630
rect 2870 -655 2875 -630
rect 2840 -675 2875 -655
rect 2840 -700 2845 -675
rect 2870 -700 2875 -675
rect 2840 -725 2875 -700
rect 2840 -750 2845 -725
rect 2870 -750 2875 -725
rect 2840 -770 2875 -750
rect 2900 -585 2935 -575
rect 2900 -610 2905 -585
rect 2930 -610 2935 -585
rect 2900 -630 2935 -610
rect 2900 -655 2905 -630
rect 2930 -655 2935 -630
rect 2900 -675 2935 -655
rect 2900 -700 2905 -675
rect 2930 -700 2935 -675
rect 2900 -725 2935 -700
rect 2900 -750 2905 -725
rect 2930 -750 2935 -725
rect 2900 -770 2935 -750
rect 2960 -585 2995 -575
rect 2960 -610 2965 -585
rect 2990 -610 2995 -585
rect 2960 -630 2995 -610
rect 2960 -655 2965 -630
rect 2990 -655 2995 -630
rect 2960 -675 2995 -655
rect 2960 -700 2965 -675
rect 2990 -700 2995 -675
rect 2960 -725 2995 -700
rect 2960 -750 2965 -725
rect 2990 -750 2995 -725
rect 2960 -770 2995 -750
rect 3020 -585 3055 -575
rect 3020 -610 3025 -585
rect 3050 -610 3055 -585
rect 3020 -630 3055 -610
rect 3020 -655 3025 -630
rect 3050 -655 3055 -630
rect 3020 -675 3055 -655
rect 3020 -700 3025 -675
rect 3050 -700 3055 -675
rect 3020 -725 3055 -700
rect 3020 -750 3025 -725
rect 3050 -750 3055 -725
rect 3020 -770 3055 -750
rect 3080 -585 3115 -575
rect 3080 -610 3085 -585
rect 3110 -610 3115 -585
rect 3080 -630 3115 -610
rect 3080 -655 3085 -630
rect 3110 -655 3115 -630
rect 3080 -675 3115 -655
rect 3080 -700 3085 -675
rect 3110 -700 3115 -675
rect 3080 -725 3115 -700
rect 3080 -750 3085 -725
rect 3110 -750 3115 -725
rect 3080 -770 3115 -750
rect 3140 -585 3175 -575
rect 3140 -610 3145 -585
rect 3170 -610 3175 -585
rect 3140 -630 3175 -610
rect 3140 -655 3145 -630
rect 3170 -655 3175 -630
rect 3140 -675 3175 -655
rect 3140 -700 3145 -675
rect 3170 -700 3175 -675
rect 3140 -725 3175 -700
rect 3140 -750 3145 -725
rect 3170 -750 3175 -725
rect 3140 -770 3175 -750
rect 3200 -585 3235 -575
rect 3200 -610 3205 -585
rect 3230 -610 3235 -585
rect 3200 -630 3235 -610
rect 3200 -655 3205 -630
rect 3230 -655 3235 -630
rect 3200 -675 3235 -655
rect 3200 -700 3205 -675
rect 3230 -700 3235 -675
rect 3200 -725 3235 -700
rect 3200 -750 3205 -725
rect 3230 -750 3235 -725
rect 3200 -770 3235 -750
rect 3260 -585 3295 -575
rect 3260 -610 3265 -585
rect 3290 -610 3295 -585
rect 3260 -630 3295 -610
rect 3260 -655 3265 -630
rect 3290 -655 3295 -630
rect 3260 -675 3295 -655
rect 3260 -700 3265 -675
rect 3290 -700 3295 -675
rect 3260 -725 3295 -700
rect 3260 -750 3265 -725
rect 3290 -750 3295 -725
rect 3260 -770 3295 -750
rect 3320 -585 3355 -575
rect 3320 -610 3325 -585
rect 3350 -610 3355 -585
rect 3320 -630 3355 -610
rect 3320 -655 3325 -630
rect 3350 -655 3355 -630
rect 3320 -675 3355 -655
rect 3320 -700 3325 -675
rect 3350 -700 3355 -675
rect 3320 -725 3355 -700
rect 3320 -750 3325 -725
rect 3350 -750 3355 -725
rect 3320 -770 3355 -750
rect 3380 -585 3415 -575
rect 3380 -610 3385 -585
rect 3410 -610 3415 -585
rect 3380 -630 3415 -610
rect 3380 -655 3385 -630
rect 3410 -655 3415 -630
rect 3380 -675 3415 -655
rect 3380 -700 3385 -675
rect 3410 -700 3415 -675
rect 3380 -725 3415 -700
rect 3380 -750 3385 -725
rect 3410 -750 3415 -725
rect 3380 -770 3415 -750
rect 3440 -585 3475 -575
rect 3440 -610 3445 -585
rect 3470 -610 3475 -585
rect 3440 -630 3475 -610
rect 3440 -655 3445 -630
rect 3470 -655 3475 -630
rect 3440 -675 3475 -655
rect 3440 -700 3445 -675
rect 3470 -700 3475 -675
rect 3440 -725 3475 -700
rect 3440 -750 3445 -725
rect 3470 -750 3475 -725
rect 3440 -770 3475 -750
rect 3500 -585 3535 -575
rect 3500 -610 3505 -585
rect 3530 -610 3535 -585
rect 3500 -630 3535 -610
rect 3500 -655 3505 -630
rect 3530 -655 3535 -630
rect 3500 -675 3535 -655
rect 3500 -700 3505 -675
rect 3530 -700 3535 -675
rect 3500 -725 3535 -700
rect 3500 -750 3505 -725
rect 3530 -750 3535 -725
rect 3500 -770 3535 -750
rect 3560 -585 3595 -575
rect 3560 -610 3565 -585
rect 3590 -610 3595 -585
rect 3560 -630 3595 -610
rect 3560 -655 3565 -630
rect 3590 -655 3595 -630
rect 3560 -675 3595 -655
rect 3560 -700 3565 -675
rect 3590 -700 3595 -675
rect 3560 -725 3595 -700
rect 3560 -750 3565 -725
rect 3590 -750 3595 -725
rect 3560 -770 3595 -750
rect 3620 -585 3655 -575
rect 3620 -610 3625 -585
rect 3650 -610 3655 -585
rect 3620 -630 3655 -610
rect 3620 -655 3625 -630
rect 3650 -655 3655 -630
rect 3620 -675 3655 -655
rect 3620 -700 3625 -675
rect 3650 -700 3655 -675
rect 3620 -725 3655 -700
rect 3620 -750 3625 -725
rect 3650 -750 3655 -725
rect 3620 -770 3655 -750
rect 3680 -585 3715 -575
rect 3680 -610 3685 -585
rect 3710 -610 3715 -585
rect 3680 -630 3715 -610
rect 3680 -655 3685 -630
rect 3710 -655 3715 -630
rect 3680 -675 3715 -655
rect 3680 -700 3685 -675
rect 3710 -700 3715 -675
rect 3680 -725 3715 -700
rect 3680 -750 3685 -725
rect 3710 -750 3715 -725
rect 3680 -770 3715 -750
rect 3740 -585 3775 -575
rect 3740 -610 3745 -585
rect 3770 -610 3775 -585
rect 3740 -630 3775 -610
rect 3740 -655 3745 -630
rect 3770 -655 3775 -630
rect 3740 -675 3775 -655
rect 3740 -700 3745 -675
rect 3770 -700 3775 -675
rect 3740 -725 3775 -700
rect 3740 -750 3745 -725
rect 3770 -750 3775 -725
rect 3740 -770 3775 -750
rect 3800 -585 3835 -575
rect 3800 -610 3805 -585
rect 3830 -610 3835 -585
rect 3800 -630 3835 -610
rect 3800 -655 3805 -630
rect 3830 -655 3835 -630
rect 3800 -675 3835 -655
rect 3800 -700 3805 -675
rect 3830 -700 3835 -675
rect 3800 -725 3835 -700
rect 3800 -750 3805 -725
rect 3830 -750 3835 -725
rect 3800 -770 3835 -750
rect 3860 -585 3895 -575
rect 3860 -610 3865 -585
rect 3890 -610 3895 -585
rect 3860 -630 3895 -610
rect 3860 -655 3865 -630
rect 3890 -655 3895 -630
rect 3860 -675 3895 -655
rect 3860 -700 3865 -675
rect 3890 -700 3895 -675
rect 3860 -725 3895 -700
rect 3860 -750 3865 -725
rect 3890 -750 3895 -725
rect 3860 -770 3895 -750
rect 3920 -585 3955 -575
rect 3920 -610 3925 -585
rect 3950 -610 3955 -585
rect 3920 -630 3955 -610
rect 3920 -655 3925 -630
rect 3950 -655 3955 -630
rect 3920 -675 3955 -655
rect 3920 -700 3925 -675
rect 3950 -700 3955 -675
rect 3920 -725 3955 -700
rect 3920 -750 3925 -725
rect 3950 -750 3955 -725
rect 3920 -770 3955 -750
rect 3980 -585 4015 -575
rect 3980 -610 3985 -585
rect 4010 -610 4015 -585
rect 3980 -630 4015 -610
rect 3980 -655 3985 -630
rect 4010 -655 4015 -630
rect 3980 -675 4015 -655
rect 3980 -700 3985 -675
rect 4010 -700 4015 -675
rect 3980 -725 4015 -700
rect 3980 -750 3985 -725
rect 4010 -750 4015 -725
rect 3980 -770 4015 -750
rect 4040 -585 4075 -575
rect 4040 -610 4045 -585
rect 4070 -610 4075 -585
rect 4040 -630 4075 -610
rect 4040 -655 4045 -630
rect 4070 -655 4075 -630
rect 4040 -675 4075 -655
rect 4040 -700 4045 -675
rect 4070 -700 4075 -675
rect 4040 -725 4075 -700
rect 4040 -750 4045 -725
rect 4070 -750 4075 -725
rect 4040 -770 4075 -750
rect 4100 -585 4135 -575
rect 4100 -610 4105 -585
rect 4130 -610 4135 -585
rect 4100 -630 4135 -610
rect 4100 -655 4105 -630
rect 4130 -655 4135 -630
rect 4100 -675 4135 -655
rect 4100 -700 4105 -675
rect 4130 -700 4135 -675
rect 4100 -725 4135 -700
rect 4100 -750 4105 -725
rect 4130 -750 4135 -725
rect 4100 -770 4135 -750
rect 4160 -585 4195 -575
rect 4160 -610 4165 -585
rect 4190 -610 4195 -585
rect 4160 -630 4195 -610
rect 4160 -655 4165 -630
rect 4190 -655 4195 -630
rect 4160 -675 4195 -655
rect 4160 -700 4165 -675
rect 4190 -700 4195 -675
rect 4160 -725 4195 -700
rect 4160 -750 4165 -725
rect 4190 -750 4195 -725
rect 4160 -770 4195 -750
rect 4220 -585 4255 -575
rect 4220 -610 4225 -585
rect 4250 -610 4255 -585
rect 4220 -630 4255 -610
rect 4220 -655 4225 -630
rect 4250 -655 4255 -630
rect 4220 -675 4255 -655
rect 4220 -700 4225 -675
rect 4250 -700 4255 -675
rect 4220 -725 4255 -700
rect 4220 -750 4225 -725
rect 4250 -750 4255 -725
rect 4220 -770 4255 -750
rect 4280 -585 4315 -575
rect 4280 -610 4285 -585
rect 4310 -610 4315 -585
rect 4280 -630 4315 -610
rect 4280 -655 4285 -630
rect 4310 -655 4315 -630
rect 4280 -675 4315 -655
rect 4280 -700 4285 -675
rect 4310 -700 4315 -675
rect 4280 -725 4315 -700
rect 4280 -750 4285 -725
rect 4310 -750 4315 -725
rect 4280 -770 4315 -750
rect 4340 -585 4375 -575
rect 4340 -610 4345 -585
rect 4370 -610 4375 -585
rect 4340 -630 4375 -610
rect 4340 -655 4345 -630
rect 4370 -655 4375 -630
rect 4340 -675 4375 -655
rect 4340 -700 4345 -675
rect 4370 -700 4375 -675
rect 4340 -725 4375 -700
rect 4340 -750 4345 -725
rect 4370 -750 4375 -725
rect 4340 -770 4375 -750
rect 4400 -585 4435 -575
rect 4400 -610 4405 -585
rect 4430 -610 4435 -585
rect 4400 -630 4435 -610
rect 4400 -655 4405 -630
rect 4430 -655 4435 -630
rect 4400 -675 4435 -655
rect 4400 -700 4405 -675
rect 4430 -700 4435 -675
rect 4400 -725 4435 -700
rect 4400 -750 4405 -725
rect 4430 -750 4435 -725
rect 4400 -770 4435 -750
rect 4460 -585 4495 -575
rect 4460 -610 4465 -585
rect 4490 -610 4495 -585
rect 4460 -630 4495 -610
rect 4460 -655 4465 -630
rect 4490 -655 4495 -630
rect 4460 -675 4495 -655
rect 4460 -700 4465 -675
rect 4490 -700 4495 -675
rect 4460 -725 4495 -700
rect 4460 -750 4465 -725
rect 4490 -750 4495 -725
rect 4460 -770 4495 -750
rect 4520 -585 4555 -575
rect 4520 -610 4525 -585
rect 4550 -610 4555 -585
rect 4520 -630 4555 -610
rect 4520 -655 4525 -630
rect 4550 -655 4555 -630
rect 4520 -675 4555 -655
rect 4520 -700 4525 -675
rect 4550 -700 4555 -675
rect 4520 -725 4555 -700
rect 4520 -750 4525 -725
rect 4550 -750 4555 -725
rect 4520 -770 4555 -750
rect 4580 -585 4615 -575
rect 4580 -610 4585 -585
rect 4610 -610 4615 -585
rect 4580 -630 4615 -610
rect 4580 -655 4585 -630
rect 4610 -655 4615 -630
rect 4580 -675 4615 -655
rect 4580 -700 4585 -675
rect 4610 -700 4615 -675
rect 4580 -725 4615 -700
rect 4580 -750 4585 -725
rect 4610 -750 4615 -725
rect 4580 -770 4615 -750
rect 4640 -585 4675 -575
rect 4640 -610 4645 -585
rect 4670 -610 4675 -585
rect 4640 -630 4675 -610
rect 4640 -655 4645 -630
rect 4670 -655 4675 -630
rect 4640 -675 4675 -655
rect 4640 -700 4645 -675
rect 4670 -700 4675 -675
rect 4640 -725 4675 -700
rect 4640 -750 4645 -725
rect 4670 -750 4675 -725
rect 4640 -770 4675 -750
rect 4700 -585 4735 -575
rect 4700 -610 4705 -585
rect 4730 -610 4735 -585
rect 4700 -630 4735 -610
rect 4700 -655 4705 -630
rect 4730 -655 4735 -630
rect 4700 -675 4735 -655
rect 4700 -700 4705 -675
rect 4730 -700 4735 -675
rect 4700 -725 4735 -700
rect 4700 -750 4705 -725
rect 4730 -750 4735 -725
rect 4700 -770 4735 -750
rect 4760 -585 4795 -575
rect 4760 -610 4765 -585
rect 4790 -610 4795 -585
rect 4760 -630 4795 -610
rect 4760 -655 4765 -630
rect 4790 -655 4795 -630
rect 4760 -675 4795 -655
rect 4760 -700 4765 -675
rect 4790 -700 4795 -675
rect 4760 -725 4795 -700
rect 4760 -750 4765 -725
rect 4790 -750 4795 -725
rect 4760 -770 4795 -750
rect 4820 -585 4855 -575
rect 4820 -610 4825 -585
rect 4850 -610 4855 -585
rect 4820 -630 4855 -610
rect 4820 -655 4825 -630
rect 4850 -655 4855 -630
rect 4820 -675 4855 -655
rect 4820 -700 4825 -675
rect 4850 -700 4855 -675
rect 4820 -725 4855 -700
rect 4820 -750 4825 -725
rect 4850 -750 4855 -725
rect 4820 -770 4855 -750
rect 4880 -585 4915 -575
rect 4880 -610 4885 -585
rect 4910 -610 4915 -585
rect 4880 -630 4915 -610
rect 4880 -655 4885 -630
rect 4910 -655 4915 -630
rect 4880 -675 4915 -655
rect 4880 -700 4885 -675
rect 4910 -700 4915 -675
rect 4880 -725 4915 -700
rect 4880 -750 4885 -725
rect 4910 -750 4915 -725
rect 4880 -770 4915 -750
rect 4940 -585 4975 -575
rect 4940 -610 4945 -585
rect 4970 -610 4975 -585
rect 4940 -630 4975 -610
rect 4940 -655 4945 -630
rect 4970 -655 4975 -630
rect 4940 -675 4975 -655
rect 4940 -700 4945 -675
rect 4970 -700 4975 -675
rect 4940 -725 4975 -700
rect 4940 -750 4945 -725
rect 4970 -750 4975 -725
rect 4940 -770 4975 -750
rect 5000 -585 5035 -575
rect 5000 -610 5005 -585
rect 5030 -610 5035 -585
rect 5000 -630 5035 -610
rect 5000 -655 5005 -630
rect 5030 -655 5035 -630
rect 5000 -675 5035 -655
rect 5000 -700 5005 -675
rect 5030 -700 5035 -675
rect 5000 -725 5035 -700
rect 5000 -750 5005 -725
rect 5030 -750 5035 -725
rect 5000 -770 5035 -750
rect 5060 -585 5095 -575
rect 5060 -610 5065 -585
rect 5090 -610 5095 -585
rect 5060 -630 5095 -610
rect 5060 -655 5065 -630
rect 5090 -655 5095 -630
rect 5060 -675 5095 -655
rect 5060 -700 5065 -675
rect 5090 -700 5095 -675
rect 5060 -725 5095 -700
rect 5060 -750 5065 -725
rect 5090 -750 5095 -725
rect 5060 -770 5095 -750
rect 5120 -585 5155 -575
rect 5120 -610 5125 -585
rect 5150 -610 5155 -585
rect 5120 -630 5155 -610
rect 5120 -655 5125 -630
rect 5150 -655 5155 -630
rect 5120 -675 5155 -655
rect 5120 -700 5125 -675
rect 5150 -700 5155 -675
rect 5120 -725 5155 -700
rect 5120 -750 5125 -725
rect 5150 -750 5155 -725
rect 5120 -770 5155 -750
rect 5180 -585 5215 -575
rect 5180 -610 5185 -585
rect 5210 -610 5215 -585
rect 5180 -630 5215 -610
rect 5180 -655 5185 -630
rect 5210 -655 5215 -630
rect 5180 -675 5215 -655
rect 5180 -700 5185 -675
rect 5210 -700 5215 -675
rect 5180 -725 5215 -700
rect 5180 -750 5185 -725
rect 5210 -750 5215 -725
rect 5180 -770 5215 -750
rect 5240 -585 5275 -575
rect 5240 -610 5245 -585
rect 5270 -610 5275 -585
rect 5240 -630 5275 -610
rect 5240 -655 5245 -630
rect 5270 -655 5275 -630
rect 5240 -675 5275 -655
rect 5240 -700 5245 -675
rect 5270 -700 5275 -675
rect 5240 -725 5275 -700
rect 5240 -750 5245 -725
rect 5270 -750 5275 -725
rect 5240 -770 5275 -750
rect 5300 -585 5335 -575
rect 5300 -610 5305 -585
rect 5330 -610 5335 -585
rect 5300 -630 5335 -610
rect 5300 -655 5305 -630
rect 5330 -655 5335 -630
rect 5300 -675 5335 -655
rect 5300 -700 5305 -675
rect 5330 -700 5335 -675
rect 5300 -725 5335 -700
rect 5300 -750 5305 -725
rect 5330 -750 5335 -725
rect 5300 -770 5335 -750
rect 5360 -585 5395 -575
rect 5360 -610 5365 -585
rect 5390 -610 5395 -585
rect 5360 -630 5395 -610
rect 5360 -655 5365 -630
rect 5390 -655 5395 -630
rect 5360 -675 5395 -655
rect 5360 -700 5365 -675
rect 5390 -700 5395 -675
rect 5360 -725 5395 -700
rect 5360 -750 5365 -725
rect 5390 -750 5395 -725
rect 5360 -770 5395 -750
rect 5420 -585 5455 -575
rect 5420 -610 5425 -585
rect 5450 -610 5455 -585
rect 5420 -630 5455 -610
rect 5420 -655 5425 -630
rect 5450 -655 5455 -630
rect 5420 -675 5455 -655
rect 5420 -700 5425 -675
rect 5450 -700 5455 -675
rect 5420 -725 5455 -700
rect 5420 -750 5425 -725
rect 5450 -750 5455 -725
rect 5420 -770 5455 -750
rect 5480 -585 5515 -575
rect 5480 -610 5485 -585
rect 5510 -610 5515 -585
rect 5480 -630 5515 -610
rect 5480 -655 5485 -630
rect 5510 -655 5515 -630
rect 5480 -675 5515 -655
rect 5480 -700 5485 -675
rect 5510 -700 5515 -675
rect 5480 -725 5515 -700
rect 5480 -750 5485 -725
rect 5510 -750 5515 -725
rect 5480 -770 5515 -750
rect 5540 -585 5575 -575
rect 5540 -610 5545 -585
rect 5570 -610 5575 -585
rect 5540 -630 5575 -610
rect 5540 -655 5545 -630
rect 5570 -655 5575 -630
rect 5540 -675 5575 -655
rect 5540 -700 5545 -675
rect 5570 -700 5575 -675
rect 5540 -725 5575 -700
rect 5540 -750 5545 -725
rect 5570 -750 5575 -725
rect 5540 -770 5575 -750
rect 5600 -585 5635 -575
rect 5600 -610 5605 -585
rect 5630 -610 5635 -585
rect 5600 -630 5635 -610
rect 5600 -655 5605 -630
rect 5630 -655 5635 -630
rect 5600 -675 5635 -655
rect 5600 -700 5605 -675
rect 5630 -700 5635 -675
rect 5600 -725 5635 -700
rect 5600 -750 5605 -725
rect 5630 -750 5635 -725
rect 5600 -770 5635 -750
rect 5660 -585 5695 -575
rect 5660 -610 5665 -585
rect 5690 -610 5695 -585
rect 5660 -630 5695 -610
rect 5660 -655 5665 -630
rect 5690 -655 5695 -630
rect 5660 -675 5695 -655
rect 5660 -700 5665 -675
rect 5690 -700 5695 -675
rect 5660 -725 5695 -700
rect 5660 -750 5665 -725
rect 5690 -750 5695 -725
rect 5660 -770 5695 -750
rect 5720 -585 5755 -575
rect 5720 -610 5725 -585
rect 5750 -610 5755 -585
rect 5720 -630 5755 -610
rect 5720 -655 5725 -630
rect 5750 -655 5755 -630
rect 5720 -675 5755 -655
rect 5720 -700 5725 -675
rect 5750 -700 5755 -675
rect 5720 -725 5755 -700
rect 5720 -750 5725 -725
rect 5750 -750 5755 -725
rect 5720 -770 5755 -750
rect 5780 -585 5815 -575
rect 5780 -610 5785 -585
rect 5810 -610 5815 -585
rect 5780 -630 5815 -610
rect 5780 -655 5785 -630
rect 5810 -655 5815 -630
rect 5780 -675 5815 -655
rect 5780 -700 5785 -675
rect 5810 -700 5815 -675
rect 5780 -725 5815 -700
rect 5780 -750 5785 -725
rect 5810 -750 5815 -725
rect 5780 -770 5815 -750
rect 5840 -585 5875 -575
rect 5840 -610 5845 -585
rect 5870 -610 5875 -585
rect 5840 -630 5875 -610
rect 5840 -655 5845 -630
rect 5870 -655 5875 -630
rect 5840 -675 5875 -655
rect 5840 -700 5845 -675
rect 5870 -700 5875 -675
rect 5840 -725 5875 -700
rect 5840 -750 5845 -725
rect 5870 -750 5875 -725
rect 5840 -770 5875 -750
rect 5900 -585 5935 -575
rect 5900 -610 5905 -585
rect 5930 -610 5935 -585
rect 5900 -630 5935 -610
rect 5900 -655 5905 -630
rect 5930 -655 5935 -630
rect 5900 -675 5935 -655
rect 5900 -700 5905 -675
rect 5930 -700 5935 -675
rect 5900 -725 5935 -700
rect 5900 -750 5905 -725
rect 5930 -750 5935 -725
rect 5900 -770 5935 -750
rect 5960 -585 5995 -575
rect 5960 -610 5965 -585
rect 5990 -610 5995 -585
rect 5960 -630 5995 -610
rect 5960 -655 5965 -630
rect 5990 -655 5995 -630
rect 5960 -675 5995 -655
rect 5960 -700 5965 -675
rect 5990 -700 5995 -675
rect 5960 -725 5995 -700
rect 5960 -750 5965 -725
rect 5990 -750 5995 -725
rect 5960 -770 5995 -750
rect 6020 -585 6055 -575
rect 6020 -610 6025 -585
rect 6050 -610 6055 -585
rect 6020 -630 6055 -610
rect 6020 -655 6025 -630
rect 6050 -655 6055 -630
rect 6020 -675 6055 -655
rect 6020 -700 6025 -675
rect 6050 -700 6055 -675
rect 6020 -725 6055 -700
rect 6020 -750 6025 -725
rect 6050 -750 6055 -725
rect 6020 -770 6055 -750
rect 6080 -585 6115 -575
rect 6080 -610 6085 -585
rect 6110 -610 6115 -585
rect 6080 -630 6115 -610
rect 6080 -655 6085 -630
rect 6110 -655 6115 -630
rect 6080 -675 6115 -655
rect 6080 -700 6085 -675
rect 6110 -700 6115 -675
rect 6080 -725 6115 -700
rect 6080 -750 6085 -725
rect 6110 -750 6115 -725
rect 6080 -770 6115 -750
rect 6140 -585 6175 -575
rect 6140 -610 6145 -585
rect 6170 -610 6175 -585
rect 6140 -630 6175 -610
rect 6140 -655 6145 -630
rect 6170 -655 6175 -630
rect 6140 -675 6175 -655
rect 6140 -700 6145 -675
rect 6170 -700 6175 -675
rect 6140 -725 6175 -700
rect 6140 -750 6145 -725
rect 6170 -750 6175 -725
rect 6140 -770 6175 -750
rect 6200 -585 6235 -575
rect 6200 -610 6205 -585
rect 6230 -610 6235 -585
rect 6200 -630 6235 -610
rect 6200 -655 6205 -630
rect 6230 -655 6235 -630
rect 6200 -675 6235 -655
rect 6200 -700 6205 -675
rect 6230 -700 6235 -675
rect 6200 -725 6235 -700
rect 6200 -750 6205 -725
rect 6230 -750 6235 -725
rect 6200 -770 6235 -750
rect 6260 -585 6295 -575
rect 6260 -610 6265 -585
rect 6290 -610 6295 -585
rect 6260 -630 6295 -610
rect 6260 -655 6265 -630
rect 6290 -655 6295 -630
rect 6260 -675 6295 -655
rect 6260 -700 6265 -675
rect 6290 -700 6295 -675
rect 6260 -725 6295 -700
rect 6260 -750 6265 -725
rect 6290 -750 6295 -725
rect 6260 -770 6295 -750
rect 6320 -585 6355 -575
rect 6320 -610 6325 -585
rect 6350 -610 6355 -585
rect 6320 -630 6355 -610
rect 6320 -655 6325 -630
rect 6350 -655 6355 -630
rect 6320 -675 6355 -655
rect 6320 -700 6325 -675
rect 6350 -700 6355 -675
rect 6320 -725 6355 -700
rect 6320 -750 6325 -725
rect 6350 -750 6355 -725
rect 6320 -770 6355 -750
rect 6380 -585 6415 -575
rect 6380 -610 6385 -585
rect 6410 -610 6415 -585
rect 6380 -630 6415 -610
rect 6380 -655 6385 -630
rect 6410 -655 6415 -630
rect 6380 -675 6415 -655
rect 6380 -700 6385 -675
rect 6410 -700 6415 -675
rect 6380 -725 6415 -700
rect 6380 -750 6385 -725
rect 6410 -750 6415 -725
rect 6380 -770 6415 -750
rect 6440 -585 6475 -575
rect 6440 -610 6445 -585
rect 6470 -610 6475 -585
rect 6440 -630 6475 -610
rect 6440 -655 6445 -630
rect 6470 -655 6475 -630
rect 6440 -675 6475 -655
rect 6440 -700 6445 -675
rect 6470 -700 6475 -675
rect 6440 -725 6475 -700
rect 6440 -750 6445 -725
rect 6470 -750 6475 -725
rect 6440 -770 6475 -750
rect 6500 -585 6535 -575
rect 6500 -610 6505 -585
rect 6530 -610 6535 -585
rect 6500 -630 6535 -610
rect 6500 -655 6505 -630
rect 6530 -655 6535 -630
rect 6500 -675 6535 -655
rect 6500 -700 6505 -675
rect 6530 -700 6535 -675
rect 6500 -725 6535 -700
rect 6500 -750 6505 -725
rect 6530 -750 6535 -725
rect 6500 -770 6535 -750
rect 6560 -585 6595 -575
rect 6560 -610 6565 -585
rect 6590 -610 6595 -585
rect 6560 -630 6595 -610
rect 6560 -655 6565 -630
rect 6590 -655 6595 -630
rect 6560 -675 6595 -655
rect 6560 -700 6565 -675
rect 6590 -700 6595 -675
rect 6560 -725 6595 -700
rect 6560 -750 6565 -725
rect 6590 -750 6595 -725
rect 6560 -770 6595 -750
rect 6620 -585 6655 -575
rect 6620 -610 6625 -585
rect 6650 -610 6655 -585
rect 6620 -630 6655 -610
rect 6620 -655 6625 -630
rect 6650 -655 6655 -630
rect 6620 -675 6655 -655
rect 6620 -700 6625 -675
rect 6650 -700 6655 -675
rect 6620 -725 6655 -700
rect 6620 -750 6625 -725
rect 6650 -750 6655 -725
rect 6620 -770 6655 -750
rect 6680 -585 6715 -575
rect 6680 -610 6685 -585
rect 6710 -610 6715 -585
rect 6680 -630 6715 -610
rect 6680 -655 6685 -630
rect 6710 -655 6715 -630
rect 6680 -675 6715 -655
rect 6680 -700 6685 -675
rect 6710 -700 6715 -675
rect 6680 -725 6715 -700
rect 6680 -750 6685 -725
rect 6710 -750 6715 -725
rect 6680 -770 6715 -750
rect 6740 -585 6775 -575
rect 6740 -610 6745 -585
rect 6770 -610 6775 -585
rect 6740 -630 6775 -610
rect 6740 -655 6745 -630
rect 6770 -655 6775 -630
rect 6740 -675 6775 -655
rect 6740 -700 6745 -675
rect 6770 -700 6775 -675
rect 6740 -725 6775 -700
rect 6740 -750 6745 -725
rect 6770 -750 6775 -725
rect 6740 -770 6775 -750
rect 6800 -585 6835 -575
rect 6800 -610 6805 -585
rect 6830 -610 6835 -585
rect 6800 -630 6835 -610
rect 6800 -655 6805 -630
rect 6830 -655 6835 -630
rect 6800 -675 6835 -655
rect 6800 -700 6805 -675
rect 6830 -700 6835 -675
rect 6800 -725 6835 -700
rect 6800 -750 6805 -725
rect 6830 -750 6835 -725
rect 6800 -770 6835 -750
rect 6860 -585 6895 -575
rect 6860 -610 6865 -585
rect 6890 -610 6895 -585
rect 6860 -630 6895 -610
rect 6860 -655 6865 -630
rect 6890 -655 6895 -630
rect 6860 -675 6895 -655
rect 6860 -700 6865 -675
rect 6890 -700 6895 -675
rect 6860 -725 6895 -700
rect 6860 -750 6865 -725
rect 6890 -750 6895 -725
rect 6860 -770 6895 -750
rect 6920 -585 6955 -575
rect 6920 -610 6925 -585
rect 6950 -610 6955 -585
rect 6920 -630 6955 -610
rect 6920 -655 6925 -630
rect 6950 -655 6955 -630
rect 6920 -675 6955 -655
rect 6920 -700 6925 -675
rect 6950 -700 6955 -675
rect 6920 -725 6955 -700
rect 6920 -750 6925 -725
rect 6950 -750 6955 -725
rect 6920 -770 6955 -750
rect 6980 -585 7015 -575
rect 6980 -610 6985 -585
rect 7010 -610 7015 -585
rect 6980 -630 7015 -610
rect 6980 -655 6985 -630
rect 7010 -655 7015 -630
rect 6980 -675 7015 -655
rect 6980 -700 6985 -675
rect 7010 -700 7015 -675
rect 6980 -725 7015 -700
rect 6980 -750 6985 -725
rect 7010 -750 7015 -725
rect 6980 -770 7015 -750
rect 7040 -585 7075 -575
rect 7040 -610 7045 -585
rect 7070 -610 7075 -585
rect 7040 -630 7075 -610
rect 7040 -655 7045 -630
rect 7070 -655 7075 -630
rect 7040 -675 7075 -655
rect 7040 -700 7045 -675
rect 7070 -700 7075 -675
rect 7040 -725 7075 -700
rect 7040 -750 7045 -725
rect 7070 -750 7075 -725
rect 7040 -770 7075 -750
rect 7100 -585 7135 -575
rect 7100 -610 7105 -585
rect 7130 -610 7135 -585
rect 7100 -630 7135 -610
rect 7100 -655 7105 -630
rect 7130 -655 7135 -630
rect 7100 -675 7135 -655
rect 7100 -700 7105 -675
rect 7130 -700 7135 -675
rect 7100 -725 7135 -700
rect 7100 -750 7105 -725
rect 7130 -750 7135 -725
rect 7100 -770 7135 -750
rect 7160 -585 7195 -575
rect 7160 -610 7165 -585
rect 7190 -610 7195 -585
rect 7160 -630 7195 -610
rect 7160 -655 7165 -630
rect 7190 -655 7195 -630
rect 7160 -675 7195 -655
rect 7160 -700 7165 -675
rect 7190 -700 7195 -675
rect 7160 -725 7195 -700
rect 7160 -750 7165 -725
rect 7190 -750 7195 -725
rect 7160 -770 7195 -750
rect 7220 -585 7255 -575
rect 7220 -610 7225 -585
rect 7250 -610 7255 -585
rect 7220 -630 7255 -610
rect 7220 -655 7225 -630
rect 7250 -655 7255 -630
rect 7220 -675 7255 -655
rect 7220 -700 7225 -675
rect 7250 -700 7255 -675
rect 7220 -725 7255 -700
rect 7220 -750 7225 -725
rect 7250 -750 7255 -725
rect 7220 -770 7255 -750
rect 7280 -585 7315 -575
rect 7280 -610 7285 -585
rect 7310 -610 7315 -585
rect 7280 -630 7315 -610
rect 7280 -655 7285 -630
rect 7310 -655 7315 -630
rect 7280 -675 7315 -655
rect 7280 -700 7285 -675
rect 7310 -700 7315 -675
rect 7280 -725 7315 -700
rect 7280 -750 7285 -725
rect 7310 -750 7315 -725
rect 7280 -770 7315 -750
rect 7340 -585 7375 -575
rect 7340 -610 7345 -585
rect 7370 -610 7375 -585
rect 7340 -630 7375 -610
rect 7340 -655 7345 -630
rect 7370 -655 7375 -630
rect 7340 -675 7375 -655
rect 7340 -700 7345 -675
rect 7370 -700 7375 -675
rect 7340 -725 7375 -700
rect 7340 -750 7345 -725
rect 7370 -750 7375 -725
rect 7340 -770 7375 -750
rect 7400 -585 7435 -575
rect 7400 -610 7405 -585
rect 7430 -610 7435 -585
rect 7400 -630 7435 -610
rect 7400 -655 7405 -630
rect 7430 -655 7435 -630
rect 7400 -675 7435 -655
rect 7400 -700 7405 -675
rect 7430 -700 7435 -675
rect 7400 -725 7435 -700
rect 7400 -750 7405 -725
rect 7430 -750 7435 -725
rect 7400 -770 7435 -750
rect 7460 -585 7495 -575
rect 7460 -610 7465 -585
rect 7490 -610 7495 -585
rect 7460 -630 7495 -610
rect 7460 -655 7465 -630
rect 7490 -655 7495 -630
rect 7460 -675 7495 -655
rect 7460 -700 7465 -675
rect 7490 -700 7495 -675
rect 7460 -725 7495 -700
rect 7460 -750 7465 -725
rect 7490 -750 7495 -725
rect 7460 -770 7495 -750
rect 7520 -585 7555 -575
rect 7520 -610 7525 -585
rect 7550 -610 7555 -585
rect 7520 -630 7555 -610
rect 7520 -655 7525 -630
rect 7550 -655 7555 -630
rect 7520 -675 7555 -655
rect 7520 -700 7525 -675
rect 7550 -700 7555 -675
rect 7520 -725 7555 -700
rect 7520 -750 7525 -725
rect 7550 -750 7555 -725
rect 7520 -770 7555 -750
rect 7580 -585 7615 -575
rect 7580 -610 7585 -585
rect 7610 -610 7615 -585
rect 7580 -630 7615 -610
rect 7580 -655 7585 -630
rect 7610 -655 7615 -630
rect 7580 -675 7615 -655
rect 7580 -700 7585 -675
rect 7610 -700 7615 -675
rect 7580 -725 7615 -700
rect 7580 -750 7585 -725
rect 7610 -750 7615 -725
rect 7580 -770 7615 -750
rect 7640 -585 7675 -575
rect 7640 -610 7645 -585
rect 7670 -610 7675 -585
rect 7640 -630 7675 -610
rect 7640 -655 7645 -630
rect 7670 -655 7675 -630
rect 7640 -675 7675 -655
rect 7640 -700 7645 -675
rect 7670 -700 7675 -675
rect 7640 -725 7675 -700
rect 7640 -750 7645 -725
rect 7670 -750 7675 -725
rect 7640 -770 7675 -750
rect 7700 -585 7735 -575
rect 7700 -610 7705 -585
rect 7730 -610 7735 -585
rect 7700 -630 7735 -610
rect 7700 -655 7705 -630
rect 7730 -655 7735 -630
rect 7700 -675 7735 -655
rect 7700 -700 7705 -675
rect 7730 -700 7735 -675
rect 7700 -725 7735 -700
rect 7700 -750 7705 -725
rect 7730 -750 7735 -725
rect 7700 -770 7735 -750
rect 7760 -585 7795 -575
rect 7760 -610 7765 -585
rect 7790 -610 7795 -585
rect 7760 -630 7795 -610
rect 7760 -655 7765 -630
rect 7790 -655 7795 -630
rect 7760 -675 7795 -655
rect 7760 -700 7765 -675
rect 7790 -700 7795 -675
rect 7760 -725 7795 -700
rect 7760 -750 7765 -725
rect 7790 -750 7795 -725
rect 7760 -770 7795 -750
rect 7820 -585 7855 -575
rect 7820 -610 7825 -585
rect 7850 -610 7855 -585
rect 7820 -630 7855 -610
rect 7820 -655 7825 -630
rect 7850 -655 7855 -630
rect 7820 -675 7855 -655
rect 7820 -700 7825 -675
rect 7850 -700 7855 -675
rect 7820 -725 7855 -700
rect 7820 -750 7825 -725
rect 7850 -750 7855 -725
rect 7820 -770 7855 -750
rect 7880 -585 7915 -575
rect 7880 -610 7885 -585
rect 7910 -610 7915 -585
rect 7880 -630 7915 -610
rect 7880 -655 7885 -630
rect 7910 -655 7915 -630
rect 7880 -675 7915 -655
rect 7880 -700 7885 -675
rect 7910 -700 7915 -675
rect 7880 -725 7915 -700
rect 7880 -750 7885 -725
rect 7910 -750 7915 -725
rect 7880 -770 7915 -750
rect 7940 -585 7975 -575
rect 7940 -610 7945 -585
rect 7970 -610 7975 -585
rect 7940 -630 7975 -610
rect 7940 -655 7945 -630
rect 7970 -655 7975 -630
rect 7940 -675 7975 -655
rect 7940 -700 7945 -675
rect 7970 -700 7975 -675
rect 7940 -725 7975 -700
rect 7940 -750 7945 -725
rect 7970 -750 7975 -725
rect 7940 -770 7975 -750
rect 8000 -585 8035 -575
rect 8000 -610 8005 -585
rect 8030 -610 8035 -585
rect 8000 -630 8035 -610
rect 8000 -655 8005 -630
rect 8030 -655 8035 -630
rect 8000 -675 8035 -655
rect 8000 -700 8005 -675
rect 8030 -700 8035 -675
rect 8000 -725 8035 -700
rect 8000 -750 8005 -725
rect 8030 -750 8035 -725
rect 8000 -770 8035 -750
rect 8060 -585 8095 -575
rect 8060 -610 8065 -585
rect 8090 -610 8095 -585
rect 8060 -630 8095 -610
rect 8060 -655 8065 -630
rect 8090 -655 8095 -630
rect 8060 -675 8095 -655
rect 8060 -700 8065 -675
rect 8090 -700 8095 -675
rect 8060 -725 8095 -700
rect 8060 -750 8065 -725
rect 8090 -750 8095 -725
rect 8060 -770 8095 -750
rect 8120 -585 8155 -575
rect 8120 -610 8125 -585
rect 8150 -610 8155 -585
rect 8120 -630 8155 -610
rect 8120 -655 8125 -630
rect 8150 -655 8155 -630
rect 8120 -675 8155 -655
rect 8120 -700 8125 -675
rect 8150 -700 8155 -675
rect 8120 -725 8155 -700
rect 8120 -750 8125 -725
rect 8150 -750 8155 -725
rect 8120 -770 8155 -750
rect 8180 -585 8215 -575
rect 8180 -610 8185 -585
rect 8210 -610 8215 -585
rect 8180 -630 8215 -610
rect 8180 -655 8185 -630
rect 8210 -655 8215 -630
rect 8180 -675 8215 -655
rect 8180 -700 8185 -675
rect 8210 -700 8215 -675
rect 8180 -725 8215 -700
rect 8180 -750 8185 -725
rect 8210 -750 8215 -725
rect 8180 -770 8215 -750
rect 8240 -585 8275 -575
rect 8240 -610 8245 -585
rect 8270 -610 8275 -585
rect 8240 -630 8275 -610
rect 8240 -655 8245 -630
rect 8270 -655 8275 -630
rect 8240 -675 8275 -655
rect 8240 -700 8245 -675
rect 8270 -700 8275 -675
rect 8240 -725 8275 -700
rect 8240 -750 8245 -725
rect 8270 -750 8275 -725
rect 8240 -770 8275 -750
rect 8300 -585 8335 -575
rect 8300 -610 8305 -585
rect 8330 -610 8335 -585
rect 8300 -630 8335 -610
rect 8300 -655 8305 -630
rect 8330 -655 8335 -630
rect 8300 -675 8335 -655
rect 8300 -700 8305 -675
rect 8330 -700 8335 -675
rect 8300 -725 8335 -700
rect 8300 -750 8305 -725
rect 8330 -750 8335 -725
rect 8300 -770 8335 -750
rect 8360 -585 8395 -575
rect 8360 -610 8365 -585
rect 8390 -610 8395 -585
rect 8360 -630 8395 -610
rect 8360 -655 8365 -630
rect 8390 -655 8395 -630
rect 8360 -675 8395 -655
rect 8360 -700 8365 -675
rect 8390 -700 8395 -675
rect 8360 -725 8395 -700
rect 8360 -750 8365 -725
rect 8390 -750 8395 -725
rect 8360 -770 8395 -750
rect 8420 -585 8455 -575
rect 8420 -610 8425 -585
rect 8450 -610 8455 -585
rect 8420 -630 8455 -610
rect 8420 -655 8425 -630
rect 8450 -655 8455 -630
rect 8420 -675 8455 -655
rect 8420 -700 8425 -675
rect 8450 -700 8455 -675
rect 8420 -725 8455 -700
rect 8420 -750 8425 -725
rect 8450 -750 8455 -725
rect 8420 -770 8455 -750
rect 8480 -585 8515 -575
rect 8480 -610 8485 -585
rect 8510 -610 8515 -585
rect 8480 -630 8515 -610
rect 8480 -655 8485 -630
rect 8510 -655 8515 -630
rect 8480 -675 8515 -655
rect 8480 -700 8485 -675
rect 8510 -700 8515 -675
rect 8480 -725 8515 -700
rect 8480 -750 8485 -725
rect 8510 -750 8515 -725
rect 8480 -770 8515 -750
rect 8540 -585 8575 -575
rect 8540 -610 8545 -585
rect 8570 -610 8575 -585
rect 8540 -630 8575 -610
rect 8540 -655 8545 -630
rect 8570 -655 8575 -630
rect 8540 -675 8575 -655
rect 8540 -700 8545 -675
rect 8570 -700 8575 -675
rect 8540 -725 8575 -700
rect 8540 -750 8545 -725
rect 8570 -750 8575 -725
rect 8540 -770 8575 -750
rect 8600 -585 8635 -575
rect 8600 -610 8605 -585
rect 8630 -610 8635 -585
rect 8600 -630 8635 -610
rect 8600 -655 8605 -630
rect 8630 -655 8635 -630
rect 8600 -675 8635 -655
rect 8600 -700 8605 -675
rect 8630 -700 8635 -675
rect 8600 -725 8635 -700
rect 8600 -750 8605 -725
rect 8630 -750 8635 -725
rect 8600 -770 8635 -750
rect 8660 -585 8695 -575
rect 8660 -610 8665 -585
rect 8690 -610 8695 -585
rect 8660 -630 8695 -610
rect 8660 -655 8665 -630
rect 8690 -655 8695 -630
rect 8660 -675 8695 -655
rect 8660 -700 8665 -675
rect 8690 -700 8695 -675
rect 8660 -725 8695 -700
rect 8660 -750 8665 -725
rect 8690 -750 8695 -725
rect 8660 -770 8695 -750
rect 8720 -585 8755 -575
rect 8720 -610 8725 -585
rect 8750 -610 8755 -585
rect 8720 -630 8755 -610
rect 8720 -655 8725 -630
rect 8750 -655 8755 -630
rect 8720 -675 8755 -655
rect 8720 -700 8725 -675
rect 8750 -700 8755 -675
rect 8720 -725 8755 -700
rect 8720 -750 8725 -725
rect 8750 -750 8755 -725
rect 8720 -770 8755 -750
rect 8780 -585 8815 -575
rect 8780 -610 8785 -585
rect 8810 -610 8815 -585
rect 8780 -630 8815 -610
rect 8780 -655 8785 -630
rect 8810 -655 8815 -630
rect 8780 -675 8815 -655
rect 8780 -700 8785 -675
rect 8810 -700 8815 -675
rect 8780 -725 8815 -700
rect 8780 -750 8785 -725
rect 8810 -750 8815 -725
rect 8780 -770 8815 -750
rect 8840 -585 8875 -575
rect 8840 -610 8845 -585
rect 8870 -610 8875 -585
rect 8840 -630 8875 -610
rect 8840 -655 8845 -630
rect 8870 -655 8875 -630
rect 8840 -675 8875 -655
rect 8840 -700 8845 -675
rect 8870 -700 8875 -675
rect 8840 -725 8875 -700
rect 8840 -750 8845 -725
rect 8870 -750 8875 -725
rect 8840 -770 8875 -750
rect 8900 -585 8935 -575
rect 8900 -610 8905 -585
rect 8930 -610 8935 -585
rect 8900 -630 8935 -610
rect 8900 -655 8905 -630
rect 8930 -655 8935 -630
rect 8900 -675 8935 -655
rect 8900 -700 8905 -675
rect 8930 -700 8935 -675
rect 8900 -725 8935 -700
rect 8900 -750 8905 -725
rect 8930 -750 8935 -725
rect 8900 -770 8935 -750
rect 8960 -585 8995 -575
rect 8960 -610 8965 -585
rect 8990 -610 8995 -585
rect 8960 -630 8995 -610
rect 8960 -655 8965 -630
rect 8990 -655 8995 -630
rect 8960 -675 8995 -655
rect 8960 -700 8965 -675
rect 8990 -700 8995 -675
rect 8960 -725 8995 -700
rect 8960 -750 8965 -725
rect 8990 -750 8995 -725
rect 8960 -770 8995 -750
rect 9020 -585 9055 -575
rect 9020 -610 9025 -585
rect 9050 -610 9055 -585
rect 9020 -630 9055 -610
rect 9020 -655 9025 -630
rect 9050 -655 9055 -630
rect 9020 -675 9055 -655
rect 9020 -700 9025 -675
rect 9050 -700 9055 -675
rect 9020 -725 9055 -700
rect 9020 -750 9025 -725
rect 9050 -750 9055 -725
rect 9020 -770 9055 -750
rect 9080 -585 9115 -575
rect 9080 -610 9085 -585
rect 9110 -610 9115 -585
rect 9080 -630 9115 -610
rect 9080 -655 9085 -630
rect 9110 -655 9115 -630
rect 9080 -675 9115 -655
rect 9080 -700 9085 -675
rect 9110 -700 9115 -675
rect 9080 -725 9115 -700
rect 9080 -750 9085 -725
rect 9110 -750 9115 -725
rect 9080 -770 9115 -750
rect 9140 -585 9175 -575
rect 9140 -610 9145 -585
rect 9170 -610 9175 -585
rect 9140 -630 9175 -610
rect 9140 -655 9145 -630
rect 9170 -655 9175 -630
rect 9140 -675 9175 -655
rect 9140 -700 9145 -675
rect 9170 -700 9175 -675
rect 9140 -725 9175 -700
rect 9140 -750 9145 -725
rect 9170 -750 9175 -725
rect 9140 -770 9175 -750
rect 9200 -585 9235 -575
rect 9200 -610 9205 -585
rect 9230 -610 9235 -585
rect 9200 -630 9235 -610
rect 9200 -655 9205 -630
rect 9230 -655 9235 -630
rect 9200 -675 9235 -655
rect 9200 -700 9205 -675
rect 9230 -700 9235 -675
rect 9200 -725 9235 -700
rect 9200 -750 9205 -725
rect 9230 -750 9235 -725
rect 9200 -770 9235 -750
rect 9260 -585 9295 -575
rect 9260 -610 9265 -585
rect 9290 -610 9295 -585
rect 9260 -630 9295 -610
rect 9260 -655 9265 -630
rect 9290 -655 9295 -630
rect 9260 -675 9295 -655
rect 9260 -700 9265 -675
rect 9290 -700 9295 -675
rect 9260 -725 9295 -700
rect 9260 -750 9265 -725
rect 9290 -750 9295 -725
rect 9260 -770 9295 -750
rect 9320 -585 9355 -575
rect 9320 -610 9325 -585
rect 9350 -610 9355 -585
rect 9320 -630 9355 -610
rect 9320 -655 9325 -630
rect 9350 -655 9355 -630
rect 9320 -675 9355 -655
rect 9320 -700 9325 -675
rect 9350 -700 9355 -675
rect 9320 -725 9355 -700
rect 9320 -750 9325 -725
rect 9350 -750 9355 -725
rect 9320 -770 9355 -750
rect 9380 -585 9415 -575
rect 9380 -610 9385 -585
rect 9410 -610 9415 -585
rect 9380 -630 9415 -610
rect 9380 -655 9385 -630
rect 9410 -655 9415 -630
rect 9380 -675 9415 -655
rect 9380 -700 9385 -675
rect 9410 -700 9415 -675
rect 9380 -725 9415 -700
rect 9380 -750 9385 -725
rect 9410 -750 9415 -725
rect 9380 -770 9415 -750
rect 9440 -585 9475 -575
rect 9440 -610 9445 -585
rect 9470 -610 9475 -585
rect 9440 -630 9475 -610
rect 9440 -655 9445 -630
rect 9470 -655 9475 -630
rect 9440 -675 9475 -655
rect 9440 -700 9445 -675
rect 9470 -700 9475 -675
rect 9440 -725 9475 -700
rect 9440 -750 9445 -725
rect 9470 -750 9475 -725
rect 9440 -770 9475 -750
rect 9500 -585 9535 -575
rect 9500 -610 9505 -585
rect 9530 -610 9535 -585
rect 9500 -630 9535 -610
rect 9500 -655 9505 -630
rect 9530 -655 9535 -630
rect 9500 -675 9535 -655
rect 9500 -700 9505 -675
rect 9530 -700 9535 -675
rect 9500 -725 9535 -700
rect 9500 -750 9505 -725
rect 9530 -750 9535 -725
rect 9500 -770 9535 -750
rect 9560 -585 9595 -575
rect 9560 -610 9565 -585
rect 9590 -610 9595 -585
rect 9560 -630 9595 -610
rect 9560 -655 9565 -630
rect 9590 -655 9595 -630
rect 9560 -675 9595 -655
rect 9560 -700 9565 -675
rect 9590 -700 9595 -675
rect 9560 -725 9595 -700
rect 9560 -750 9565 -725
rect 9590 -750 9595 -725
rect 9560 -770 9595 -750
rect 9620 -585 9655 -575
rect 9620 -610 9625 -585
rect 9650 -610 9655 -585
rect 9620 -630 9655 -610
rect 9620 -655 9625 -630
rect 9650 -655 9655 -630
rect 9620 -675 9655 -655
rect 9620 -700 9625 -675
rect 9650 -700 9655 -675
rect 9620 -725 9655 -700
rect 9620 -750 9625 -725
rect 9650 -750 9655 -725
rect 9620 -770 9655 -750
rect 9680 -585 9715 -575
rect 9680 -610 9685 -585
rect 9710 -610 9715 -585
rect 9680 -630 9715 -610
rect 9680 -655 9685 -630
rect 9710 -655 9715 -630
rect 9680 -675 9715 -655
rect 9680 -700 9685 -675
rect 9710 -700 9715 -675
rect 9680 -725 9715 -700
rect 9680 -750 9685 -725
rect 9710 -750 9715 -725
rect 9680 -770 9715 -750
rect 9740 -585 9775 -575
rect 9740 -610 9745 -585
rect 9770 -610 9775 -585
rect 9740 -630 9775 -610
rect 9740 -655 9745 -630
rect 9770 -655 9775 -630
rect 9740 -675 9775 -655
rect 9740 -700 9745 -675
rect 9770 -700 9775 -675
rect 9740 -725 9775 -700
rect 9740 -750 9745 -725
rect 9770 -750 9775 -725
rect 9740 -770 9775 -750
rect 9800 -585 9835 -575
rect 9800 -610 9805 -585
rect 9830 -610 9835 -585
rect 9800 -630 9835 -610
rect 9800 -655 9805 -630
rect 9830 -655 9835 -630
rect 9800 -675 9835 -655
rect 9800 -700 9805 -675
rect 9830 -700 9835 -675
rect 9800 -725 9835 -700
rect 9800 -750 9805 -725
rect 9830 -750 9835 -725
rect 9800 -770 9835 -750
rect 9860 -585 9895 -575
rect 9860 -610 9865 -585
rect 9890 -610 9895 -585
rect 9860 -630 9895 -610
rect 9860 -655 9865 -630
rect 9890 -655 9895 -630
rect 9860 -675 9895 -655
rect 9860 -700 9865 -675
rect 9890 -700 9895 -675
rect 9860 -725 9895 -700
rect 9860 -750 9865 -725
rect 9890 -750 9895 -725
rect 9860 -770 9895 -750
rect 9920 -585 9955 -575
rect 9920 -610 9925 -585
rect 9950 -610 9955 -585
rect 9920 -630 9955 -610
rect 9920 -655 9925 -630
rect 9950 -655 9955 -630
rect 9920 -675 9955 -655
rect 9920 -700 9925 -675
rect 9950 -700 9955 -675
rect 9920 -725 9955 -700
rect 9920 -750 9925 -725
rect 9950 -750 9955 -725
rect 9920 -770 9955 -750
rect 9980 -585 10015 -575
rect 9980 -610 9985 -585
rect 10010 -610 10015 -585
rect 9980 -630 10015 -610
rect 9980 -655 9985 -630
rect 10010 -655 10015 -630
rect 9980 -675 10015 -655
rect 9980 -700 9985 -675
rect 10010 -700 10015 -675
rect 9980 -725 10015 -700
rect 9980 -750 9985 -725
rect 10010 -750 10015 -725
rect 9980 -770 10015 -750
rect 10040 -585 10075 -575
rect 10040 -610 10045 -585
rect 10070 -610 10075 -585
rect 10040 -630 10075 -610
rect 10040 -655 10045 -630
rect 10070 -655 10075 -630
rect 10040 -675 10075 -655
rect 10040 -700 10045 -675
rect 10070 -700 10075 -675
rect 10040 -725 10075 -700
rect 10040 -750 10045 -725
rect 10070 -750 10075 -725
rect 10040 -770 10075 -750
rect 10100 -585 10135 -575
rect 10100 -610 10105 -585
rect 10130 -610 10135 -585
rect 10100 -630 10135 -610
rect 10100 -655 10105 -630
rect 10130 -655 10135 -630
rect 10100 -675 10135 -655
rect 10100 -700 10105 -675
rect 10130 -700 10135 -675
rect 10100 -725 10135 -700
rect 10100 -750 10105 -725
rect 10130 -750 10135 -725
rect 10100 -770 10135 -750
rect 10160 -585 10195 -575
rect 10160 -610 10165 -585
rect 10190 -610 10195 -585
rect 10160 -630 10195 -610
rect 10160 -655 10165 -630
rect 10190 -655 10195 -630
rect 10160 -675 10195 -655
rect 10160 -700 10165 -675
rect 10190 -700 10195 -675
rect 10160 -725 10195 -700
rect 10160 -750 10165 -725
rect 10190 -750 10195 -725
rect 10160 -770 10195 -750
rect 10220 -585 10255 -575
rect 10220 -610 10225 -585
rect 10250 -610 10255 -585
rect 10220 -630 10255 -610
rect 10220 -655 10225 -630
rect 10250 -655 10255 -630
rect 10220 -675 10255 -655
rect 10220 -700 10225 -675
rect 10250 -700 10255 -675
rect 10220 -725 10255 -700
rect 10220 -750 10225 -725
rect 10250 -750 10255 -725
rect 10220 -770 10255 -750
rect 10280 -585 10315 -575
rect 10280 -610 10285 -585
rect 10310 -610 10315 -585
rect 10280 -630 10315 -610
rect 10280 -655 10285 -630
rect 10310 -655 10315 -630
rect 10280 -675 10315 -655
rect 10280 -700 10285 -675
rect 10310 -700 10315 -675
rect 10280 -725 10315 -700
rect 10280 -750 10285 -725
rect 10310 -750 10315 -725
rect 10280 -770 10315 -750
rect 10340 -585 10375 -575
rect 10340 -610 10345 -585
rect 10370 -610 10375 -585
rect 10340 -630 10375 -610
rect 10340 -655 10345 -630
rect 10370 -655 10375 -630
rect 10340 -675 10375 -655
rect 10340 -700 10345 -675
rect 10370 -700 10375 -675
rect 10340 -725 10375 -700
rect 10340 -750 10345 -725
rect 10370 -750 10375 -725
rect 10340 -770 10375 -750
rect 10400 -585 10435 -575
rect 10400 -610 10405 -585
rect 10430 -610 10435 -585
rect 10400 -630 10435 -610
rect 10400 -655 10405 -630
rect 10430 -655 10435 -630
rect 10400 -675 10435 -655
rect 10400 -700 10405 -675
rect 10430 -700 10435 -675
rect 10400 -725 10435 -700
rect 10400 -750 10405 -725
rect 10430 -750 10435 -725
rect 10400 -770 10435 -750
rect 10460 -585 10495 -575
rect 10460 -610 10465 -585
rect 10490 -610 10495 -585
rect 10460 -630 10495 -610
rect 10460 -655 10465 -630
rect 10490 -655 10495 -630
rect 10460 -675 10495 -655
rect 10460 -700 10465 -675
rect 10490 -700 10495 -675
rect 10460 -725 10495 -700
rect 10460 -750 10465 -725
rect 10490 -750 10495 -725
rect 10460 -770 10495 -750
rect 10520 -585 10555 -575
rect 10520 -610 10525 -585
rect 10550 -610 10555 -585
rect 10520 -630 10555 -610
rect 10520 -655 10525 -630
rect 10550 -655 10555 -630
rect 10520 -675 10555 -655
rect 10520 -700 10525 -675
rect 10550 -700 10555 -675
rect 10520 -725 10555 -700
rect 10520 -750 10525 -725
rect 10550 -750 10555 -725
rect 10520 -770 10555 -750
rect 10580 -585 10615 -575
rect 10580 -610 10585 -585
rect 10610 -610 10615 -585
rect 10580 -630 10615 -610
rect 10580 -655 10585 -630
rect 10610 -655 10615 -630
rect 10580 -675 10615 -655
rect 10580 -700 10585 -675
rect 10610 -700 10615 -675
rect 10580 -725 10615 -700
rect 10580 -750 10585 -725
rect 10610 -750 10615 -725
rect 10580 -770 10615 -750
rect 10640 -585 10675 -575
rect 10640 -610 10645 -585
rect 10670 -610 10675 -585
rect 10640 -630 10675 -610
rect 10640 -655 10645 -630
rect 10670 -655 10675 -630
rect 10640 -675 10675 -655
rect 10640 -700 10645 -675
rect 10670 -700 10675 -675
rect 10640 -725 10675 -700
rect 10640 -750 10645 -725
rect 10670 -750 10675 -725
rect 10640 -770 10675 -750
rect 10700 -585 10735 -575
rect 10700 -610 10705 -585
rect 10730 -610 10735 -585
rect 10700 -630 10735 -610
rect 10700 -655 10705 -630
rect 10730 -655 10735 -630
rect 10700 -675 10735 -655
rect 10700 -700 10705 -675
rect 10730 -700 10735 -675
rect 10700 -725 10735 -700
rect 10700 -750 10705 -725
rect 10730 -750 10735 -725
rect 10700 -770 10735 -750
rect 10760 -585 10795 -575
rect 10760 -610 10765 -585
rect 10790 -610 10795 -585
rect 10760 -630 10795 -610
rect 10760 -655 10765 -630
rect 10790 -655 10795 -630
rect 10760 -675 10795 -655
rect 10760 -700 10765 -675
rect 10790 -700 10795 -675
rect 10760 -725 10795 -700
rect 10760 -750 10765 -725
rect 10790 -750 10795 -725
rect 10760 -770 10795 -750
rect 10820 -585 10855 -575
rect 10820 -610 10825 -585
rect 10850 -610 10855 -585
rect 10820 -630 10855 -610
rect 10820 -655 10825 -630
rect 10850 -655 10855 -630
rect 10820 -675 10855 -655
rect 10820 -700 10825 -675
rect 10850 -700 10855 -675
rect 10820 -725 10855 -700
rect 10820 -750 10825 -725
rect 10850 -750 10855 -725
rect 10820 -770 10855 -750
rect 10880 -585 10915 -575
rect 10880 -610 10885 -585
rect 10910 -610 10915 -585
rect 10880 -630 10915 -610
rect 10880 -655 10885 -630
rect 10910 -655 10915 -630
rect 10880 -675 10915 -655
rect 10880 -700 10885 -675
rect 10910 -700 10915 -675
rect 10880 -725 10915 -700
rect 10880 -750 10885 -725
rect 10910 -750 10915 -725
rect 10880 -770 10915 -750
rect 10940 -585 10975 -575
rect 10940 -610 10945 -585
rect 10970 -610 10975 -585
rect 10940 -630 10975 -610
rect 10940 -655 10945 -630
rect 10970 -655 10975 -630
rect 10940 -675 10975 -655
rect 10940 -700 10945 -675
rect 10970 -700 10975 -675
rect 10940 -725 10975 -700
rect 10940 -750 10945 -725
rect 10970 -750 10975 -725
rect 10940 -770 10975 -750
rect 11000 -585 11035 -575
rect 11000 -610 11005 -585
rect 11030 -610 11035 -585
rect 11000 -630 11035 -610
rect 11000 -655 11005 -630
rect 11030 -655 11035 -630
rect 11000 -675 11035 -655
rect 11000 -700 11005 -675
rect 11030 -700 11035 -675
rect 11000 -725 11035 -700
rect 11000 -750 11005 -725
rect 11030 -750 11035 -725
rect 11000 -770 11035 -750
rect 11060 -585 11095 -575
rect 11060 -610 11065 -585
rect 11090 -610 11095 -585
rect 11060 -630 11095 -610
rect 11060 -655 11065 -630
rect 11090 -655 11095 -630
rect 11060 -675 11095 -655
rect 11060 -700 11065 -675
rect 11090 -700 11095 -675
rect 11060 -725 11095 -700
rect 11060 -750 11065 -725
rect 11090 -750 11095 -725
rect 11060 -770 11095 -750
rect 11120 -585 11155 -575
rect 11120 -610 11125 -585
rect 11150 -610 11155 -585
rect 11120 -630 11155 -610
rect 11120 -655 11125 -630
rect 11150 -655 11155 -630
rect 11120 -675 11155 -655
rect 11120 -700 11125 -675
rect 11150 -700 11155 -675
rect 11120 -725 11155 -700
rect 11120 -750 11125 -725
rect 11150 -750 11155 -725
rect 11120 -770 11155 -750
rect 11180 -585 11215 -575
rect 11180 -610 11185 -585
rect 11210 -610 11215 -585
rect 11180 -630 11215 -610
rect 11180 -655 11185 -630
rect 11210 -655 11215 -630
rect 11180 -675 11215 -655
rect 11180 -700 11185 -675
rect 11210 -700 11215 -675
rect 11180 -725 11215 -700
rect 11180 -750 11185 -725
rect 11210 -750 11215 -725
rect 11180 -770 11215 -750
rect 11240 -585 11275 -575
rect 11240 -610 11245 -585
rect 11270 -610 11275 -585
rect 11240 -630 11275 -610
rect 11240 -655 11245 -630
rect 11270 -655 11275 -630
rect 11240 -675 11275 -655
rect 11240 -700 11245 -675
rect 11270 -700 11275 -675
rect 11240 -725 11275 -700
rect 11240 -750 11245 -725
rect 11270 -750 11275 -725
rect 11240 -770 11275 -750
rect 11300 -585 11335 -575
rect 11300 -610 11305 -585
rect 11330 -610 11335 -585
rect 11300 -630 11335 -610
rect 11300 -655 11305 -630
rect 11330 -655 11335 -630
rect 11300 -675 11335 -655
rect 11300 -700 11305 -675
rect 11330 -700 11335 -675
rect 11300 -725 11335 -700
rect 11300 -750 11305 -725
rect 11330 -750 11335 -725
rect 11300 -770 11335 -750
rect 11360 -585 11395 -575
rect 11360 -610 11365 -585
rect 11390 -610 11395 -585
rect 11360 -630 11395 -610
rect 11360 -655 11365 -630
rect 11390 -655 11395 -630
rect 11360 -675 11395 -655
rect 11360 -700 11365 -675
rect 11390 -700 11395 -675
rect 11360 -725 11395 -700
rect 11360 -750 11365 -725
rect 11390 -750 11395 -725
rect 11360 -770 11395 -750
rect 11420 -585 11455 -575
rect 11420 -610 11425 -585
rect 11450 -610 11455 -585
rect 11420 -630 11455 -610
rect 11420 -655 11425 -630
rect 11450 -655 11455 -630
rect 11420 -675 11455 -655
rect 11420 -700 11425 -675
rect 11450 -700 11455 -675
rect 11420 -725 11455 -700
rect 11420 -750 11425 -725
rect 11450 -750 11455 -725
rect 11420 -770 11455 -750
rect 11480 -585 11515 -575
rect 11480 -610 11485 -585
rect 11510 -610 11515 -585
rect 11480 -630 11515 -610
rect 11480 -655 11485 -630
rect 11510 -655 11515 -630
rect 11480 -675 11515 -655
rect 11480 -700 11485 -675
rect 11510 -700 11515 -675
rect 11480 -725 11515 -700
rect 11480 -750 11485 -725
rect 11510 -750 11515 -725
rect 11480 -770 11515 -750
rect 11540 -585 11575 -575
rect 11540 -610 11545 -585
rect 11570 -610 11575 -585
rect 11540 -630 11575 -610
rect 11540 -655 11545 -630
rect 11570 -655 11575 -630
rect 11540 -675 11575 -655
rect 11540 -700 11545 -675
rect 11570 -700 11575 -675
rect 11540 -725 11575 -700
rect 11540 -750 11545 -725
rect 11570 -750 11575 -725
rect 11540 -770 11575 -750
rect 11600 -585 11635 -575
rect 11600 -610 11605 -585
rect 11630 -610 11635 -585
rect 11600 -630 11635 -610
rect 11600 -655 11605 -630
rect 11630 -655 11635 -630
rect 11600 -675 11635 -655
rect 11600 -700 11605 -675
rect 11630 -700 11635 -675
rect 11600 -725 11635 -700
rect 11600 -750 11605 -725
rect 11630 -750 11635 -725
rect 11600 -770 11635 -750
rect 11660 -585 11695 -575
rect 11660 -610 11665 -585
rect 11690 -610 11695 -585
rect 11660 -630 11695 -610
rect 11660 -655 11665 -630
rect 11690 -655 11695 -630
rect 11660 -675 11695 -655
rect 11660 -700 11665 -675
rect 11690 -700 11695 -675
rect 11660 -725 11695 -700
rect 11660 -750 11665 -725
rect 11690 -750 11695 -725
rect 11660 -770 11695 -750
rect 11720 -585 11755 -575
rect 11720 -610 11725 -585
rect 11750 -610 11755 -585
rect 11720 -630 11755 -610
rect 11720 -655 11725 -630
rect 11750 -655 11755 -630
rect 11720 -675 11755 -655
rect 11720 -700 11725 -675
rect 11750 -700 11755 -675
rect 11720 -725 11755 -700
rect 11720 -750 11725 -725
rect 11750 -750 11755 -725
rect 11720 -770 11755 -750
rect 11780 -585 11815 -575
rect 11780 -610 11785 -585
rect 11810 -610 11815 -585
rect 11780 -630 11815 -610
rect 11780 -655 11785 -630
rect 11810 -655 11815 -630
rect 11780 -675 11815 -655
rect 11780 -700 11785 -675
rect 11810 -700 11815 -675
rect 11780 -725 11815 -700
rect 11780 -750 11785 -725
rect 11810 -750 11815 -725
rect 11780 -770 11815 -750
rect 11840 -585 11875 -575
rect 11840 -610 11845 -585
rect 11870 -610 11875 -585
rect 11840 -630 11875 -610
rect 11840 -655 11845 -630
rect 11870 -655 11875 -630
rect 11840 -675 11875 -655
rect 11840 -700 11845 -675
rect 11870 -700 11875 -675
rect 11840 -725 11875 -700
rect 11840 -750 11845 -725
rect 11870 -750 11875 -725
rect 11840 -770 11875 -750
rect 11900 -585 11935 -575
rect 11900 -610 11905 -585
rect 11930 -610 11935 -585
rect 11900 -630 11935 -610
rect 11900 -655 11905 -630
rect 11930 -655 11935 -630
rect 11900 -675 11935 -655
rect 11900 -700 11905 -675
rect 11930 -700 11935 -675
rect 11900 -725 11935 -700
rect 11900 -750 11905 -725
rect 11930 -750 11935 -725
rect 11900 -770 11935 -750
rect 11960 -585 11995 -575
rect 11960 -610 11965 -585
rect 11990 -610 11995 -585
rect 11960 -630 11995 -610
rect 11960 -655 11965 -630
rect 11990 -655 11995 -630
rect 11960 -675 11995 -655
rect 11960 -700 11965 -675
rect 11990 -700 11995 -675
rect 11960 -725 11995 -700
rect 11960 -750 11965 -725
rect 11990 -750 11995 -725
rect 11960 -770 11995 -750
rect 12020 -585 12055 -575
rect 12020 -610 12025 -585
rect 12050 -610 12055 -585
rect 12020 -630 12055 -610
rect 12020 -655 12025 -630
rect 12050 -655 12055 -630
rect 12020 -675 12055 -655
rect 12020 -700 12025 -675
rect 12050 -700 12055 -675
rect 12020 -725 12055 -700
rect 12020 -750 12025 -725
rect 12050 -750 12055 -725
rect 12020 -770 12055 -750
rect 12080 -585 12115 -575
rect 12080 -610 12085 -585
rect 12110 -610 12115 -585
rect 12080 -630 12115 -610
rect 12080 -655 12085 -630
rect 12110 -655 12115 -630
rect 12080 -675 12115 -655
rect 12080 -700 12085 -675
rect 12110 -700 12115 -675
rect 12080 -725 12115 -700
rect 12080 -750 12085 -725
rect 12110 -750 12115 -725
rect 12080 -770 12115 -750
rect 12140 -585 12175 -575
rect 12140 -610 12145 -585
rect 12170 -610 12175 -585
rect 12140 -630 12175 -610
rect 12140 -655 12145 -630
rect 12170 -655 12175 -630
rect 12140 -675 12175 -655
rect 12140 -700 12145 -675
rect 12170 -700 12175 -675
rect 12140 -725 12175 -700
rect 12140 -750 12145 -725
rect 12170 -750 12175 -725
rect 12140 -770 12175 -750
rect 12200 -585 12235 -575
rect 12200 -610 12205 -585
rect 12230 -610 12235 -585
rect 12200 -630 12235 -610
rect 12200 -655 12205 -630
rect 12230 -655 12235 -630
rect 12200 -675 12235 -655
rect 12200 -700 12205 -675
rect 12230 -700 12235 -675
rect 12200 -725 12235 -700
rect 12200 -750 12205 -725
rect 12230 -750 12235 -725
rect 12200 -770 12235 -750
rect 12260 -585 12295 -575
rect 12260 -610 12265 -585
rect 12290 -610 12295 -585
rect 12260 -630 12295 -610
rect 12260 -655 12265 -630
rect 12290 -655 12295 -630
rect 12260 -675 12295 -655
rect 12260 -700 12265 -675
rect 12290 -700 12295 -675
rect 12260 -725 12295 -700
rect 12260 -750 12265 -725
rect 12290 -750 12295 -725
rect 12260 -770 12295 -750
rect 12320 -585 12355 -575
rect 12320 -610 12325 -585
rect 12350 -610 12355 -585
rect 12320 -630 12355 -610
rect 12320 -655 12325 -630
rect 12350 -655 12355 -630
rect 12320 -675 12355 -655
rect 12320 -700 12325 -675
rect 12350 -700 12355 -675
rect 12320 -725 12355 -700
rect 12320 -750 12325 -725
rect 12350 -750 12355 -725
rect 12320 -770 12355 -750
rect 12380 -585 12415 -575
rect 12380 -610 12385 -585
rect 12410 -610 12415 -585
rect 12380 -630 12415 -610
rect 12380 -655 12385 -630
rect 12410 -655 12415 -630
rect 12380 -675 12415 -655
rect 12380 -700 12385 -675
rect 12410 -700 12415 -675
rect 12380 -725 12415 -700
rect 12380 -750 12385 -725
rect 12410 -750 12415 -725
rect 12380 -770 12415 -750
rect 12440 -585 12475 -575
rect 12440 -610 12445 -585
rect 12470 -610 12475 -585
rect 12440 -630 12475 -610
rect 12440 -655 12445 -630
rect 12470 -655 12475 -630
rect 12440 -675 12475 -655
rect 12440 -700 12445 -675
rect 12470 -700 12475 -675
rect 12440 -725 12475 -700
rect 12440 -750 12445 -725
rect 12470 -750 12475 -725
rect 12440 -770 12475 -750
rect 12500 -585 12535 -575
rect 12500 -610 12505 -585
rect 12530 -610 12535 -585
rect 12500 -630 12535 -610
rect 12500 -655 12505 -630
rect 12530 -655 12535 -630
rect 12500 -675 12535 -655
rect 12500 -700 12505 -675
rect 12530 -700 12535 -675
rect 12500 -725 12535 -700
rect 12500 -750 12505 -725
rect 12530 -750 12535 -725
rect 12500 -770 12535 -750
rect 12560 -585 12595 -575
rect 12560 -610 12565 -585
rect 12590 -610 12595 -585
rect 12560 -630 12595 -610
rect 12560 -655 12565 -630
rect 12590 -655 12595 -630
rect 12560 -675 12595 -655
rect 12560 -700 12565 -675
rect 12590 -700 12595 -675
rect 12560 -725 12595 -700
rect 12560 -750 12565 -725
rect 12590 -750 12595 -725
rect 12560 -770 12595 -750
rect 12620 -585 12655 -575
rect 12620 -610 12625 -585
rect 12650 -610 12655 -585
rect 12620 -630 12655 -610
rect 12620 -655 12625 -630
rect 12650 -655 12655 -630
rect 12620 -675 12655 -655
rect 12620 -700 12625 -675
rect 12650 -700 12655 -675
rect 12620 -725 12655 -700
rect 12620 -750 12625 -725
rect 12650 -750 12655 -725
rect 12620 -770 12655 -750
rect 12680 -585 12715 -575
rect 12680 -610 12685 -585
rect 12710 -610 12715 -585
rect 12680 -630 12715 -610
rect 12680 -655 12685 -630
rect 12710 -655 12715 -630
rect 12680 -675 12715 -655
rect 12680 -700 12685 -675
rect 12710 -700 12715 -675
rect 12680 -725 12715 -700
rect 12680 -750 12685 -725
rect 12710 -750 12715 -725
rect 12680 -770 12715 -750
rect 12740 -585 12775 -575
rect 12740 -610 12745 -585
rect 12770 -610 12775 -585
rect 12740 -630 12775 -610
rect 12740 -655 12745 -630
rect 12770 -655 12775 -630
rect 12740 -675 12775 -655
rect 12740 -700 12745 -675
rect 12770 -700 12775 -675
rect 12740 -725 12775 -700
rect 12740 -750 12745 -725
rect 12770 -750 12775 -725
rect 12740 -770 12775 -750
rect 12800 -585 12835 -575
rect 12800 -610 12805 -585
rect 12830 -610 12835 -585
rect 12800 -630 12835 -610
rect 12800 -655 12805 -630
rect 12830 -655 12835 -630
rect 12800 -675 12835 -655
rect 12800 -700 12805 -675
rect 12830 -700 12835 -675
rect 12800 -725 12835 -700
rect 12800 -750 12805 -725
rect 12830 -750 12835 -725
rect 12800 -770 12835 -750
rect 12860 -585 12895 -575
rect 12860 -610 12865 -585
rect 12890 -610 12895 -585
rect 12860 -630 12895 -610
rect 12860 -655 12865 -630
rect 12890 -655 12895 -630
rect 12860 -675 12895 -655
rect 12860 -700 12865 -675
rect 12890 -700 12895 -675
rect 12860 -725 12895 -700
rect 12860 -750 12865 -725
rect 12890 -750 12895 -725
rect 12860 -770 12895 -750
rect 12920 -585 12955 -575
rect 12920 -610 12925 -585
rect 12950 -610 12955 -585
rect 12920 -630 12955 -610
rect 12920 -655 12925 -630
rect 12950 -655 12955 -630
rect 12920 -675 12955 -655
rect 12920 -700 12925 -675
rect 12950 -700 12955 -675
rect 12920 -725 12955 -700
rect 12920 -750 12925 -725
rect 12950 -750 12955 -725
rect 12920 -770 12955 -750
rect 12980 -585 13015 -575
rect 12980 -610 12985 -585
rect 13010 -610 13015 -585
rect 12980 -630 13015 -610
rect 12980 -655 12985 -630
rect 13010 -655 13015 -630
rect 12980 -675 13015 -655
rect 12980 -700 12985 -675
rect 13010 -700 13015 -675
rect 12980 -725 13015 -700
rect 12980 -750 12985 -725
rect 13010 -750 13015 -725
rect 12980 -770 13015 -750
rect 13040 -585 13075 -575
rect 13040 -610 13045 -585
rect 13070 -610 13075 -585
rect 13040 -630 13075 -610
rect 13040 -655 13045 -630
rect 13070 -655 13075 -630
rect 13040 -675 13075 -655
rect 13040 -700 13045 -675
rect 13070 -700 13075 -675
rect 13040 -725 13075 -700
rect 13040 -750 13045 -725
rect 13070 -750 13075 -725
rect 13040 -770 13075 -750
rect 13100 -585 13135 -575
rect 13100 -610 13105 -585
rect 13130 -610 13135 -585
rect 13100 -630 13135 -610
rect 13100 -655 13105 -630
rect 13130 -655 13135 -630
rect 13100 -675 13135 -655
rect 13100 -700 13105 -675
rect 13130 -700 13135 -675
rect 13100 -725 13135 -700
rect 13100 -750 13105 -725
rect 13130 -750 13135 -725
rect 13100 -770 13135 -750
rect 13160 -585 13195 -575
rect 13160 -610 13165 -585
rect 13190 -610 13195 -585
rect 13160 -630 13195 -610
rect 13160 -655 13165 -630
rect 13190 -655 13195 -630
rect 13160 -675 13195 -655
rect 13160 -700 13165 -675
rect 13190 -700 13195 -675
rect 13160 -725 13195 -700
rect 13160 -750 13165 -725
rect 13190 -750 13195 -725
rect 13160 -770 13195 -750
rect 13220 -585 13255 -575
rect 13220 -610 13225 -585
rect 13250 -610 13255 -585
rect 13220 -630 13255 -610
rect 13220 -655 13225 -630
rect 13250 -655 13255 -630
rect 13220 -675 13255 -655
rect 13220 -700 13225 -675
rect 13250 -700 13255 -675
rect 13220 -725 13255 -700
rect 13220 -750 13225 -725
rect 13250 -750 13255 -725
rect 13220 -770 13255 -750
rect 13280 -585 13315 -575
rect 13280 -610 13285 -585
rect 13310 -610 13315 -585
rect 13280 -630 13315 -610
rect 13280 -655 13285 -630
rect 13310 -655 13315 -630
rect 13280 -675 13315 -655
rect 13280 -700 13285 -675
rect 13310 -700 13315 -675
rect 13280 -725 13315 -700
rect 13280 -750 13285 -725
rect 13310 -750 13315 -725
rect 13280 -770 13315 -750
rect 13340 -585 13375 -575
rect 13340 -610 13345 -585
rect 13370 -610 13375 -585
rect 13340 -630 13375 -610
rect 13340 -655 13345 -630
rect 13370 -655 13375 -630
rect 13340 -675 13375 -655
rect 13340 -700 13345 -675
rect 13370 -700 13375 -675
rect 13340 -725 13375 -700
rect 13340 -750 13345 -725
rect 13370 -750 13375 -725
rect 13340 -770 13375 -750
rect 13400 -585 13435 -575
rect 13400 -610 13405 -585
rect 13430 -610 13435 -585
rect 13400 -630 13435 -610
rect 13400 -655 13405 -630
rect 13430 -655 13435 -630
rect 13400 -675 13435 -655
rect 13400 -700 13405 -675
rect 13430 -700 13435 -675
rect 13400 -725 13435 -700
rect 13400 -750 13405 -725
rect 13430 -750 13435 -725
rect 13400 -770 13435 -750
rect 13460 -585 13495 -575
rect 13460 -610 13465 -585
rect 13490 -610 13495 -585
rect 13460 -630 13495 -610
rect 13460 -655 13465 -630
rect 13490 -655 13495 -630
rect 13460 -675 13495 -655
rect 13460 -700 13465 -675
rect 13490 -700 13495 -675
rect 13460 -725 13495 -700
rect 13460 -750 13465 -725
rect 13490 -750 13495 -725
rect 13460 -770 13495 -750
rect 13520 -585 13555 -575
rect 13520 -610 13525 -585
rect 13550 -610 13555 -585
rect 13520 -630 13555 -610
rect 13520 -655 13525 -630
rect 13550 -655 13555 -630
rect 13520 -675 13555 -655
rect 13520 -700 13525 -675
rect 13550 -700 13555 -675
rect 13520 -725 13555 -700
rect 13520 -750 13525 -725
rect 13550 -750 13555 -725
rect 13520 -770 13555 -750
rect 13580 -585 13615 -575
rect 13580 -610 13585 -585
rect 13610 -610 13615 -585
rect 13580 -630 13615 -610
rect 13580 -655 13585 -630
rect 13610 -655 13615 -630
rect 13580 -675 13615 -655
rect 13580 -700 13585 -675
rect 13610 -700 13615 -675
rect 13580 -725 13615 -700
rect 13580 -750 13585 -725
rect 13610 -750 13615 -725
rect 13580 -770 13615 -750
rect 13640 -585 13675 -575
rect 13640 -610 13645 -585
rect 13670 -610 13675 -585
rect 13640 -630 13675 -610
rect 13640 -655 13645 -630
rect 13670 -655 13675 -630
rect 13640 -675 13675 -655
rect 13640 -700 13645 -675
rect 13670 -700 13675 -675
rect 13640 -725 13675 -700
rect 13640 -750 13645 -725
rect 13670 -750 13675 -725
rect 13640 -770 13675 -750
rect 13700 -585 13735 -575
rect 13700 -610 13705 -585
rect 13730 -610 13735 -585
rect 13700 -630 13735 -610
rect 13700 -655 13705 -630
rect 13730 -655 13735 -630
rect 13700 -675 13735 -655
rect 13700 -700 13705 -675
rect 13730 -700 13735 -675
rect 13700 -725 13735 -700
rect 13700 -750 13705 -725
rect 13730 -750 13735 -725
rect 13700 -770 13735 -750
rect 13760 -585 13795 -575
rect 13760 -610 13765 -585
rect 13790 -610 13795 -585
rect 13760 -630 13795 -610
rect 13760 -655 13765 -630
rect 13790 -655 13795 -630
rect 13760 -675 13795 -655
rect 13760 -700 13765 -675
rect 13790 -700 13795 -675
rect 13760 -725 13795 -700
rect 13760 -750 13765 -725
rect 13790 -750 13795 -725
rect 13760 -770 13795 -750
rect 13820 -585 13855 -575
rect 13820 -610 13825 -585
rect 13850 -610 13855 -585
rect 13820 -630 13855 -610
rect 13820 -655 13825 -630
rect 13850 -655 13855 -630
rect 13820 -675 13855 -655
rect 13820 -700 13825 -675
rect 13850 -700 13855 -675
rect 13820 -725 13855 -700
rect 13820 -750 13825 -725
rect 13850 -750 13855 -725
rect 13820 -770 13855 -750
rect 13880 -585 13915 -575
rect 13880 -610 13885 -585
rect 13910 -610 13915 -585
rect 13880 -630 13915 -610
rect 13880 -655 13885 -630
rect 13910 -655 13915 -630
rect 13880 -675 13915 -655
rect 13880 -700 13885 -675
rect 13910 -700 13915 -675
rect 13880 -725 13915 -700
rect 13880 -750 13885 -725
rect 13910 -750 13915 -725
rect 13880 -770 13915 -750
rect 13940 -585 13975 -575
rect 13940 -610 13945 -585
rect 13970 -610 13975 -585
rect 13940 -630 13975 -610
rect 13940 -655 13945 -630
rect 13970 -655 13975 -630
rect 13940 -675 13975 -655
rect 13940 -700 13945 -675
rect 13970 -700 13975 -675
rect 13940 -725 13975 -700
rect 13940 -750 13945 -725
rect 13970 -750 13975 -725
rect 13940 -770 13975 -750
rect 14000 -585 14035 -575
rect 14000 -610 14005 -585
rect 14030 -610 14035 -585
rect 14000 -630 14035 -610
rect 14000 -655 14005 -630
rect 14030 -655 14035 -630
rect 14000 -675 14035 -655
rect 14000 -700 14005 -675
rect 14030 -700 14035 -675
rect 14000 -725 14035 -700
rect 14000 -750 14005 -725
rect 14030 -750 14035 -725
rect 14000 -770 14035 -750
rect 14060 -585 14095 -575
rect 14060 -610 14065 -585
rect 14090 -610 14095 -585
rect 14060 -630 14095 -610
rect 14060 -655 14065 -630
rect 14090 -655 14095 -630
rect 14060 -675 14095 -655
rect 14060 -700 14065 -675
rect 14090 -700 14095 -675
rect 14060 -725 14095 -700
rect 14060 -750 14065 -725
rect 14090 -750 14095 -725
rect 14060 -770 14095 -750
rect 14120 -585 14155 -575
rect 14120 -610 14125 -585
rect 14150 -610 14155 -585
rect 14120 -630 14155 -610
rect 14120 -655 14125 -630
rect 14150 -655 14155 -630
rect 14120 -675 14155 -655
rect 14120 -700 14125 -675
rect 14150 -700 14155 -675
rect 14120 -725 14155 -700
rect 14120 -750 14125 -725
rect 14150 -750 14155 -725
rect 14120 -770 14155 -750
rect 14180 -585 14215 -575
rect 14180 -610 14185 -585
rect 14210 -610 14215 -585
rect 14180 -630 14215 -610
rect 14180 -655 14185 -630
rect 14210 -655 14215 -630
rect 14180 -675 14215 -655
rect 14180 -700 14185 -675
rect 14210 -700 14215 -675
rect 14180 -725 14215 -700
rect 14180 -750 14185 -725
rect 14210 -750 14215 -725
rect 14180 -770 14215 -750
rect 14240 -585 14275 -575
rect 14240 -610 14245 -585
rect 14270 -610 14275 -585
rect 14240 -630 14275 -610
rect 14240 -655 14245 -630
rect 14270 -655 14275 -630
rect 14240 -675 14275 -655
rect 14240 -700 14245 -675
rect 14270 -700 14275 -675
rect 14240 -725 14275 -700
rect 14240 -750 14245 -725
rect 14270 -750 14275 -725
rect 14240 -770 14275 -750
rect 14300 -585 14335 -575
rect 14300 -610 14305 -585
rect 14330 -610 14335 -585
rect 14300 -630 14335 -610
rect 14300 -655 14305 -630
rect 14330 -655 14335 -630
rect 14300 -675 14335 -655
rect 14300 -700 14305 -675
rect 14330 -700 14335 -675
rect 14300 -725 14335 -700
rect 14300 -750 14305 -725
rect 14330 -750 14335 -725
rect 14300 -770 14335 -750
rect 14360 -585 14395 -575
rect 14360 -610 14365 -585
rect 14390 -610 14395 -585
rect 14360 -630 14395 -610
rect 14360 -655 14365 -630
rect 14390 -655 14395 -630
rect 14360 -675 14395 -655
rect 14360 -700 14365 -675
rect 14390 -700 14395 -675
rect 14360 -725 14395 -700
rect 14360 -750 14365 -725
rect 14390 -750 14395 -725
rect 14360 -770 14395 -750
rect 14420 -585 14455 -575
rect 14420 -610 14425 -585
rect 14450 -610 14455 -585
rect 14420 -630 14455 -610
rect 14420 -655 14425 -630
rect 14450 -655 14455 -630
rect 14420 -675 14455 -655
rect 14420 -700 14425 -675
rect 14450 -700 14455 -675
rect 14420 -725 14455 -700
rect 14420 -750 14425 -725
rect 14450 -750 14455 -725
rect 14420 -770 14455 -750
rect 14480 -585 14515 -575
rect 14480 -610 14485 -585
rect 14510 -610 14515 -585
rect 14480 -630 14515 -610
rect 14480 -655 14485 -630
rect 14510 -655 14515 -630
rect 14480 -675 14515 -655
rect 14480 -700 14485 -675
rect 14510 -700 14515 -675
rect 14480 -725 14515 -700
rect 14480 -750 14485 -725
rect 14510 -750 14515 -725
rect 14480 -770 14515 -750
rect 14540 -585 14575 -575
rect 14540 -610 14545 -585
rect 14570 -610 14575 -585
rect 14540 -630 14575 -610
rect 14540 -655 14545 -630
rect 14570 -655 14575 -630
rect 14540 -675 14575 -655
rect 14540 -700 14545 -675
rect 14570 -700 14575 -675
rect 14540 -725 14575 -700
rect 14540 -750 14545 -725
rect 14570 -750 14575 -725
rect 14540 -770 14575 -750
rect 14600 -585 14635 -575
rect 14600 -610 14605 -585
rect 14630 -610 14635 -585
rect 14600 -630 14635 -610
rect 14600 -655 14605 -630
rect 14630 -655 14635 -630
rect 14600 -675 14635 -655
rect 14600 -700 14605 -675
rect 14630 -700 14635 -675
rect 14600 -725 14635 -700
rect 14600 -750 14605 -725
rect 14630 -750 14635 -725
rect 14600 -770 14635 -750
rect 14660 -585 14695 -575
rect 14660 -610 14665 -585
rect 14690 -610 14695 -585
rect 14660 -630 14695 -610
rect 14660 -655 14665 -630
rect 14690 -655 14695 -630
rect 14660 -675 14695 -655
rect 14660 -700 14665 -675
rect 14690 -700 14695 -675
rect 14660 -725 14695 -700
rect 14660 -750 14665 -725
rect 14690 -750 14695 -725
rect 14660 -770 14695 -750
rect 14720 -585 14755 -575
rect 14720 -610 14725 -585
rect 14750 -610 14755 -585
rect 14720 -630 14755 -610
rect 14720 -655 14725 -630
rect 14750 -655 14755 -630
rect 14720 -675 14755 -655
rect 14720 -700 14725 -675
rect 14750 -700 14755 -675
rect 14720 -725 14755 -700
rect 14720 -750 14725 -725
rect 14750 -750 14755 -725
rect 14720 -770 14755 -750
rect 14780 -585 14815 -575
rect 14780 -610 14785 -585
rect 14810 -610 14815 -585
rect 14780 -630 14815 -610
rect 14780 -655 14785 -630
rect 14810 -655 14815 -630
rect 14780 -675 14815 -655
rect 14780 -700 14785 -675
rect 14810 -700 14815 -675
rect 14780 -725 14815 -700
rect 14780 -750 14785 -725
rect 14810 -750 14815 -725
rect 14780 -770 14815 -750
rect 14840 -585 14875 -575
rect 14840 -610 14845 -585
rect 14870 -610 14875 -585
rect 14840 -630 14875 -610
rect 14840 -655 14845 -630
rect 14870 -655 14875 -630
rect 14840 -675 14875 -655
rect 14840 -700 14845 -675
rect 14870 -700 14875 -675
rect 14840 -725 14875 -700
rect 14840 -750 14845 -725
rect 14870 -750 14875 -725
rect 14840 -770 14875 -750
rect 14900 -585 14935 -575
rect 14900 -610 14905 -585
rect 14930 -610 14935 -585
rect 14900 -630 14935 -610
rect 14900 -655 14905 -630
rect 14930 -655 14935 -630
rect 14900 -675 14935 -655
rect 14900 -700 14905 -675
rect 14930 -700 14935 -675
rect 14900 -725 14935 -700
rect 14900 -750 14905 -725
rect 14930 -750 14935 -725
rect 14900 -770 14935 -750
rect 14960 -585 14995 -575
rect 14960 -610 14965 -585
rect 14990 -610 14995 -585
rect 14960 -630 14995 -610
rect 14960 -655 14965 -630
rect 14990 -655 14995 -630
rect 14960 -675 14995 -655
rect 14960 -700 14965 -675
rect 14990 -700 14995 -675
rect 14960 -725 14995 -700
rect 14960 -750 14965 -725
rect 14990 -750 14995 -725
rect 14960 -770 14995 -750
rect 15020 -585 15055 -575
rect 15020 -610 15025 -585
rect 15050 -610 15055 -585
rect 15020 -630 15055 -610
rect 15020 -655 15025 -630
rect 15050 -655 15055 -630
rect 15020 -675 15055 -655
rect 15020 -700 15025 -675
rect 15050 -700 15055 -675
rect 15020 -725 15055 -700
rect 15020 -750 15025 -725
rect 15050 -750 15055 -725
rect 15020 -770 15055 -750
rect 15080 -585 15115 -575
rect 15080 -610 15085 -585
rect 15110 -610 15115 -585
rect 15080 -630 15115 -610
rect 15080 -655 15085 -630
rect 15110 -655 15115 -630
rect 15080 -675 15115 -655
rect 15080 -700 15085 -675
rect 15110 -700 15115 -675
rect 15080 -725 15115 -700
rect 15080 -750 15085 -725
rect 15110 -750 15115 -725
rect 15080 -770 15115 -750
rect 15140 -585 15175 -575
rect 15140 -610 15145 -585
rect 15170 -610 15175 -585
rect 15140 -630 15175 -610
rect 15140 -655 15145 -630
rect 15170 -655 15175 -630
rect 15140 -675 15175 -655
rect 15140 -700 15145 -675
rect 15170 -700 15175 -675
rect 15140 -725 15175 -700
rect 15140 -750 15145 -725
rect 15170 -750 15175 -725
rect 15140 -770 15175 -750
rect 15200 -585 15235 -575
rect 15200 -610 15205 -585
rect 15230 -610 15235 -585
rect 15200 -630 15235 -610
rect 15200 -655 15205 -630
rect 15230 -655 15235 -630
rect 15200 -675 15235 -655
rect 15200 -700 15205 -675
rect 15230 -700 15235 -675
rect 15200 -725 15235 -700
rect 15200 -750 15205 -725
rect 15230 -750 15235 -725
rect 15200 -770 15235 -750
rect 15260 -585 15295 -575
rect 15260 -610 15265 -585
rect 15290 -610 15295 -585
rect 15260 -630 15295 -610
rect 15260 -655 15265 -630
rect 15290 -655 15295 -630
rect 15260 -675 15295 -655
rect 15260 -700 15265 -675
rect 15290 -700 15295 -675
rect 15260 -725 15295 -700
rect 15260 -750 15265 -725
rect 15290 -750 15295 -725
rect 15260 -770 15295 -750
rect 15320 -585 15355 -575
rect 15320 -610 15325 -585
rect 15350 -610 15355 -585
rect 15320 -630 15355 -610
rect 15320 -655 15325 -630
rect 15350 -655 15355 -630
rect 15320 -675 15355 -655
rect 15320 -700 15325 -675
rect 15350 -700 15355 -675
rect 15320 -725 15355 -700
rect 15320 -750 15325 -725
rect 15350 -750 15355 -725
rect 15320 -770 15355 -750
rect 15380 -585 15415 -575
rect 15380 -610 15385 -585
rect 15410 -610 15415 -585
rect 15380 -630 15415 -610
rect 15380 -655 15385 -630
rect 15410 -655 15415 -630
rect 15380 -675 15415 -655
rect 15380 -700 15385 -675
rect 15410 -700 15415 -675
rect 15380 -725 15415 -700
rect 15380 -750 15385 -725
rect 15410 -750 15415 -725
rect 15380 -770 15415 -750
rect 15440 -585 15475 -575
rect 15440 -610 15445 -585
rect 15470 -610 15475 -585
rect 15440 -630 15475 -610
rect 15440 -655 15445 -630
rect 15470 -655 15475 -630
rect 15440 -675 15475 -655
rect 15440 -700 15445 -675
rect 15470 -700 15475 -675
rect 15440 -725 15475 -700
rect 15440 -750 15445 -725
rect 15470 -750 15475 -725
rect 15440 -770 15475 -750
rect 15500 -585 15535 -575
rect 15500 -610 15505 -585
rect 15530 -610 15535 -585
rect 15500 -630 15535 -610
rect 15500 -655 15505 -630
rect 15530 -655 15535 -630
rect 15500 -675 15535 -655
rect 15500 -700 15505 -675
rect 15530 -700 15535 -675
rect 15500 -725 15535 -700
rect 15500 -750 15505 -725
rect 15530 -750 15535 -725
rect 15500 -770 15535 -750
rect 15560 -585 15595 -575
rect 15560 -610 15565 -585
rect 15590 -610 15595 -585
rect 15560 -630 15595 -610
rect 15560 -655 15565 -630
rect 15590 -655 15595 -630
rect 15560 -675 15595 -655
rect 15560 -700 15565 -675
rect 15590 -700 15595 -675
rect 15560 -725 15595 -700
rect 15560 -750 15565 -725
rect 15590 -750 15595 -725
rect 15560 -770 15595 -750
rect 15620 -585 15655 -575
rect 15620 -610 15625 -585
rect 15650 -610 15655 -585
rect 15620 -630 15655 -610
rect 15620 -655 15625 -630
rect 15650 -655 15655 -630
rect 15620 -675 15655 -655
rect 15620 -700 15625 -675
rect 15650 -700 15655 -675
rect 15620 -725 15655 -700
rect 15620 -750 15625 -725
rect 15650 -750 15655 -725
rect 15620 -770 15655 -750
rect 15680 -585 15715 -575
rect 15680 -610 15685 -585
rect 15710 -610 15715 -585
rect 15680 -630 15715 -610
rect 15680 -655 15685 -630
rect 15710 -655 15715 -630
rect 15680 -675 15715 -655
rect 15680 -700 15685 -675
rect 15710 -700 15715 -675
rect 15680 -725 15715 -700
rect 15680 -750 15685 -725
rect 15710 -750 15715 -725
rect 15680 -770 15715 -750
rect 15740 -585 15775 -575
rect 15740 -610 15745 -585
rect 15770 -610 15775 -585
rect 15740 -630 15775 -610
rect 15740 -655 15745 -630
rect 15770 -655 15775 -630
rect 15740 -675 15775 -655
rect 15740 -700 15745 -675
rect 15770 -700 15775 -675
rect 15740 -725 15775 -700
rect 15740 -750 15745 -725
rect 15770 -750 15775 -725
rect 15740 -770 15775 -750
rect 15800 -585 15835 -575
rect 15800 -610 15805 -585
rect 15830 -610 15835 -585
rect 15800 -630 15835 -610
rect 15800 -655 15805 -630
rect 15830 -655 15835 -630
rect 15800 -675 15835 -655
rect 15800 -700 15805 -675
rect 15830 -700 15835 -675
rect 15800 -725 15835 -700
rect 15800 -750 15805 -725
rect 15830 -750 15835 -725
rect 15800 -770 15835 -750
rect 15860 -585 15895 -575
rect 15860 -610 15865 -585
rect 15890 -610 15895 -585
rect 15860 -630 15895 -610
rect 15860 -655 15865 -630
rect 15890 -655 15895 -630
rect 15860 -675 15895 -655
rect 15860 -700 15865 -675
rect 15890 -700 15895 -675
rect 15860 -725 15895 -700
rect 15860 -750 15865 -725
rect 15890 -750 15895 -725
rect 15860 -770 15895 -750
rect 15920 -585 15955 -575
rect 15920 -610 15925 -585
rect 15950 -610 15955 -585
rect 15920 -630 15955 -610
rect 15920 -655 15925 -630
rect 15950 -655 15955 -630
rect 15920 -675 15955 -655
rect 15920 -700 15925 -675
rect 15950 -700 15955 -675
rect 15920 -725 15955 -700
rect 15920 -750 15925 -725
rect 15950 -750 15955 -725
rect 15920 -770 15955 -750
rect 15980 -585 16015 -575
rect 15980 -610 15985 -585
rect 16010 -610 16015 -585
rect 15980 -630 16015 -610
rect 15980 -655 15985 -630
rect 16010 -655 16015 -630
rect 15980 -675 16015 -655
rect 15980 -700 15985 -675
rect 16010 -700 16015 -675
rect 15980 -725 16015 -700
rect 15980 -750 15985 -725
rect 16010 -750 16015 -725
rect 15980 -770 16015 -750
rect 16040 -585 16075 -575
rect 16040 -610 16045 -585
rect 16070 -610 16075 -585
rect 16040 -630 16075 -610
rect 16040 -655 16045 -630
rect 16070 -655 16075 -630
rect 16040 -675 16075 -655
rect 16040 -700 16045 -675
rect 16070 -700 16075 -675
rect 16040 -725 16075 -700
rect 16040 -750 16045 -725
rect 16070 -750 16075 -725
rect 16040 -770 16075 -750
rect 16100 -585 16135 -575
rect 16100 -610 16105 -585
rect 16130 -610 16135 -585
rect 16100 -630 16135 -610
rect 16100 -655 16105 -630
rect 16130 -655 16135 -630
rect 16100 -675 16135 -655
rect 16100 -700 16105 -675
rect 16130 -700 16135 -675
rect 16100 -725 16135 -700
rect 16100 -750 16105 -725
rect 16130 -750 16135 -725
rect 16100 -770 16135 -750
rect 16160 -585 16195 -575
rect 16160 -610 16165 -585
rect 16190 -610 16195 -585
rect 16160 -630 16195 -610
rect 16160 -655 16165 -630
rect 16190 -655 16195 -630
rect 16160 -675 16195 -655
rect 16160 -700 16165 -675
rect 16190 -700 16195 -675
rect 16160 -725 16195 -700
rect 16160 -750 16165 -725
rect 16190 -750 16195 -725
rect 16160 -770 16195 -750
rect 16220 -585 16255 -575
rect 16220 -610 16225 -585
rect 16250 -610 16255 -585
rect 16220 -630 16255 -610
rect 16220 -655 16225 -630
rect 16250 -655 16255 -630
rect 16220 -675 16255 -655
rect 16220 -700 16225 -675
rect 16250 -700 16255 -675
rect 16220 -725 16255 -700
rect 16220 -750 16225 -725
rect 16250 -750 16255 -725
rect 16220 -770 16255 -750
rect 16280 -585 16315 -575
rect 16280 -610 16285 -585
rect 16310 -610 16315 -585
rect 16280 -630 16315 -610
rect 16280 -655 16285 -630
rect 16310 -655 16315 -630
rect 16280 -675 16315 -655
rect 16280 -700 16285 -675
rect 16310 -700 16315 -675
rect 16280 -725 16315 -700
rect 16280 -750 16285 -725
rect 16310 -750 16315 -725
rect 16280 -770 16315 -750
rect 16340 -585 16375 -575
rect 16340 -610 16345 -585
rect 16370 -610 16375 -585
rect 16340 -630 16375 -610
rect 16340 -655 16345 -630
rect 16370 -655 16375 -630
rect 16340 -675 16375 -655
rect 16340 -700 16345 -675
rect 16370 -700 16375 -675
rect 16340 -725 16375 -700
rect 16340 -750 16345 -725
rect 16370 -750 16375 -725
rect 16340 -770 16375 -750
rect 16400 -585 16435 -575
rect 16400 -610 16405 -585
rect 16430 -610 16435 -585
rect 16400 -630 16435 -610
rect 16400 -655 16405 -630
rect 16430 -655 16435 -630
rect 16400 -675 16435 -655
rect 16400 -700 16405 -675
rect 16430 -700 16435 -675
rect 16400 -725 16435 -700
rect 16400 -750 16405 -725
rect 16430 -750 16435 -725
rect 16400 -770 16435 -750
rect 16460 -585 16495 -575
rect 16460 -610 16465 -585
rect 16490 -610 16495 -585
rect 16460 -630 16495 -610
rect 16460 -655 16465 -630
rect 16490 -655 16495 -630
rect 16460 -675 16495 -655
rect 16460 -700 16465 -675
rect 16490 -700 16495 -675
rect 16460 -725 16495 -700
rect 16460 -750 16465 -725
rect 16490 -750 16495 -725
rect 16460 -770 16495 -750
rect 16520 -585 16555 -575
rect 16520 -610 16525 -585
rect 16550 -610 16555 -585
rect 16520 -630 16555 -610
rect 16520 -655 16525 -630
rect 16550 -655 16555 -630
rect 16520 -675 16555 -655
rect 16520 -700 16525 -675
rect 16550 -700 16555 -675
rect 16520 -725 16555 -700
rect 16520 -750 16525 -725
rect 16550 -750 16555 -725
rect 16520 -770 16555 -750
rect 16580 -585 16615 -575
rect 16580 -610 16585 -585
rect 16610 -610 16615 -585
rect 16580 -630 16615 -610
rect 16580 -655 16585 -630
rect 16610 -655 16615 -630
rect 16580 -675 16615 -655
rect 16580 -700 16585 -675
rect 16610 -700 16615 -675
rect 16580 -725 16615 -700
rect 16580 -750 16585 -725
rect 16610 -750 16615 -725
rect 16580 -770 16615 -750
rect 16640 -585 16675 -575
rect 16640 -610 16645 -585
rect 16670 -610 16675 -585
rect 16640 -630 16675 -610
rect 16640 -655 16645 -630
rect 16670 -655 16675 -630
rect 16640 -675 16675 -655
rect 16640 -700 16645 -675
rect 16670 -700 16675 -675
rect 16640 -725 16675 -700
rect 16640 -750 16645 -725
rect 16670 -750 16675 -725
rect 16640 -770 16675 -750
rect 16700 -585 16735 -575
rect 16700 -610 16705 -585
rect 16730 -610 16735 -585
rect 16700 -630 16735 -610
rect 16700 -655 16705 -630
rect 16730 -655 16735 -630
rect 16700 -675 16735 -655
rect 16700 -700 16705 -675
rect 16730 -700 16735 -675
rect 16700 -725 16735 -700
rect 16700 -750 16705 -725
rect 16730 -750 16735 -725
rect 16700 -770 16735 -750
rect 16760 -585 16795 -575
rect 16760 -610 16765 -585
rect 16790 -610 16795 -585
rect 16760 -630 16795 -610
rect 16760 -655 16765 -630
rect 16790 -655 16795 -630
rect 16760 -675 16795 -655
rect 16760 -700 16765 -675
rect 16790 -700 16795 -675
rect 16760 -725 16795 -700
rect 16760 -750 16765 -725
rect 16790 -750 16795 -725
rect 16760 -770 16795 -750
rect 16820 -585 16855 -575
rect 16820 -610 16825 -585
rect 16850 -610 16855 -585
rect 16820 -630 16855 -610
rect 16820 -655 16825 -630
rect 16850 -655 16855 -630
rect 16820 -675 16855 -655
rect 16820 -700 16825 -675
rect 16850 -700 16855 -675
rect 16820 -725 16855 -700
rect 16820 -750 16825 -725
rect 16850 -750 16855 -725
rect 16820 -770 16855 -750
rect 16880 -585 16915 -575
rect 16880 -610 16885 -585
rect 16910 -610 16915 -585
rect 16880 -630 16915 -610
rect 16880 -655 16885 -630
rect 16910 -655 16915 -630
rect 16880 -675 16915 -655
rect 16880 -700 16885 -675
rect 16910 -700 16915 -675
rect 16880 -725 16915 -700
rect 16880 -750 16885 -725
rect 16910 -750 16915 -725
rect 16880 -770 16915 -750
rect 16940 -585 16975 -575
rect 16940 -610 16945 -585
rect 16970 -610 16975 -585
rect 16940 -630 16975 -610
rect 16940 -655 16945 -630
rect 16970 -655 16975 -630
rect 16940 -675 16975 -655
rect 16940 -700 16945 -675
rect 16970 -700 16975 -675
rect 16940 -725 16975 -700
rect 16940 -750 16945 -725
rect 16970 -750 16975 -725
rect 16940 -770 16975 -750
rect 17000 -585 17035 -575
rect 17000 -610 17005 -585
rect 17030 -610 17035 -585
rect 17000 -630 17035 -610
rect 17000 -655 17005 -630
rect 17030 -655 17035 -630
rect 17000 -675 17035 -655
rect 17000 -700 17005 -675
rect 17030 -700 17035 -675
rect 17000 -725 17035 -700
rect 17000 -750 17005 -725
rect 17030 -750 17035 -725
rect 17000 -770 17035 -750
rect 17060 -585 17095 -575
rect 17060 -610 17065 -585
rect 17090 -610 17095 -585
rect 17060 -630 17095 -610
rect 17060 -655 17065 -630
rect 17090 -655 17095 -630
rect 17060 -675 17095 -655
rect 17060 -700 17065 -675
rect 17090 -700 17095 -675
rect 17060 -725 17095 -700
rect 17060 -750 17065 -725
rect 17090 -750 17095 -725
rect 17060 -770 17095 -750
rect 17120 -585 17155 -575
rect 17120 -610 17125 -585
rect 17150 -610 17155 -585
rect 17120 -630 17155 -610
rect 17120 -655 17125 -630
rect 17150 -655 17155 -630
rect 17120 -675 17155 -655
rect 17120 -700 17125 -675
rect 17150 -700 17155 -675
rect 17120 -725 17155 -700
rect 17120 -750 17125 -725
rect 17150 -750 17155 -725
rect 17120 -770 17155 -750
rect 17180 -585 17215 -575
rect 17180 -610 17185 -585
rect 17210 -610 17215 -585
rect 17180 -630 17215 -610
rect 17180 -655 17185 -630
rect 17210 -655 17215 -630
rect 17180 -675 17215 -655
rect 17180 -700 17185 -675
rect 17210 -700 17215 -675
rect 17180 -725 17215 -700
rect 17180 -750 17185 -725
rect 17210 -750 17215 -725
rect 17180 -770 17215 -750
rect 17240 -585 17275 -575
rect 17240 -610 17245 -585
rect 17270 -610 17275 -585
rect 17240 -630 17275 -610
rect 17240 -655 17245 -630
rect 17270 -655 17275 -630
rect 17240 -675 17275 -655
rect 17240 -700 17245 -675
rect 17270 -700 17275 -675
rect 17240 -725 17275 -700
rect 17240 -750 17245 -725
rect 17270 -750 17275 -725
rect 17240 -770 17275 -750
rect 17300 -585 17335 -575
rect 17300 -610 17305 -585
rect 17330 -610 17335 -585
rect 17300 -630 17335 -610
rect 17300 -655 17305 -630
rect 17330 -655 17335 -630
rect 17300 -675 17335 -655
rect 17300 -700 17305 -675
rect 17330 -700 17335 -675
rect 17300 -725 17335 -700
rect 17300 -750 17305 -725
rect 17330 -750 17335 -725
rect 17300 -770 17335 -750
rect 17360 -585 17395 -575
rect 17360 -610 17365 -585
rect 17390 -610 17395 -585
rect 17360 -630 17395 -610
rect 17360 -655 17365 -630
rect 17390 -655 17395 -630
rect 17360 -675 17395 -655
rect 17360 -700 17365 -675
rect 17390 -700 17395 -675
rect 17360 -725 17395 -700
rect 17360 -750 17365 -725
rect 17390 -750 17395 -725
rect 17360 -770 17395 -750
rect 17420 -585 17455 -575
rect 17420 -610 17425 -585
rect 17450 -610 17455 -585
rect 17420 -630 17455 -610
rect 17420 -655 17425 -630
rect 17450 -655 17455 -630
rect 17420 -675 17455 -655
rect 17420 -700 17425 -675
rect 17450 -700 17455 -675
rect 17420 -725 17455 -700
rect 17420 -750 17425 -725
rect 17450 -750 17455 -725
rect 17420 -770 17455 -750
rect 17480 -585 17515 -575
rect 17480 -610 17485 -585
rect 17510 -610 17515 -585
rect 17480 -630 17515 -610
rect 17480 -655 17485 -630
rect 17510 -655 17515 -630
rect 17480 -675 17515 -655
rect 17480 -700 17485 -675
rect 17510 -700 17515 -675
rect 17480 -725 17515 -700
rect 17480 -750 17485 -725
rect 17510 -750 17515 -725
rect 17480 -770 17515 -750
rect 17540 -585 17575 -575
rect 17540 -610 17545 -585
rect 17570 -610 17575 -585
rect 17540 -630 17575 -610
rect 17540 -655 17545 -630
rect 17570 -655 17575 -630
rect 17540 -675 17575 -655
rect 17540 -700 17545 -675
rect 17570 -700 17575 -675
rect 17540 -725 17575 -700
rect 17540 -750 17545 -725
rect 17570 -750 17575 -725
rect 17540 -770 17575 -750
rect 17600 -585 17635 -575
rect 17600 -610 17605 -585
rect 17630 -610 17635 -585
rect 17600 -630 17635 -610
rect 17600 -655 17605 -630
rect 17630 -655 17635 -630
rect 17600 -675 17635 -655
rect 17600 -700 17605 -675
rect 17630 -700 17635 -675
rect 17600 -725 17635 -700
rect 17600 -750 17605 -725
rect 17630 -750 17635 -725
rect 17600 -770 17635 -750
rect 17660 -585 17695 -575
rect 17660 -610 17665 -585
rect 17690 -610 17695 -585
rect 17660 -630 17695 -610
rect 17660 -655 17665 -630
rect 17690 -655 17695 -630
rect 17660 -675 17695 -655
rect 17660 -700 17665 -675
rect 17690 -700 17695 -675
rect 17660 -725 17695 -700
rect 17660 -750 17665 -725
rect 17690 -750 17695 -725
rect 17660 -770 17695 -750
rect 17720 -585 17755 -575
rect 17720 -610 17725 -585
rect 17750 -610 17755 -585
rect 17720 -630 17755 -610
rect 17720 -655 17725 -630
rect 17750 -655 17755 -630
rect 17720 -675 17755 -655
rect 17720 -700 17725 -675
rect 17750 -700 17755 -675
rect 17720 -725 17755 -700
rect 17720 -750 17725 -725
rect 17750 -750 17755 -725
rect 17720 -770 17755 -750
rect 17780 -585 17815 -575
rect 17780 -610 17785 -585
rect 17810 -610 17815 -585
rect 17780 -630 17815 -610
rect 17780 -655 17785 -630
rect 17810 -655 17815 -630
rect 17780 -675 17815 -655
rect 17780 -700 17785 -675
rect 17810 -700 17815 -675
rect 17780 -725 17815 -700
rect 17780 -750 17785 -725
rect 17810 -750 17815 -725
rect 17780 -770 17815 -750
rect 17840 -585 17875 -575
rect 17840 -610 17845 -585
rect 17870 -610 17875 -585
rect 17840 -630 17875 -610
rect 17840 -655 17845 -630
rect 17870 -655 17875 -630
rect 17840 -675 17875 -655
rect 17840 -700 17845 -675
rect 17870 -700 17875 -675
rect 17840 -725 17875 -700
rect 17840 -750 17845 -725
rect 17870 -750 17875 -725
rect 17840 -770 17875 -750
rect 17900 -585 17935 -575
rect 17900 -610 17905 -585
rect 17930 -610 17935 -585
rect 17900 -630 17935 -610
rect 17900 -655 17905 -630
rect 17930 -655 17935 -630
rect 17900 -675 17935 -655
rect 17900 -700 17905 -675
rect 17930 -700 17935 -675
rect 17900 -725 17935 -700
rect 17900 -750 17905 -725
rect 17930 -750 17935 -725
rect 17900 -770 17935 -750
rect 17960 -585 17995 -575
rect 17960 -610 17965 -585
rect 17990 -610 17995 -585
rect 17960 -630 17995 -610
rect 17960 -655 17965 -630
rect 17990 -655 17995 -630
rect 17960 -675 17995 -655
rect 17960 -700 17965 -675
rect 17990 -700 17995 -675
rect 17960 -725 17995 -700
rect 17960 -750 17965 -725
rect 17990 -750 17995 -725
rect 17960 -770 17995 -750
rect 18020 -585 18055 -575
rect 18020 -610 18025 -585
rect 18050 -610 18055 -585
rect 18020 -630 18055 -610
rect 18020 -655 18025 -630
rect 18050 -655 18055 -630
rect 18020 -675 18055 -655
rect 18020 -700 18025 -675
rect 18050 -700 18055 -675
rect 18020 -725 18055 -700
rect 18020 -750 18025 -725
rect 18050 -750 18055 -725
rect 18020 -770 18055 -750
rect 18080 -585 18115 -575
rect 18080 -610 18085 -585
rect 18110 -610 18115 -585
rect 18080 -630 18115 -610
rect 18080 -655 18085 -630
rect 18110 -655 18115 -630
rect 18080 -675 18115 -655
rect 18080 -700 18085 -675
rect 18110 -700 18115 -675
rect 18080 -725 18115 -700
rect 18080 -750 18085 -725
rect 18110 -750 18115 -725
rect 18080 -770 18115 -750
rect 18140 -585 18175 -575
rect 18140 -610 18145 -585
rect 18170 -610 18175 -585
rect 18140 -630 18175 -610
rect 18140 -655 18145 -630
rect 18170 -655 18175 -630
rect 18140 -675 18175 -655
rect 18140 -700 18145 -675
rect 18170 -700 18175 -675
rect 18140 -725 18175 -700
rect 18140 -750 18145 -725
rect 18170 -750 18175 -725
rect 18140 -770 18175 -750
rect 18200 -585 18235 -575
rect 18200 -610 18205 -585
rect 18230 -610 18235 -585
rect 18200 -630 18235 -610
rect 18200 -655 18205 -630
rect 18230 -655 18235 -630
rect 18200 -675 18235 -655
rect 18200 -700 18205 -675
rect 18230 -700 18235 -675
rect 18200 -725 18235 -700
rect 18200 -750 18205 -725
rect 18230 -750 18235 -725
rect 18200 -770 18235 -750
rect 18260 -585 18295 -575
rect 18260 -610 18265 -585
rect 18290 -610 18295 -585
rect 18260 -630 18295 -610
rect 18260 -655 18265 -630
rect 18290 -655 18295 -630
rect 18260 -675 18295 -655
rect 18260 -700 18265 -675
rect 18290 -700 18295 -675
rect 18260 -725 18295 -700
rect 18260 -750 18265 -725
rect 18290 -750 18295 -725
rect 18260 -770 18295 -750
rect 18320 -585 18355 -575
rect 18320 -610 18325 -585
rect 18350 -610 18355 -585
rect 18320 -630 18355 -610
rect 18320 -655 18325 -630
rect 18350 -655 18355 -630
rect 18320 -675 18355 -655
rect 18320 -700 18325 -675
rect 18350 -700 18355 -675
rect 18320 -725 18355 -700
rect 18320 -750 18325 -725
rect 18350 -750 18355 -725
rect 18320 -770 18355 -750
rect 18380 -585 18415 -575
rect 18380 -610 18385 -585
rect 18410 -610 18415 -585
rect 18380 -630 18415 -610
rect 18380 -655 18385 -630
rect 18410 -655 18415 -630
rect 18380 -675 18415 -655
rect 18380 -700 18385 -675
rect 18410 -700 18415 -675
rect 18380 -725 18415 -700
rect 18380 -750 18385 -725
rect 18410 -750 18415 -725
rect 18380 -770 18415 -750
rect 18440 -585 18475 -575
rect 18440 -610 18445 -585
rect 18470 -610 18475 -585
rect 18440 -630 18475 -610
rect 18440 -655 18445 -630
rect 18470 -655 18475 -630
rect 18440 -675 18475 -655
rect 18440 -700 18445 -675
rect 18470 -700 18475 -675
rect 18440 -725 18475 -700
rect 18440 -750 18445 -725
rect 18470 -750 18475 -725
rect 18440 -770 18475 -750
rect 18500 -585 18535 -575
rect 18500 -610 18505 -585
rect 18530 -610 18535 -585
rect 18500 -630 18535 -610
rect 18500 -655 18505 -630
rect 18530 -655 18535 -630
rect 18500 -675 18535 -655
rect 18500 -700 18505 -675
rect 18530 -700 18535 -675
rect 18500 -725 18535 -700
rect 18500 -750 18505 -725
rect 18530 -750 18535 -725
rect 18500 -770 18535 -750
rect 18560 -585 18595 -575
rect 18560 -610 18565 -585
rect 18590 -610 18595 -585
rect 18560 -630 18595 -610
rect 18560 -655 18565 -630
rect 18590 -655 18595 -630
rect 18560 -675 18595 -655
rect 18560 -700 18565 -675
rect 18590 -700 18595 -675
rect 18560 -725 18595 -700
rect 18560 -750 18565 -725
rect 18590 -750 18595 -725
rect 18560 -770 18595 -750
rect 18620 -585 18655 -575
rect 18620 -610 18625 -585
rect 18650 -610 18655 -585
rect 18620 -630 18655 -610
rect 18620 -655 18625 -630
rect 18650 -655 18655 -630
rect 18620 -675 18655 -655
rect 18620 -700 18625 -675
rect 18650 -700 18655 -675
rect 18620 -725 18655 -700
rect 18620 -750 18625 -725
rect 18650 -750 18655 -725
rect 18620 -770 18655 -750
rect 18680 -585 18715 -575
rect 18680 -610 18685 -585
rect 18710 -610 18715 -585
rect 18680 -630 18715 -610
rect 18680 -655 18685 -630
rect 18710 -655 18715 -630
rect 18680 -675 18715 -655
rect 18680 -700 18685 -675
rect 18710 -700 18715 -675
rect 18680 -725 18715 -700
rect 18680 -750 18685 -725
rect 18710 -750 18715 -725
rect 18680 -770 18715 -750
rect 18740 -585 18775 -575
rect 18740 -610 18745 -585
rect 18770 -610 18775 -585
rect 18740 -630 18775 -610
rect 18740 -655 18745 -630
rect 18770 -655 18775 -630
rect 18740 -675 18775 -655
rect 18740 -700 18745 -675
rect 18770 -700 18775 -675
rect 18740 -725 18775 -700
rect 18740 -750 18745 -725
rect 18770 -750 18775 -725
rect 18740 -770 18775 -750
rect 18800 -585 18835 -575
rect 18800 -610 18805 -585
rect 18830 -610 18835 -585
rect 18800 -630 18835 -610
rect 18800 -655 18805 -630
rect 18830 -655 18835 -630
rect 18800 -675 18835 -655
rect 18800 -700 18805 -675
rect 18830 -700 18835 -675
rect 18800 -725 18835 -700
rect 18800 -750 18805 -725
rect 18830 -750 18835 -725
rect 18800 -770 18835 -750
rect 18860 -585 18895 -575
rect 18860 -610 18865 -585
rect 18890 -610 18895 -585
rect 18860 -630 18895 -610
rect 18860 -655 18865 -630
rect 18890 -655 18895 -630
rect 18860 -675 18895 -655
rect 18860 -700 18865 -675
rect 18890 -700 18895 -675
rect 18860 -725 18895 -700
rect 18860 -750 18865 -725
rect 18890 -750 18895 -725
rect 18860 -770 18895 -750
rect 18920 -585 18955 -575
rect 18920 -610 18925 -585
rect 18950 -610 18955 -585
rect 18920 -630 18955 -610
rect 18920 -655 18925 -630
rect 18950 -655 18955 -630
rect 18920 -675 18955 -655
rect 18920 -700 18925 -675
rect 18950 -700 18955 -675
rect 18920 -725 18955 -700
rect 18920 -750 18925 -725
rect 18950 -750 18955 -725
rect 18920 -770 18955 -750
rect 18980 -585 19015 -575
rect 18980 -610 18985 -585
rect 19010 -610 19015 -585
rect 18980 -630 19015 -610
rect 18980 -655 18985 -630
rect 19010 -655 19015 -630
rect 18980 -675 19015 -655
rect 18980 -700 18985 -675
rect 19010 -700 19015 -675
rect 18980 -725 19015 -700
rect 18980 -750 18985 -725
rect 19010 -750 19015 -725
rect 18980 -770 19015 -750
rect 19040 -585 19075 -575
rect 19040 -610 19045 -585
rect 19070 -610 19075 -585
rect 19040 -630 19075 -610
rect 19040 -655 19045 -630
rect 19070 -655 19075 -630
rect 19040 -675 19075 -655
rect 19040 -700 19045 -675
rect 19070 -700 19075 -675
rect 19040 -725 19075 -700
rect 19040 -750 19045 -725
rect 19070 -750 19075 -725
rect 19040 -770 19075 -750
rect 19100 -585 19135 -575
rect 19100 -610 19105 -585
rect 19130 -610 19135 -585
rect 19100 -630 19135 -610
rect 19100 -655 19105 -630
rect 19130 -655 19135 -630
rect 19100 -675 19135 -655
rect 19100 -700 19105 -675
rect 19130 -700 19135 -675
rect 19100 -725 19135 -700
rect 19100 -750 19105 -725
rect 19130 -750 19135 -725
rect 19100 -770 19135 -750
rect 19160 -585 19195 -575
rect 19160 -610 19165 -585
rect 19190 -610 19195 -585
rect 19160 -630 19195 -610
rect 19160 -655 19165 -630
rect 19190 -655 19195 -630
rect 19160 -675 19195 -655
rect 19160 -700 19165 -675
rect 19190 -700 19195 -675
rect 19160 -725 19195 -700
rect 19160 -750 19165 -725
rect 19190 -750 19195 -725
rect 19160 -770 19195 -750
rect 19220 -585 19255 -575
rect 19220 -610 19225 -585
rect 19250 -610 19255 -585
rect 19220 -630 19255 -610
rect 19220 -655 19225 -630
rect 19250 -655 19255 -630
rect 19220 -675 19255 -655
rect 19220 -700 19225 -675
rect 19250 -700 19255 -675
rect 19220 -725 19255 -700
rect 19220 -750 19225 -725
rect 19250 -750 19255 -725
rect 19220 -770 19255 -750
rect 19280 -585 19315 -575
rect 19280 -610 19285 -585
rect 19310 -610 19315 -585
rect 19280 -630 19315 -610
rect 19280 -655 19285 -630
rect 19310 -655 19315 -630
rect 19280 -675 19315 -655
rect 19280 -700 19285 -675
rect 19310 -700 19315 -675
rect 19280 -725 19315 -700
rect 19280 -750 19285 -725
rect 19310 -750 19315 -725
rect 19280 -770 19315 -750
rect 19340 -585 19375 -575
rect 19340 -610 19345 -585
rect 19370 -610 19375 -585
rect 19340 -630 19375 -610
rect 19340 -655 19345 -630
rect 19370 -655 19375 -630
rect 19340 -675 19375 -655
rect 19340 -700 19345 -675
rect 19370 -700 19375 -675
rect 19340 -725 19375 -700
rect 19340 -750 19345 -725
rect 19370 -750 19375 -725
rect 19340 -770 19375 -750
rect 19400 -585 19435 -575
rect 19400 -610 19405 -585
rect 19430 -610 19435 -585
rect 19400 -630 19435 -610
rect 19400 -655 19405 -630
rect 19430 -655 19435 -630
rect 19400 -675 19435 -655
rect 19400 -700 19405 -675
rect 19430 -700 19435 -675
rect 19400 -725 19435 -700
rect 19400 -750 19405 -725
rect 19430 -750 19435 -725
rect 19400 -770 19435 -750
rect 19460 -585 19495 -575
rect 19460 -610 19465 -585
rect 19490 -610 19495 -585
rect 19460 -630 19495 -610
rect 19460 -655 19465 -630
rect 19490 -655 19495 -630
rect 19460 -675 19495 -655
rect 19460 -700 19465 -675
rect 19490 -700 19495 -675
rect 19460 -725 19495 -700
rect 19460 -750 19465 -725
rect 19490 -750 19495 -725
rect 19460 -770 19495 -750
rect 19520 -585 19555 -575
rect 19520 -610 19525 -585
rect 19550 -610 19555 -585
rect 19520 -630 19555 -610
rect 19520 -655 19525 -630
rect 19550 -655 19555 -630
rect 19520 -675 19555 -655
rect 19520 -700 19525 -675
rect 19550 -700 19555 -675
rect 19520 -725 19555 -700
rect 19520 -750 19525 -725
rect 19550 -750 19555 -725
rect 19520 -770 19555 -750
rect 19580 -585 19615 -575
rect 19580 -610 19585 -585
rect 19610 -610 19615 -585
rect 19580 -630 19615 -610
rect 19580 -655 19585 -630
rect 19610 -655 19615 -630
rect 19580 -675 19615 -655
rect 19580 -700 19585 -675
rect 19610 -700 19615 -675
rect 19580 -725 19615 -700
rect 19580 -750 19585 -725
rect 19610 -750 19615 -725
rect 19580 -770 19615 -750
rect 19640 -585 19675 -575
rect 19640 -610 19645 -585
rect 19670 -610 19675 -585
rect 19640 -630 19675 -610
rect 19640 -655 19645 -630
rect 19670 -655 19675 -630
rect 19640 -675 19675 -655
rect 19640 -700 19645 -675
rect 19670 -700 19675 -675
rect 19640 -725 19675 -700
rect 19640 -750 19645 -725
rect 19670 -750 19675 -725
rect 19640 -770 19675 -750
rect 19700 -585 19735 -575
rect 19700 -610 19705 -585
rect 19730 -610 19735 -585
rect 19700 -630 19735 -610
rect 19700 -655 19705 -630
rect 19730 -655 19735 -630
rect 19700 -675 19735 -655
rect 19700 -700 19705 -675
rect 19730 -700 19735 -675
rect 19700 -725 19735 -700
rect 19700 -750 19705 -725
rect 19730 -750 19735 -725
rect 19700 -770 19735 -750
rect 19760 -585 19795 -575
rect 19760 -610 19765 -585
rect 19790 -610 19795 -585
rect 19760 -630 19795 -610
rect 19760 -655 19765 -630
rect 19790 -655 19795 -630
rect 19760 -675 19795 -655
rect 19760 -700 19765 -675
rect 19790 -700 19795 -675
rect 19760 -725 19795 -700
rect 19760 -750 19765 -725
rect 19790 -750 19795 -725
rect 19760 -770 19795 -750
rect 19820 -585 19855 -575
rect 19820 -610 19825 -585
rect 19850 -610 19855 -585
rect 19820 -630 19855 -610
rect 19820 -655 19825 -630
rect 19850 -655 19855 -630
rect 19820 -675 19855 -655
rect 19820 -700 19825 -675
rect 19850 -700 19855 -675
rect 19820 -725 19855 -700
rect 19820 -750 19825 -725
rect 19850 -750 19855 -725
rect 19820 -770 19855 -750
rect 19880 -585 19915 -575
rect 19880 -610 19885 -585
rect 19910 -610 19915 -585
rect 19880 -630 19915 -610
rect 19880 -655 19885 -630
rect 19910 -655 19915 -630
rect 19880 -675 19915 -655
rect 19880 -700 19885 -675
rect 19910 -700 19915 -675
rect 19880 -725 19915 -700
rect 19880 -750 19885 -725
rect 19910 -750 19915 -725
rect 19880 -770 19915 -750
rect 19940 -585 19975 -575
rect 19940 -610 19945 -585
rect 19970 -610 19975 -585
rect 19940 -630 19975 -610
rect 19940 -655 19945 -630
rect 19970 -655 19975 -630
rect 19940 -675 19975 -655
rect 19940 -700 19945 -675
rect 19970 -700 19975 -675
rect 19940 -725 19975 -700
rect 19940 -750 19945 -725
rect 19970 -750 19975 -725
rect 19940 -770 19975 -750
rect 20000 -585 20035 -575
rect 20000 -610 20005 -585
rect 20030 -610 20035 -585
rect 20000 -630 20035 -610
rect 20000 -655 20005 -630
rect 20030 -655 20035 -630
rect 20000 -675 20035 -655
rect 20000 -700 20005 -675
rect 20030 -700 20035 -675
rect 20000 -725 20035 -700
rect 20000 -750 20005 -725
rect 20030 -750 20035 -725
rect 20000 -770 20035 -750
rect 20060 -585 20095 -575
rect 20060 -610 20065 -585
rect 20090 -610 20095 -585
rect 20060 -630 20095 -610
rect 20060 -655 20065 -630
rect 20090 -655 20095 -630
rect 20060 -675 20095 -655
rect 20060 -700 20065 -675
rect 20090 -700 20095 -675
rect 20060 -725 20095 -700
rect 20060 -750 20065 -725
rect 20090 -750 20095 -725
rect 20060 -770 20095 -750
rect 20120 -585 20155 -575
rect 20120 -610 20125 -585
rect 20150 -610 20155 -585
rect 20120 -630 20155 -610
rect 20120 -655 20125 -630
rect 20150 -655 20155 -630
rect 20120 -675 20155 -655
rect 20120 -700 20125 -675
rect 20150 -700 20155 -675
rect 20120 -725 20155 -700
rect 20120 -750 20125 -725
rect 20150 -750 20155 -725
rect 20120 -770 20155 -750
rect 20180 -585 20215 -575
rect 20180 -610 20185 -585
rect 20210 -610 20215 -585
rect 20180 -630 20215 -610
rect 20180 -655 20185 -630
rect 20210 -655 20215 -630
rect 20180 -675 20215 -655
rect 20180 -700 20185 -675
rect 20210 -700 20215 -675
rect 20180 -725 20215 -700
rect 20180 -750 20185 -725
rect 20210 -750 20215 -725
rect 20180 -770 20215 -750
rect 20240 -585 20275 -575
rect 20240 -610 20245 -585
rect 20270 -610 20275 -585
rect 20240 -630 20275 -610
rect 20240 -655 20245 -630
rect 20270 -655 20275 -630
rect 20240 -675 20275 -655
rect 20240 -700 20245 -675
rect 20270 -700 20275 -675
rect 20240 -725 20275 -700
rect 20240 -750 20245 -725
rect 20270 -750 20275 -725
rect 20240 -770 20275 -750
rect 20300 -585 20335 -575
rect 20300 -610 20305 -585
rect 20330 -610 20335 -585
rect 20300 -630 20335 -610
rect 20300 -655 20305 -630
rect 20330 -655 20335 -630
rect 20300 -675 20335 -655
rect 20300 -700 20305 -675
rect 20330 -700 20335 -675
rect 20300 -725 20335 -700
rect 20300 -750 20305 -725
rect 20330 -750 20335 -725
rect 20300 -770 20335 -750
rect 20360 -585 20395 -575
rect 20360 -610 20365 -585
rect 20390 -610 20395 -585
rect 20360 -630 20395 -610
rect 20360 -655 20365 -630
rect 20390 -655 20395 -630
rect 20360 -675 20395 -655
rect 20360 -700 20365 -675
rect 20390 -700 20395 -675
rect 20360 -725 20395 -700
rect 20360 -750 20365 -725
rect 20390 -750 20395 -725
rect 20360 -770 20395 -750
rect 20420 -585 20455 -575
rect 20420 -610 20425 -585
rect 20450 -610 20455 -585
rect 20420 -630 20455 -610
rect 20420 -655 20425 -630
rect 20450 -655 20455 -630
rect 20420 -675 20455 -655
rect 20420 -700 20425 -675
rect 20450 -700 20455 -675
rect 20420 -725 20455 -700
rect 20420 -750 20425 -725
rect 20450 -750 20455 -725
rect 20420 -770 20455 -750
rect 20480 -585 20515 -575
rect 20480 -610 20485 -585
rect 20510 -610 20515 -585
rect 20480 -630 20515 -610
rect 20480 -655 20485 -630
rect 20510 -655 20515 -630
rect 20480 -675 20515 -655
rect 20480 -700 20485 -675
rect 20510 -700 20515 -675
rect 20480 -725 20515 -700
rect 20480 -750 20485 -725
rect 20510 -750 20515 -725
rect 20480 -770 20515 -750
rect 20540 -585 20575 -575
rect 20540 -610 20545 -585
rect 20570 -610 20575 -585
rect 20540 -630 20575 -610
rect 20540 -655 20545 -630
rect 20570 -655 20575 -630
rect 20540 -675 20575 -655
rect 20540 -700 20545 -675
rect 20570 -700 20575 -675
rect 20540 -725 20575 -700
rect 20540 -750 20545 -725
rect 20570 -750 20575 -725
rect 20540 -770 20575 -750
rect 20600 -585 20635 -575
rect 20600 -610 20605 -585
rect 20630 -610 20635 -585
rect 20600 -630 20635 -610
rect 20600 -655 20605 -630
rect 20630 -655 20635 -630
rect 20600 -675 20635 -655
rect 20600 -700 20605 -675
rect 20630 -700 20635 -675
rect 20600 -725 20635 -700
rect 20600 -750 20605 -725
rect 20630 -750 20635 -725
rect 20600 -770 20635 -750
rect 20660 -585 20695 -575
rect 20660 -610 20665 -585
rect 20690 -610 20695 -585
rect 20660 -630 20695 -610
rect 20660 -655 20665 -630
rect 20690 -655 20695 -630
rect 20660 -675 20695 -655
rect 20660 -700 20665 -675
rect 20690 -700 20695 -675
rect 20660 -725 20695 -700
rect 20660 -750 20665 -725
rect 20690 -750 20695 -725
rect 20660 -770 20695 -750
rect 20720 -585 20755 -575
rect 20720 -610 20725 -585
rect 20750 -610 20755 -585
rect 20720 -630 20755 -610
rect 20720 -655 20725 -630
rect 20750 -655 20755 -630
rect 20720 -675 20755 -655
rect 20720 -700 20725 -675
rect 20750 -700 20755 -675
rect 20720 -725 20755 -700
rect 20720 -750 20725 -725
rect 20750 -750 20755 -725
rect 20720 -770 20755 -750
rect 20780 -585 20815 -575
rect 20780 -610 20785 -585
rect 20810 -610 20815 -585
rect 20780 -630 20815 -610
rect 20780 -655 20785 -630
rect 20810 -655 20815 -630
rect 20780 -675 20815 -655
rect 20780 -700 20785 -675
rect 20810 -700 20815 -675
rect 20780 -725 20815 -700
rect 20780 -750 20785 -725
rect 20810 -750 20815 -725
rect 20780 -770 20815 -750
rect 20840 -585 20875 -575
rect 20840 -610 20845 -585
rect 20870 -610 20875 -585
rect 20840 -630 20875 -610
rect 20840 -655 20845 -630
rect 20870 -655 20875 -630
rect 20840 -675 20875 -655
rect 20840 -700 20845 -675
rect 20870 -700 20875 -675
rect 20840 -725 20875 -700
rect 20840 -750 20845 -725
rect 20870 -750 20875 -725
rect 20840 -770 20875 -750
rect 20900 -585 20935 -575
rect 20900 -610 20905 -585
rect 20930 -610 20935 -585
rect 20900 -630 20935 -610
rect 20900 -655 20905 -630
rect 20930 -655 20935 -630
rect 20900 -675 20935 -655
rect 20900 -700 20905 -675
rect 20930 -700 20935 -675
rect 20900 -725 20935 -700
rect 20900 -750 20905 -725
rect 20930 -750 20935 -725
rect 20900 -770 20935 -750
rect 20960 -585 20995 -575
rect 20960 -610 20965 -585
rect 20990 -610 20995 -585
rect 20960 -630 20995 -610
rect 20960 -655 20965 -630
rect 20990 -655 20995 -630
rect 20960 -675 20995 -655
rect 20960 -700 20965 -675
rect 20990 -700 20995 -675
rect 20960 -725 20995 -700
rect 20960 -750 20965 -725
rect 20990 -750 20995 -725
rect 20960 -770 20995 -750
rect 21020 -585 21055 -575
rect 21020 -610 21025 -585
rect 21050 -610 21055 -585
rect 21020 -630 21055 -610
rect 21020 -655 21025 -630
rect 21050 -655 21055 -630
rect 21020 -675 21055 -655
rect 21020 -700 21025 -675
rect 21050 -700 21055 -675
rect 21020 -725 21055 -700
rect 21020 -750 21025 -725
rect 21050 -750 21055 -725
rect 21020 -770 21055 -750
rect 21080 -585 21115 -575
rect 21080 -610 21085 -585
rect 21110 -610 21115 -585
rect 21080 -630 21115 -610
rect 21080 -655 21085 -630
rect 21110 -655 21115 -630
rect 21080 -675 21115 -655
rect 21080 -700 21085 -675
rect 21110 -700 21115 -675
rect 21080 -725 21115 -700
rect 21080 -750 21085 -725
rect 21110 -750 21115 -725
rect 21080 -770 21115 -750
rect 21140 -585 21175 -575
rect 21140 -610 21145 -585
rect 21170 -610 21175 -585
rect 21140 -630 21175 -610
rect 21140 -655 21145 -630
rect 21170 -655 21175 -630
rect 21140 -675 21175 -655
rect 21140 -700 21145 -675
rect 21170 -700 21175 -675
rect 21140 -725 21175 -700
rect 21140 -750 21145 -725
rect 21170 -750 21175 -725
rect 21140 -770 21175 -750
rect 21200 -585 21235 -575
rect 21200 -610 21205 -585
rect 21230 -610 21235 -585
rect 21200 -630 21235 -610
rect 21200 -655 21205 -630
rect 21230 -655 21235 -630
rect 21200 -675 21235 -655
rect 21200 -700 21205 -675
rect 21230 -700 21235 -675
rect 21200 -725 21235 -700
rect 21200 -750 21205 -725
rect 21230 -750 21235 -725
rect 21200 -770 21235 -750
rect 21260 -585 21295 -575
rect 21260 -610 21265 -585
rect 21290 -610 21295 -585
rect 21260 -630 21295 -610
rect 21260 -655 21265 -630
rect 21290 -655 21295 -630
rect 21260 -675 21295 -655
rect 21260 -700 21265 -675
rect 21290 -700 21295 -675
rect 21260 -725 21295 -700
rect 21260 -750 21265 -725
rect 21290 -750 21295 -725
rect 21260 -770 21295 -750
rect 21320 -585 21355 -575
rect 21320 -610 21325 -585
rect 21350 -610 21355 -585
rect 21320 -630 21355 -610
rect 21320 -655 21325 -630
rect 21350 -655 21355 -630
rect 21320 -675 21355 -655
rect 21320 -700 21325 -675
rect 21350 -700 21355 -675
rect 21320 -725 21355 -700
rect 21320 -750 21325 -725
rect 21350 -750 21355 -725
rect 21320 -770 21355 -750
rect 21380 -585 21415 -575
rect 21380 -610 21385 -585
rect 21410 -610 21415 -585
rect 21380 -630 21415 -610
rect 21380 -655 21385 -630
rect 21410 -655 21415 -630
rect 21380 -675 21415 -655
rect 21380 -700 21385 -675
rect 21410 -700 21415 -675
rect 21380 -725 21415 -700
rect 21380 -750 21385 -725
rect 21410 -750 21415 -725
rect 21380 -770 21415 -750
rect 21440 -585 21475 -575
rect 21440 -610 21445 -585
rect 21470 -610 21475 -585
rect 21440 -630 21475 -610
rect 21440 -655 21445 -630
rect 21470 -655 21475 -630
rect 21440 -675 21475 -655
rect 21440 -700 21445 -675
rect 21470 -700 21475 -675
rect 21440 -725 21475 -700
rect 21440 -750 21445 -725
rect 21470 -750 21475 -725
rect 21440 -770 21475 -750
rect 21500 -585 21535 -575
rect 21500 -610 21505 -585
rect 21530 -610 21535 -585
rect 21500 -630 21535 -610
rect 21500 -655 21505 -630
rect 21530 -655 21535 -630
rect 21500 -675 21535 -655
rect 21500 -700 21505 -675
rect 21530 -700 21535 -675
rect 21500 -725 21535 -700
rect 21500 -750 21505 -725
rect 21530 -750 21535 -725
rect 21500 -770 21535 -750
rect 21560 -585 21595 -575
rect 21560 -610 21565 -585
rect 21590 -610 21595 -585
rect 21560 -630 21595 -610
rect 21560 -655 21565 -630
rect 21590 -655 21595 -630
rect 21560 -675 21595 -655
rect 21560 -700 21565 -675
rect 21590 -700 21595 -675
rect 21560 -725 21595 -700
rect 21560 -750 21565 -725
rect 21590 -750 21595 -725
rect 21560 -770 21595 -750
rect 21620 -585 21655 -575
rect 21620 -610 21625 -585
rect 21650 -610 21655 -585
rect 21620 -630 21655 -610
rect 21620 -655 21625 -630
rect 21650 -655 21655 -630
rect 21620 -675 21655 -655
rect 21620 -700 21625 -675
rect 21650 -700 21655 -675
rect 21620 -725 21655 -700
rect 21620 -750 21625 -725
rect 21650 -750 21655 -725
rect 21620 -770 21655 -750
rect 21680 -585 21715 -575
rect 21680 -610 21685 -585
rect 21710 -610 21715 -585
rect 21680 -630 21715 -610
rect 21680 -655 21685 -630
rect 21710 -655 21715 -630
rect 21680 -675 21715 -655
rect 21680 -700 21685 -675
rect 21710 -700 21715 -675
rect 21680 -725 21715 -700
rect 21680 -750 21685 -725
rect 21710 -750 21715 -725
rect 21680 -770 21715 -750
rect 21740 -585 21775 -575
rect 21740 -610 21745 -585
rect 21770 -610 21775 -585
rect 21740 -630 21775 -610
rect 21740 -655 21745 -630
rect 21770 -655 21775 -630
rect 21740 -675 21775 -655
rect 21740 -700 21745 -675
rect 21770 -700 21775 -675
rect 21740 -725 21775 -700
rect 21740 -750 21745 -725
rect 21770 -750 21775 -725
rect 21740 -770 21775 -750
rect 21800 -585 21835 -575
rect 21800 -610 21805 -585
rect 21830 -610 21835 -585
rect 21800 -630 21835 -610
rect 21800 -655 21805 -630
rect 21830 -655 21835 -630
rect 21800 -675 21835 -655
rect 21800 -700 21805 -675
rect 21830 -700 21835 -675
rect 21800 -725 21835 -700
rect 21800 -750 21805 -725
rect 21830 -750 21835 -725
rect 21800 -770 21835 -750
rect 21860 -585 21895 -575
rect 21860 -610 21865 -585
rect 21890 -610 21895 -585
rect 21860 -630 21895 -610
rect 21860 -655 21865 -630
rect 21890 -655 21895 -630
rect 21860 -675 21895 -655
rect 21860 -700 21865 -675
rect 21890 -700 21895 -675
rect 21860 -725 21895 -700
rect 21860 -750 21865 -725
rect 21890 -750 21895 -725
rect 21860 -770 21895 -750
rect 21920 -585 21955 -575
rect 21920 -610 21925 -585
rect 21950 -610 21955 -585
rect 21920 -630 21955 -610
rect 21920 -655 21925 -630
rect 21950 -655 21955 -630
rect 21920 -675 21955 -655
rect 21920 -700 21925 -675
rect 21950 -700 21955 -675
rect 21920 -725 21955 -700
rect 21920 -750 21925 -725
rect 21950 -750 21955 -725
rect 21920 -770 21955 -750
rect 21980 -585 22015 -575
rect 21980 -610 21985 -585
rect 22010 -610 22015 -585
rect 21980 -630 22015 -610
rect 21980 -655 21985 -630
rect 22010 -655 22015 -630
rect 21980 -675 22015 -655
rect 21980 -700 21985 -675
rect 22010 -700 22015 -675
rect 21980 -725 22015 -700
rect 21980 -750 21985 -725
rect 22010 -750 22015 -725
rect 21980 -770 22015 -750
rect 22040 -585 22075 -575
rect 22040 -610 22045 -585
rect 22070 -610 22075 -585
rect 22040 -630 22075 -610
rect 22040 -655 22045 -630
rect 22070 -655 22075 -630
rect 22040 -675 22075 -655
rect 22040 -700 22045 -675
rect 22070 -700 22075 -675
rect 22040 -725 22075 -700
rect 22040 -750 22045 -725
rect 22070 -750 22075 -725
rect 22040 -770 22075 -750
rect 22100 -585 22135 -575
rect 22100 -610 22105 -585
rect 22130 -610 22135 -585
rect 22100 -630 22135 -610
rect 22100 -655 22105 -630
rect 22130 -655 22135 -630
rect 22100 -675 22135 -655
rect 22100 -700 22105 -675
rect 22130 -700 22135 -675
rect 22100 -725 22135 -700
rect 22100 -750 22105 -725
rect 22130 -750 22135 -725
rect 22100 -770 22135 -750
rect 22160 -585 22195 -575
rect 22160 -610 22165 -585
rect 22190 -610 22195 -585
rect 22160 -630 22195 -610
rect 22160 -655 22165 -630
rect 22190 -655 22195 -630
rect 22160 -675 22195 -655
rect 22160 -700 22165 -675
rect 22190 -700 22195 -675
rect 22160 -725 22195 -700
rect 22160 -750 22165 -725
rect 22190 -750 22195 -725
rect 22160 -770 22195 -750
rect 22220 -585 22255 -575
rect 22220 -610 22225 -585
rect 22250 -610 22255 -585
rect 22220 -630 22255 -610
rect 22220 -655 22225 -630
rect 22250 -655 22255 -630
rect 22220 -675 22255 -655
rect 22220 -700 22225 -675
rect 22250 -700 22255 -675
rect 22220 -725 22255 -700
rect 22220 -750 22225 -725
rect 22250 -750 22255 -725
rect 22220 -770 22255 -750
rect 22280 -585 22315 -575
rect 22280 -610 22285 -585
rect 22310 -610 22315 -585
rect 22280 -630 22315 -610
rect 22280 -655 22285 -630
rect 22310 -655 22315 -630
rect 22280 -675 22315 -655
rect 22280 -700 22285 -675
rect 22310 -700 22315 -675
rect 22280 -725 22315 -700
rect 22280 -750 22285 -725
rect 22310 -750 22315 -725
rect 22280 -770 22315 -750
rect 22340 -585 22375 -575
rect 22340 -610 22345 -585
rect 22370 -610 22375 -585
rect 22340 -630 22375 -610
rect 22340 -655 22345 -630
rect 22370 -655 22375 -630
rect 22340 -675 22375 -655
rect 22340 -700 22345 -675
rect 22370 -700 22375 -675
rect 22340 -725 22375 -700
rect 22340 -750 22345 -725
rect 22370 -750 22375 -725
rect 22340 -770 22375 -750
rect 22400 -585 22435 -575
rect 22400 -610 22405 -585
rect 22430 -610 22435 -585
rect 22400 -630 22435 -610
rect 22400 -655 22405 -630
rect 22430 -655 22435 -630
rect 22400 -675 22435 -655
rect 22400 -700 22405 -675
rect 22430 -700 22435 -675
rect 22400 -725 22435 -700
rect 22400 -750 22405 -725
rect 22430 -750 22435 -725
rect 22400 -770 22435 -750
rect 22460 -585 22495 -575
rect 22460 -610 22465 -585
rect 22490 -610 22495 -585
rect 22460 -630 22495 -610
rect 22460 -655 22465 -630
rect 22490 -655 22495 -630
rect 22460 -675 22495 -655
rect 22460 -700 22465 -675
rect 22490 -700 22495 -675
rect 22460 -725 22495 -700
rect 22460 -750 22465 -725
rect 22490 -750 22495 -725
rect 22460 -770 22495 -750
rect 22520 -585 22555 -575
rect 22520 -610 22525 -585
rect 22550 -610 22555 -585
rect 22520 -630 22555 -610
rect 22520 -655 22525 -630
rect 22550 -655 22555 -630
rect 22520 -675 22555 -655
rect 22520 -700 22525 -675
rect 22550 -700 22555 -675
rect 22520 -725 22555 -700
rect 22520 -750 22525 -725
rect 22550 -750 22555 -725
rect 22520 -770 22555 -750
rect 22580 -585 22615 -575
rect 22580 -610 22585 -585
rect 22610 -610 22615 -585
rect 22580 -630 22615 -610
rect 22580 -655 22585 -630
rect 22610 -655 22615 -630
rect 22580 -675 22615 -655
rect 22580 -700 22585 -675
rect 22610 -700 22615 -675
rect 22580 -725 22615 -700
rect 22580 -750 22585 -725
rect 22610 -750 22615 -725
rect 22580 -770 22615 -750
rect 22640 -585 22675 -575
rect 22640 -610 22645 -585
rect 22670 -610 22675 -585
rect 22640 -630 22675 -610
rect 22640 -655 22645 -630
rect 22670 -655 22675 -630
rect 22640 -675 22675 -655
rect 22640 -700 22645 -675
rect 22670 -700 22675 -675
rect 22640 -725 22675 -700
rect 22640 -750 22645 -725
rect 22670 -750 22675 -725
rect 22640 -770 22675 -750
rect 22700 -585 22735 -575
rect 22700 -610 22705 -585
rect 22730 -610 22735 -585
rect 22700 -630 22735 -610
rect 22700 -655 22705 -630
rect 22730 -655 22735 -630
rect 22700 -675 22735 -655
rect 22700 -700 22705 -675
rect 22730 -700 22735 -675
rect 22700 -725 22735 -700
rect 22700 -750 22705 -725
rect 22730 -750 22735 -725
rect 22700 -770 22735 -750
rect 22760 -585 22795 -575
rect 22760 -610 22765 -585
rect 22790 -610 22795 -585
rect 22760 -630 22795 -610
rect 22760 -655 22765 -630
rect 22790 -655 22795 -630
rect 22760 -675 22795 -655
rect 22760 -700 22765 -675
rect 22790 -700 22795 -675
rect 22760 -725 22795 -700
rect 22760 -750 22765 -725
rect 22790 -750 22795 -725
rect 22760 -770 22795 -750
rect 22820 -585 22855 -575
rect 22820 -610 22825 -585
rect 22850 -610 22855 -585
rect 22820 -630 22855 -610
rect 22820 -655 22825 -630
rect 22850 -655 22855 -630
rect 22820 -675 22855 -655
rect 22820 -700 22825 -675
rect 22850 -700 22855 -675
rect 22820 -725 22855 -700
rect 22820 -750 22825 -725
rect 22850 -750 22855 -725
rect 22820 -770 22855 -750
rect 22880 -585 22915 -575
rect 22880 -610 22885 -585
rect 22910 -610 22915 -585
rect 22880 -630 22915 -610
rect 22880 -655 22885 -630
rect 22910 -655 22915 -630
rect 22880 -675 22915 -655
rect 22880 -700 22885 -675
rect 22910 -700 22915 -675
rect 22880 -725 22915 -700
rect 22880 -750 22885 -725
rect 22910 -750 22915 -725
rect 22880 -770 22915 -750
rect 22940 -585 22975 -575
rect 22940 -610 22945 -585
rect 22970 -610 22975 -585
rect 22940 -630 22975 -610
rect 22940 -655 22945 -630
rect 22970 -655 22975 -630
rect 22940 -675 22975 -655
rect 22940 -700 22945 -675
rect 22970 -700 22975 -675
rect 22940 -725 22975 -700
rect 22940 -750 22945 -725
rect 22970 -750 22975 -725
rect 22940 -770 22975 -750
rect 23000 -585 23035 -575
rect 23000 -610 23005 -585
rect 23030 -610 23035 -585
rect 23000 -630 23035 -610
rect 23000 -655 23005 -630
rect 23030 -655 23035 -630
rect 23000 -675 23035 -655
rect 23000 -700 23005 -675
rect 23030 -700 23035 -675
rect 23000 -725 23035 -700
rect 23000 -750 23005 -725
rect 23030 -750 23035 -725
rect 23000 -770 23035 -750
rect 23060 -585 23095 -575
rect 23060 -610 23065 -585
rect 23090 -610 23095 -585
rect 23060 -630 23095 -610
rect 23060 -655 23065 -630
rect 23090 -655 23095 -630
rect 23060 -675 23095 -655
rect 23060 -700 23065 -675
rect 23090 -700 23095 -675
rect 23060 -725 23095 -700
rect 23060 -750 23065 -725
rect 23090 -750 23095 -725
rect 23060 -770 23095 -750
rect 23120 -585 23155 -575
rect 23120 -610 23125 -585
rect 23150 -610 23155 -585
rect 23120 -630 23155 -610
rect 23120 -655 23125 -630
rect 23150 -655 23155 -630
rect 23120 -675 23155 -655
rect 23120 -700 23125 -675
rect 23150 -700 23155 -675
rect 23120 -725 23155 -700
rect 23120 -750 23125 -725
rect 23150 -750 23155 -725
rect 23120 -770 23155 -750
rect 23180 -585 23215 -575
rect 23180 -610 23185 -585
rect 23210 -610 23215 -585
rect 23180 -630 23215 -610
rect 23180 -655 23185 -630
rect 23210 -655 23215 -630
rect 23180 -675 23215 -655
rect 23180 -700 23185 -675
rect 23210 -700 23215 -675
rect 23180 -725 23215 -700
rect 23180 -750 23185 -725
rect 23210 -750 23215 -725
rect 23180 -770 23215 -750
rect 23240 -585 23275 -575
rect 23240 -610 23245 -585
rect 23270 -610 23275 -585
rect 23240 -630 23275 -610
rect 23240 -655 23245 -630
rect 23270 -655 23275 -630
rect 23240 -675 23275 -655
rect 23240 -700 23245 -675
rect 23270 -700 23275 -675
rect 23240 -725 23275 -700
rect 23240 -750 23245 -725
rect 23270 -750 23275 -725
rect 23240 -770 23275 -750
rect 23300 -585 23335 -575
rect 23300 -610 23305 -585
rect 23330 -610 23335 -585
rect 23300 -630 23335 -610
rect 23300 -655 23305 -630
rect 23330 -655 23335 -630
rect 23300 -675 23335 -655
rect 23300 -700 23305 -675
rect 23330 -700 23335 -675
rect 23300 -725 23335 -700
rect 23300 -750 23305 -725
rect 23330 -750 23335 -725
rect 23300 -770 23335 -750
rect 23360 -585 23395 -575
rect 23360 -610 23365 -585
rect 23390 -610 23395 -585
rect 23360 -630 23395 -610
rect 23360 -655 23365 -630
rect 23390 -655 23395 -630
rect 23360 -675 23395 -655
rect 23360 -700 23365 -675
rect 23390 -700 23395 -675
rect 23360 -725 23395 -700
rect 23360 -750 23365 -725
rect 23390 -750 23395 -725
rect 23360 -770 23395 -750
rect 23420 -585 23455 -575
rect 23420 -610 23425 -585
rect 23450 -610 23455 -585
rect 23420 -630 23455 -610
rect 23420 -655 23425 -630
rect 23450 -655 23455 -630
rect 23420 -675 23455 -655
rect 23420 -700 23425 -675
rect 23450 -700 23455 -675
rect 23420 -725 23455 -700
rect 23420 -750 23425 -725
rect 23450 -750 23455 -725
rect 23420 -770 23455 -750
rect 23480 -585 23515 -575
rect 23480 -610 23485 -585
rect 23510 -610 23515 -585
rect 23480 -630 23515 -610
rect 23480 -655 23485 -630
rect 23510 -655 23515 -630
rect 23480 -675 23515 -655
rect 23480 -700 23485 -675
rect 23510 -700 23515 -675
rect 23480 -725 23515 -700
rect 23480 -750 23485 -725
rect 23510 -750 23515 -725
rect 23480 -770 23515 -750
rect 23540 -585 23575 -575
rect 23540 -610 23545 -585
rect 23570 -610 23575 -585
rect 23540 -630 23575 -610
rect 23540 -655 23545 -630
rect 23570 -655 23575 -630
rect 23540 -675 23575 -655
rect 23540 -700 23545 -675
rect 23570 -700 23575 -675
rect 23540 -725 23575 -700
rect 23540 -750 23545 -725
rect 23570 -750 23575 -725
rect 23540 -770 23575 -750
rect 23600 -585 23635 -575
rect 23600 -610 23605 -585
rect 23630 -610 23635 -585
rect 23600 -630 23635 -610
rect 23600 -655 23605 -630
rect 23630 -655 23635 -630
rect 23600 -675 23635 -655
rect 23600 -700 23605 -675
rect 23630 -700 23635 -675
rect 23600 -725 23635 -700
rect 23600 -750 23605 -725
rect 23630 -750 23635 -725
rect 23600 -770 23635 -750
rect 23660 -585 23695 -575
rect 23660 -610 23665 -585
rect 23690 -610 23695 -585
rect 23660 -630 23695 -610
rect 23660 -655 23665 -630
rect 23690 -655 23695 -630
rect 23660 -675 23695 -655
rect 23660 -700 23665 -675
rect 23690 -700 23695 -675
rect 23660 -725 23695 -700
rect 23660 -750 23665 -725
rect 23690 -750 23695 -725
rect 23660 -770 23695 -750
rect 23720 -585 23755 -575
rect 23720 -610 23725 -585
rect 23750 -610 23755 -585
rect 23720 -630 23755 -610
rect 23720 -655 23725 -630
rect 23750 -655 23755 -630
rect 23720 -675 23755 -655
rect 23720 -700 23725 -675
rect 23750 -700 23755 -675
rect 23720 -725 23755 -700
rect 23720 -750 23725 -725
rect 23750 -750 23755 -725
rect 23720 -770 23755 -750
rect 23780 -585 23815 -575
rect 23780 -610 23785 -585
rect 23810 -610 23815 -585
rect 23780 -630 23815 -610
rect 23780 -655 23785 -630
rect 23810 -655 23815 -630
rect 23780 -675 23815 -655
rect 23780 -700 23785 -675
rect 23810 -700 23815 -675
rect 23780 -725 23815 -700
rect 23780 -750 23785 -725
rect 23810 -750 23815 -725
rect 23780 -770 23815 -750
rect 23840 -585 23875 -575
rect 23840 -610 23845 -585
rect 23870 -610 23875 -585
rect 23840 -630 23875 -610
rect 23840 -655 23845 -630
rect 23870 -655 23875 -630
rect 23840 -675 23875 -655
rect 23840 -700 23845 -675
rect 23870 -700 23875 -675
rect 23840 -725 23875 -700
rect 23840 -750 23845 -725
rect 23870 -750 23875 -725
rect 23840 -770 23875 -750
rect 23900 -585 23935 -575
rect 23900 -610 23905 -585
rect 23930 -610 23935 -585
rect 23900 -630 23935 -610
rect 23900 -655 23905 -630
rect 23930 -655 23935 -630
rect 23900 -675 23935 -655
rect 23900 -700 23905 -675
rect 23930 -700 23935 -675
rect 23900 -725 23935 -700
rect 23900 -750 23905 -725
rect 23930 -750 23935 -725
rect 23900 -770 23935 -750
rect 23960 -585 23995 -575
rect 23960 -610 23965 -585
rect 23990 -610 23995 -585
rect 23960 -630 23995 -610
rect 23960 -655 23965 -630
rect 23990 -655 23995 -630
rect 23960 -675 23995 -655
rect 23960 -700 23965 -675
rect 23990 -700 23995 -675
rect 23960 -725 23995 -700
rect 23960 -750 23965 -725
rect 23990 -750 23995 -725
rect 23960 -770 23995 -750
rect 24020 -585 24055 -575
rect 24020 -610 24025 -585
rect 24050 -610 24055 -585
rect 24020 -630 24055 -610
rect 24020 -655 24025 -630
rect 24050 -655 24055 -630
rect 24020 -675 24055 -655
rect 24020 -700 24025 -675
rect 24050 -700 24055 -675
rect 24020 -725 24055 -700
rect 24020 -750 24025 -725
rect 24050 -750 24055 -725
rect 24020 -770 24055 -750
rect 24080 -585 24115 -575
rect 24080 -610 24085 -585
rect 24110 -610 24115 -585
rect 24080 -630 24115 -610
rect 24080 -655 24085 -630
rect 24110 -655 24115 -630
rect 24080 -675 24115 -655
rect 24080 -700 24085 -675
rect 24110 -700 24115 -675
rect 24080 -725 24115 -700
rect 24080 -750 24085 -725
rect 24110 -750 24115 -725
rect 24080 -770 24115 -750
rect 24140 -585 24175 -575
rect 24140 -610 24145 -585
rect 24170 -610 24175 -585
rect 24140 -630 24175 -610
rect 24140 -655 24145 -630
rect 24170 -655 24175 -630
rect 24140 -675 24175 -655
rect 24140 -700 24145 -675
rect 24170 -700 24175 -675
rect 24140 -725 24175 -700
rect 24140 -750 24145 -725
rect 24170 -750 24175 -725
rect 24140 -770 24175 -750
rect 24200 -585 24235 -575
rect 24200 -610 24205 -585
rect 24230 -610 24235 -585
rect 24200 -630 24235 -610
rect 24200 -655 24205 -630
rect 24230 -655 24235 -630
rect 24200 -675 24235 -655
rect 24200 -700 24205 -675
rect 24230 -700 24235 -675
rect 24200 -725 24235 -700
rect 24200 -750 24205 -725
rect 24230 -750 24235 -725
rect 24200 -770 24235 -750
rect 24260 -585 24295 -575
rect 24260 -610 24265 -585
rect 24290 -610 24295 -585
rect 24260 -630 24295 -610
rect 24260 -655 24265 -630
rect 24290 -655 24295 -630
rect 24260 -675 24295 -655
rect 24260 -700 24265 -675
rect 24290 -700 24295 -675
rect 24260 -725 24295 -700
rect 24260 -750 24265 -725
rect 24290 -750 24295 -725
rect 24260 -770 24295 -750
rect 24320 -585 24355 -575
rect 24320 -610 24325 -585
rect 24350 -610 24355 -585
rect 24320 -630 24355 -610
rect 24320 -655 24325 -630
rect 24350 -655 24355 -630
rect 24320 -675 24355 -655
rect 24320 -700 24325 -675
rect 24350 -700 24355 -675
rect 24320 -725 24355 -700
rect 24320 -750 24325 -725
rect 24350 -750 24355 -725
rect 24320 -770 24355 -750
rect 24380 -585 24415 -575
rect 24380 -610 24385 -585
rect 24410 -610 24415 -585
rect 24380 -630 24415 -610
rect 24380 -655 24385 -630
rect 24410 -655 24415 -630
rect 24380 -675 24415 -655
rect 24380 -700 24385 -675
rect 24410 -700 24415 -675
rect 24380 -725 24415 -700
rect 24380 -750 24385 -725
rect 24410 -750 24415 -725
rect 24380 -770 24415 -750
rect 24440 -585 24475 -575
rect 24440 -610 24445 -585
rect 24470 -610 24475 -585
rect 24440 -630 24475 -610
rect 24440 -655 24445 -630
rect 24470 -655 24475 -630
rect 24440 -675 24475 -655
rect 24440 -700 24445 -675
rect 24470 -700 24475 -675
rect 24440 -725 24475 -700
rect 24440 -750 24445 -725
rect 24470 -750 24475 -725
rect 24440 -770 24475 -750
rect 24500 -585 24535 -575
rect 24500 -610 24505 -585
rect 24530 -610 24535 -585
rect 24500 -630 24535 -610
rect 24500 -655 24505 -630
rect 24530 -655 24535 -630
rect 24500 -675 24535 -655
rect 24500 -700 24505 -675
rect 24530 -700 24535 -675
rect 24500 -725 24535 -700
rect 24500 -750 24505 -725
rect 24530 -750 24535 -725
rect 24500 -770 24535 -750
rect 24560 -585 24595 -575
rect 24560 -610 24565 -585
rect 24590 -610 24595 -585
rect 24560 -630 24595 -610
rect 24560 -655 24565 -630
rect 24590 -655 24595 -630
rect 24560 -675 24595 -655
rect 24560 -700 24565 -675
rect 24590 -700 24595 -675
rect 24560 -725 24595 -700
rect 24560 -750 24565 -725
rect 24590 -750 24595 -725
rect 24560 -770 24595 -750
rect 24620 -585 24655 -575
rect 24620 -610 24625 -585
rect 24650 -610 24655 -585
rect 24620 -630 24655 -610
rect 24620 -655 24625 -630
rect 24650 -655 24655 -630
rect 24620 -675 24655 -655
rect 24620 -700 24625 -675
rect 24650 -700 24655 -675
rect 24620 -725 24655 -700
rect 24620 -750 24625 -725
rect 24650 -750 24655 -725
rect 24620 -770 24655 -750
rect 24680 -585 24715 -575
rect 24680 -610 24685 -585
rect 24710 -610 24715 -585
rect 24680 -630 24715 -610
rect 24680 -655 24685 -630
rect 24710 -655 24715 -630
rect 24680 -675 24715 -655
rect 24680 -700 24685 -675
rect 24710 -700 24715 -675
rect 24680 -725 24715 -700
rect 24680 -750 24685 -725
rect 24710 -750 24715 -725
rect 24680 -770 24715 -750
rect 24740 -585 24775 -575
rect 24740 -610 24745 -585
rect 24770 -610 24775 -585
rect 24740 -630 24775 -610
rect 24740 -655 24745 -630
rect 24770 -655 24775 -630
rect 24740 -675 24775 -655
rect 24740 -700 24745 -675
rect 24770 -700 24775 -675
rect 24740 -725 24775 -700
rect 24740 -750 24745 -725
rect 24770 -750 24775 -725
rect 24740 -770 24775 -750
rect 24800 -585 24835 -575
rect 24800 -610 24805 -585
rect 24830 -610 24835 -585
rect 24800 -630 24835 -610
rect 24800 -655 24805 -630
rect 24830 -655 24835 -630
rect 24800 -675 24835 -655
rect 24800 -700 24805 -675
rect 24830 -700 24835 -675
rect 24800 -725 24835 -700
rect 24800 -750 24805 -725
rect 24830 -750 24835 -725
rect 24800 -770 24835 -750
rect 24860 -585 24895 -575
rect 24860 -610 24865 -585
rect 24890 -610 24895 -585
rect 24860 -630 24895 -610
rect 24860 -655 24865 -630
rect 24890 -655 24895 -630
rect 24860 -675 24895 -655
rect 24860 -700 24865 -675
rect 24890 -700 24895 -675
rect 24860 -725 24895 -700
rect 24860 -750 24865 -725
rect 24890 -750 24895 -725
rect 24860 -770 24895 -750
rect 24920 -585 24955 -575
rect 24920 -610 24925 -585
rect 24950 -610 24955 -585
rect 24920 -630 24955 -610
rect 24920 -655 24925 -630
rect 24950 -655 24955 -630
rect 24920 -675 24955 -655
rect 24920 -700 24925 -675
rect 24950 -700 24955 -675
rect 24920 -725 24955 -700
rect 24920 -750 24925 -725
rect 24950 -750 24955 -725
rect 24920 -770 24955 -750
rect 24980 -585 25015 -575
rect 24980 -610 24985 -585
rect 25010 -610 25015 -585
rect 24980 -630 25015 -610
rect 24980 -655 24985 -630
rect 25010 -655 25015 -630
rect 24980 -675 25015 -655
rect 24980 -700 24985 -675
rect 25010 -700 25015 -675
rect 24980 -725 25015 -700
rect 24980 -750 24985 -725
rect 25010 -750 25015 -725
rect 24980 -770 25015 -750
rect 25040 -585 25075 -575
rect 25040 -610 25045 -585
rect 25070 -610 25075 -585
rect 25040 -630 25075 -610
rect 25040 -655 25045 -630
rect 25070 -655 25075 -630
rect 25040 -675 25075 -655
rect 25040 -700 25045 -675
rect 25070 -700 25075 -675
rect 25040 -725 25075 -700
rect 25040 -750 25045 -725
rect 25070 -750 25075 -725
rect 25040 -770 25075 -750
rect 25100 -585 25135 -575
rect 25100 -610 25105 -585
rect 25130 -610 25135 -585
rect 25100 -630 25135 -610
rect 25100 -655 25105 -630
rect 25130 -655 25135 -630
rect 25100 -675 25135 -655
rect 25100 -700 25105 -675
rect 25130 -700 25135 -675
rect 25100 -725 25135 -700
rect 25100 -750 25105 -725
rect 25130 -750 25135 -725
rect 25100 -770 25135 -750
rect 25160 -585 25195 -575
rect 25160 -610 25165 -585
rect 25190 -610 25195 -585
rect 25160 -630 25195 -610
rect 25160 -655 25165 -630
rect 25190 -655 25195 -630
rect 25160 -675 25195 -655
rect 25160 -700 25165 -675
rect 25190 -700 25195 -675
rect 25160 -725 25195 -700
rect 25160 -750 25165 -725
rect 25190 -750 25195 -725
rect 25160 -770 25195 -750
rect 25220 -585 25255 -575
rect 25220 -610 25225 -585
rect 25250 -610 25255 -585
rect 25220 -630 25255 -610
rect 25220 -655 25225 -630
rect 25250 -655 25255 -630
rect 25220 -675 25255 -655
rect 25220 -700 25225 -675
rect 25250 -700 25255 -675
rect 25220 -725 25255 -700
rect 25220 -750 25225 -725
rect 25250 -750 25255 -725
rect 25220 -770 25255 -750
rect 25280 -585 25315 -575
rect 25280 -610 25285 -585
rect 25310 -610 25315 -585
rect 25280 -630 25315 -610
rect 25280 -655 25285 -630
rect 25310 -655 25315 -630
rect 25280 -675 25315 -655
rect 25280 -700 25285 -675
rect 25310 -700 25315 -675
rect 25280 -725 25315 -700
rect 25280 -750 25285 -725
rect 25310 -750 25315 -725
rect 25280 -770 25315 -750
rect 25340 -585 25375 -575
rect 25340 -610 25345 -585
rect 25370 -610 25375 -585
rect 25340 -630 25375 -610
rect 25340 -655 25345 -630
rect 25370 -655 25375 -630
rect 25340 -675 25375 -655
rect 25340 -700 25345 -675
rect 25370 -700 25375 -675
rect 25340 -725 25375 -700
rect 25340 -750 25345 -725
rect 25370 -750 25375 -725
rect 25340 -770 25375 -750
rect 25400 -585 25435 -575
rect 25400 -610 25405 -585
rect 25430 -610 25435 -585
rect 25400 -630 25435 -610
rect 25400 -655 25405 -630
rect 25430 -655 25435 -630
rect 25400 -675 25435 -655
rect 25400 -700 25405 -675
rect 25430 -700 25435 -675
rect 25400 -725 25435 -700
rect 25400 -750 25405 -725
rect 25430 -750 25435 -725
rect 25400 -770 25435 -750
rect 25460 -585 25495 -575
rect 25460 -610 25465 -585
rect 25490 -610 25495 -585
rect 25460 -630 25495 -610
rect 25460 -655 25465 -630
rect 25490 -655 25495 -630
rect 25460 -675 25495 -655
rect 25460 -700 25465 -675
rect 25490 -700 25495 -675
rect 25460 -725 25495 -700
rect 25460 -750 25465 -725
rect 25490 -750 25495 -725
rect 25460 -770 25495 -750
rect 25520 -585 25555 -575
rect 25520 -610 25525 -585
rect 25550 -610 25555 -585
rect 25520 -630 25555 -610
rect 25520 -655 25525 -630
rect 25550 -655 25555 -630
rect 25520 -675 25555 -655
rect 25520 -700 25525 -675
rect 25550 -700 25555 -675
rect 25520 -725 25555 -700
rect 25520 -750 25525 -725
rect 25550 -750 25555 -725
rect 25520 -770 25555 -750
rect 25580 -585 25615 -575
rect 25580 -610 25585 -585
rect 25610 -610 25615 -585
rect 25580 -630 25615 -610
rect 25580 -655 25585 -630
rect 25610 -655 25615 -630
rect 25580 -675 25615 -655
rect 25580 -700 25585 -675
rect 25610 -700 25615 -675
rect 25580 -725 25615 -700
rect 25580 -750 25585 -725
rect 25610 -750 25615 -725
rect 25580 -770 25615 -750
rect 25640 -585 25675 -575
rect 25640 -610 25645 -585
rect 25670 -610 25675 -585
rect 25640 -630 25675 -610
rect 25640 -655 25645 -630
rect 25670 -655 25675 -630
rect 25640 -675 25675 -655
rect 25640 -700 25645 -675
rect 25670 -700 25675 -675
rect 25640 -725 25675 -700
rect 25640 -750 25645 -725
rect 25670 -750 25675 -725
rect 25640 -770 25675 -750
rect 25700 -585 25735 -575
rect 25700 -610 25705 -585
rect 25730 -610 25735 -585
rect 25700 -630 25735 -610
rect 25700 -655 25705 -630
rect 25730 -655 25735 -630
rect 25700 -675 25735 -655
rect 25700 -700 25705 -675
rect 25730 -700 25735 -675
rect 25700 -725 25735 -700
rect 25700 -750 25705 -725
rect 25730 -750 25735 -725
rect 25700 -770 25735 -750
rect 25760 -585 25795 -575
rect 25760 -610 25765 -585
rect 25790 -610 25795 -585
rect 25760 -630 25795 -610
rect 25760 -655 25765 -630
rect 25790 -655 25795 -630
rect 25760 -675 25795 -655
rect 25760 -700 25765 -675
rect 25790 -700 25795 -675
rect 25760 -725 25795 -700
rect 25760 -750 25765 -725
rect 25790 -750 25795 -725
rect 25760 -770 25795 -750
rect 25820 -585 25855 -575
rect 25820 -610 25825 -585
rect 25850 -610 25855 -585
rect 25820 -630 25855 -610
rect 25820 -655 25825 -630
rect 25850 -655 25855 -630
rect 25820 -675 25855 -655
rect 25820 -700 25825 -675
rect 25850 -700 25855 -675
rect 25820 -725 25855 -700
rect 25820 -750 25825 -725
rect 25850 -750 25855 -725
rect 25820 -770 25855 -750
rect 25880 -585 25915 -575
rect 25880 -610 25885 -585
rect 25910 -610 25915 -585
rect 25880 -630 25915 -610
rect 25880 -655 25885 -630
rect 25910 -655 25915 -630
rect 25880 -675 25915 -655
rect 25880 -700 25885 -675
rect 25910 -700 25915 -675
rect 25880 -725 25915 -700
rect 25880 -750 25885 -725
rect 25910 -750 25915 -725
rect 25880 -770 25915 -750
rect 25940 -585 25975 -575
rect 25940 -610 25945 -585
rect 25970 -610 25975 -585
rect 25940 -630 25975 -610
rect 25940 -655 25945 -630
rect 25970 -655 25975 -630
rect 25940 -675 25975 -655
rect 25940 -700 25945 -675
rect 25970 -700 25975 -675
rect 25940 -725 25975 -700
rect 25940 -750 25945 -725
rect 25970 -750 25975 -725
rect 25940 -770 25975 -750
rect 26000 -585 26035 -575
rect 26000 -610 26005 -585
rect 26030 -610 26035 -585
rect 26000 -630 26035 -610
rect 26000 -655 26005 -630
rect 26030 -655 26035 -630
rect 26000 -675 26035 -655
rect 26000 -700 26005 -675
rect 26030 -700 26035 -675
rect 26000 -725 26035 -700
rect 26000 -750 26005 -725
rect 26030 -750 26035 -725
rect 26000 -770 26035 -750
rect 26060 -585 26095 -575
rect 26060 -610 26065 -585
rect 26090 -610 26095 -585
rect 26060 -630 26095 -610
rect 26060 -655 26065 -630
rect 26090 -655 26095 -630
rect 26060 -675 26095 -655
rect 26060 -700 26065 -675
rect 26090 -700 26095 -675
rect 26060 -725 26095 -700
rect 26060 -750 26065 -725
rect 26090 -750 26095 -725
rect 26060 -770 26095 -750
rect 26120 -585 26155 -575
rect 26120 -610 26125 -585
rect 26150 -610 26155 -585
rect 26120 -630 26155 -610
rect 26120 -655 26125 -630
rect 26150 -655 26155 -630
rect 26120 -675 26155 -655
rect 26120 -700 26125 -675
rect 26150 -700 26155 -675
rect 26120 -725 26155 -700
rect 26120 -750 26125 -725
rect 26150 -750 26155 -725
rect 26120 -770 26155 -750
rect 26180 -585 26215 -575
rect 26180 -610 26185 -585
rect 26210 -610 26215 -585
rect 26180 -630 26215 -610
rect 26180 -655 26185 -630
rect 26210 -655 26215 -630
rect 26180 -675 26215 -655
rect 26180 -700 26185 -675
rect 26210 -700 26215 -675
rect 26180 -725 26215 -700
rect 26180 -750 26185 -725
rect 26210 -750 26215 -725
rect 26180 -770 26215 -750
rect 26240 -585 26275 -575
rect 26240 -610 26245 -585
rect 26270 -610 26275 -585
rect 26240 -630 26275 -610
rect 26240 -655 26245 -630
rect 26270 -655 26275 -630
rect 26240 -675 26275 -655
rect 26240 -700 26245 -675
rect 26270 -700 26275 -675
rect 26240 -725 26275 -700
rect 26240 -750 26245 -725
rect 26270 -750 26275 -725
rect 26240 -770 26275 -750
rect 26300 -585 26335 -575
rect 26300 -610 26305 -585
rect 26330 -610 26335 -585
rect 26300 -630 26335 -610
rect 26300 -655 26305 -630
rect 26330 -655 26335 -630
rect 26300 -675 26335 -655
rect 26300 -700 26305 -675
rect 26330 -700 26335 -675
rect 26300 -725 26335 -700
rect 26300 -750 26305 -725
rect 26330 -750 26335 -725
rect 26300 -770 26335 -750
rect 26360 -585 26395 -575
rect 26360 -610 26365 -585
rect 26390 -610 26395 -585
rect 26360 -630 26395 -610
rect 26360 -655 26365 -630
rect 26390 -655 26395 -630
rect 26360 -675 26395 -655
rect 26360 -700 26365 -675
rect 26390 -700 26395 -675
rect 26360 -725 26395 -700
rect 26360 -750 26365 -725
rect 26390 -750 26395 -725
rect 26360 -770 26395 -750
rect 26420 -585 26455 -575
rect 26420 -610 26425 -585
rect 26450 -610 26455 -585
rect 26420 -630 26455 -610
rect 26420 -655 26425 -630
rect 26450 -655 26455 -630
rect 26420 -675 26455 -655
rect 26420 -700 26425 -675
rect 26450 -700 26455 -675
rect 26420 -725 26455 -700
rect 26420 -750 26425 -725
rect 26450 -750 26455 -725
rect 26420 -770 26455 -750
rect 26480 -585 26515 -575
rect 26480 -610 26485 -585
rect 26510 -610 26515 -585
rect 26480 -630 26515 -610
rect 26480 -655 26485 -630
rect 26510 -655 26515 -630
rect 26480 -675 26515 -655
rect 26480 -700 26485 -675
rect 26510 -700 26515 -675
rect 26480 -725 26515 -700
rect 26480 -750 26485 -725
rect 26510 -750 26515 -725
rect 26480 -770 26515 -750
rect 26540 -585 26575 -575
rect 26540 -610 26545 -585
rect 26570 -610 26575 -585
rect 26540 -630 26575 -610
rect 26540 -655 26545 -630
rect 26570 -655 26575 -630
rect 26540 -675 26575 -655
rect 26540 -700 26545 -675
rect 26570 -700 26575 -675
rect 26540 -725 26575 -700
rect 26540 -750 26545 -725
rect 26570 -750 26575 -725
rect 26540 -770 26575 -750
rect 26600 -585 26635 -575
rect 26600 -610 26605 -585
rect 26630 -610 26635 -585
rect 26600 -630 26635 -610
rect 26600 -655 26605 -630
rect 26630 -655 26635 -630
rect 26600 -675 26635 -655
rect 26600 -700 26605 -675
rect 26630 -700 26635 -675
rect 26600 -725 26635 -700
rect 26600 -750 26605 -725
rect 26630 -750 26635 -725
rect 26600 -770 26635 -750
rect 26660 -585 26695 -575
rect 26660 -610 26665 -585
rect 26690 -610 26695 -585
rect 26660 -630 26695 -610
rect 26660 -655 26665 -630
rect 26690 -655 26695 -630
rect 26660 -675 26695 -655
rect 26660 -700 26665 -675
rect 26690 -700 26695 -675
rect 26660 -725 26695 -700
rect 26660 -750 26665 -725
rect 26690 -750 26695 -725
rect 26660 -770 26695 -750
rect 26720 -585 26755 -575
rect 26720 -610 26725 -585
rect 26750 -610 26755 -585
rect 26720 -630 26755 -610
rect 26720 -655 26725 -630
rect 26750 -655 26755 -630
rect 26720 -675 26755 -655
rect 26720 -700 26725 -675
rect 26750 -700 26755 -675
rect 26720 -725 26755 -700
rect 26720 -750 26725 -725
rect 26750 -750 26755 -725
rect 26720 -770 26755 -750
rect 26780 -585 26815 -575
rect 26780 -610 26785 -585
rect 26810 -610 26815 -585
rect 26780 -630 26815 -610
rect 26780 -655 26785 -630
rect 26810 -655 26815 -630
rect 26780 -675 26815 -655
rect 26780 -700 26785 -675
rect 26810 -700 26815 -675
rect 26780 -725 26815 -700
rect 26780 -750 26785 -725
rect 26810 -750 26815 -725
rect 26780 -770 26815 -750
rect 26840 -585 26875 -575
rect 26840 -610 26845 -585
rect 26870 -610 26875 -585
rect 26840 -630 26875 -610
rect 26840 -655 26845 -630
rect 26870 -655 26875 -630
rect 26840 -675 26875 -655
rect 26840 -700 26845 -675
rect 26870 -700 26875 -675
rect 26840 -725 26875 -700
rect 26840 -750 26845 -725
rect 26870 -750 26875 -725
rect 26840 -770 26875 -750
rect 26900 -585 26935 -575
rect 26900 -610 26905 -585
rect 26930 -610 26935 -585
rect 26900 -630 26935 -610
rect 26900 -655 26905 -630
rect 26930 -655 26935 -630
rect 26900 -675 26935 -655
rect 26900 -700 26905 -675
rect 26930 -700 26935 -675
rect 26900 -725 26935 -700
rect 26900 -750 26905 -725
rect 26930 -750 26935 -725
rect 26900 -770 26935 -750
rect 26960 -585 26995 -575
rect 26960 -610 26965 -585
rect 26990 -610 26995 -585
rect 26960 -630 26995 -610
rect 26960 -655 26965 -630
rect 26990 -655 26995 -630
rect 26960 -675 26995 -655
rect 26960 -700 26965 -675
rect 26990 -700 26995 -675
rect 26960 -725 26995 -700
rect 26960 -750 26965 -725
rect 26990 -750 26995 -725
rect 26960 -770 26995 -750
rect 27020 -585 27055 -575
rect 27020 -610 27025 -585
rect 27050 -610 27055 -585
rect 27020 -630 27055 -610
rect 27020 -655 27025 -630
rect 27050 -655 27055 -630
rect 27020 -675 27055 -655
rect 27020 -700 27025 -675
rect 27050 -700 27055 -675
rect 27020 -725 27055 -700
rect 27020 -750 27025 -725
rect 27050 -750 27055 -725
rect 27020 -770 27055 -750
rect 27080 -585 27115 -575
rect 27080 -610 27085 -585
rect 27110 -610 27115 -585
rect 27080 -630 27115 -610
rect 27080 -655 27085 -630
rect 27110 -655 27115 -630
rect 27080 -675 27115 -655
rect 27080 -700 27085 -675
rect 27110 -700 27115 -675
rect 27080 -725 27115 -700
rect 27080 -750 27085 -725
rect 27110 -750 27115 -725
rect 27080 -770 27115 -750
rect 27140 -585 27175 -575
rect 27140 -610 27145 -585
rect 27170 -610 27175 -585
rect 27140 -630 27175 -610
rect 27140 -655 27145 -630
rect 27170 -655 27175 -630
rect 27140 -675 27175 -655
rect 27140 -700 27145 -675
rect 27170 -700 27175 -675
rect 27140 -725 27175 -700
rect 27140 -750 27145 -725
rect 27170 -750 27175 -725
rect 27140 -770 27175 -750
rect 27200 -585 27235 -575
rect 27200 -610 27205 -585
rect 27230 -610 27235 -585
rect 27200 -630 27235 -610
rect 27200 -655 27205 -630
rect 27230 -655 27235 -630
rect 27200 -675 27235 -655
rect 27200 -700 27205 -675
rect 27230 -700 27235 -675
rect 27200 -725 27235 -700
rect 27200 -750 27205 -725
rect 27230 -750 27235 -725
rect 27200 -770 27235 -750
rect 27260 -585 27295 -575
rect 27260 -610 27265 -585
rect 27290 -610 27295 -585
rect 27260 -630 27295 -610
rect 27260 -655 27265 -630
rect 27290 -655 27295 -630
rect 27260 -675 27295 -655
rect 27260 -700 27265 -675
rect 27290 -700 27295 -675
rect 27260 -725 27295 -700
rect 27260 -750 27265 -725
rect 27290 -750 27295 -725
rect 27260 -770 27295 -750
rect 27320 -585 27355 -575
rect 27320 -610 27325 -585
rect 27350 -610 27355 -585
rect 27320 -630 27355 -610
rect 27320 -655 27325 -630
rect 27350 -655 27355 -630
rect 27320 -675 27355 -655
rect 27320 -700 27325 -675
rect 27350 -700 27355 -675
rect 27320 -725 27355 -700
rect 27320 -750 27325 -725
rect 27350 -750 27355 -725
rect 27320 -770 27355 -750
rect 27380 -585 27415 -575
rect 27380 -610 27385 -585
rect 27410 -610 27415 -585
rect 27380 -630 27415 -610
rect 27380 -655 27385 -630
rect 27410 -655 27415 -630
rect 27380 -675 27415 -655
rect 27380 -700 27385 -675
rect 27410 -700 27415 -675
rect 27380 -725 27415 -700
rect 27380 -750 27385 -725
rect 27410 -750 27415 -725
rect 27380 -770 27415 -750
rect 27440 -585 27475 -575
rect 27440 -610 27445 -585
rect 27470 -610 27475 -585
rect 27440 -630 27475 -610
rect 27440 -655 27445 -630
rect 27470 -655 27475 -630
rect 27440 -675 27475 -655
rect 27440 -700 27445 -675
rect 27470 -700 27475 -675
rect 27440 -725 27475 -700
rect 27440 -750 27445 -725
rect 27470 -750 27475 -725
rect 27440 -770 27475 -750
rect 27500 -585 27535 -575
rect 27500 -610 27505 -585
rect 27530 -610 27535 -585
rect 27500 -630 27535 -610
rect 27500 -655 27505 -630
rect 27530 -655 27535 -630
rect 27500 -675 27535 -655
rect 27500 -700 27505 -675
rect 27530 -700 27535 -675
rect 27500 -725 27535 -700
rect 27500 -750 27505 -725
rect 27530 -750 27535 -725
rect 27500 -770 27535 -750
rect 27560 -585 27595 -575
rect 27560 -610 27565 -585
rect 27590 -610 27595 -585
rect 27560 -630 27595 -610
rect 27560 -655 27565 -630
rect 27590 -655 27595 -630
rect 27560 -675 27595 -655
rect 27560 -700 27565 -675
rect 27590 -700 27595 -675
rect 27560 -725 27595 -700
rect 27560 -750 27565 -725
rect 27590 -750 27595 -725
rect 27560 -770 27595 -750
rect 27620 -585 27655 -575
rect 27620 -610 27625 -585
rect 27650 -610 27655 -585
rect 27620 -630 27655 -610
rect 27620 -655 27625 -630
rect 27650 -655 27655 -630
rect 27620 -675 27655 -655
rect 27620 -700 27625 -675
rect 27650 -700 27655 -675
rect 27620 -725 27655 -700
rect 27620 -750 27625 -725
rect 27650 -750 27655 -725
rect 27620 -770 27655 -750
rect 27680 -585 27715 -575
rect 27680 -610 27685 -585
rect 27710 -610 27715 -585
rect 27680 -630 27715 -610
rect 27680 -655 27685 -630
rect 27710 -655 27715 -630
rect 27680 -675 27715 -655
rect 27680 -700 27685 -675
rect 27710 -700 27715 -675
rect 27680 -725 27715 -700
rect 27680 -750 27685 -725
rect 27710 -750 27715 -725
rect 27680 -770 27715 -750
rect 27740 -585 27775 -575
rect 27740 -610 27745 -585
rect 27770 -610 27775 -585
rect 27740 -630 27775 -610
rect 27740 -655 27745 -630
rect 27770 -655 27775 -630
rect 27740 -675 27775 -655
rect 27740 -700 27745 -675
rect 27770 -700 27775 -675
rect 27740 -725 27775 -700
rect 27740 -750 27745 -725
rect 27770 -750 27775 -725
rect 27740 -770 27775 -750
rect 27800 -585 27835 -575
rect 27800 -610 27805 -585
rect 27830 -610 27835 -585
rect 27800 -630 27835 -610
rect 27800 -655 27805 -630
rect 27830 -655 27835 -630
rect 27800 -675 27835 -655
rect 27800 -700 27805 -675
rect 27830 -700 27835 -675
rect 27800 -725 27835 -700
rect 27800 -750 27805 -725
rect 27830 -750 27835 -725
rect 27800 -770 27835 -750
rect 27860 -585 27895 -575
rect 27860 -610 27865 -585
rect 27890 -610 27895 -585
rect 27860 -630 27895 -610
rect 27860 -655 27865 -630
rect 27890 -655 27895 -630
rect 27860 -675 27895 -655
rect 27860 -700 27865 -675
rect 27890 -700 27895 -675
rect 27860 -725 27895 -700
rect 27860 -750 27865 -725
rect 27890 -750 27895 -725
rect 27860 -770 27895 -750
rect 27920 -585 27955 -575
rect 27920 -610 27925 -585
rect 27950 -610 27955 -585
rect 27920 -630 27955 -610
rect 27920 -655 27925 -630
rect 27950 -655 27955 -630
rect 27920 -675 27955 -655
rect 27920 -700 27925 -675
rect 27950 -700 27955 -675
rect 27920 -725 27955 -700
rect 27920 -750 27925 -725
rect 27950 -750 27955 -725
rect 27920 -770 27955 -750
rect 27980 -585 28015 -575
rect 27980 -610 27985 -585
rect 28010 -610 28015 -585
rect 27980 -630 28015 -610
rect 27980 -655 27985 -630
rect 28010 -655 28015 -630
rect 27980 -675 28015 -655
rect 27980 -700 27985 -675
rect 28010 -700 28015 -675
rect 27980 -725 28015 -700
rect 27980 -750 27985 -725
rect 28010 -750 28015 -725
rect 27980 -770 28015 -750
rect 28040 -585 28075 -575
rect 28040 -610 28045 -585
rect 28070 -610 28075 -585
rect 28040 -630 28075 -610
rect 28040 -655 28045 -630
rect 28070 -655 28075 -630
rect 28040 -675 28075 -655
rect 28040 -700 28045 -675
rect 28070 -700 28075 -675
rect 28040 -725 28075 -700
rect 28040 -750 28045 -725
rect 28070 -750 28075 -725
rect 28040 -770 28075 -750
rect 28100 -585 28135 -575
rect 28100 -610 28105 -585
rect 28130 -610 28135 -585
rect 28100 -630 28135 -610
rect 28100 -655 28105 -630
rect 28130 -655 28135 -630
rect 28100 -675 28135 -655
rect 28100 -700 28105 -675
rect 28130 -700 28135 -675
rect 28100 -725 28135 -700
rect 28100 -750 28105 -725
rect 28130 -750 28135 -725
rect 28100 -770 28135 -750
rect 28160 -585 28195 -575
rect 28160 -610 28165 -585
rect 28190 -610 28195 -585
rect 28160 -630 28195 -610
rect 28160 -655 28165 -630
rect 28190 -655 28195 -630
rect 28160 -675 28195 -655
rect 28160 -700 28165 -675
rect 28190 -700 28195 -675
rect 28160 -725 28195 -700
rect 28160 -750 28165 -725
rect 28190 -750 28195 -725
rect 28160 -770 28195 -750
rect 28220 -585 28255 -575
rect 28220 -610 28225 -585
rect 28250 -610 28255 -585
rect 28220 -630 28255 -610
rect 28220 -655 28225 -630
rect 28250 -655 28255 -630
rect 28220 -675 28255 -655
rect 28220 -700 28225 -675
rect 28250 -700 28255 -675
rect 28220 -725 28255 -700
rect 28220 -750 28225 -725
rect 28250 -750 28255 -725
rect 28220 -770 28255 -750
rect 28280 -585 28315 -575
rect 28280 -610 28285 -585
rect 28310 -610 28315 -585
rect 28280 -630 28315 -610
rect 28280 -655 28285 -630
rect 28310 -655 28315 -630
rect 28280 -675 28315 -655
rect 28280 -700 28285 -675
rect 28310 -700 28315 -675
rect 28280 -725 28315 -700
rect 28280 -750 28285 -725
rect 28310 -750 28315 -725
rect 28280 -770 28315 -750
rect 28340 -585 28375 -575
rect 28340 -610 28345 -585
rect 28370 -610 28375 -585
rect 28340 -630 28375 -610
rect 28340 -655 28345 -630
rect 28370 -655 28375 -630
rect 28340 -675 28375 -655
rect 28340 -700 28345 -675
rect 28370 -700 28375 -675
rect 28340 -725 28375 -700
rect 28340 -750 28345 -725
rect 28370 -750 28375 -725
rect 28340 -770 28375 -750
rect 28400 -585 28435 -575
rect 28400 -610 28405 -585
rect 28430 -610 28435 -585
rect 28400 -630 28435 -610
rect 28400 -655 28405 -630
rect 28430 -655 28435 -630
rect 28400 -675 28435 -655
rect 28400 -700 28405 -675
rect 28430 -700 28435 -675
rect 28400 -725 28435 -700
rect 28400 -750 28405 -725
rect 28430 -750 28435 -725
rect 28400 -770 28435 -750
rect 28460 -585 28495 -575
rect 28460 -610 28465 -585
rect 28490 -610 28495 -585
rect 28460 -630 28495 -610
rect 28460 -655 28465 -630
rect 28490 -655 28495 -630
rect 28460 -675 28495 -655
rect 28460 -700 28465 -675
rect 28490 -700 28495 -675
rect 28460 -725 28495 -700
rect 28460 -750 28465 -725
rect 28490 -750 28495 -725
rect 28460 -770 28495 -750
rect 28520 -585 28555 -575
rect 28520 -610 28525 -585
rect 28550 -610 28555 -585
rect 28520 -630 28555 -610
rect 28520 -655 28525 -630
rect 28550 -655 28555 -630
rect 28520 -675 28555 -655
rect 28520 -700 28525 -675
rect 28550 -700 28555 -675
rect 28520 -725 28555 -700
rect 28520 -750 28525 -725
rect 28550 -750 28555 -725
rect 28520 -770 28555 -750
rect 28580 -585 28615 -575
rect 28580 -610 28585 -585
rect 28610 -610 28615 -585
rect 28580 -630 28615 -610
rect 28580 -655 28585 -630
rect 28610 -655 28615 -630
rect 28580 -675 28615 -655
rect 28580 -700 28585 -675
rect 28610 -700 28615 -675
rect 28580 -725 28615 -700
rect 28580 -750 28585 -725
rect 28610 -750 28615 -725
rect 28580 -770 28615 -750
rect 28640 -585 28675 -575
rect 28640 -610 28645 -585
rect 28670 -610 28675 -585
rect 28640 -630 28675 -610
rect 28640 -655 28645 -630
rect 28670 -655 28675 -630
rect 28640 -675 28675 -655
rect 28640 -700 28645 -675
rect 28670 -700 28675 -675
rect 28640 -725 28675 -700
rect 28640 -750 28645 -725
rect 28670 -750 28675 -725
rect 28640 -770 28675 -750
rect 28700 -585 28735 -575
rect 28700 -610 28705 -585
rect 28730 -610 28735 -585
rect 28700 -630 28735 -610
rect 28700 -655 28705 -630
rect 28730 -655 28735 -630
rect 28700 -675 28735 -655
rect 28700 -700 28705 -675
rect 28730 -700 28735 -675
rect 28700 -725 28735 -700
rect 28700 -750 28705 -725
rect 28730 -750 28735 -725
rect 28700 -770 28735 -750
rect 28760 -585 28795 -575
rect 28760 -610 28765 -585
rect 28790 -610 28795 -585
rect 28760 -630 28795 -610
rect 28760 -655 28765 -630
rect 28790 -655 28795 -630
rect 28760 -675 28795 -655
rect 28760 -700 28765 -675
rect 28790 -700 28795 -675
rect 28760 -725 28795 -700
rect 28760 -750 28765 -725
rect 28790 -750 28795 -725
rect 28760 -770 28795 -750
rect 28820 -585 28855 -575
rect 28820 -610 28825 -585
rect 28850 -610 28855 -585
rect 28820 -630 28855 -610
rect 28820 -655 28825 -630
rect 28850 -655 28855 -630
rect 28820 -675 28855 -655
rect 28820 -700 28825 -675
rect 28850 -700 28855 -675
rect 28820 -725 28855 -700
rect 28820 -750 28825 -725
rect 28850 -750 28855 -725
rect 28820 -770 28855 -750
rect 28880 -585 28915 -575
rect 28880 -610 28885 -585
rect 28910 -610 28915 -585
rect 28880 -630 28915 -610
rect 28880 -655 28885 -630
rect 28910 -655 28915 -630
rect 28880 -675 28915 -655
rect 28880 -700 28885 -675
rect 28910 -700 28915 -675
rect 28880 -725 28915 -700
rect 28880 -750 28885 -725
rect 28910 -750 28915 -725
rect 28880 -770 28915 -750
rect 28940 -585 28975 -575
rect 28940 -610 28945 -585
rect 28970 -610 28975 -585
rect 28940 -630 28975 -610
rect 28940 -655 28945 -630
rect 28970 -655 28975 -630
rect 28940 -675 28975 -655
rect 28940 -700 28945 -675
rect 28970 -700 28975 -675
rect 28940 -725 28975 -700
rect 28940 -750 28945 -725
rect 28970 -750 28975 -725
rect 28940 -770 28975 -750
rect 29000 -585 29035 -575
rect 29000 -610 29005 -585
rect 29030 -610 29035 -585
rect 29000 -630 29035 -610
rect 29000 -655 29005 -630
rect 29030 -655 29035 -630
rect 29000 -675 29035 -655
rect 29000 -700 29005 -675
rect 29030 -700 29035 -675
rect 29000 -725 29035 -700
rect 29000 -750 29005 -725
rect 29030 -750 29035 -725
rect 29000 -770 29035 -750
rect 29060 -585 29095 -575
rect 29060 -610 29065 -585
rect 29090 -610 29095 -585
rect 29060 -630 29095 -610
rect 29060 -655 29065 -630
rect 29090 -655 29095 -630
rect 29060 -675 29095 -655
rect 29060 -700 29065 -675
rect 29090 -700 29095 -675
rect 29060 -725 29095 -700
rect 29060 -750 29065 -725
rect 29090 -750 29095 -725
rect 29060 -770 29095 -750
rect 29120 -585 29155 -575
rect 29120 -610 29125 -585
rect 29150 -610 29155 -585
rect 29120 -630 29155 -610
rect 29120 -655 29125 -630
rect 29150 -655 29155 -630
rect 29120 -675 29155 -655
rect 29120 -700 29125 -675
rect 29150 -700 29155 -675
rect 29120 -725 29155 -700
rect 29120 -750 29125 -725
rect 29150 -750 29155 -725
rect 29120 -770 29155 -750
rect 29180 -585 29215 -575
rect 29180 -610 29185 -585
rect 29210 -610 29215 -585
rect 29180 -630 29215 -610
rect 29180 -655 29185 -630
rect 29210 -655 29215 -630
rect 29180 -675 29215 -655
rect 29180 -700 29185 -675
rect 29210 -700 29215 -675
rect 29180 -725 29215 -700
rect 29180 -750 29185 -725
rect 29210 -750 29215 -725
rect 29180 -770 29215 -750
rect 29240 -585 29275 -575
rect 29240 -610 29245 -585
rect 29270 -610 29275 -585
rect 29240 -630 29275 -610
rect 29240 -655 29245 -630
rect 29270 -655 29275 -630
rect 29240 -675 29275 -655
rect 29240 -700 29245 -675
rect 29270 -700 29275 -675
rect 29240 -725 29275 -700
rect 29240 -750 29245 -725
rect 29270 -750 29275 -725
rect 29240 -770 29275 -750
rect 29300 -585 29335 -575
rect 29300 -610 29305 -585
rect 29330 -610 29335 -585
rect 29300 -630 29335 -610
rect 29300 -655 29305 -630
rect 29330 -655 29335 -630
rect 29300 -675 29335 -655
rect 29300 -700 29305 -675
rect 29330 -700 29335 -675
rect 29300 -725 29335 -700
rect 29300 -750 29305 -725
rect 29330 -750 29335 -725
rect 29300 -770 29335 -750
rect 29360 -585 29395 -575
rect 29360 -610 29365 -585
rect 29390 -610 29395 -585
rect 29360 -630 29395 -610
rect 29360 -655 29365 -630
rect 29390 -655 29395 -630
rect 29360 -675 29395 -655
rect 29360 -700 29365 -675
rect 29390 -700 29395 -675
rect 29360 -725 29395 -700
rect 29360 -750 29365 -725
rect 29390 -750 29395 -725
rect 29360 -770 29395 -750
rect 29420 -585 29455 -575
rect 29420 -610 29425 -585
rect 29450 -610 29455 -585
rect 29420 -630 29455 -610
rect 29420 -655 29425 -630
rect 29450 -655 29455 -630
rect 29420 -675 29455 -655
rect 29420 -700 29425 -675
rect 29450 -700 29455 -675
rect 29420 -725 29455 -700
rect 29420 -750 29425 -725
rect 29450 -750 29455 -725
rect 29420 -770 29455 -750
rect 29480 -585 29515 -575
rect 29480 -610 29485 -585
rect 29510 -610 29515 -585
rect 29480 -630 29515 -610
rect 29480 -655 29485 -630
rect 29510 -655 29515 -630
rect 29480 -675 29515 -655
rect 29480 -700 29485 -675
rect 29510 -700 29515 -675
rect 29480 -725 29515 -700
rect 29480 -750 29485 -725
rect 29510 -750 29515 -725
rect 29480 -770 29515 -750
rect 29540 -585 29575 -575
rect 29540 -610 29545 -585
rect 29570 -610 29575 -585
rect 29540 -630 29575 -610
rect 29540 -655 29545 -630
rect 29570 -655 29575 -630
rect 29540 -675 29575 -655
rect 29540 -700 29545 -675
rect 29570 -700 29575 -675
rect 29540 -725 29575 -700
rect 29540 -750 29545 -725
rect 29570 -750 29575 -725
rect 29540 -770 29575 -750
rect 29600 -585 29635 -575
rect 29600 -610 29605 -585
rect 29630 -610 29635 -585
rect 29600 -630 29635 -610
rect 29600 -655 29605 -630
rect 29630 -655 29635 -630
rect 29600 -675 29635 -655
rect 29600 -700 29605 -675
rect 29630 -700 29635 -675
rect 29600 -725 29635 -700
rect 29600 -750 29605 -725
rect 29630 -750 29635 -725
rect 29600 -770 29635 -750
rect 29660 -585 29695 -575
rect 29660 -610 29665 -585
rect 29690 -610 29695 -585
rect 29660 -630 29695 -610
rect 29660 -655 29665 -630
rect 29690 -655 29695 -630
rect 29660 -675 29695 -655
rect 29660 -700 29665 -675
rect 29690 -700 29695 -675
rect 29660 -725 29695 -700
rect 29660 -750 29665 -725
rect 29690 -750 29695 -725
rect 29660 -770 29695 -750
rect 29720 -585 29755 -575
rect 29720 -610 29725 -585
rect 29750 -610 29755 -585
rect 29720 -630 29755 -610
rect 29720 -655 29725 -630
rect 29750 -655 29755 -630
rect 29720 -675 29755 -655
rect 29720 -700 29725 -675
rect 29750 -700 29755 -675
rect 29720 -725 29755 -700
rect 29720 -750 29725 -725
rect 29750 -750 29755 -725
rect 29720 -770 29755 -750
rect 29780 -585 29815 -575
rect 29780 -610 29785 -585
rect 29810 -610 29815 -585
rect 29780 -630 29815 -610
rect 29780 -655 29785 -630
rect 29810 -655 29815 -630
rect 29780 -675 29815 -655
rect 29780 -700 29785 -675
rect 29810 -700 29815 -675
rect 29780 -725 29815 -700
rect 29780 -750 29785 -725
rect 29810 -750 29815 -725
rect 29780 -770 29815 -750
rect 29840 -585 29875 -575
rect 29840 -610 29845 -585
rect 29870 -610 29875 -585
rect 29840 -630 29875 -610
rect 29840 -655 29845 -630
rect 29870 -655 29875 -630
rect 29840 -675 29875 -655
rect 29840 -700 29845 -675
rect 29870 -700 29875 -675
rect 29840 -725 29875 -700
rect 29840 -750 29845 -725
rect 29870 -750 29875 -725
rect 29840 -770 29875 -750
rect 29900 -585 29935 -575
rect 29900 -610 29905 -585
rect 29930 -610 29935 -585
rect 29900 -630 29935 -610
rect 29900 -655 29905 -630
rect 29930 -655 29935 -630
rect 29900 -675 29935 -655
rect 29900 -700 29905 -675
rect 29930 -700 29935 -675
rect 29900 -725 29935 -700
rect 29900 -750 29905 -725
rect 29930 -750 29935 -725
rect 29900 -770 29935 -750
rect 29960 -585 29995 -575
rect 29960 -610 29965 -585
rect 29990 -610 29995 -585
rect 29960 -630 29995 -610
rect 29960 -655 29965 -630
rect 29990 -655 29995 -630
rect 29960 -675 29995 -655
rect 29960 -700 29965 -675
rect 29990 -700 29995 -675
rect 29960 -725 29995 -700
rect 29960 -750 29965 -725
rect 29990 -750 29995 -725
rect 29960 -770 29995 -750
rect 30020 -585 30055 -575
rect 30020 -610 30025 -585
rect 30050 -610 30055 -585
rect 30020 -630 30055 -610
rect 30020 -655 30025 -630
rect 30050 -655 30055 -630
rect 30020 -675 30055 -655
rect 30020 -700 30025 -675
rect 30050 -700 30055 -675
rect 30020 -725 30055 -700
rect 30020 -750 30025 -725
rect 30050 -750 30055 -725
rect 30020 -770 30055 -750
rect 30080 -585 30115 -575
rect 30080 -610 30085 -585
rect 30110 -610 30115 -585
rect 30080 -630 30115 -610
rect 30080 -655 30085 -630
rect 30110 -655 30115 -630
rect 30080 -675 30115 -655
rect 30080 -700 30085 -675
rect 30110 -700 30115 -675
rect 30080 -725 30115 -700
rect 30080 -750 30085 -725
rect 30110 -750 30115 -725
rect 30080 -770 30115 -750
rect 30140 -585 30175 -575
rect 30140 -610 30145 -585
rect 30170 -610 30175 -585
rect 30140 -630 30175 -610
rect 30140 -655 30145 -630
rect 30170 -655 30175 -630
rect 30140 -675 30175 -655
rect 30140 -700 30145 -675
rect 30170 -700 30175 -675
rect 30140 -725 30175 -700
rect 30140 -750 30145 -725
rect 30170 -750 30175 -725
rect 30140 -770 30175 -750
rect 30200 -585 30235 -575
rect 30200 -610 30205 -585
rect 30230 -610 30235 -585
rect 30200 -630 30235 -610
rect 30200 -655 30205 -630
rect 30230 -655 30235 -630
rect 30200 -675 30235 -655
rect 30200 -700 30205 -675
rect 30230 -700 30235 -675
rect 30200 -725 30235 -700
rect 30200 -750 30205 -725
rect 30230 -750 30235 -725
rect 30200 -770 30235 -750
rect 30260 -585 30295 -575
rect 30260 -610 30265 -585
rect 30290 -610 30295 -585
rect 30260 -630 30295 -610
rect 30260 -655 30265 -630
rect 30290 -655 30295 -630
rect 30260 -675 30295 -655
rect 30260 -700 30265 -675
rect 30290 -700 30295 -675
rect 30260 -725 30295 -700
rect 30260 -750 30265 -725
rect 30290 -750 30295 -725
rect 30260 -770 30295 -750
rect 30320 -585 30355 -575
rect 30320 -610 30325 -585
rect 30350 -610 30355 -585
rect 30320 -630 30355 -610
rect 30320 -655 30325 -630
rect 30350 -655 30355 -630
rect 30320 -675 30355 -655
rect 30320 -700 30325 -675
rect 30350 -700 30355 -675
rect 30320 -725 30355 -700
rect 30320 -750 30325 -725
rect 30350 -750 30355 -725
rect 30320 -770 30355 -750
rect 30380 -585 30415 -575
rect 30380 -610 30385 -585
rect 30410 -610 30415 -585
rect 30380 -630 30415 -610
rect 30380 -655 30385 -630
rect 30410 -655 30415 -630
rect 30380 -675 30415 -655
rect 30380 -700 30385 -675
rect 30410 -700 30415 -675
rect 30380 -725 30415 -700
rect 30380 -750 30385 -725
rect 30410 -750 30415 -725
rect 30380 -770 30415 -750
rect 30440 -585 30475 -575
rect 30440 -610 30445 -585
rect 30470 -610 30475 -585
rect 30440 -630 30475 -610
rect 30440 -655 30445 -630
rect 30470 -655 30475 -630
rect 30440 -675 30475 -655
rect 30440 -700 30445 -675
rect 30470 -700 30475 -675
rect 30440 -725 30475 -700
rect 30440 -750 30445 -725
rect 30470 -750 30475 -725
rect 30440 -770 30475 -750
rect 30500 -585 30535 -575
rect 30500 -610 30505 -585
rect 30530 -610 30535 -585
rect 30500 -630 30535 -610
rect 30500 -655 30505 -630
rect 30530 -655 30535 -630
rect 30500 -675 30535 -655
rect 30500 -700 30505 -675
rect 30530 -700 30535 -675
rect 30500 -725 30535 -700
rect 30500 -750 30505 -725
rect 30530 -750 30535 -725
rect 30500 -770 30535 -750
rect 30560 -585 30595 -575
rect 30560 -610 30565 -585
rect 30590 -610 30595 -585
rect 30560 -630 30595 -610
rect 30560 -655 30565 -630
rect 30590 -655 30595 -630
rect 30560 -675 30595 -655
rect 30560 -700 30565 -675
rect 30590 -700 30595 -675
rect 30560 -725 30595 -700
rect 30560 -750 30565 -725
rect 30590 -750 30595 -725
rect 30560 -770 30595 -750
rect 30620 -585 30655 -575
rect 30620 -610 30625 -585
rect 30650 -610 30655 -585
rect 30620 -630 30655 -610
rect 30620 -655 30625 -630
rect 30650 -655 30655 -630
rect 30620 -675 30655 -655
rect 30620 -700 30625 -675
rect 30650 -700 30655 -675
rect 30620 -725 30655 -700
rect 30620 -750 30625 -725
rect 30650 -750 30655 -725
rect 30620 -770 30655 -750
rect 30680 -585 30715 -575
rect 30680 -610 30685 -585
rect 30710 -610 30715 -585
rect 30680 -630 30715 -610
rect 30680 -655 30685 -630
rect 30710 -655 30715 -630
rect 30680 -675 30715 -655
rect 30680 -700 30685 -675
rect 30710 -700 30715 -675
rect 30680 -725 30715 -700
rect 30680 -750 30685 -725
rect 30710 -750 30715 -725
rect 30680 -770 30715 -750
rect 31060 -770 31200 -320
rect 25 -785 45 -770
rect 85 -810 110 -770
rect 145 -785 165 -770
rect 265 -785 285 -770
rect 325 -810 350 -770
rect 385 -785 405 -770
rect 505 -785 525 -770
rect 565 -810 590 -770
rect 625 -785 645 -770
rect 745 -785 765 -770
rect 80 -825 115 -810
rect 80 -850 85 -825
rect 110 -850 115 -825
rect 80 -860 115 -850
rect 320 -825 355 -810
rect 320 -850 325 -825
rect 350 -850 355 -825
rect 320 -860 355 -850
rect 560 -825 595 -810
rect 805 -825 830 -770
rect 865 -785 885 -770
rect 985 -785 1005 -770
rect 1045 -810 1070 -770
rect 1105 -785 1125 -770
rect 1225 -785 1245 -770
rect 1285 -810 1310 -770
rect 1345 -785 1365 -770
rect 1465 -785 1485 -770
rect 1525 -810 1550 -770
rect 1585 -785 1605 -770
rect 1705 -785 1725 -770
rect 1765 -810 1790 -770
rect 1825 -785 1845 -770
rect 1945 -785 1965 -770
rect 2005 -810 2030 -770
rect 2065 -785 2085 -770
rect 2185 -785 2205 -770
rect 2245 -810 2270 -770
rect 2305 -785 2325 -770
rect 2425 -785 2445 -770
rect 2485 -810 2510 -770
rect 2545 -785 2565 -770
rect 2665 -785 2685 -770
rect 2725 -810 2750 -770
rect 2785 -785 2805 -770
rect 2905 -785 2925 -770
rect 1040 -825 1075 -810
rect 560 -850 565 -825
rect 590 -850 595 -825
rect 560 -860 595 -850
rect 790 -835 845 -825
rect 790 -870 800 -835
rect 835 -870 845 -835
rect 1040 -850 1045 -825
rect 1070 -850 1075 -825
rect 1040 -860 1075 -850
rect 1280 -825 1315 -810
rect 1280 -850 1285 -825
rect 1310 -850 1315 -825
rect 1280 -860 1315 -850
rect 1520 -825 1555 -810
rect 1520 -850 1525 -825
rect 1550 -850 1555 -825
rect 1520 -860 1555 -850
rect 1760 -825 1795 -810
rect 1760 -850 1765 -825
rect 1790 -850 1795 -825
rect 1760 -860 1795 -850
rect 2000 -825 2035 -810
rect 2000 -850 2005 -825
rect 2030 -850 2035 -825
rect 2000 -860 2035 -850
rect 2240 -825 2275 -810
rect 2240 -850 2245 -825
rect 2270 -850 2275 -825
rect 2240 -860 2275 -850
rect 2480 -825 2515 -810
rect 2480 -850 2485 -825
rect 2510 -850 2515 -825
rect 2480 -860 2515 -850
rect 2720 -825 2755 -810
rect 2965 -825 2990 -770
rect 3025 -785 3045 -770
rect 3145 -785 3165 -770
rect 3205 -810 3230 -770
rect 3265 -785 3285 -770
rect 3385 -785 3405 -770
rect 3445 -810 3470 -770
rect 3505 -785 3525 -770
rect 3625 -785 3645 -770
rect 3685 -810 3710 -770
rect 3745 -785 3765 -770
rect 3865 -785 3885 -770
rect 3925 -810 3950 -770
rect 3985 -785 4005 -770
rect 4105 -785 4125 -770
rect 4165 -810 4190 -770
rect 4225 -785 4245 -770
rect 4345 -785 4365 -770
rect 4405 -810 4430 -770
rect 4465 -785 4485 -770
rect 4585 -785 4605 -770
rect 4645 -810 4670 -770
rect 4705 -785 4725 -770
rect 4825 -785 4845 -770
rect 4885 -810 4910 -770
rect 4945 -785 4965 -770
rect 5065 -785 5085 -770
rect 3200 -825 3235 -810
rect 2720 -850 2725 -825
rect 2750 -850 2755 -825
rect 2720 -860 2755 -850
rect 2950 -835 3005 -825
rect 790 -880 845 -870
rect 2950 -870 2960 -835
rect 2995 -870 3005 -835
rect 3200 -850 3205 -825
rect 3230 -850 3235 -825
rect 3200 -860 3235 -850
rect 3440 -825 3475 -810
rect 3440 -850 3445 -825
rect 3470 -850 3475 -825
rect 3440 -860 3475 -850
rect 3680 -825 3715 -810
rect 3680 -850 3685 -825
rect 3710 -850 3715 -825
rect 3680 -860 3715 -850
rect 3920 -825 3955 -810
rect 3920 -850 3925 -825
rect 3950 -850 3955 -825
rect 3920 -860 3955 -850
rect 4160 -825 4195 -810
rect 4160 -850 4165 -825
rect 4190 -850 4195 -825
rect 4160 -860 4195 -850
rect 4400 -825 4435 -810
rect 4400 -850 4405 -825
rect 4430 -850 4435 -825
rect 4400 -860 4435 -850
rect 4640 -825 4675 -810
rect 4640 -850 4645 -825
rect 4670 -850 4675 -825
rect 4640 -860 4675 -850
rect 4880 -825 4915 -810
rect 5125 -825 5150 -770
rect 5185 -785 5205 -770
rect 5305 -785 5325 -770
rect 5365 -810 5390 -770
rect 5425 -785 5445 -770
rect 5545 -785 5565 -770
rect 5605 -810 5630 -770
rect 5665 -785 5685 -770
rect 5785 -785 5805 -770
rect 5845 -810 5870 -770
rect 5905 -785 5925 -770
rect 6025 -785 6045 -770
rect 6085 -810 6110 -770
rect 6145 -785 6165 -770
rect 6265 -785 6285 -770
rect 6325 -810 6350 -770
rect 6385 -785 6405 -770
rect 6505 -785 6525 -770
rect 6565 -810 6590 -770
rect 6625 -785 6645 -770
rect 6745 -785 6765 -770
rect 6805 -810 6830 -770
rect 6865 -785 6885 -770
rect 6985 -785 7005 -770
rect 7045 -810 7070 -770
rect 7105 -785 7125 -770
rect 7225 -785 7245 -770
rect 5360 -825 5395 -810
rect 4880 -850 4885 -825
rect 4910 -850 4915 -825
rect 4880 -860 4915 -850
rect 5110 -835 5165 -825
rect 2950 -880 3005 -870
rect 5110 -870 5120 -835
rect 5155 -870 5165 -835
rect 5360 -850 5365 -825
rect 5390 -850 5395 -825
rect 5360 -860 5395 -850
rect 5600 -825 5635 -810
rect 5600 -850 5605 -825
rect 5630 -850 5635 -825
rect 5600 -860 5635 -850
rect 5840 -825 5875 -810
rect 5840 -850 5845 -825
rect 5870 -850 5875 -825
rect 5840 -860 5875 -850
rect 6080 -825 6115 -810
rect 6080 -850 6085 -825
rect 6110 -850 6115 -825
rect 6080 -860 6115 -850
rect 6320 -825 6355 -810
rect 6320 -850 6325 -825
rect 6350 -850 6355 -825
rect 6320 -860 6355 -850
rect 6560 -825 6595 -810
rect 6560 -850 6565 -825
rect 6590 -850 6595 -825
rect 6560 -860 6595 -850
rect 6800 -825 6835 -810
rect 6800 -850 6805 -825
rect 6830 -850 6835 -825
rect 6800 -860 6835 -850
rect 7040 -825 7075 -810
rect 7285 -825 7310 -770
rect 7345 -785 7365 -770
rect 7465 -785 7485 -770
rect 7525 -810 7550 -770
rect 7585 -785 7605 -770
rect 7705 -785 7725 -770
rect 7765 -810 7790 -770
rect 7825 -785 7845 -770
rect 7945 -785 7965 -770
rect 8005 -810 8030 -770
rect 8065 -785 8085 -770
rect 8185 -785 8205 -770
rect 8245 -810 8270 -770
rect 8305 -785 8325 -770
rect 8425 -785 8445 -770
rect 8485 -810 8510 -770
rect 8545 -785 8565 -770
rect 8665 -785 8685 -770
rect 8725 -810 8750 -770
rect 8785 -785 8805 -770
rect 8905 -785 8925 -770
rect 8965 -810 8990 -770
rect 9025 -785 9045 -770
rect 9145 -785 9165 -770
rect 9205 -810 9230 -770
rect 9265 -785 9285 -770
rect 9385 -785 9405 -770
rect 7520 -825 7555 -810
rect 7040 -850 7045 -825
rect 7070 -850 7075 -825
rect 7040 -860 7075 -850
rect 7270 -835 7325 -825
rect 5110 -880 5165 -870
rect 7270 -870 7280 -835
rect 7315 -870 7325 -835
rect 7520 -850 7525 -825
rect 7550 -850 7555 -825
rect 7520 -860 7555 -850
rect 7760 -825 7795 -810
rect 7760 -850 7765 -825
rect 7790 -850 7795 -825
rect 7760 -860 7795 -850
rect 8000 -825 8035 -810
rect 8000 -850 8005 -825
rect 8030 -850 8035 -825
rect 8000 -860 8035 -850
rect 8240 -825 8275 -810
rect 8240 -850 8245 -825
rect 8270 -850 8275 -825
rect 8240 -860 8275 -850
rect 8480 -825 8515 -810
rect 8480 -850 8485 -825
rect 8510 -850 8515 -825
rect 8480 -860 8515 -850
rect 8720 -825 8755 -810
rect 8720 -850 8725 -825
rect 8750 -850 8755 -825
rect 8720 -860 8755 -850
rect 8960 -825 8995 -810
rect 8960 -850 8965 -825
rect 8990 -850 8995 -825
rect 8960 -860 8995 -850
rect 9200 -825 9235 -810
rect 9445 -825 9470 -770
rect 9505 -785 9525 -770
rect 9625 -785 9645 -770
rect 9685 -810 9710 -770
rect 9745 -785 9765 -770
rect 9865 -785 9885 -770
rect 9925 -810 9950 -770
rect 9985 -785 10005 -770
rect 10105 -785 10125 -770
rect 10165 -810 10190 -770
rect 10225 -785 10245 -770
rect 10345 -785 10365 -770
rect 10405 -810 10430 -770
rect 10465 -785 10485 -770
rect 10585 -785 10605 -770
rect 10645 -810 10670 -770
rect 10705 -785 10725 -770
rect 10825 -785 10845 -770
rect 10885 -810 10910 -770
rect 10945 -785 10965 -770
rect 11065 -785 11085 -770
rect 11125 -810 11150 -770
rect 11185 -785 11205 -770
rect 11305 -785 11325 -770
rect 11365 -810 11390 -770
rect 11425 -785 11445 -770
rect 11545 -785 11565 -770
rect 9680 -825 9715 -810
rect 9200 -850 9205 -825
rect 9230 -850 9235 -825
rect 9200 -860 9235 -850
rect 9430 -835 9485 -825
rect 7270 -880 7325 -870
rect 9430 -870 9440 -835
rect 9475 -870 9485 -835
rect 9680 -850 9685 -825
rect 9710 -850 9715 -825
rect 9680 -860 9715 -850
rect 9920 -825 9955 -810
rect 9920 -850 9925 -825
rect 9950 -850 9955 -825
rect 9920 -860 9955 -850
rect 10160 -825 10195 -810
rect 10160 -850 10165 -825
rect 10190 -850 10195 -825
rect 10160 -860 10195 -850
rect 10400 -825 10435 -810
rect 10400 -850 10405 -825
rect 10430 -850 10435 -825
rect 10400 -860 10435 -850
rect 10640 -825 10675 -810
rect 10640 -850 10645 -825
rect 10670 -850 10675 -825
rect 10640 -860 10675 -850
rect 10880 -825 10915 -810
rect 10880 -850 10885 -825
rect 10910 -850 10915 -825
rect 10880 -860 10915 -850
rect 11120 -825 11155 -810
rect 11120 -850 11125 -825
rect 11150 -850 11155 -825
rect 11120 -860 11155 -850
rect 11360 -825 11395 -810
rect 11605 -825 11630 -770
rect 11665 -785 11685 -770
rect 11785 -785 11805 -770
rect 11845 -810 11870 -770
rect 11905 -785 11925 -770
rect 12025 -785 12045 -770
rect 12085 -810 12110 -770
rect 12145 -785 12165 -770
rect 12265 -785 12285 -770
rect 12325 -810 12350 -770
rect 12385 -785 12405 -770
rect 12505 -785 12525 -770
rect 12565 -810 12590 -770
rect 12625 -785 12645 -770
rect 12745 -785 12765 -770
rect 12805 -810 12830 -770
rect 12865 -785 12885 -770
rect 12985 -785 13005 -770
rect 13045 -810 13070 -770
rect 13105 -785 13125 -770
rect 13225 -785 13245 -770
rect 13285 -810 13310 -770
rect 13345 -785 13365 -770
rect 13465 -785 13485 -770
rect 13525 -810 13550 -770
rect 13585 -785 13605 -770
rect 13705 -785 13725 -770
rect 11840 -825 11875 -810
rect 11360 -850 11365 -825
rect 11390 -850 11395 -825
rect 11360 -860 11395 -850
rect 11590 -835 11645 -825
rect 9430 -880 9485 -870
rect 11590 -870 11600 -835
rect 11635 -870 11645 -835
rect 11840 -850 11845 -825
rect 11870 -850 11875 -825
rect 11840 -860 11875 -850
rect 12080 -825 12115 -810
rect 12080 -850 12085 -825
rect 12110 -850 12115 -825
rect 12080 -860 12115 -850
rect 12320 -825 12355 -810
rect 12320 -850 12325 -825
rect 12350 -850 12355 -825
rect 12320 -860 12355 -850
rect 12560 -825 12595 -810
rect 12560 -850 12565 -825
rect 12590 -850 12595 -825
rect 12560 -860 12595 -850
rect 12800 -825 12835 -810
rect 12800 -850 12805 -825
rect 12830 -850 12835 -825
rect 12800 -860 12835 -850
rect 13040 -825 13075 -810
rect 13040 -850 13045 -825
rect 13070 -850 13075 -825
rect 13040 -860 13075 -850
rect 13280 -825 13315 -810
rect 13280 -850 13285 -825
rect 13310 -850 13315 -825
rect 13280 -860 13315 -850
rect 13520 -825 13555 -810
rect 13765 -825 13790 -770
rect 13825 -785 13845 -770
rect 13945 -785 13965 -770
rect 14005 -810 14030 -770
rect 14065 -785 14085 -770
rect 14185 -785 14205 -770
rect 14245 -810 14270 -770
rect 14305 -785 14325 -770
rect 14425 -785 14445 -770
rect 14485 -810 14510 -770
rect 14545 -785 14565 -770
rect 14665 -785 14685 -770
rect 14725 -810 14750 -770
rect 14785 -785 14805 -770
rect 14905 -785 14925 -770
rect 14965 -810 14990 -770
rect 15025 -785 15045 -770
rect 15145 -785 15165 -770
rect 15205 -810 15230 -770
rect 15265 -785 15285 -770
rect 15385 -785 15405 -770
rect 15445 -810 15470 -770
rect 15505 -785 15525 -770
rect 15625 -785 15645 -770
rect 15685 -810 15710 -770
rect 15745 -785 15765 -770
rect 15865 -785 15885 -770
rect 14000 -825 14035 -810
rect 13520 -850 13525 -825
rect 13550 -850 13555 -825
rect 13520 -860 13555 -850
rect 13750 -835 13805 -825
rect 11590 -880 11645 -870
rect 13750 -870 13760 -835
rect 13795 -870 13805 -835
rect 14000 -850 14005 -825
rect 14030 -850 14035 -825
rect 14000 -860 14035 -850
rect 14240 -825 14275 -810
rect 14240 -850 14245 -825
rect 14270 -850 14275 -825
rect 14240 -860 14275 -850
rect 14480 -825 14515 -810
rect 14480 -850 14485 -825
rect 14510 -850 14515 -825
rect 14480 -860 14515 -850
rect 14720 -825 14755 -810
rect 14720 -850 14725 -825
rect 14750 -850 14755 -825
rect 14720 -860 14755 -850
rect 14960 -825 14995 -810
rect 14960 -850 14965 -825
rect 14990 -850 14995 -825
rect 14960 -860 14995 -850
rect 15200 -825 15235 -810
rect 15200 -850 15205 -825
rect 15230 -850 15235 -825
rect 15200 -860 15235 -850
rect 15440 -825 15475 -810
rect 15440 -850 15445 -825
rect 15470 -850 15475 -825
rect 15440 -860 15475 -850
rect 15680 -825 15715 -810
rect 15925 -825 15950 -770
rect 15985 -785 16005 -770
rect 16105 -785 16125 -770
rect 16165 -810 16190 -770
rect 16225 -785 16245 -770
rect 16345 -785 16365 -770
rect 16405 -810 16430 -770
rect 16465 -785 16485 -770
rect 16585 -785 16605 -770
rect 16645 -810 16670 -770
rect 16705 -785 16725 -770
rect 16825 -785 16845 -770
rect 16885 -810 16910 -770
rect 16945 -785 16965 -770
rect 17065 -785 17085 -770
rect 17125 -810 17150 -770
rect 17185 -785 17205 -770
rect 17305 -785 17325 -770
rect 17365 -810 17390 -770
rect 17425 -785 17445 -770
rect 17545 -785 17565 -770
rect 17605 -810 17630 -770
rect 17665 -785 17685 -770
rect 17785 -785 17805 -770
rect 17845 -810 17870 -770
rect 17905 -785 17925 -770
rect 18025 -785 18045 -770
rect 16160 -825 16195 -810
rect 15680 -850 15685 -825
rect 15710 -850 15715 -825
rect 15680 -860 15715 -850
rect 15910 -835 15965 -825
rect 13750 -880 13805 -870
rect 15910 -870 15920 -835
rect 15955 -870 15965 -835
rect 16160 -850 16165 -825
rect 16190 -850 16195 -825
rect 16160 -860 16195 -850
rect 16400 -825 16435 -810
rect 16400 -850 16405 -825
rect 16430 -850 16435 -825
rect 16400 -860 16435 -850
rect 16640 -825 16675 -810
rect 16640 -850 16645 -825
rect 16670 -850 16675 -825
rect 16640 -860 16675 -850
rect 16880 -825 16915 -810
rect 16880 -850 16885 -825
rect 16910 -850 16915 -825
rect 16880 -860 16915 -850
rect 17120 -825 17155 -810
rect 17120 -850 17125 -825
rect 17150 -850 17155 -825
rect 17120 -860 17155 -850
rect 17360 -825 17395 -810
rect 17360 -850 17365 -825
rect 17390 -850 17395 -825
rect 17360 -860 17395 -850
rect 17600 -825 17635 -810
rect 17600 -850 17605 -825
rect 17630 -850 17635 -825
rect 17600 -860 17635 -850
rect 17840 -825 17875 -810
rect 18085 -825 18110 -770
rect 18145 -785 18165 -770
rect 18265 -785 18285 -770
rect 18325 -810 18350 -770
rect 18385 -785 18405 -770
rect 18505 -785 18525 -770
rect 18565 -810 18590 -770
rect 18625 -785 18645 -770
rect 18745 -785 18765 -770
rect 18805 -810 18830 -770
rect 18865 -785 18885 -770
rect 18985 -785 19005 -770
rect 19045 -810 19070 -770
rect 19105 -785 19125 -770
rect 19225 -785 19245 -770
rect 19285 -810 19310 -770
rect 19345 -785 19365 -770
rect 19465 -785 19485 -770
rect 19525 -810 19550 -770
rect 19585 -785 19605 -770
rect 19705 -785 19725 -770
rect 19765 -810 19790 -770
rect 19825 -785 19845 -770
rect 19945 -785 19965 -770
rect 20005 -810 20030 -770
rect 20065 -785 20085 -770
rect 20185 -785 20205 -770
rect 18320 -825 18355 -810
rect 17840 -850 17845 -825
rect 17870 -850 17875 -825
rect 17840 -860 17875 -850
rect 18070 -835 18125 -825
rect 15910 -880 15965 -870
rect 18070 -870 18080 -835
rect 18115 -870 18125 -835
rect 18320 -850 18325 -825
rect 18350 -850 18355 -825
rect 18320 -860 18355 -850
rect 18560 -825 18595 -810
rect 18560 -850 18565 -825
rect 18590 -850 18595 -825
rect 18560 -860 18595 -850
rect 18800 -825 18835 -810
rect 18800 -850 18805 -825
rect 18830 -850 18835 -825
rect 18800 -860 18835 -850
rect 19040 -825 19075 -810
rect 19040 -850 19045 -825
rect 19070 -850 19075 -825
rect 19040 -860 19075 -850
rect 19280 -825 19315 -810
rect 19280 -850 19285 -825
rect 19310 -850 19315 -825
rect 19280 -860 19315 -850
rect 19520 -825 19555 -810
rect 19520 -850 19525 -825
rect 19550 -850 19555 -825
rect 19520 -860 19555 -850
rect 19760 -825 19795 -810
rect 19760 -850 19765 -825
rect 19790 -850 19795 -825
rect 19760 -860 19795 -850
rect 20000 -825 20035 -810
rect 20245 -825 20270 -770
rect 20305 -785 20325 -770
rect 20425 -785 20445 -770
rect 20485 -810 20510 -770
rect 20545 -785 20565 -770
rect 20665 -785 20685 -770
rect 20725 -810 20750 -770
rect 20785 -785 20805 -770
rect 20905 -785 20925 -770
rect 20965 -810 20990 -770
rect 21025 -785 21045 -770
rect 21145 -785 21165 -770
rect 21205 -810 21230 -770
rect 21265 -785 21285 -770
rect 21385 -785 21405 -770
rect 21445 -810 21470 -770
rect 21505 -785 21525 -770
rect 21625 -785 21645 -770
rect 21685 -810 21710 -770
rect 21745 -785 21765 -770
rect 21865 -785 21885 -770
rect 21925 -810 21950 -770
rect 21985 -785 22005 -770
rect 22105 -785 22125 -770
rect 22165 -810 22190 -770
rect 22225 -785 22245 -770
rect 22345 -785 22365 -770
rect 20480 -825 20515 -810
rect 20000 -850 20005 -825
rect 20030 -850 20035 -825
rect 20000 -860 20035 -850
rect 20230 -835 20285 -825
rect 18070 -880 18125 -870
rect 20230 -870 20240 -835
rect 20275 -870 20285 -835
rect 20480 -850 20485 -825
rect 20510 -850 20515 -825
rect 20480 -860 20515 -850
rect 20720 -825 20755 -810
rect 20720 -850 20725 -825
rect 20750 -850 20755 -825
rect 20720 -860 20755 -850
rect 20960 -825 20995 -810
rect 20960 -850 20965 -825
rect 20990 -850 20995 -825
rect 20960 -860 20995 -850
rect 21200 -825 21235 -810
rect 21200 -850 21205 -825
rect 21230 -850 21235 -825
rect 21200 -860 21235 -850
rect 21440 -825 21475 -810
rect 21440 -850 21445 -825
rect 21470 -850 21475 -825
rect 21440 -860 21475 -850
rect 21680 -825 21715 -810
rect 21680 -850 21685 -825
rect 21710 -850 21715 -825
rect 21680 -860 21715 -850
rect 21920 -825 21955 -810
rect 21920 -850 21925 -825
rect 21950 -850 21955 -825
rect 21920 -860 21955 -850
rect 22160 -825 22195 -810
rect 22405 -825 22430 -770
rect 22465 -785 22485 -770
rect 22585 -785 22605 -770
rect 22645 -810 22670 -770
rect 22705 -785 22725 -770
rect 22825 -785 22845 -770
rect 22885 -810 22910 -770
rect 22945 -785 22965 -770
rect 23065 -785 23085 -770
rect 23125 -810 23150 -770
rect 23185 -785 23205 -770
rect 23305 -785 23325 -770
rect 23365 -810 23390 -770
rect 23425 -785 23445 -770
rect 23545 -785 23565 -770
rect 23605 -810 23630 -770
rect 23665 -785 23685 -770
rect 23785 -785 23805 -770
rect 23845 -810 23870 -770
rect 23905 -785 23925 -770
rect 24025 -785 24045 -770
rect 24085 -810 24110 -770
rect 24145 -785 24165 -770
rect 24265 -785 24285 -770
rect 22640 -825 22675 -810
rect 22160 -850 22165 -825
rect 22190 -850 22195 -825
rect 22160 -860 22195 -850
rect 22390 -835 22445 -825
rect 20230 -880 20285 -870
rect 22390 -870 22400 -835
rect 22435 -870 22445 -835
rect 22640 -850 22645 -825
rect 22670 -850 22675 -825
rect 22640 -860 22675 -850
rect 22880 -825 22915 -810
rect 22880 -850 22885 -825
rect 22910 -850 22915 -825
rect 22880 -860 22915 -850
rect 23120 -825 23155 -810
rect 23120 -850 23125 -825
rect 23150 -850 23155 -825
rect 23120 -860 23155 -850
rect 23360 -825 23395 -810
rect 23360 -850 23365 -825
rect 23390 -850 23395 -825
rect 23360 -860 23395 -850
rect 23600 -825 23635 -810
rect 23600 -850 23605 -825
rect 23630 -850 23635 -825
rect 23600 -860 23635 -850
rect 23840 -825 23875 -810
rect 23840 -850 23845 -825
rect 23870 -850 23875 -825
rect 23840 -860 23875 -850
rect 24080 -825 24115 -810
rect 24325 -825 24350 -770
rect 24385 -785 24405 -770
rect 24505 -785 24525 -770
rect 24565 -810 24590 -770
rect 24625 -785 24645 -770
rect 24745 -785 24765 -770
rect 24805 -810 24830 -770
rect 24865 -785 24885 -770
rect 24985 -785 25005 -770
rect 25045 -810 25070 -770
rect 25105 -785 25125 -770
rect 25225 -785 25245 -770
rect 25285 -810 25310 -770
rect 25345 -785 25365 -770
rect 25465 -785 25485 -770
rect 25525 -810 25550 -770
rect 25585 -785 25605 -770
rect 25705 -785 25725 -770
rect 25765 -810 25790 -770
rect 25825 -785 25845 -770
rect 25945 -785 25965 -770
rect 26005 -810 26030 -770
rect 26065 -785 26085 -770
rect 26185 -785 26205 -770
rect 24560 -825 24595 -810
rect 24080 -850 24085 -825
rect 24110 -850 24115 -825
rect 24080 -860 24115 -850
rect 24310 -835 24365 -825
rect 22390 -880 22445 -870
rect 24310 -870 24320 -835
rect 24355 -870 24365 -835
rect 24560 -850 24565 -825
rect 24590 -850 24595 -825
rect 24560 -860 24595 -850
rect 24800 -825 24835 -810
rect 24800 -850 24805 -825
rect 24830 -850 24835 -825
rect 24800 -860 24835 -850
rect 25040 -825 25075 -810
rect 25040 -850 25045 -825
rect 25070 -850 25075 -825
rect 25040 -860 25075 -850
rect 25280 -825 25315 -810
rect 25280 -850 25285 -825
rect 25310 -850 25315 -825
rect 25280 -860 25315 -850
rect 25520 -825 25555 -810
rect 25520 -850 25525 -825
rect 25550 -850 25555 -825
rect 25520 -860 25555 -850
rect 25760 -825 25795 -810
rect 25760 -850 25765 -825
rect 25790 -850 25795 -825
rect 25760 -860 25795 -850
rect 26000 -825 26035 -810
rect 26245 -825 26270 -770
rect 26305 -785 26325 -770
rect 26425 -785 26445 -770
rect 26485 -810 26510 -770
rect 26545 -785 26565 -770
rect 26665 -785 26685 -770
rect 26725 -810 26750 -770
rect 26785 -785 26805 -770
rect 26905 -785 26925 -770
rect 26965 -810 26990 -770
rect 27025 -785 27045 -770
rect 27145 -785 27165 -770
rect 27205 -810 27230 -770
rect 27265 -785 27285 -770
rect 27385 -785 27405 -770
rect 27445 -810 27470 -770
rect 27505 -785 27525 -770
rect 27625 -785 27645 -770
rect 27685 -810 27710 -770
rect 27745 -785 27765 -770
rect 27865 -785 27885 -770
rect 27925 -810 27950 -770
rect 27985 -785 28005 -770
rect 28105 -785 28125 -770
rect 26480 -825 26515 -810
rect 26000 -850 26005 -825
rect 26030 -850 26035 -825
rect 26000 -860 26035 -850
rect 26230 -835 26285 -825
rect 24310 -880 24365 -870
rect 26230 -870 26240 -835
rect 26275 -870 26285 -835
rect 26480 -850 26485 -825
rect 26510 -850 26515 -825
rect 26480 -860 26515 -850
rect 26720 -825 26755 -810
rect 26720 -850 26725 -825
rect 26750 -850 26755 -825
rect 26720 -860 26755 -850
rect 26960 -825 26995 -810
rect 26960 -850 26965 -825
rect 26990 -850 26995 -825
rect 26960 -860 26995 -850
rect 27200 -825 27235 -810
rect 27200 -850 27205 -825
rect 27230 -850 27235 -825
rect 27200 -860 27235 -850
rect 27440 -825 27475 -810
rect 27440 -850 27445 -825
rect 27470 -850 27475 -825
rect 27440 -860 27475 -850
rect 27680 -825 27715 -810
rect 27680 -850 27685 -825
rect 27710 -850 27715 -825
rect 27680 -860 27715 -850
rect 27920 -825 27955 -810
rect 28165 -825 28190 -770
rect 28225 -785 28245 -770
rect 28345 -785 28365 -770
rect 28405 -810 28430 -770
rect 28465 -785 28485 -770
rect 28585 -785 28605 -770
rect 28645 -810 28670 -770
rect 28705 -785 28725 -770
rect 28825 -785 28845 -770
rect 28885 -810 28910 -770
rect 28945 -785 28965 -770
rect 29065 -785 29085 -770
rect 29125 -810 29150 -770
rect 29185 -785 29205 -770
rect 29305 -785 29325 -770
rect 29365 -810 29390 -770
rect 29425 -785 29445 -770
rect 29545 -785 29565 -770
rect 29605 -810 29630 -770
rect 29665 -785 29685 -770
rect 29785 -785 29805 -770
rect 28400 -825 28435 -810
rect 27920 -850 27925 -825
rect 27950 -850 27955 -825
rect 27920 -860 27955 -850
rect 28150 -835 28205 -825
rect 26230 -880 26285 -870
rect 28150 -870 28160 -835
rect 28195 -870 28205 -835
rect 28400 -850 28405 -825
rect 28430 -850 28435 -825
rect 28400 -860 28435 -850
rect 28640 -825 28675 -810
rect 28640 -850 28645 -825
rect 28670 -850 28675 -825
rect 28640 -860 28675 -850
rect 28880 -825 28915 -810
rect 28880 -850 28885 -825
rect 28910 -850 28915 -825
rect 28880 -860 28915 -850
rect 29120 -825 29155 -810
rect 29120 -850 29125 -825
rect 29150 -850 29155 -825
rect 29120 -860 29155 -850
rect 29360 -825 29395 -810
rect 29360 -850 29365 -825
rect 29390 -850 29395 -825
rect 29360 -860 29395 -850
rect 29600 -825 29635 -810
rect 29845 -825 29870 -770
rect 29905 -785 29925 -770
rect 30025 -785 30045 -770
rect 30085 -810 30110 -770
rect 30145 -785 30165 -770
rect 30265 -785 30285 -770
rect 30325 -810 30350 -770
rect 30385 -785 30405 -770
rect 30505 -785 30525 -770
rect 30565 -810 30590 -770
rect 30625 -785 30645 -770
rect 30080 -825 30115 -810
rect 29600 -850 29605 -825
rect 29630 -850 29635 -825
rect 29600 -860 29635 -850
rect 29830 -835 29885 -825
rect 28150 -880 28205 -870
rect 29830 -870 29840 -835
rect 29875 -870 29885 -835
rect 30080 -850 30085 -825
rect 30110 -850 30115 -825
rect 30080 -860 30115 -850
rect 30320 -825 30355 -810
rect 30320 -850 30325 -825
rect 30350 -850 30355 -825
rect 30320 -860 30355 -850
rect 30560 -825 30595 -810
rect 30560 -850 30565 -825
rect 30590 -850 30595 -825
rect 30560 -860 30595 -850
rect 29830 -880 29885 -870
rect 31060 -870 31080 -770
rect 31180 -870 31200 -770
rect 31060 -945 31200 -870
rect -460 -965 31200 -945
rect -460 -1065 -275 -965
rect -175 -1065 275 -965
rect 375 -1065 825 -965
rect 925 -1065 1375 -965
rect 1475 -1065 1925 -965
rect 2025 -1065 2475 -965
rect 2575 -1065 3025 -965
rect 3125 -1065 3575 -965
rect 3675 -1065 4125 -965
rect 4225 -1065 4675 -965
rect 4775 -1065 5225 -965
rect 5325 -1065 5775 -965
rect 5875 -1065 6325 -965
rect 6425 -1065 6875 -965
rect 6975 -1065 7425 -965
rect 7525 -1065 7975 -965
rect 8075 -1065 8525 -965
rect 8625 -1065 9075 -965
rect 9175 -1065 9625 -965
rect 9725 -1065 10175 -965
rect 10275 -1065 10725 -965
rect 10825 -1065 11275 -965
rect 11375 -1065 11825 -965
rect 11925 -1065 12375 -965
rect 12475 -1065 12925 -965
rect 13025 -1065 13475 -965
rect 13575 -1065 14025 -965
rect 14125 -1065 14575 -965
rect 14675 -1065 15125 -965
rect 15225 -1065 15675 -965
rect 15775 -1065 16225 -965
rect 16325 -1065 16775 -965
rect 16875 -1065 17325 -965
rect 17425 -1065 17875 -965
rect 17975 -1065 18425 -965
rect 18525 -1065 18975 -965
rect 19075 -1065 19525 -965
rect 19625 -1065 20075 -965
rect 20175 -1065 20625 -965
rect 20725 -1065 21175 -965
rect 21275 -1065 22065 -965
rect 22165 -1065 22615 -965
rect 22715 -1065 23165 -965
rect 23265 -1065 23715 -965
rect 23815 -1065 24265 -965
rect 24365 -1065 24815 -965
rect 24915 -1065 25365 -965
rect 25465 -1065 25915 -965
rect 26015 -1065 26465 -965
rect 26565 -1065 27015 -965
rect 27115 -1065 27565 -965
rect 27665 -1065 28115 -965
rect 28215 -1065 28665 -965
rect 28765 -1065 29215 -965
rect 29315 -1065 29765 -965
rect 29865 -1065 30315 -965
rect 30415 -1065 30865 -965
rect 30965 -1065 31200 -965
rect -460 -1085 31200 -1065
<< viali >>
rect 195 240 230 275
rect 441 240 461 260
rect 746 240 766 260
rect 991 240 1011 260
rect 1231 240 1251 260
rect 1476 240 1496 260
rect 1781 240 1801 260
rect 2026 240 2046 260
rect 2265 270 2300 305
rect 2511 240 2531 260
rect 2751 240 2771 260
rect 2996 240 3016 260
rect 3236 240 3256 260
rect 3481 240 3501 260
rect 3721 240 3741 260
rect 3966 240 3986 260
rect 4205 270 4240 305
rect 386 200 406 220
rect 506 200 526 220
rect 691 200 711 220
rect 811 200 831 220
rect 936 200 956 220
rect 1056 200 1076 220
rect 1176 200 1196 220
rect 1296 200 1316 220
rect 1421 200 1441 220
rect 1541 200 1561 220
rect 1726 200 1746 220
rect 1846 200 1866 220
rect 1971 200 1991 220
rect 2091 200 2111 220
rect 2211 200 2231 220
rect 2331 200 2351 220
rect 2456 200 2476 220
rect 2576 200 2596 220
rect 2696 200 2716 220
rect 2816 200 2836 220
rect 2941 200 2961 220
rect 3061 200 3081 220
rect 3181 200 3201 220
rect 3301 200 3321 220
rect 3426 200 3446 220
rect 3546 200 3566 220
rect 3666 200 3686 220
rect 3786 200 3806 220
rect 3911 200 3931 220
rect 4451 240 4471 260
rect 4691 240 4711 260
rect 4936 240 4956 260
rect 5176 240 5196 260
rect 5421 240 5441 260
rect 5726 240 5746 260
rect 5971 240 5991 260
rect 6211 240 6231 260
rect 6455 270 6490 305
rect 6696 240 6716 260
rect 6941 240 6961 260
rect 7181 240 7201 260
rect 7421 240 7441 260
rect 7661 240 7681 260
rect 7906 240 7926 260
rect 8146 240 8166 260
rect 8391 240 8411 260
rect 8631 240 8651 260
rect 8876 240 8896 260
rect 9116 240 9136 260
rect 9360 270 9395 305
rect 4031 200 4051 220
rect 4151 200 4171 220
rect 4271 200 4291 220
rect 4396 200 4416 220
rect 4516 200 4536 220
rect 4636 200 4656 220
rect 4756 200 4776 220
rect 4881 200 4901 220
rect 5001 200 5021 220
rect 5121 200 5141 220
rect 5241 200 5261 220
rect 5366 200 5386 220
rect 5486 200 5506 220
rect 5671 200 5691 220
rect 5791 200 5811 220
rect 5916 200 5936 220
rect 6036 200 6056 220
rect 6156 200 6176 220
rect 6276 200 6296 220
rect 6401 200 6421 220
rect 6521 200 6541 220
rect 6641 200 6661 220
rect 6761 200 6781 220
rect 6886 200 6906 220
rect 7006 200 7026 220
rect 7126 200 7146 220
rect 7246 200 7266 220
rect 7366 200 7386 220
rect 7486 200 7506 220
rect 7606 200 7626 220
rect 7726 200 7746 220
rect 7851 200 7871 220
rect 7971 200 7991 220
rect 8091 200 8111 220
rect 8211 200 8231 220
rect 8336 200 8356 220
rect 8456 200 8476 220
rect 8576 200 8596 220
rect 8696 200 8716 220
rect 8821 200 8841 220
rect 8941 200 8961 220
rect 9061 200 9081 220
rect 9606 240 9626 260
rect 9851 240 9871 260
rect 10091 240 10111 260
rect 10336 240 10356 260
rect 10576 240 10596 260
rect 10821 240 10841 260
rect 11061 240 11081 260
rect 11305 270 11340 305
rect 11546 240 11566 260
rect 11791 240 11811 260
rect 12031 240 12051 260
rect 12276 240 12296 260
rect 12516 240 12536 260
rect 12761 240 12781 260
rect 13000 270 13035 305
rect 13246 240 13266 260
rect 13486 240 13506 260
rect 13731 240 13751 260
rect 13971 240 13991 260
rect 14216 240 14236 260
rect 14456 240 14476 260
rect 14701 240 14721 260
rect 14941 240 14961 260
rect 15185 270 15220 305
rect 15426 240 15446 260
rect 15671 240 15691 260
rect 15911 240 15931 260
rect 16156 240 16176 260
rect 16396 240 16416 260
rect 16641 240 16661 260
rect 16881 240 16901 260
rect 17126 240 17146 260
rect 17365 270 17400 305
rect 17611 240 17631 260
rect 17851 240 17871 260
rect 18096 240 18116 260
rect 18336 240 18356 260
rect 18581 240 18601 260
rect 18821 240 18841 260
rect 19066 240 19086 260
rect 19306 240 19326 260
rect 19550 270 19585 305
rect 19791 240 19811 260
rect 20036 240 20056 260
rect 20276 240 20296 260
rect 20521 240 20541 260
rect 20760 270 20795 305
rect 21006 240 21026 260
rect 9181 200 9201 220
rect 9306 200 9326 220
rect 9426 200 9446 220
rect 9551 200 9571 220
rect 9671 200 9691 220
rect 9796 200 9816 220
rect 9916 200 9936 220
rect 10036 200 10056 220
rect 10156 200 10176 220
rect 10281 200 10301 220
rect 10401 200 10421 220
rect 10521 200 10541 220
rect 10641 200 10661 220
rect 10766 200 10786 220
rect 10886 200 10906 220
rect 11006 200 11026 220
rect 11126 200 11146 220
rect 11251 200 11271 220
rect 11371 200 11391 220
rect 11491 200 11511 220
rect 11611 200 11631 220
rect 11736 200 11756 220
rect 11856 200 11876 220
rect 11976 200 11996 220
rect 12096 200 12116 220
rect 12221 200 12241 220
rect 12341 200 12361 220
rect 12461 200 12481 220
rect 12581 200 12601 220
rect 12706 200 12726 220
rect 12826 200 12846 220
rect 12946 200 12966 220
rect 13066 200 13086 220
rect 13191 200 13211 220
rect 13311 200 13331 220
rect 13431 200 13451 220
rect 13551 200 13571 220
rect 13676 200 13696 220
rect 13796 200 13816 220
rect 13916 200 13936 220
rect 14036 200 14056 220
rect 14161 200 14181 220
rect 14281 200 14301 220
rect 14401 200 14421 220
rect 14521 200 14541 220
rect 14646 200 14666 220
rect 14766 200 14786 220
rect 14886 200 14906 220
rect 15006 200 15026 220
rect 15131 200 15151 220
rect 15251 200 15271 220
rect 15371 200 15391 220
rect 15491 200 15511 220
rect 15616 200 15636 220
rect 15736 200 15756 220
rect 15856 200 15876 220
rect 15976 200 15996 220
rect 16101 200 16121 220
rect 16221 200 16241 220
rect 16341 200 16361 220
rect 16461 200 16481 220
rect 16586 200 16606 220
rect 16706 200 16726 220
rect 16826 200 16846 220
rect 16946 200 16966 220
rect 17071 200 17091 220
rect 17191 200 17211 220
rect 17311 200 17331 220
rect 17431 200 17451 220
rect 17556 200 17576 220
rect 17676 200 17696 220
rect 17796 200 17816 220
rect 17916 200 17936 220
rect 18041 200 18061 220
rect 18161 200 18181 220
rect 18281 200 18301 220
rect 18401 200 18421 220
rect 18526 200 18546 220
rect 18646 200 18666 220
rect 18766 200 18786 220
rect 18886 200 18906 220
rect 19011 200 19031 220
rect 19131 200 19151 220
rect 19251 200 19271 220
rect 19371 200 19391 220
rect 19496 200 19516 220
rect 19616 200 19636 220
rect 19736 200 19756 220
rect 19856 200 19876 220
rect 19981 200 20001 220
rect 20101 200 20121 220
rect 20221 200 20241 220
rect 20341 200 20361 220
rect 20466 200 20486 220
rect 20586 200 20606 220
rect 20706 200 20726 220
rect 20826 200 20846 220
rect 20951 200 20971 220
rect 21071 200 21091 220
rect 326 55 346 75
rect 441 55 461 75
rect 561 55 581 75
rect 631 55 651 75
rect 746 55 766 75
rect 876 55 896 75
rect 991 55 1011 75
rect 1116 55 1136 75
rect 1231 55 1251 75
rect 1361 55 1381 75
rect 1476 55 1496 75
rect 326 -65 346 -45
rect 446 -70 466 -50
rect 1596 55 1616 75
rect 1666 55 1686 75
rect 1781 55 1801 75
rect 1911 55 1931 75
rect 2026 55 2046 75
rect 2151 55 2171 75
rect 2266 55 2286 75
rect 2396 55 2416 75
rect 2511 55 2531 75
rect 2636 55 2656 75
rect 2751 55 2771 75
rect 2881 55 2901 75
rect 2996 55 3016 75
rect 3121 55 3141 75
rect 3236 55 3256 75
rect 3366 55 3386 75
rect 3481 55 3501 75
rect 3606 55 3626 75
rect 3721 55 3741 75
rect 3851 55 3871 75
rect 3966 55 3986 75
rect 4091 55 4111 75
rect 4206 55 4226 75
rect 4336 55 4356 75
rect 4451 55 4471 75
rect 4576 55 4596 75
rect 4691 55 4711 75
rect 4821 55 4841 75
rect 4936 55 4956 75
rect 5061 55 5081 75
rect 5176 55 5196 75
rect 5306 55 5326 75
rect 5421 55 5441 75
rect 561 -70 581 -50
rect 631 -65 651 -45
rect 751 -70 771 -50
rect 876 -65 896 -45
rect 996 -70 1016 -50
rect 1116 -65 1136 -45
rect 1236 -70 1256 -50
rect 1361 -65 1381 -45
rect 1481 -70 1501 -50
rect 5541 55 5561 75
rect 5611 55 5631 75
rect 5726 55 5746 75
rect 5856 55 5876 75
rect 5971 55 5991 75
rect 6096 55 6116 75
rect 6211 55 6231 75
rect 6341 55 6361 75
rect 6456 55 6476 75
rect 6581 55 6601 75
rect 6696 55 6716 75
rect 6826 55 6846 75
rect 6941 55 6961 75
rect 7066 55 7086 75
rect 7181 55 7201 75
rect 7306 55 7326 75
rect 7421 55 7441 75
rect 7546 55 7566 75
rect 7661 55 7681 75
rect 7791 55 7811 75
rect 7906 55 7926 75
rect 8031 55 8051 75
rect 8146 55 8166 75
rect 8276 55 8296 75
rect 8391 55 8411 75
rect 8516 55 8536 75
rect 8631 55 8651 75
rect 8761 55 8781 75
rect 8876 55 8896 75
rect 9001 55 9021 75
rect 9116 55 9136 75
rect 9246 55 9266 75
rect 9361 55 9381 75
rect 9491 55 9511 75
rect 9606 55 9626 75
rect 9736 55 9756 75
rect 9851 55 9871 75
rect 9976 55 9996 75
rect 10091 55 10111 75
rect 10221 55 10241 75
rect 10336 55 10356 75
rect 10461 55 10481 75
rect 10576 55 10596 75
rect 10706 55 10726 75
rect 10821 55 10841 75
rect 10946 55 10966 75
rect 11061 55 11081 75
rect 11191 55 11211 75
rect 11306 55 11326 75
rect 11431 55 11451 75
rect 11546 55 11566 75
rect 11676 55 11696 75
rect 11791 55 11811 75
rect 11916 55 11936 75
rect 12031 55 12051 75
rect 12161 55 12181 75
rect 12276 55 12296 75
rect 12401 55 12421 75
rect 12516 55 12536 75
rect 12646 55 12666 75
rect 12761 55 12781 75
rect 12886 55 12906 75
rect 13001 55 13021 75
rect 13131 55 13151 75
rect 13246 55 13266 75
rect 13371 55 13391 75
rect 13486 55 13506 75
rect 13616 55 13636 75
rect 13731 55 13751 75
rect 13856 55 13876 75
rect 13971 55 13991 75
rect 14101 55 14121 75
rect 14216 55 14236 75
rect 14341 55 14361 75
rect 14456 55 14476 75
rect 14586 55 14606 75
rect 14701 55 14721 75
rect 14826 55 14846 75
rect 14941 55 14961 75
rect 15071 55 15091 75
rect 15186 55 15206 75
rect 15311 55 15331 75
rect 15426 55 15446 75
rect 15556 55 15576 75
rect 15671 55 15691 75
rect 15796 55 15816 75
rect 15911 55 15931 75
rect 16041 55 16061 75
rect 16156 55 16176 75
rect 16281 55 16301 75
rect 16396 55 16416 75
rect 16526 55 16546 75
rect 16641 55 16661 75
rect 16766 55 16786 75
rect 16881 55 16901 75
rect 17011 55 17031 75
rect 17126 55 17146 75
rect 17251 55 17271 75
rect 17366 55 17386 75
rect 17496 55 17516 75
rect 17611 55 17631 75
rect 17736 55 17756 75
rect 17851 55 17871 75
rect 17981 55 18001 75
rect 18096 55 18116 75
rect 18221 55 18241 75
rect 18336 55 18356 75
rect 18466 55 18486 75
rect 18581 55 18601 75
rect 18706 55 18726 75
rect 18821 55 18841 75
rect 18951 55 18971 75
rect 19066 55 19086 75
rect 19191 55 19211 75
rect 19306 55 19326 75
rect 19436 55 19456 75
rect 19551 55 19571 75
rect 19676 55 19696 75
rect 19791 55 19811 75
rect 19921 55 19941 75
rect 20036 55 20056 75
rect 20161 55 20181 75
rect 20276 55 20296 75
rect 20406 55 20426 75
rect 20521 55 20541 75
rect 20646 55 20666 75
rect 20761 55 20781 75
rect 20891 55 20911 75
rect 21006 55 21026 75
rect 21126 55 21146 75
rect 1596 -70 1616 -50
rect 1666 -65 1686 -45
rect 1786 -70 1806 -50
rect 1911 -65 1931 -45
rect 2031 -70 2051 -50
rect 2151 -65 2171 -45
rect 2271 -70 2291 -50
rect 2396 -65 2416 -45
rect 2516 -70 2536 -50
rect 2636 -65 2656 -45
rect 2756 -70 2776 -50
rect 2881 -65 2901 -45
rect 3001 -70 3021 -50
rect 3121 -65 3141 -45
rect 3241 -70 3261 -50
rect 3366 -65 3386 -45
rect 3486 -70 3506 -50
rect 3606 -65 3626 -45
rect 3726 -70 3746 -50
rect 3851 -65 3871 -45
rect 3971 -70 3991 -50
rect 4091 -65 4111 -45
rect 4211 -70 4231 -50
rect 4336 -65 4356 -45
rect 4456 -70 4476 -50
rect 4576 -65 4596 -45
rect 4696 -70 4716 -50
rect 4821 -65 4841 -45
rect 4941 -70 4961 -50
rect 5061 -65 5081 -45
rect 5181 -70 5201 -50
rect 5306 -65 5326 -45
rect 5426 -70 5446 -50
rect 21160 -10 21180 10
rect 5541 -70 5561 -50
rect 5611 -65 5631 -45
rect 5731 -70 5751 -50
rect 5856 -65 5876 -45
rect 5976 -70 5996 -50
rect 6096 -65 6116 -45
rect 6216 -70 6236 -50
rect 6341 -65 6361 -45
rect 6461 -70 6481 -50
rect 6581 -65 6601 -45
rect 6701 -70 6721 -50
rect 6826 -65 6846 -45
rect 6946 -70 6966 -50
rect 7066 -65 7086 -45
rect 7186 -70 7206 -50
rect 7306 -65 7326 -45
rect 7426 -70 7446 -50
rect 7546 -65 7566 -45
rect 7666 -70 7686 -50
rect 7791 -65 7811 -45
rect 7911 -70 7931 -50
rect 8031 -65 8051 -45
rect 8151 -70 8171 -50
rect 8276 -65 8296 -45
rect 8396 -70 8416 -50
rect 8516 -65 8536 -45
rect 8636 -70 8656 -50
rect 8761 -65 8781 -45
rect 8881 -70 8901 -50
rect 9001 -65 9021 -45
rect 9121 -70 9141 -50
rect 9246 -65 9266 -45
rect 9366 -70 9386 -50
rect 9491 -65 9511 -45
rect 9611 -70 9631 -50
rect 9736 -65 9756 -45
rect 9856 -70 9876 -50
rect 9976 -65 9996 -45
rect 10096 -70 10116 -50
rect 10221 -65 10241 -45
rect 10341 -70 10361 -50
rect 10461 -65 10481 -45
rect 10581 -70 10601 -50
rect 10706 -65 10726 -45
rect 10826 -70 10846 -50
rect 10946 -65 10966 -45
rect 11066 -70 11086 -50
rect 11191 -65 11211 -45
rect 11311 -70 11331 -50
rect 11431 -65 11451 -45
rect 11551 -70 11571 -50
rect 11676 -65 11696 -45
rect 11796 -70 11816 -50
rect 11916 -65 11936 -45
rect 12036 -70 12056 -50
rect 12161 -65 12181 -45
rect 12281 -70 12301 -50
rect 12401 -65 12421 -45
rect 12521 -70 12541 -50
rect 12646 -65 12666 -45
rect 12766 -70 12786 -50
rect 12886 -65 12906 -45
rect 13006 -70 13026 -50
rect 13131 -65 13151 -45
rect 13251 -70 13271 -50
rect 13371 -65 13391 -45
rect 13491 -70 13511 -50
rect 13616 -65 13636 -45
rect 13736 -70 13756 -50
rect 13856 -65 13876 -45
rect 13976 -70 13996 -50
rect 14101 -65 14121 -45
rect 14221 -70 14241 -50
rect 14341 -65 14361 -45
rect 14461 -70 14481 -50
rect 14586 -65 14606 -45
rect 14706 -70 14726 -50
rect 14826 -65 14846 -45
rect 14946 -70 14966 -50
rect 15071 -65 15091 -45
rect 15191 -70 15211 -50
rect 15311 -65 15331 -45
rect 15431 -70 15451 -50
rect 15556 -65 15576 -45
rect 15676 -70 15696 -50
rect 15796 -65 15816 -45
rect 15916 -70 15936 -50
rect 16041 -65 16061 -45
rect 16161 -70 16181 -50
rect 16281 -65 16301 -45
rect 16401 -70 16421 -50
rect 16526 -65 16546 -45
rect 16646 -70 16666 -50
rect 16766 -65 16786 -45
rect 16886 -70 16906 -50
rect 17011 -65 17031 -45
rect 17131 -70 17151 -50
rect 17251 -65 17271 -45
rect 17371 -70 17391 -50
rect 17496 -65 17516 -45
rect 17616 -70 17636 -50
rect 17736 -65 17756 -45
rect 17856 -70 17876 -50
rect 17981 -65 18001 -45
rect 18101 -70 18121 -50
rect 18221 -65 18241 -45
rect 18341 -70 18361 -50
rect 18466 -65 18486 -45
rect 18586 -70 18606 -50
rect 18706 -65 18726 -45
rect 18826 -70 18846 -50
rect 18951 -65 18971 -45
rect 19071 -70 19091 -50
rect 19191 -65 19211 -45
rect 19311 -70 19331 -50
rect 19436 -65 19456 -45
rect 19556 -70 19576 -50
rect 19676 -65 19696 -45
rect 19796 -70 19816 -50
rect 19921 -65 19941 -45
rect 20041 -70 20061 -50
rect 20161 -65 20181 -45
rect 20281 -70 20301 -50
rect 20406 -65 20426 -45
rect 20526 -70 20546 -50
rect 20646 -65 20666 -45
rect 20766 -70 20786 -50
rect 20891 -65 20911 -45
rect 21011 -70 21031 -50
rect 21126 -70 21146 -50
rect 386 -145 406 -125
rect 191 -190 211 -170
rect 506 -145 526 -125
rect 691 -145 711 -125
rect 436 -190 456 -170
rect 811 -145 831 -125
rect 936 -145 956 -125
rect 741 -190 761 -170
rect 1056 -145 1076 -125
rect 1176 -145 1196 -125
rect 986 -190 1006 -170
rect 1296 -145 1316 -125
rect 1421 -145 1441 -125
rect 1226 -190 1246 -170
rect 1541 -145 1561 -125
rect 1726 -145 1746 -125
rect 1471 -190 1491 -170
rect 1846 -145 1866 -125
rect 1971 -145 1991 -125
rect 1776 -190 1796 -170
rect 2091 -145 2111 -125
rect 2211 -145 2231 -125
rect 2021 -190 2041 -170
rect 2331 -145 2351 -125
rect 2456 -145 2476 -125
rect 2261 -190 2281 -170
rect 2576 -145 2596 -125
rect 2696 -145 2716 -125
rect 2506 -190 2526 -170
rect 2816 -145 2836 -125
rect 2941 -145 2961 -125
rect 2746 -190 2766 -170
rect 3061 -145 3081 -125
rect 3181 -145 3201 -125
rect 2991 -190 3011 -170
rect 3301 -145 3321 -125
rect 3426 -145 3446 -125
rect 3231 -190 3251 -170
rect 3546 -145 3566 -125
rect 3666 -145 3686 -125
rect 3476 -190 3496 -170
rect 3786 -145 3806 -125
rect 3911 -145 3931 -125
rect 3716 -190 3736 -170
rect 4031 -145 4051 -125
rect 4151 -145 4171 -125
rect 3961 -190 3981 -170
rect 4271 -145 4291 -125
rect 4396 -145 4416 -125
rect -415 -240 -365 -190
rect 1635 -240 1675 -200
rect 4201 -190 4221 -170
rect 4516 -145 4536 -125
rect 4636 -145 4656 -125
rect 4446 -190 4466 -170
rect 4756 -145 4776 -125
rect 4881 -145 4901 -125
rect 4686 -190 4706 -170
rect 5001 -145 5021 -125
rect 5121 -145 5141 -125
rect 4931 -190 4951 -170
rect 5241 -145 5261 -125
rect 5366 -145 5386 -125
rect 5171 -190 5191 -170
rect 5486 -145 5506 -125
rect 5671 -145 5691 -125
rect 5416 -190 5436 -170
rect 5791 -145 5811 -125
rect 5916 -145 5936 -125
rect 5721 -190 5741 -170
rect 6036 -145 6056 -125
rect 6156 -145 6176 -125
rect 5966 -190 5986 -170
rect 6276 -145 6296 -125
rect 6401 -140 6421 -120
rect 6521 -145 6541 -125
rect 6641 -145 6661 -125
rect 6206 -190 6226 -170
rect 6761 -145 6781 -125
rect 6886 -145 6906 -125
rect 4060 -235 4100 -195
rect 6691 -190 6711 -170
rect 7006 -145 7026 -125
rect 7126 -145 7146 -125
rect 6936 -190 6956 -170
rect 7246 -145 7266 -125
rect 7366 -145 7386 -125
rect 7176 -190 7196 -170
rect 7486 -145 7506 -125
rect 7606 -145 7626 -125
rect 7416 -190 7436 -170
rect 7726 -145 7746 -125
rect 7851 -145 7871 -125
rect 7971 -145 7991 -125
rect 8091 -145 8111 -125
rect 7656 -190 7676 -170
rect 8211 -145 8231 -125
rect 8336 -145 8356 -125
rect 95 -270 115 -250
rect 25 -315 45 -295
rect 335 -270 355 -250
rect 145 -315 165 -295
rect 265 -315 285 -295
rect 575 -270 595 -250
rect 385 -315 405 -295
rect 505 -315 525 -295
rect 815 -270 835 -250
rect 625 -315 645 -295
rect 745 -315 765 -295
rect 1055 -270 1075 -250
rect 865 -315 885 -295
rect 985 -315 1005 -295
rect 1295 -270 1315 -250
rect 1105 -315 1125 -295
rect 1225 -315 1245 -295
rect 1535 -270 1555 -250
rect 1345 -315 1365 -295
rect 1465 -315 1485 -295
rect 1775 -270 1795 -250
rect 1585 -315 1605 -295
rect 1705 -315 1725 -295
rect 2015 -270 2035 -250
rect 1825 -315 1845 -295
rect 1945 -315 1965 -295
rect 2255 -270 2275 -250
rect 2065 -315 2085 -295
rect 2185 -315 2205 -295
rect 2495 -270 2515 -250
rect 2305 -315 2325 -295
rect 2425 -315 2445 -295
rect 2735 -270 2755 -250
rect 2545 -315 2565 -295
rect 2665 -315 2685 -295
rect 2975 -270 2995 -250
rect 2785 -315 2805 -295
rect 2905 -315 2925 -295
rect 3215 -270 3235 -250
rect 3025 -315 3045 -295
rect 3145 -315 3165 -295
rect 3455 -270 3475 -250
rect 3265 -315 3285 -295
rect 3385 -315 3405 -295
rect 3695 -270 3715 -250
rect 3505 -315 3525 -295
rect 3625 -315 3645 -295
rect 3935 -270 3955 -250
rect 3745 -315 3765 -295
rect 3865 -315 3885 -295
rect 4175 -270 4195 -250
rect 3985 -315 4005 -295
rect 4105 -315 4125 -295
rect 4415 -270 4435 -250
rect 4225 -315 4245 -295
rect 4345 -315 4365 -295
rect 4655 -270 4675 -250
rect 4465 -315 4485 -295
rect 4585 -315 4605 -295
rect 4895 -270 4915 -250
rect 4705 -315 4725 -295
rect 4825 -315 4845 -295
rect 5135 -270 5155 -250
rect 4945 -315 4965 -295
rect 5065 -315 5085 -295
rect 5375 -270 5395 -250
rect 5185 -315 5205 -295
rect 5305 -315 5325 -295
rect 5615 -270 5635 -250
rect 5425 -315 5445 -295
rect 5545 -315 5565 -295
rect 5855 -270 5875 -250
rect 5665 -315 5685 -295
rect 5785 -315 5805 -295
rect 6095 -270 6115 -250
rect 5905 -315 5925 -295
rect 6025 -315 6045 -295
rect 6335 -270 6355 -250
rect 6455 -260 6495 -220
rect 8141 -190 8161 -170
rect 8456 -145 8476 -125
rect 8576 -145 8596 -125
rect 8386 -190 8406 -170
rect 8696 -145 8716 -125
rect 8821 -145 8841 -125
rect 8626 -190 8646 -170
rect 8941 -145 8961 -125
rect 9061 -145 9081 -125
rect 8871 -190 8891 -170
rect 9181 -145 9201 -125
rect 9306 -145 9326 -125
rect 9111 -190 9131 -170
rect 9426 -145 9446 -125
rect 9551 -140 9571 -120
rect 9671 -145 9691 -125
rect 9796 -145 9816 -125
rect 9356 -190 9376 -170
rect 9916 -145 9936 -125
rect 10036 -145 10056 -125
rect 6575 -270 6595 -250
rect 6145 -315 6165 -295
rect 6265 -315 6285 -295
rect 6385 -315 6405 -295
rect 6505 -315 6525 -295
rect 6815 -270 6835 -250
rect 6625 -315 6645 -295
rect 6745 -315 6765 -295
rect 7055 -270 7075 -250
rect 6865 -315 6885 -295
rect 6985 -315 7005 -295
rect 7295 -270 7315 -250
rect 7105 -315 7125 -295
rect 7225 -315 7245 -295
rect 7535 -270 7555 -250
rect 7345 -315 7365 -295
rect 7465 -315 7485 -295
rect 7775 -270 7795 -250
rect 7880 -260 7920 -220
rect 9846 -190 9866 -170
rect 10156 -145 10176 -125
rect 10281 -145 10301 -125
rect 10086 -190 10106 -170
rect 10401 -145 10421 -125
rect 10521 -145 10541 -125
rect 10331 -190 10351 -170
rect 10641 -145 10661 -125
rect 10766 -145 10786 -125
rect 10571 -190 10591 -170
rect 10886 -145 10906 -125
rect 11006 -145 11026 -125
rect 10816 -190 10836 -170
rect 11126 -145 11146 -125
rect 11251 -145 11271 -125
rect 11056 -190 11076 -170
rect 11371 -145 11391 -125
rect 11491 -145 11511 -125
rect 11301 -190 11321 -170
rect 11611 -145 11631 -125
rect 11736 -145 11756 -125
rect 11541 -190 11561 -170
rect 11856 -145 11876 -125
rect 11976 -145 11996 -125
rect 12096 -145 12116 -125
rect 12221 -145 12241 -125
rect 11786 -190 11806 -170
rect 12341 -145 12361 -125
rect 12461 -145 12481 -125
rect 12271 -190 12291 -170
rect 12581 -145 12601 -125
rect 12706 -145 12726 -125
rect 12511 -190 12531 -170
rect 12826 -145 12846 -125
rect 12946 -145 12966 -125
rect 12756 -190 12776 -170
rect 13066 -145 13086 -125
rect 13191 -145 13211 -125
rect 12996 -190 13016 -170
rect 13311 -145 13331 -125
rect 13431 -145 13451 -125
rect 13241 -190 13261 -170
rect 13551 -145 13571 -125
rect 13676 -145 13696 -125
rect 13481 -190 13501 -170
rect 13796 -145 13816 -125
rect 13916 -145 13936 -125
rect 14036 -145 14056 -125
rect 14161 -145 14181 -125
rect 13726 -190 13746 -170
rect 14281 -145 14301 -125
rect 14401 -145 14421 -125
rect 14211 -190 14231 -170
rect 14521 -145 14541 -125
rect 14646 -145 14666 -125
rect 14451 -190 14471 -170
rect 14766 -145 14786 -125
rect 14886 -145 14906 -125
rect 14696 -190 14716 -170
rect 15006 -145 15026 -125
rect 15131 -145 15151 -125
rect 14936 -190 14956 -170
rect 15251 -145 15271 -125
rect 15371 -145 15391 -125
rect 15181 -190 15201 -170
rect 15491 -145 15511 -125
rect 15616 -145 15636 -125
rect 15421 -190 15441 -170
rect 15736 -145 15756 -125
rect 15856 -145 15876 -125
rect 15976 -145 15996 -125
rect 16101 -145 16121 -125
rect 15666 -190 15686 -170
rect 16221 -145 16241 -125
rect 16341 -145 16361 -125
rect 8015 -270 8035 -250
rect 7585 -315 7605 -295
rect 7705 -315 7725 -295
rect 7825 -315 7845 -295
rect 7945 -315 7965 -295
rect 8255 -270 8275 -250
rect 8065 -315 8085 -295
rect 8185 -315 8205 -295
rect 8495 -270 8515 -250
rect 8305 -315 8325 -295
rect 8425 -315 8445 -295
rect 8735 -270 8755 -250
rect 8545 -315 8565 -295
rect 8665 -315 8685 -295
rect 8975 -270 8995 -250
rect 8785 -315 8805 -295
rect 8905 -315 8925 -295
rect 9215 -270 9235 -250
rect 9025 -315 9045 -295
rect 9145 -315 9165 -295
rect 9455 -270 9475 -250
rect 9570 -250 9610 -210
rect 9265 -315 9285 -295
rect 9385 -315 9405 -295
rect 9695 -270 9715 -250
rect 9505 -315 9525 -295
rect 9625 -315 9645 -295
rect 9935 -270 9955 -250
rect 9745 -315 9765 -295
rect 9865 -315 9885 -295
rect 10175 -270 10195 -250
rect 9985 -315 10005 -295
rect 10105 -315 10125 -295
rect 10415 -270 10435 -250
rect 10225 -315 10245 -295
rect 10345 -315 10365 -295
rect 10655 -270 10675 -250
rect 10465 -315 10485 -295
rect 10585 -315 10605 -295
rect 10895 -270 10915 -250
rect 10705 -315 10725 -295
rect 10825 -315 10845 -295
rect 11135 -270 11155 -250
rect 10945 -315 10965 -295
rect 11065 -315 11085 -295
rect 11375 -270 11395 -250
rect 11185 -315 11205 -295
rect 11305 -315 11325 -295
rect 11615 -270 11635 -250
rect 11425 -315 11445 -295
rect 11545 -315 11565 -295
rect 11855 -270 11875 -250
rect 11950 -260 11990 -220
rect 12095 -270 12115 -250
rect 11665 -315 11685 -295
rect 11785 -315 11805 -295
rect 11905 -315 11925 -295
rect 12025 -315 12045 -295
rect 12335 -270 12355 -250
rect 12145 -315 12165 -295
rect 12265 -315 12285 -295
rect 12575 -270 12595 -250
rect 12385 -315 12405 -295
rect 12505 -315 12525 -295
rect 12815 -270 12835 -250
rect 12625 -315 12645 -295
rect 12745 -315 12765 -295
rect 13055 -270 13075 -250
rect 12865 -315 12885 -295
rect 12985 -315 13005 -295
rect 13295 -270 13315 -250
rect 13105 -315 13125 -295
rect 13225 -315 13245 -295
rect 13535 -270 13555 -250
rect 13345 -315 13365 -295
rect 13465 -315 13485 -295
rect 13775 -270 13795 -250
rect 13870 -260 13910 -220
rect 16151 -190 16171 -170
rect 16461 -145 16481 -125
rect 16586 -145 16606 -125
rect 16391 -190 16411 -170
rect 16706 -145 16726 -125
rect 16826 -145 16846 -125
rect 16636 -190 16656 -170
rect 16946 -145 16966 -125
rect 17071 -145 17091 -125
rect 16876 -190 16896 -170
rect 17191 -145 17211 -125
rect 17311 -145 17331 -125
rect 17121 -190 17141 -170
rect 17431 -145 17451 -125
rect 17556 -145 17576 -125
rect 17361 -190 17381 -170
rect 17676 -145 17696 -125
rect 17796 -145 17816 -125
rect 17606 -190 17626 -170
rect 17916 -145 17936 -125
rect 18041 -145 18061 -125
rect 17846 -190 17866 -170
rect 18161 -145 18181 -125
rect 18281 -145 18301 -125
rect 18091 -190 18111 -170
rect 18401 -145 18421 -125
rect 18526 -145 18546 -125
rect 18331 -190 18351 -170
rect 18646 -145 18666 -125
rect 18766 -145 18786 -125
rect 18576 -190 18596 -170
rect 18886 -145 18906 -125
rect 19011 -145 19031 -125
rect 18816 -190 18836 -170
rect 19131 -145 19151 -125
rect 19251 -145 19271 -125
rect 19061 -190 19081 -170
rect 19371 -145 19391 -125
rect 19496 -145 19516 -125
rect 19301 -190 19321 -170
rect 19616 -145 19636 -125
rect 19736 -145 19756 -125
rect 19546 -190 19566 -170
rect 19856 -145 19876 -125
rect 19981 -145 20001 -125
rect 19786 -190 19806 -170
rect 20101 -145 20121 -125
rect 20221 -145 20241 -125
rect 20031 -190 20051 -170
rect 20341 -145 20361 -125
rect 20466 -145 20486 -125
rect 20271 -190 20291 -170
rect 20586 -145 20606 -125
rect 20706 -145 20726 -125
rect 20516 -190 20536 -170
rect 20826 -145 20846 -125
rect 20951 -145 20971 -125
rect 20756 -190 20776 -170
rect 21071 -145 21091 -125
rect 21001 -190 21021 -170
rect 14015 -270 14035 -250
rect 13585 -315 13605 -295
rect 13705 -315 13725 -295
rect 13825 -315 13845 -295
rect 13945 -315 13965 -295
rect 14255 -270 14275 -250
rect 14065 -315 14085 -295
rect 14185 -315 14205 -295
rect 14495 -270 14515 -250
rect 14305 -315 14325 -295
rect 14425 -315 14445 -295
rect 14735 -270 14755 -250
rect 14545 -315 14565 -295
rect 14665 -315 14685 -295
rect 14975 -270 14995 -250
rect 14785 -315 14805 -295
rect 14905 -315 14925 -295
rect 15215 -270 15235 -250
rect 15025 -315 15045 -295
rect 15145 -315 15165 -295
rect 15455 -270 15475 -250
rect 15265 -315 15285 -295
rect 15385 -315 15405 -295
rect 15695 -270 15715 -250
rect 15815 -260 15855 -220
rect 17705 -250 17745 -210
rect 19645 -250 19685 -210
rect 15935 -270 15955 -250
rect 15505 -315 15525 -295
rect 15625 -315 15645 -295
rect 15745 -315 15765 -295
rect 15865 -315 15885 -295
rect 16175 -270 16195 -250
rect 15985 -315 16005 -295
rect 16105 -315 16125 -295
rect 16415 -270 16435 -250
rect 16225 -315 16245 -295
rect 16345 -315 16365 -295
rect 16655 -270 16675 -250
rect 16465 -315 16485 -295
rect 16585 -315 16605 -295
rect 16895 -270 16915 -250
rect 16705 -315 16725 -295
rect 16825 -315 16845 -295
rect 17135 -270 17155 -250
rect 16945 -315 16965 -295
rect 17065 -315 17085 -295
rect 17375 -270 17395 -250
rect 17185 -315 17205 -295
rect 17305 -315 17325 -295
rect 17615 -270 17635 -250
rect 17425 -315 17445 -295
rect 17545 -315 17565 -295
rect 17855 -270 17875 -250
rect 17665 -315 17685 -295
rect 17785 -315 17805 -295
rect 18095 -270 18115 -250
rect 17905 -315 17925 -295
rect 18025 -315 18045 -295
rect 18335 -270 18355 -250
rect 18145 -315 18165 -295
rect 18265 -315 18285 -295
rect 18575 -270 18595 -250
rect 18385 -315 18405 -295
rect 18505 -315 18525 -295
rect 18815 -270 18835 -250
rect 18625 -315 18645 -295
rect 18745 -315 18765 -295
rect 19055 -270 19075 -250
rect 18865 -315 18885 -295
rect 18985 -315 19005 -295
rect 19295 -270 19315 -250
rect 19105 -315 19125 -295
rect 19225 -315 19245 -295
rect 19535 -270 19555 -250
rect 19345 -315 19365 -295
rect 19465 -315 19485 -295
rect 19775 -270 19795 -250
rect 19585 -315 19605 -295
rect 19705 -315 19725 -295
rect 20015 -270 20035 -250
rect 19825 -315 19845 -295
rect 19945 -315 19965 -295
rect 20255 -270 20275 -250
rect 20065 -315 20085 -295
rect 20185 -315 20205 -295
rect 20495 -270 20515 -250
rect 20305 -315 20325 -295
rect 20425 -315 20445 -295
rect 20735 -270 20755 -250
rect 20545 -315 20565 -295
rect 20665 -315 20685 -295
rect 20975 -270 20995 -250
rect 20785 -315 20805 -295
rect 20905 -315 20925 -295
rect 21215 -270 21235 -250
rect 21025 -315 21045 -295
rect 21145 -315 21165 -295
rect 21455 -270 21475 -250
rect 21265 -315 21285 -295
rect 21385 -315 21405 -295
rect 21695 -270 21715 -250
rect 21505 -315 21525 -295
rect 21625 -315 21645 -295
rect 21935 -270 21955 -250
rect 21745 -315 21765 -295
rect 21865 -315 21885 -295
rect 22175 -270 22195 -250
rect 21985 -315 22005 -295
rect 22105 -315 22125 -295
rect 22415 -270 22435 -250
rect 22225 -315 22245 -295
rect 22345 -315 22365 -295
rect 22655 -270 22675 -250
rect 22465 -315 22485 -295
rect 22585 -315 22605 -295
rect 22895 -270 22915 -250
rect 22705 -315 22725 -295
rect 22825 -315 22845 -295
rect 23135 -270 23155 -250
rect 22945 -315 22965 -295
rect 23065 -315 23085 -295
rect 23375 -270 23395 -250
rect 23185 -315 23205 -295
rect 23305 -315 23325 -295
rect 23615 -270 23635 -250
rect 23425 -315 23445 -295
rect 23545 -315 23565 -295
rect 23855 -270 23875 -250
rect 23665 -315 23685 -295
rect 23785 -315 23805 -295
rect 24095 -270 24115 -250
rect 23905 -315 23925 -295
rect 24025 -315 24045 -295
rect 24335 -270 24355 -250
rect 24145 -315 24165 -295
rect 24265 -315 24285 -295
rect 24575 -270 24595 -250
rect 24385 -315 24405 -295
rect 24505 -315 24525 -295
rect 24815 -270 24835 -250
rect 24625 -315 24645 -295
rect 24745 -315 24765 -295
rect 25055 -270 25075 -250
rect 24865 -315 24885 -295
rect 24985 -315 25005 -295
rect 25295 -270 25315 -250
rect 25105 -315 25125 -295
rect 25225 -315 25245 -295
rect 25535 -270 25555 -250
rect 25345 -315 25365 -295
rect 25465 -315 25485 -295
rect 25775 -270 25795 -250
rect 25585 -315 25605 -295
rect 25705 -315 25725 -295
rect 26015 -270 26035 -250
rect 25825 -315 25845 -295
rect 25945 -315 25965 -295
rect 26255 -270 26275 -250
rect 26065 -315 26085 -295
rect 26185 -315 26205 -295
rect 26495 -270 26515 -250
rect 26305 -315 26325 -295
rect 26425 -315 26445 -295
rect 26735 -270 26755 -250
rect 26545 -315 26565 -295
rect 26665 -315 26685 -295
rect 26975 -270 26995 -250
rect 26785 -315 26805 -295
rect 26905 -315 26925 -295
rect 27215 -270 27235 -250
rect 27025 -315 27045 -295
rect 27145 -315 27165 -295
rect 27455 -270 27475 -250
rect 27265 -315 27285 -295
rect 27385 -315 27405 -295
rect 27695 -270 27715 -250
rect 27505 -315 27525 -295
rect 27625 -315 27645 -295
rect 27935 -270 27955 -250
rect 27745 -315 27765 -295
rect 27865 -315 27885 -295
rect 28175 -270 28195 -250
rect 27985 -315 28005 -295
rect 28105 -315 28125 -295
rect 28415 -270 28435 -250
rect 28225 -315 28245 -295
rect 28345 -315 28365 -295
rect 28655 -270 28675 -250
rect 28465 -315 28485 -295
rect 28585 -315 28605 -295
rect 28895 -270 28915 -250
rect 28705 -315 28725 -295
rect 28825 -315 28845 -295
rect 29135 -270 29155 -250
rect 28945 -315 28965 -295
rect 29065 -315 29085 -295
rect 29375 -270 29395 -250
rect 29185 -315 29205 -295
rect 29305 -315 29325 -295
rect 29615 -270 29635 -250
rect 29425 -315 29445 -295
rect 29545 -315 29565 -295
rect 29855 -270 29875 -250
rect 29665 -315 29685 -295
rect 29785 -315 29805 -295
rect 30095 -270 30115 -250
rect 29905 -315 29925 -295
rect 30025 -315 30045 -295
rect 30335 -270 30355 -250
rect 30145 -315 30165 -295
rect 30265 -315 30285 -295
rect 30575 -270 30595 -250
rect 30385 -315 30405 -295
rect 30505 -315 30525 -295
rect 30625 -315 30645 -295
rect -30 -440 -10 -420
rect 85 -440 105 -420
rect 210 -440 230 -420
rect 325 -440 345 -420
rect 450 -440 470 -420
rect 565 -440 585 -420
rect 690 -440 710 -420
rect 805 -440 825 -420
rect 930 -440 950 -420
rect 1045 -440 1065 -420
rect 1170 -440 1190 -420
rect 1285 -440 1305 -420
rect 1410 -440 1430 -420
rect 1525 -440 1545 -420
rect 1650 -440 1670 -420
rect 1765 -440 1785 -420
rect 1890 -440 1910 -420
rect 2005 -440 2025 -420
rect 2130 -440 2150 -420
rect 2245 -440 2265 -420
rect 2370 -440 2390 -420
rect 2485 -440 2505 -420
rect 2610 -440 2630 -420
rect 2725 -440 2745 -420
rect 2850 -440 2870 -420
rect 2965 -440 2985 -420
rect 3090 -440 3110 -420
rect 3205 -440 3225 -420
rect 3330 -440 3350 -420
rect 3445 -440 3465 -420
rect 3570 -440 3590 -420
rect 3685 -440 3705 -420
rect 3810 -440 3830 -420
rect 3925 -440 3945 -420
rect 4050 -440 4070 -420
rect 4165 -440 4185 -420
rect 4290 -440 4310 -420
rect 4405 -440 4425 -420
rect 4530 -440 4550 -420
rect 4645 -440 4665 -420
rect 4770 -440 4790 -420
rect 4885 -440 4905 -420
rect 5010 -440 5030 -420
rect 5125 -440 5145 -420
rect 5250 -440 5270 -420
rect 5365 -440 5385 -420
rect 5490 -440 5510 -420
rect 5605 -440 5625 -420
rect 5730 -440 5750 -420
rect 5845 -440 5865 -420
rect 5970 -440 5990 -420
rect 6085 -440 6105 -420
rect 6210 -440 6230 -420
rect 6325 -440 6345 -420
rect 6450 -440 6470 -420
rect 6565 -440 6585 -420
rect 6690 -440 6710 -420
rect 6805 -440 6825 -420
rect 6930 -440 6950 -420
rect 7045 -440 7065 -420
rect 7170 -440 7190 -420
rect 7285 -440 7305 -420
rect 7410 -440 7430 -420
rect 7525 -440 7545 -420
rect 7650 -440 7670 -420
rect 7765 -440 7785 -420
rect 7890 -440 7910 -420
rect 8005 -440 8025 -420
rect 8130 -440 8150 -420
rect 8245 -440 8265 -420
rect 8370 -440 8390 -420
rect 8485 -440 8505 -420
rect 8610 -440 8630 -420
rect 8725 -440 8745 -420
rect 8850 -440 8870 -420
rect 8965 -440 8985 -420
rect 9090 -440 9110 -420
rect 9205 -440 9225 -420
rect 9330 -440 9350 -420
rect 9445 -440 9465 -420
rect 9570 -440 9590 -420
rect 9685 -440 9705 -420
rect 9810 -440 9830 -420
rect 9925 -440 9945 -420
rect 10050 -440 10070 -420
rect 10165 -440 10185 -420
rect 10290 -440 10310 -420
rect 10405 -440 10425 -420
rect 10530 -440 10550 -420
rect 10645 -440 10665 -420
rect 10770 -440 10790 -420
rect 10885 -440 10905 -420
rect 11010 -440 11030 -420
rect 11125 -440 11145 -420
rect 11250 -440 11270 -420
rect 11365 -440 11385 -420
rect 11490 -440 11510 -420
rect 11605 -440 11625 -420
rect 11730 -440 11750 -420
rect 11845 -440 11865 -420
rect 11970 -440 11990 -420
rect 12085 -440 12105 -420
rect 12210 -440 12230 -420
rect 12325 -440 12345 -420
rect 12450 -440 12470 -420
rect 12565 -440 12585 -420
rect 12690 -440 12710 -420
rect 12805 -440 12825 -420
rect 12930 -440 12950 -420
rect 13045 -440 13065 -420
rect 13170 -440 13190 -420
rect 13285 -440 13305 -420
rect 13410 -440 13430 -420
rect 13525 -440 13545 -420
rect 13650 -440 13670 -420
rect 13765 -440 13785 -420
rect 13890 -440 13910 -420
rect 14005 -440 14025 -420
rect 14130 -440 14150 -420
rect 14245 -440 14265 -420
rect 14370 -440 14390 -420
rect 14485 -440 14505 -420
rect 14610 -440 14630 -420
rect 14725 -440 14745 -420
rect 14850 -440 14870 -420
rect 14965 -440 14985 -420
rect 15090 -440 15110 -420
rect 15205 -440 15225 -420
rect 15330 -440 15350 -420
rect 15445 -440 15465 -420
rect 15570 -440 15590 -420
rect 15685 -440 15705 -420
rect 15810 -440 15830 -420
rect 15925 -440 15945 -420
rect 16050 -440 16070 -420
rect 16165 -440 16185 -420
rect 16290 -440 16310 -420
rect 16405 -440 16425 -420
rect 16530 -440 16550 -420
rect 16645 -440 16665 -420
rect 16770 -440 16790 -420
rect 16885 -440 16905 -420
rect 17010 -440 17030 -420
rect 17125 -440 17145 -420
rect 17250 -440 17270 -420
rect 17365 -440 17385 -420
rect 17490 -440 17510 -420
rect 17605 -440 17625 -420
rect 17730 -440 17750 -420
rect 17845 -440 17865 -420
rect 17970 -440 17990 -420
rect 18085 -440 18105 -420
rect 18210 -440 18230 -420
rect 18325 -440 18345 -420
rect 18450 -440 18470 -420
rect 18565 -440 18585 -420
rect 18690 -440 18710 -420
rect 18805 -440 18825 -420
rect 18930 -440 18950 -420
rect 19045 -440 19065 -420
rect 19170 -440 19190 -420
rect 19285 -440 19305 -420
rect 19410 -440 19430 -420
rect 19525 -440 19545 -420
rect 19650 -440 19670 -420
rect 19765 -440 19785 -420
rect 19890 -440 19910 -420
rect 20005 -440 20025 -420
rect 20130 -440 20150 -420
rect 20245 -440 20265 -420
rect 20370 -440 20390 -420
rect 20485 -440 20505 -420
rect 20610 -440 20630 -420
rect 20725 -440 20745 -420
rect 20850 -440 20870 -420
rect 20965 -440 20985 -420
rect 21090 -440 21110 -420
rect 21205 -440 21225 -420
rect 21330 -440 21350 -420
rect 21445 -440 21465 -420
rect 21570 -440 21590 -420
rect 21685 -440 21705 -420
rect 21810 -440 21830 -420
rect 21925 -440 21945 -420
rect 22050 -440 22070 -420
rect 22165 -440 22185 -420
rect 22290 -440 22310 -420
rect 22405 -440 22425 -420
rect 22530 -440 22550 -420
rect 22645 -440 22665 -420
rect 22770 -440 22790 -420
rect 22885 -440 22905 -420
rect 23010 -440 23030 -420
rect 23125 -440 23145 -420
rect 23250 -440 23270 -420
rect 23365 -440 23385 -420
rect 23490 -440 23510 -420
rect 23605 -440 23625 -420
rect 23730 -440 23750 -420
rect 23845 -440 23865 -420
rect 23970 -440 23990 -420
rect 24085 -440 24105 -420
rect 24210 -440 24230 -420
rect 24325 -440 24345 -420
rect 24450 -440 24470 -420
rect 24565 -440 24585 -420
rect 24690 -440 24710 -420
rect 24805 -440 24825 -420
rect 24930 -440 24950 -420
rect 25045 -440 25065 -420
rect 25170 -440 25190 -420
rect 25285 -440 25305 -420
rect 25410 -440 25430 -420
rect 25525 -440 25545 -420
rect 25650 -440 25670 -420
rect 25765 -440 25785 -420
rect 25890 -440 25910 -420
rect 26005 -440 26025 -420
rect 26130 -440 26150 -420
rect 26245 -440 26265 -420
rect 26370 -440 26390 -420
rect 26485 -440 26505 -420
rect 26610 -440 26630 -420
rect 26725 -440 26745 -420
rect 26850 -440 26870 -420
rect 26965 -440 26985 -420
rect 27090 -440 27110 -420
rect 27205 -440 27225 -420
rect 27330 -440 27350 -420
rect 27445 -440 27465 -420
rect 27570 -440 27590 -420
rect 27685 -440 27705 -420
rect 27810 -440 27830 -420
rect 27925 -440 27945 -420
rect 28050 -440 28070 -420
rect 28165 -440 28185 -420
rect 28290 -440 28310 -420
rect 28405 -440 28425 -420
rect 28530 -440 28550 -420
rect 28645 -440 28665 -420
rect 28770 -440 28790 -420
rect 28885 -440 28905 -420
rect 29010 -440 29030 -420
rect 29125 -440 29145 -420
rect 29250 -440 29270 -420
rect 29365 -440 29385 -420
rect 29490 -440 29510 -420
rect 29605 -440 29625 -420
rect 29730 -440 29750 -420
rect 29845 -440 29865 -420
rect 29970 -440 29990 -420
rect 30085 -440 30105 -420
rect 30210 -440 30230 -420
rect 30325 -440 30345 -420
rect 30450 -440 30470 -420
rect 30565 -440 30585 -420
rect 30685 -445 30705 -425
rect 30740 -505 30760 -485
rect -30 -565 -10 -545
rect 90 -565 110 -545
rect 210 -565 230 -545
rect 330 -565 350 -545
rect 450 -565 470 -545
rect 570 -565 590 -545
rect 690 -565 710 -545
rect 810 -565 830 -545
rect 930 -565 950 -545
rect 1050 -565 1070 -545
rect 1170 -565 1190 -545
rect 1290 -565 1310 -545
rect 1410 -565 1430 -545
rect 1530 -565 1550 -545
rect 1650 -565 1670 -545
rect 1770 -565 1790 -545
rect 1890 -565 1910 -545
rect 2010 -565 2030 -545
rect 2130 -565 2150 -545
rect 2250 -565 2270 -545
rect 2370 -565 2390 -545
rect 2490 -565 2510 -545
rect 2610 -565 2630 -545
rect 2730 -565 2750 -545
rect 2850 -565 2870 -545
rect 2970 -565 2990 -545
rect 3090 -565 3110 -545
rect 3210 -565 3230 -545
rect 3330 -565 3350 -545
rect 3450 -565 3470 -545
rect 3570 -565 3590 -545
rect 3690 -565 3710 -545
rect 3810 -565 3830 -545
rect 3930 -565 3950 -545
rect 4050 -565 4070 -545
rect 4170 -565 4190 -545
rect 4290 -565 4310 -545
rect 4410 -565 4430 -545
rect 4530 -565 4550 -545
rect 4650 -565 4670 -545
rect 4770 -565 4790 -545
rect 4890 -565 4910 -545
rect 5010 -565 5030 -545
rect 5130 -565 5150 -545
rect 5250 -565 5270 -545
rect 5370 -565 5390 -545
rect 5490 -565 5510 -545
rect 5610 -565 5630 -545
rect 5730 -565 5750 -545
rect 5850 -565 5870 -545
rect 5970 -565 5990 -545
rect 6090 -565 6110 -545
rect 6210 -565 6230 -545
rect 6330 -565 6350 -545
rect 6450 -565 6470 -545
rect 6570 -565 6590 -545
rect 6690 -565 6710 -545
rect 6810 -565 6830 -545
rect 6930 -565 6950 -545
rect 7050 -565 7070 -545
rect 7170 -565 7190 -545
rect 7290 -565 7310 -545
rect 7410 -565 7430 -545
rect 7530 -565 7550 -545
rect 7650 -565 7670 -545
rect 7770 -565 7790 -545
rect 7890 -565 7910 -545
rect 8010 -565 8030 -545
rect 8130 -565 8150 -545
rect 8250 -565 8270 -545
rect 8370 -565 8390 -545
rect 8490 -565 8510 -545
rect 8610 -565 8630 -545
rect 8730 -565 8750 -545
rect 8850 -565 8870 -545
rect 8970 -565 8990 -545
rect 9090 -565 9110 -545
rect 9210 -565 9230 -545
rect 9330 -565 9350 -545
rect 9450 -565 9470 -545
rect 9570 -565 9590 -545
rect 9690 -565 9710 -545
rect 9810 -565 9830 -545
rect 9930 -565 9950 -545
rect 10050 -565 10070 -545
rect 10170 -565 10190 -545
rect 10290 -565 10310 -545
rect 10410 -565 10430 -545
rect 10530 -565 10550 -545
rect 10650 -565 10670 -545
rect 10770 -565 10790 -545
rect 10890 -565 10910 -545
rect 11010 -565 11030 -545
rect 11130 -565 11150 -545
rect 11250 -565 11270 -545
rect 11370 -565 11390 -545
rect 11490 -565 11510 -545
rect 11610 -565 11630 -545
rect 11730 -565 11750 -545
rect 11850 -565 11870 -545
rect 11970 -565 11990 -545
rect 12090 -565 12110 -545
rect 12210 -565 12230 -545
rect 12330 -565 12350 -545
rect 12450 -565 12470 -545
rect 12570 -565 12590 -545
rect 12690 -565 12710 -545
rect 12810 -565 12830 -545
rect 12930 -565 12950 -545
rect 13050 -565 13070 -545
rect 13170 -565 13190 -545
rect 13290 -565 13310 -545
rect 13410 -565 13430 -545
rect 13530 -565 13550 -545
rect 13650 -565 13670 -545
rect 13770 -565 13790 -545
rect 13890 -565 13910 -545
rect 14010 -565 14030 -545
rect 14130 -565 14150 -545
rect 14250 -565 14270 -545
rect 14370 -565 14390 -545
rect 14490 -565 14510 -545
rect 14610 -565 14630 -545
rect 14730 -565 14750 -545
rect 14850 -565 14870 -545
rect 14970 -565 14990 -545
rect 15090 -565 15110 -545
rect 15210 -565 15230 -545
rect 15330 -565 15350 -545
rect 15450 -565 15470 -545
rect 15570 -565 15590 -545
rect 15690 -565 15710 -545
rect 15810 -565 15830 -545
rect 15930 -565 15950 -545
rect 16050 -565 16070 -545
rect 16170 -565 16190 -545
rect 16290 -565 16310 -545
rect 16410 -565 16430 -545
rect 16530 -565 16550 -545
rect 16650 -565 16670 -545
rect 16770 -565 16790 -545
rect 16890 -565 16910 -545
rect 17010 -565 17030 -545
rect 17130 -565 17150 -545
rect 17250 -565 17270 -545
rect 17370 -565 17390 -545
rect 17490 -565 17510 -545
rect 17610 -565 17630 -545
rect 17730 -565 17750 -545
rect 17850 -565 17870 -545
rect 17970 -565 17990 -545
rect 18090 -565 18110 -545
rect 18210 -565 18230 -545
rect 18330 -565 18350 -545
rect 18450 -565 18470 -545
rect 18570 -565 18590 -545
rect 18690 -565 18710 -545
rect 18810 -565 18830 -545
rect 18930 -565 18950 -545
rect 19050 -565 19070 -545
rect 19170 -565 19190 -545
rect 19290 -565 19310 -545
rect 19410 -565 19430 -545
rect 19530 -565 19550 -545
rect 19650 -565 19670 -545
rect 19770 -565 19790 -545
rect 19890 -565 19910 -545
rect 20010 -565 20030 -545
rect 20130 -565 20150 -545
rect 20250 -565 20270 -545
rect 20370 -565 20390 -545
rect 20490 -565 20510 -545
rect 20610 -565 20630 -545
rect 20730 -565 20750 -545
rect 20850 -565 20870 -545
rect 20970 -565 20990 -545
rect 21090 -565 21110 -545
rect 21210 -565 21230 -545
rect 21330 -565 21350 -545
rect 21450 -565 21470 -545
rect 21570 -565 21590 -545
rect 21690 -565 21710 -545
rect 21810 -565 21830 -545
rect 21930 -565 21950 -545
rect 22050 -565 22070 -545
rect 22170 -565 22190 -545
rect 22290 -565 22310 -545
rect 22410 -565 22430 -545
rect 22530 -565 22550 -545
rect 22650 -565 22670 -545
rect 22770 -565 22790 -545
rect 22890 -565 22910 -545
rect 23010 -565 23030 -545
rect 23130 -565 23150 -545
rect 23250 -565 23270 -545
rect 23370 -565 23390 -545
rect 23490 -565 23510 -545
rect 23610 -565 23630 -545
rect 23730 -565 23750 -545
rect 23850 -565 23870 -545
rect 23970 -565 23990 -545
rect 24090 -565 24110 -545
rect 24210 -565 24230 -545
rect 24330 -565 24350 -545
rect 24450 -565 24470 -545
rect 24570 -565 24590 -545
rect 24690 -565 24710 -545
rect 24810 -565 24830 -545
rect 24930 -565 24950 -545
rect 25050 -565 25070 -545
rect 25170 -565 25190 -545
rect 25290 -565 25310 -545
rect 25410 -565 25430 -545
rect 25530 -565 25550 -545
rect 25650 -565 25670 -545
rect 25770 -565 25790 -545
rect 25890 -565 25910 -545
rect 26010 -565 26030 -545
rect 26130 -565 26150 -545
rect 26250 -565 26270 -545
rect 26370 -565 26390 -545
rect 26490 -565 26510 -545
rect 26610 -565 26630 -545
rect 26730 -565 26750 -545
rect 26850 -565 26870 -545
rect 26970 -565 26990 -545
rect 27090 -565 27110 -545
rect 27210 -565 27230 -545
rect 27330 -565 27350 -545
rect 27450 -565 27470 -545
rect 27570 -565 27590 -545
rect 27690 -565 27710 -545
rect 27810 -565 27830 -545
rect 27930 -565 27950 -545
rect 28050 -565 28070 -545
rect 28170 -565 28190 -545
rect 28290 -565 28310 -545
rect 28410 -565 28430 -545
rect 28530 -565 28550 -545
rect 28650 -565 28670 -545
rect 28770 -565 28790 -545
rect 28890 -565 28910 -545
rect 29010 -565 29030 -545
rect 29130 -565 29150 -545
rect 29250 -565 29270 -545
rect 29370 -565 29390 -545
rect 29490 -565 29510 -545
rect 29610 -565 29630 -545
rect 29730 -565 29750 -545
rect 29850 -565 29870 -545
rect 29970 -565 29990 -545
rect 30090 -565 30110 -545
rect 30210 -565 30230 -545
rect 30330 -565 30350 -545
rect 30450 -565 30470 -545
rect 30570 -565 30590 -545
rect 30685 -565 30705 -545
rect 25 -805 45 -785
rect 145 -805 165 -785
rect 265 -805 285 -785
rect 385 -805 405 -785
rect 505 -805 525 -785
rect 625 -805 645 -785
rect 745 -805 765 -785
rect 90 -845 110 -825
rect 330 -845 350 -825
rect 865 -805 885 -785
rect 985 -805 1005 -785
rect 1105 -805 1125 -785
rect 1225 -805 1245 -785
rect 1345 -805 1365 -785
rect 1465 -805 1485 -785
rect 1585 -805 1605 -785
rect 1705 -805 1725 -785
rect 1825 -805 1845 -785
rect 1945 -805 1965 -785
rect 2065 -805 2085 -785
rect 2185 -805 2205 -785
rect 2305 -805 2325 -785
rect 2425 -805 2445 -785
rect 2545 -805 2565 -785
rect 2665 -805 2685 -785
rect 2785 -805 2805 -785
rect 2905 -805 2925 -785
rect 570 -845 590 -825
rect 800 -870 835 -835
rect 1050 -845 1070 -825
rect 1290 -845 1310 -825
rect 1530 -845 1550 -825
rect 1770 -845 1790 -825
rect 2010 -845 2030 -825
rect 2250 -845 2270 -825
rect 2490 -845 2510 -825
rect 3025 -805 3045 -785
rect 3145 -805 3165 -785
rect 3265 -805 3285 -785
rect 3385 -805 3405 -785
rect 3505 -805 3525 -785
rect 3625 -805 3645 -785
rect 3745 -805 3765 -785
rect 3865 -805 3885 -785
rect 3985 -805 4005 -785
rect 4105 -805 4125 -785
rect 4225 -805 4245 -785
rect 4345 -805 4365 -785
rect 4465 -805 4485 -785
rect 4585 -805 4605 -785
rect 4705 -805 4725 -785
rect 4825 -805 4845 -785
rect 4945 -805 4965 -785
rect 5065 -805 5085 -785
rect 2730 -845 2750 -825
rect 2960 -870 2995 -835
rect 3210 -845 3230 -825
rect 3450 -845 3470 -825
rect 3690 -845 3710 -825
rect 3930 -845 3950 -825
rect 4170 -845 4190 -825
rect 4410 -845 4430 -825
rect 4650 -845 4670 -825
rect 5185 -805 5205 -785
rect 5305 -805 5325 -785
rect 5425 -805 5445 -785
rect 5545 -805 5565 -785
rect 5665 -805 5685 -785
rect 5785 -805 5805 -785
rect 5905 -805 5925 -785
rect 6025 -805 6045 -785
rect 6145 -805 6165 -785
rect 6265 -805 6285 -785
rect 6385 -805 6405 -785
rect 6505 -805 6525 -785
rect 6625 -805 6645 -785
rect 6745 -805 6765 -785
rect 6865 -805 6885 -785
rect 6985 -805 7005 -785
rect 7105 -805 7125 -785
rect 7225 -805 7245 -785
rect 4890 -845 4910 -825
rect 5120 -870 5155 -835
rect 5370 -845 5390 -825
rect 5610 -845 5630 -825
rect 5850 -845 5870 -825
rect 6090 -845 6110 -825
rect 6330 -845 6350 -825
rect 6570 -845 6590 -825
rect 6810 -845 6830 -825
rect 7345 -805 7365 -785
rect 7465 -805 7485 -785
rect 7585 -805 7605 -785
rect 7705 -805 7725 -785
rect 7825 -805 7845 -785
rect 7945 -805 7965 -785
rect 8065 -805 8085 -785
rect 8185 -805 8205 -785
rect 8305 -805 8325 -785
rect 8425 -805 8445 -785
rect 8545 -805 8565 -785
rect 8665 -805 8685 -785
rect 8785 -805 8805 -785
rect 8905 -805 8925 -785
rect 9025 -805 9045 -785
rect 9145 -805 9165 -785
rect 9265 -805 9285 -785
rect 9385 -805 9405 -785
rect 7050 -845 7070 -825
rect 7280 -870 7315 -835
rect 7530 -845 7550 -825
rect 7770 -845 7790 -825
rect 8010 -845 8030 -825
rect 8250 -845 8270 -825
rect 8490 -845 8510 -825
rect 8730 -845 8750 -825
rect 8970 -845 8990 -825
rect 9505 -805 9525 -785
rect 9625 -805 9645 -785
rect 9745 -805 9765 -785
rect 9865 -805 9885 -785
rect 9985 -805 10005 -785
rect 10105 -805 10125 -785
rect 10225 -805 10245 -785
rect 10345 -805 10365 -785
rect 10465 -805 10485 -785
rect 10585 -805 10605 -785
rect 10705 -805 10725 -785
rect 10825 -805 10845 -785
rect 10945 -805 10965 -785
rect 11065 -805 11085 -785
rect 11185 -805 11205 -785
rect 11305 -805 11325 -785
rect 11425 -805 11445 -785
rect 11545 -805 11565 -785
rect 9210 -845 9230 -825
rect 9440 -870 9475 -835
rect 9690 -845 9710 -825
rect 9930 -845 9950 -825
rect 10170 -845 10190 -825
rect 10410 -845 10430 -825
rect 10650 -845 10670 -825
rect 10890 -845 10910 -825
rect 11130 -845 11150 -825
rect 11665 -805 11685 -785
rect 11785 -805 11805 -785
rect 11905 -805 11925 -785
rect 12025 -805 12045 -785
rect 12145 -805 12165 -785
rect 12265 -805 12285 -785
rect 12385 -805 12405 -785
rect 12505 -805 12525 -785
rect 12625 -805 12645 -785
rect 12745 -805 12765 -785
rect 12865 -805 12885 -785
rect 12985 -805 13005 -785
rect 13105 -805 13125 -785
rect 13225 -805 13245 -785
rect 13345 -805 13365 -785
rect 13465 -805 13485 -785
rect 13585 -805 13605 -785
rect 13705 -805 13725 -785
rect 11370 -845 11390 -825
rect 11600 -870 11635 -835
rect 11850 -845 11870 -825
rect 12090 -845 12110 -825
rect 12330 -845 12350 -825
rect 12570 -845 12590 -825
rect 12810 -845 12830 -825
rect 13050 -845 13070 -825
rect 13290 -845 13310 -825
rect 13825 -805 13845 -785
rect 13945 -805 13965 -785
rect 14065 -805 14085 -785
rect 14185 -805 14205 -785
rect 14305 -805 14325 -785
rect 14425 -805 14445 -785
rect 14545 -805 14565 -785
rect 14665 -805 14685 -785
rect 14785 -805 14805 -785
rect 14905 -805 14925 -785
rect 15025 -805 15045 -785
rect 15145 -805 15165 -785
rect 15265 -805 15285 -785
rect 15385 -805 15405 -785
rect 15505 -805 15525 -785
rect 15625 -805 15645 -785
rect 15745 -805 15765 -785
rect 15865 -805 15885 -785
rect 13530 -845 13550 -825
rect 13760 -870 13795 -835
rect 14010 -845 14030 -825
rect 14250 -845 14270 -825
rect 14490 -845 14510 -825
rect 14730 -845 14750 -825
rect 14970 -845 14990 -825
rect 15210 -845 15230 -825
rect 15450 -845 15470 -825
rect 15985 -805 16005 -785
rect 16105 -805 16125 -785
rect 16225 -805 16245 -785
rect 16345 -805 16365 -785
rect 16465 -805 16485 -785
rect 16585 -805 16605 -785
rect 16705 -805 16725 -785
rect 16825 -805 16845 -785
rect 16945 -805 16965 -785
rect 17065 -805 17085 -785
rect 17185 -805 17205 -785
rect 17305 -805 17325 -785
rect 17425 -805 17445 -785
rect 17545 -805 17565 -785
rect 17665 -805 17685 -785
rect 17785 -805 17805 -785
rect 17905 -805 17925 -785
rect 18025 -805 18045 -785
rect 15690 -845 15710 -825
rect 15920 -870 15955 -835
rect 16170 -845 16190 -825
rect 16410 -845 16430 -825
rect 16650 -845 16670 -825
rect 16890 -845 16910 -825
rect 17130 -845 17150 -825
rect 17370 -845 17390 -825
rect 17610 -845 17630 -825
rect 18145 -805 18165 -785
rect 18265 -805 18285 -785
rect 18385 -805 18405 -785
rect 18505 -805 18525 -785
rect 18625 -805 18645 -785
rect 18745 -805 18765 -785
rect 18865 -805 18885 -785
rect 18985 -805 19005 -785
rect 19105 -805 19125 -785
rect 19225 -805 19245 -785
rect 19345 -805 19365 -785
rect 19465 -805 19485 -785
rect 19585 -805 19605 -785
rect 19705 -805 19725 -785
rect 19825 -805 19845 -785
rect 19945 -805 19965 -785
rect 20065 -805 20085 -785
rect 20185 -805 20205 -785
rect 17850 -845 17870 -825
rect 18080 -870 18115 -835
rect 18330 -845 18350 -825
rect 18570 -845 18590 -825
rect 18810 -845 18830 -825
rect 19050 -845 19070 -825
rect 19290 -845 19310 -825
rect 19530 -845 19550 -825
rect 19770 -845 19790 -825
rect 20305 -805 20325 -785
rect 20425 -805 20445 -785
rect 20545 -805 20565 -785
rect 20665 -805 20685 -785
rect 20785 -805 20805 -785
rect 20905 -805 20925 -785
rect 21025 -805 21045 -785
rect 21145 -805 21165 -785
rect 21265 -805 21285 -785
rect 21385 -805 21405 -785
rect 21505 -805 21525 -785
rect 21625 -805 21645 -785
rect 21745 -805 21765 -785
rect 21865 -805 21885 -785
rect 21985 -805 22005 -785
rect 22105 -805 22125 -785
rect 22225 -805 22245 -785
rect 22345 -805 22365 -785
rect 20010 -845 20030 -825
rect 20240 -870 20275 -835
rect 20490 -845 20510 -825
rect 20730 -845 20750 -825
rect 20970 -845 20990 -825
rect 21210 -845 21230 -825
rect 21450 -845 21470 -825
rect 21690 -845 21710 -825
rect 21930 -845 21950 -825
rect 22465 -805 22485 -785
rect 22585 -805 22605 -785
rect 22705 -805 22725 -785
rect 22825 -805 22845 -785
rect 22945 -805 22965 -785
rect 23065 -805 23085 -785
rect 23185 -805 23205 -785
rect 23305 -805 23325 -785
rect 23425 -805 23445 -785
rect 23545 -805 23565 -785
rect 23665 -805 23685 -785
rect 23785 -805 23805 -785
rect 23905 -805 23925 -785
rect 24025 -805 24045 -785
rect 24145 -805 24165 -785
rect 24265 -805 24285 -785
rect 22170 -845 22190 -825
rect 22400 -870 22435 -835
rect 22650 -845 22670 -825
rect 22890 -845 22910 -825
rect 23130 -845 23150 -825
rect 23370 -845 23390 -825
rect 23610 -845 23630 -825
rect 23850 -845 23870 -825
rect 24385 -805 24405 -785
rect 24505 -805 24525 -785
rect 24625 -805 24645 -785
rect 24745 -805 24765 -785
rect 24865 -805 24885 -785
rect 24985 -805 25005 -785
rect 25105 -805 25125 -785
rect 25225 -805 25245 -785
rect 25345 -805 25365 -785
rect 25465 -805 25485 -785
rect 25585 -805 25605 -785
rect 25705 -805 25725 -785
rect 25825 -805 25845 -785
rect 25945 -805 25965 -785
rect 26065 -805 26085 -785
rect 26185 -805 26205 -785
rect 24090 -845 24110 -825
rect 24320 -870 24355 -835
rect 24570 -845 24590 -825
rect 24810 -845 24830 -825
rect 25050 -845 25070 -825
rect 25290 -845 25310 -825
rect 25530 -845 25550 -825
rect 25770 -845 25790 -825
rect 26305 -805 26325 -785
rect 26425 -805 26445 -785
rect 26545 -805 26565 -785
rect 26665 -805 26685 -785
rect 26785 -805 26805 -785
rect 26905 -805 26925 -785
rect 27025 -805 27045 -785
rect 27145 -805 27165 -785
rect 27265 -805 27285 -785
rect 27385 -805 27405 -785
rect 27505 -805 27525 -785
rect 27625 -805 27645 -785
rect 27745 -805 27765 -785
rect 27865 -805 27885 -785
rect 27985 -805 28005 -785
rect 28105 -805 28125 -785
rect 26010 -845 26030 -825
rect 26240 -870 26275 -835
rect 26490 -845 26510 -825
rect 26730 -845 26750 -825
rect 26970 -845 26990 -825
rect 27210 -845 27230 -825
rect 27450 -845 27470 -825
rect 27690 -845 27710 -825
rect 28225 -805 28245 -785
rect 28345 -805 28365 -785
rect 28465 -805 28485 -785
rect 28585 -805 28605 -785
rect 28705 -805 28725 -785
rect 28825 -805 28845 -785
rect 28945 -805 28965 -785
rect 29065 -805 29085 -785
rect 29185 -805 29205 -785
rect 29305 -805 29325 -785
rect 29425 -805 29445 -785
rect 29545 -805 29565 -785
rect 29665 -805 29685 -785
rect 29785 -805 29805 -785
rect 27930 -845 27950 -825
rect 28160 -870 28195 -835
rect 28410 -845 28430 -825
rect 28650 -845 28670 -825
rect 28890 -845 28910 -825
rect 29130 -845 29150 -825
rect 29370 -845 29390 -825
rect 29905 -805 29925 -785
rect 30025 -805 30045 -785
rect 30145 -805 30165 -785
rect 30265 -805 30285 -785
rect 30385 -805 30405 -785
rect 30505 -805 30525 -785
rect 30625 -805 30645 -785
rect 29610 -845 29630 -825
rect 29840 -870 29875 -835
rect 30090 -845 30110 -825
rect 30330 -845 30350 -825
rect 30570 -845 30590 -825
<< metal1 >>
rect 2255 305 2310 315
rect 185 275 240 285
rect 185 240 195 275
rect 230 240 240 275
rect 2255 270 2265 305
rect 2300 270 2310 305
rect 4195 305 4250 315
rect 4195 270 4205 305
rect 4240 270 4250 305
rect 6445 305 6500 315
rect 6445 270 6455 305
rect 6490 270 6500 305
rect 9350 305 9405 315
rect 9350 270 9360 305
rect 9395 270 9405 305
rect 11295 305 11350 315
rect 11295 270 11305 305
rect 11340 270 11350 305
rect 12990 305 13045 315
rect 12990 270 13000 305
rect 13035 270 13045 305
rect 15175 305 15230 315
rect 15175 270 15185 305
rect 15220 270 15230 305
rect 17355 305 17410 315
rect 17355 270 17365 305
rect 17400 270 17410 305
rect 19540 305 19595 315
rect 19540 270 19550 305
rect 19585 270 19595 305
rect 20750 305 20805 315
rect 20750 270 20760 305
rect 20795 270 20805 305
rect 185 230 240 240
rect 431 265 471 270
rect 431 235 436 265
rect 466 235 471 265
rect 431 230 471 235
rect 736 265 776 270
rect 736 235 741 265
rect 771 235 776 265
rect 736 230 776 235
rect 981 265 1021 270
rect 981 235 986 265
rect 1016 235 1021 265
rect 981 230 1021 235
rect 1221 265 1261 270
rect 1221 235 1226 265
rect 1256 235 1261 265
rect 1221 230 1261 235
rect 1466 265 1506 270
rect 1466 235 1471 265
rect 1501 235 1506 265
rect 1466 230 1506 235
rect 1771 265 1811 270
rect 1771 235 1776 265
rect 1806 235 1811 265
rect 1771 230 1811 235
rect 2016 265 2056 270
rect 2016 235 2021 265
rect 2051 235 2056 265
rect 2255 260 2310 270
rect 2501 265 2541 270
rect 2016 230 2056 235
rect 2501 235 2506 265
rect 2536 235 2541 265
rect 2501 230 2541 235
rect 2741 265 2781 270
rect 2741 235 2746 265
rect 2776 235 2781 265
rect 2741 230 2781 235
rect 2986 265 3026 270
rect 2986 235 2991 265
rect 3021 235 3026 265
rect 2986 230 3026 235
rect 3226 265 3266 270
rect 3226 235 3231 265
rect 3261 235 3266 265
rect 3226 230 3266 235
rect 3471 265 3511 270
rect 3471 235 3476 265
rect 3506 235 3511 265
rect 3471 230 3511 235
rect 3711 265 3751 270
rect 3711 235 3716 265
rect 3746 235 3751 265
rect 3711 230 3751 235
rect 3956 265 3996 270
rect 3956 235 3961 265
rect 3991 235 3996 265
rect 4195 260 4250 270
rect 4441 265 4481 270
rect 3956 230 3996 235
rect 4441 235 4446 265
rect 4476 235 4481 265
rect 4441 230 4481 235
rect 4681 265 4721 270
rect 4681 235 4686 265
rect 4716 235 4721 265
rect 4681 230 4721 235
rect 4926 265 4966 270
rect 4926 235 4931 265
rect 4961 235 4966 265
rect 4926 230 4966 235
rect 5166 265 5206 270
rect 5166 235 5171 265
rect 5201 235 5206 265
rect 5166 230 5206 235
rect 5411 265 5451 270
rect 5411 235 5416 265
rect 5446 235 5451 265
rect 5411 230 5451 235
rect 5716 265 5756 270
rect 5716 235 5721 265
rect 5751 235 5756 265
rect 5716 230 5756 235
rect 5961 265 6001 270
rect 5961 235 5966 265
rect 5996 235 6001 265
rect 5961 230 6001 235
rect 6201 265 6241 270
rect 6201 235 6206 265
rect 6236 235 6241 265
rect 6445 260 6500 270
rect 6686 265 6726 270
rect 6201 230 6241 235
rect 6686 235 6691 265
rect 6721 235 6726 265
rect 6686 230 6726 235
rect 6931 265 6971 270
rect 6931 235 6936 265
rect 6966 235 6971 265
rect 6931 230 6971 235
rect 7171 265 7211 270
rect 7171 235 7176 265
rect 7206 235 7211 265
rect 7171 230 7211 235
rect 7411 265 7451 270
rect 7411 235 7416 265
rect 7446 235 7451 265
rect 7411 230 7451 235
rect 7651 265 7691 270
rect 7651 235 7656 265
rect 7686 235 7691 265
rect 7651 230 7691 235
rect 7896 265 7936 270
rect 7896 235 7901 265
rect 7931 235 7936 265
rect 7896 230 7936 235
rect 8136 265 8176 270
rect 8136 235 8141 265
rect 8171 235 8176 265
rect 8136 230 8176 235
rect 8381 265 8421 270
rect 8381 235 8386 265
rect 8416 235 8421 265
rect 8381 230 8421 235
rect 8621 265 8661 270
rect 8621 235 8626 265
rect 8656 235 8661 265
rect 8621 230 8661 235
rect 8866 265 8906 270
rect 8866 235 8871 265
rect 8901 235 8906 265
rect 8866 230 8906 235
rect 9106 265 9146 270
rect 9106 235 9111 265
rect 9141 235 9146 265
rect 9350 260 9405 270
rect 9596 265 9636 270
rect 9106 230 9146 235
rect 9596 235 9601 265
rect 9631 235 9636 265
rect 9596 230 9636 235
rect 9841 265 9881 270
rect 9841 235 9846 265
rect 9876 235 9881 265
rect 9841 230 9881 235
rect 10081 265 10121 270
rect 10081 235 10086 265
rect 10116 235 10121 265
rect 10081 230 10121 235
rect 10326 265 10366 270
rect 10326 235 10331 265
rect 10361 235 10366 265
rect 10326 230 10366 235
rect 10566 265 10606 270
rect 10566 235 10571 265
rect 10601 235 10606 265
rect 10566 230 10606 235
rect 10811 265 10851 270
rect 10811 235 10816 265
rect 10846 235 10851 265
rect 10811 230 10851 235
rect 11051 265 11091 270
rect 11051 235 11056 265
rect 11086 235 11091 265
rect 11295 260 11350 270
rect 11536 265 11576 270
rect 11051 230 11091 235
rect 11536 235 11541 265
rect 11571 235 11576 265
rect 11536 230 11576 235
rect 11781 265 11821 270
rect 11781 235 11786 265
rect 11816 235 11821 265
rect 11781 230 11821 235
rect 12021 265 12061 270
rect 12021 235 12026 265
rect 12056 235 12061 265
rect 12021 230 12061 235
rect 12266 265 12306 270
rect 12266 235 12271 265
rect 12301 235 12306 265
rect 12266 230 12306 235
rect 12506 265 12546 270
rect 12506 235 12511 265
rect 12541 235 12546 265
rect 12506 230 12546 235
rect 12751 265 12791 270
rect 12751 235 12756 265
rect 12786 235 12791 265
rect 12990 260 13045 270
rect 13236 265 13276 270
rect 12751 230 12791 235
rect 13236 235 13241 265
rect 13271 235 13276 265
rect 13236 230 13276 235
rect 13476 265 13516 270
rect 13476 235 13481 265
rect 13511 235 13516 265
rect 13476 230 13516 235
rect 13721 265 13761 270
rect 13721 235 13726 265
rect 13756 235 13761 265
rect 13721 230 13761 235
rect 13961 265 14001 270
rect 13961 235 13966 265
rect 13996 235 14001 265
rect 13961 230 14001 235
rect 14206 265 14246 270
rect 14206 235 14211 265
rect 14241 235 14246 265
rect 14206 230 14246 235
rect 14446 265 14486 270
rect 14446 235 14451 265
rect 14481 235 14486 265
rect 14446 230 14486 235
rect 14691 265 14731 270
rect 14691 235 14696 265
rect 14726 235 14731 265
rect 14691 230 14731 235
rect 14931 265 14971 270
rect 14931 235 14936 265
rect 14966 235 14971 265
rect 15175 260 15230 270
rect 15416 265 15456 270
rect 14931 230 14971 235
rect 15416 235 15421 265
rect 15451 235 15456 265
rect 15416 230 15456 235
rect 15661 265 15701 270
rect 15661 235 15666 265
rect 15696 235 15701 265
rect 15661 230 15701 235
rect 15901 265 15941 270
rect 15901 235 15906 265
rect 15936 235 15941 265
rect 15901 230 15941 235
rect 16146 265 16186 270
rect 16146 235 16151 265
rect 16181 235 16186 265
rect 16146 230 16186 235
rect 16386 265 16426 270
rect 16386 235 16391 265
rect 16421 235 16426 265
rect 16386 230 16426 235
rect 16631 265 16671 270
rect 16631 235 16636 265
rect 16666 235 16671 265
rect 16631 230 16671 235
rect 16871 265 16911 270
rect 16871 235 16876 265
rect 16906 235 16911 265
rect 16871 230 16911 235
rect 17116 265 17156 270
rect 17116 235 17121 265
rect 17151 235 17156 265
rect 17355 260 17410 270
rect 17601 265 17641 270
rect 17116 230 17156 235
rect 17601 235 17606 265
rect 17636 235 17641 265
rect 17601 230 17641 235
rect 17841 265 17881 270
rect 17841 235 17846 265
rect 17876 235 17881 265
rect 17841 230 17881 235
rect 18086 265 18126 270
rect 18086 235 18091 265
rect 18121 235 18126 265
rect 18086 230 18126 235
rect 18326 265 18366 270
rect 18326 235 18331 265
rect 18361 235 18366 265
rect 18326 230 18366 235
rect 18571 265 18611 270
rect 18571 235 18576 265
rect 18606 235 18611 265
rect 18571 230 18611 235
rect 18811 265 18851 270
rect 18811 235 18816 265
rect 18846 235 18851 265
rect 18811 230 18851 235
rect 19056 265 19096 270
rect 19056 235 19061 265
rect 19091 235 19096 265
rect 19056 230 19096 235
rect 19296 265 19336 270
rect 19296 235 19301 265
rect 19331 235 19336 265
rect 19540 260 19595 270
rect 19781 265 19821 270
rect 19296 230 19336 235
rect 19781 235 19786 265
rect 19816 235 19821 265
rect 19781 230 19821 235
rect 20026 265 20066 270
rect 20026 235 20031 265
rect 20061 235 20066 265
rect 20026 230 20066 235
rect 20266 265 20306 270
rect 20266 235 20271 265
rect 20301 235 20306 265
rect 20266 230 20306 235
rect 20511 265 20551 270
rect 20511 235 20516 265
rect 20546 235 20551 265
rect 20750 260 20805 270
rect 20996 265 21036 270
rect 20511 230 20551 235
rect 20996 235 21001 265
rect 21031 235 21036 265
rect 20996 230 21036 235
rect 376 220 416 230
rect 376 200 386 220
rect 406 205 416 220
rect 496 220 536 230
rect 496 205 506 220
rect 406 200 506 205
rect 526 200 536 220
rect 376 190 536 200
rect 681 220 721 230
rect 681 200 691 220
rect 711 205 721 220
rect 801 220 841 230
rect 801 205 811 220
rect 711 200 811 205
rect 831 205 841 220
rect 926 220 966 230
rect 926 205 936 220
rect 831 200 936 205
rect 956 205 966 220
rect 1046 220 1086 230
rect 1046 205 1056 220
rect 956 200 1056 205
rect 1076 205 1086 220
rect 1166 220 1206 230
rect 1166 205 1176 220
rect 1076 200 1176 205
rect 1196 205 1206 220
rect 1286 220 1326 230
rect 1286 205 1296 220
rect 1196 200 1296 205
rect 1316 205 1326 220
rect 1411 220 1451 230
rect 1411 205 1421 220
rect 1316 200 1421 205
rect 1441 205 1451 220
rect 1531 220 1571 230
rect 1531 205 1541 220
rect 1441 200 1541 205
rect 1561 200 1571 220
rect 1716 220 1756 230
rect 1716 205 1726 220
rect 681 190 1571 200
rect 1715 200 1726 205
rect 1746 205 1756 220
rect 1836 220 1876 230
rect 1836 205 1846 220
rect 1746 200 1846 205
rect 1866 205 1876 220
rect 1961 220 2001 230
rect 1961 205 1971 220
rect 1866 200 1971 205
rect 1991 205 2001 220
rect 2081 220 2121 230
rect 2081 205 2091 220
rect 1991 200 2091 205
rect 2111 205 2121 220
rect 2201 220 2241 230
rect 2201 205 2211 220
rect 2111 200 2211 205
rect 2231 205 2241 220
rect 2321 220 2361 230
rect 2321 205 2331 220
rect 2231 200 2331 205
rect 2351 205 2361 220
rect 2446 220 2486 230
rect 2446 205 2456 220
rect 2351 200 2456 205
rect 2476 205 2486 220
rect 2566 220 2606 230
rect 2566 205 2576 220
rect 2476 200 2576 205
rect 2596 205 2606 220
rect 2686 220 2726 230
rect 2686 205 2696 220
rect 2596 200 2696 205
rect 2716 205 2726 220
rect 2806 220 2846 230
rect 2806 205 2816 220
rect 2716 200 2816 205
rect 2836 205 2846 220
rect 2931 220 2971 230
rect 2931 205 2941 220
rect 2836 200 2941 205
rect 2961 205 2971 220
rect 3051 220 3091 230
rect 3051 205 3061 220
rect 2961 200 3061 205
rect 3081 205 3091 220
rect 3171 220 3211 230
rect 3171 205 3181 220
rect 3081 200 3181 205
rect 3201 205 3211 220
rect 3291 220 3331 230
rect 3291 205 3301 220
rect 3201 200 3301 205
rect 3321 205 3331 220
rect 3416 220 3456 230
rect 3416 205 3426 220
rect 3321 200 3426 205
rect 3446 205 3456 220
rect 3536 220 3576 230
rect 3536 205 3546 220
rect 3446 200 3546 205
rect 3566 205 3576 220
rect 3656 220 3696 230
rect 3656 205 3666 220
rect 3566 200 3666 205
rect 3686 205 3696 220
rect 3776 220 3816 230
rect 3776 205 3786 220
rect 3686 200 3786 205
rect 3806 205 3816 220
rect 3901 220 3941 230
rect 3901 205 3911 220
rect 3806 200 3911 205
rect 3931 205 3941 220
rect 4021 220 4061 230
rect 4021 205 4031 220
rect 3931 200 4031 205
rect 4051 205 4061 220
rect 4141 220 4181 230
rect 4141 205 4151 220
rect 4051 200 4151 205
rect 4171 205 4181 220
rect 4261 220 4301 230
rect 4261 205 4271 220
rect 4171 200 4271 205
rect 4291 205 4301 220
rect 4386 220 4426 230
rect 4386 205 4396 220
rect 4291 200 4396 205
rect 4416 205 4426 220
rect 4506 220 4546 230
rect 4506 205 4516 220
rect 4416 200 4516 205
rect 4536 205 4546 220
rect 4626 220 4666 230
rect 4626 205 4636 220
rect 4536 200 4636 205
rect 4656 205 4666 220
rect 4746 220 4786 230
rect 4746 205 4756 220
rect 4656 200 4756 205
rect 4776 205 4786 220
rect 4871 220 4911 230
rect 4871 205 4881 220
rect 4776 200 4881 205
rect 4901 205 4911 220
rect 4991 220 5031 230
rect 4991 205 5001 220
rect 4901 200 5001 205
rect 5021 205 5031 220
rect 5111 220 5151 230
rect 5111 205 5121 220
rect 5021 200 5121 205
rect 5141 205 5151 220
rect 5231 220 5271 230
rect 5231 205 5241 220
rect 5141 200 5241 205
rect 5261 205 5271 220
rect 5356 220 5396 230
rect 5356 205 5366 220
rect 5261 200 5366 205
rect 5386 205 5396 220
rect 5476 220 5516 230
rect 5476 205 5486 220
rect 5386 200 5486 205
rect 5506 205 5516 220
rect 5661 220 5701 230
rect 5661 205 5671 220
rect 5506 200 5520 205
rect 1715 190 5520 200
rect 5660 200 5671 205
rect 5691 205 5701 220
rect 5781 220 5821 230
rect 5781 205 5791 220
rect 5691 200 5791 205
rect 5811 205 5821 220
rect 5906 220 5946 230
rect 5906 205 5916 220
rect 5811 200 5916 205
rect 5936 205 5946 220
rect 6026 220 6066 230
rect 6026 205 6036 220
rect 5936 200 6036 205
rect 6056 205 6066 220
rect 6146 220 6186 230
rect 6146 205 6156 220
rect 6056 200 6156 205
rect 6176 205 6186 220
rect 6266 220 6306 230
rect 6266 205 6276 220
rect 6176 200 6276 205
rect 6296 205 6306 220
rect 6391 220 6431 230
rect 6391 205 6401 220
rect 6296 200 6401 205
rect 6421 205 6431 220
rect 6511 220 6551 230
rect 6511 205 6521 220
rect 6421 200 6521 205
rect 6541 205 6551 220
rect 6631 220 6671 230
rect 6631 205 6641 220
rect 6541 200 6641 205
rect 6661 205 6671 220
rect 6751 220 6791 230
rect 6751 205 6761 220
rect 6661 200 6761 205
rect 6781 205 6791 220
rect 6876 220 6916 230
rect 6876 205 6886 220
rect 6781 200 6886 205
rect 6906 205 6916 220
rect 6996 220 7036 230
rect 6996 205 7006 220
rect 6906 200 7006 205
rect 7026 205 7036 220
rect 7116 220 7156 230
rect 7116 205 7126 220
rect 7026 200 7126 205
rect 7146 205 7156 220
rect 7236 220 7276 230
rect 7236 205 7246 220
rect 7146 200 7246 205
rect 7266 205 7276 220
rect 7356 220 7396 230
rect 7356 205 7366 220
rect 7266 200 7366 205
rect 7386 205 7396 220
rect 7476 220 7516 230
rect 7476 205 7486 220
rect 7386 200 7486 205
rect 7506 205 7516 220
rect 7596 220 7636 230
rect 7596 205 7606 220
rect 7506 200 7606 205
rect 7626 205 7636 220
rect 7716 220 7756 230
rect 7716 205 7726 220
rect 7626 200 7726 205
rect 7746 205 7756 220
rect 7841 220 7881 230
rect 7841 205 7851 220
rect 7746 200 7851 205
rect 7871 205 7881 220
rect 7961 220 8001 230
rect 7961 205 7971 220
rect 7871 200 7971 205
rect 7991 205 8001 220
rect 8081 220 8121 230
rect 8081 205 8091 220
rect 7991 200 8091 205
rect 8111 205 8121 220
rect 8201 220 8241 230
rect 8201 205 8211 220
rect 8111 200 8211 205
rect 8231 205 8241 220
rect 8326 220 8366 230
rect 8326 205 8336 220
rect 8231 200 8336 205
rect 8356 205 8366 220
rect 8446 220 8486 230
rect 8446 205 8456 220
rect 8356 200 8456 205
rect 8476 205 8486 220
rect 8566 220 8606 230
rect 8566 205 8576 220
rect 8476 200 8576 205
rect 8596 205 8606 220
rect 8686 220 8726 230
rect 8686 205 8696 220
rect 8596 200 8696 205
rect 8716 205 8726 220
rect 8811 220 8851 230
rect 8811 205 8821 220
rect 8716 200 8821 205
rect 8841 205 8851 220
rect 8931 220 8971 230
rect 8931 205 8941 220
rect 8841 200 8941 205
rect 8961 205 8971 220
rect 9051 220 9091 230
rect 9051 205 9061 220
rect 8961 200 9061 205
rect 9081 205 9091 220
rect 9171 220 9211 230
rect 9171 205 9181 220
rect 9081 200 9181 205
rect 9201 205 9211 220
rect 9296 220 9336 230
rect 9296 205 9306 220
rect 9201 200 9306 205
rect 9326 205 9336 220
rect 9416 220 9456 230
rect 9416 205 9426 220
rect 9326 200 9426 205
rect 9446 205 9456 220
rect 9541 220 9581 230
rect 9541 205 9551 220
rect 9446 200 9551 205
rect 9571 205 9581 220
rect 9661 220 9701 230
rect 9661 205 9671 220
rect 9571 200 9671 205
rect 9691 205 9701 220
rect 9786 220 9826 230
rect 9786 205 9796 220
rect 9691 200 9796 205
rect 9816 205 9826 220
rect 9906 220 9946 230
rect 9906 205 9916 220
rect 9816 200 9916 205
rect 9936 205 9946 220
rect 10026 220 10066 230
rect 10026 205 10036 220
rect 9936 200 10036 205
rect 10056 205 10066 220
rect 10146 220 10186 230
rect 10146 205 10156 220
rect 10056 200 10156 205
rect 10176 205 10186 220
rect 10271 220 10311 230
rect 10271 205 10281 220
rect 10176 200 10281 205
rect 10301 205 10311 220
rect 10391 220 10431 230
rect 10391 205 10401 220
rect 10301 200 10401 205
rect 10421 205 10431 220
rect 10511 220 10551 230
rect 10511 205 10521 220
rect 10421 200 10521 205
rect 10541 205 10551 220
rect 10631 220 10671 230
rect 10631 205 10641 220
rect 10541 200 10641 205
rect 10661 205 10671 220
rect 10756 220 10796 230
rect 10756 205 10766 220
rect 10661 200 10766 205
rect 10786 205 10796 220
rect 10876 220 10916 230
rect 10876 205 10886 220
rect 10786 200 10886 205
rect 10906 205 10916 220
rect 10996 220 11036 230
rect 10996 205 11006 220
rect 10906 200 11006 205
rect 11026 205 11036 220
rect 11116 220 11156 230
rect 11116 205 11126 220
rect 11026 200 11126 205
rect 11146 205 11156 220
rect 11241 220 11281 230
rect 11241 205 11251 220
rect 11146 200 11251 205
rect 11271 205 11281 220
rect 11361 220 11401 230
rect 11361 205 11371 220
rect 11271 200 11371 205
rect 11391 205 11401 220
rect 11481 220 11521 230
rect 11481 205 11491 220
rect 11391 200 11491 205
rect 11511 205 11521 220
rect 11601 220 11641 230
rect 11601 205 11611 220
rect 11511 200 11611 205
rect 11631 205 11641 220
rect 11726 220 11766 230
rect 11726 205 11736 220
rect 11631 200 11736 205
rect 11756 205 11766 220
rect 11846 220 11886 230
rect 11846 205 11856 220
rect 11756 200 11856 205
rect 11876 205 11886 220
rect 11966 220 12006 230
rect 11966 205 11976 220
rect 11876 200 11976 205
rect 11996 205 12006 220
rect 12086 220 12126 230
rect 12086 205 12096 220
rect 11996 200 12096 205
rect 12116 205 12126 220
rect 12211 220 12251 230
rect 12211 205 12221 220
rect 12116 200 12221 205
rect 12241 205 12251 220
rect 12331 220 12371 230
rect 12331 205 12341 220
rect 12241 200 12341 205
rect 12361 205 12371 220
rect 12451 220 12491 230
rect 12451 205 12461 220
rect 12361 200 12461 205
rect 12481 205 12491 220
rect 12571 220 12611 230
rect 12571 205 12581 220
rect 12481 200 12581 205
rect 12601 205 12611 220
rect 12696 220 12736 230
rect 12696 205 12706 220
rect 12601 200 12706 205
rect 12726 205 12736 220
rect 12816 220 12856 230
rect 12816 205 12826 220
rect 12726 200 12826 205
rect 12846 205 12856 220
rect 12936 220 12976 230
rect 12936 205 12946 220
rect 12846 200 12946 205
rect 12966 205 12976 220
rect 13056 220 13096 230
rect 13056 205 13066 220
rect 12966 200 13066 205
rect 13086 205 13096 220
rect 13181 220 13221 230
rect 13181 205 13191 220
rect 13086 200 13191 205
rect 13211 205 13221 220
rect 13301 220 13341 230
rect 13301 205 13311 220
rect 13211 200 13311 205
rect 13331 205 13341 220
rect 13421 220 13461 230
rect 13421 205 13431 220
rect 13331 200 13431 205
rect 13451 205 13461 220
rect 13541 220 13581 230
rect 13541 205 13551 220
rect 13451 200 13551 205
rect 13571 205 13581 220
rect 13666 220 13706 230
rect 13666 205 13676 220
rect 13571 200 13676 205
rect 13696 205 13706 220
rect 13786 220 13826 230
rect 13786 205 13796 220
rect 13696 200 13796 205
rect 13816 205 13826 220
rect 13906 220 13946 230
rect 13906 205 13916 220
rect 13816 200 13916 205
rect 13936 205 13946 220
rect 14026 220 14066 230
rect 14026 205 14036 220
rect 13936 200 14036 205
rect 14056 205 14066 220
rect 14151 220 14191 230
rect 14151 205 14161 220
rect 14056 200 14161 205
rect 14181 205 14191 220
rect 14271 220 14311 230
rect 14271 205 14281 220
rect 14181 200 14281 205
rect 14301 205 14311 220
rect 14391 220 14431 230
rect 14391 205 14401 220
rect 14301 200 14401 205
rect 14421 205 14431 220
rect 14511 220 14551 230
rect 14511 205 14521 220
rect 14421 200 14521 205
rect 14541 205 14551 220
rect 14636 220 14676 230
rect 14636 205 14646 220
rect 14541 200 14646 205
rect 14666 205 14676 220
rect 14756 220 14796 230
rect 14756 205 14766 220
rect 14666 200 14766 205
rect 14786 205 14796 220
rect 14876 220 14916 230
rect 14876 205 14886 220
rect 14786 200 14886 205
rect 14906 205 14916 220
rect 14996 220 15036 230
rect 14996 205 15006 220
rect 14906 200 15006 205
rect 15026 205 15036 220
rect 15121 220 15161 230
rect 15121 205 15131 220
rect 15026 200 15131 205
rect 15151 205 15161 220
rect 15241 220 15281 230
rect 15241 205 15251 220
rect 15151 200 15251 205
rect 15271 205 15281 220
rect 15361 220 15401 230
rect 15361 205 15371 220
rect 15271 200 15371 205
rect 15391 205 15401 220
rect 15481 220 15521 230
rect 15481 205 15491 220
rect 15391 200 15491 205
rect 15511 205 15521 220
rect 15606 220 15646 230
rect 15606 205 15616 220
rect 15511 200 15616 205
rect 15636 205 15646 220
rect 15726 220 15766 230
rect 15726 205 15736 220
rect 15636 200 15736 205
rect 15756 205 15766 220
rect 15846 220 15886 230
rect 15846 205 15856 220
rect 15756 200 15856 205
rect 15876 205 15886 220
rect 15966 220 16006 230
rect 15966 205 15976 220
rect 15876 200 15976 205
rect 15996 205 16006 220
rect 16091 220 16131 230
rect 16091 205 16101 220
rect 15996 200 16101 205
rect 16121 205 16131 220
rect 16211 220 16251 230
rect 16211 205 16221 220
rect 16121 200 16221 205
rect 16241 205 16251 220
rect 16331 220 16371 230
rect 16331 205 16341 220
rect 16241 200 16341 205
rect 16361 205 16371 220
rect 16451 220 16491 230
rect 16451 205 16461 220
rect 16361 200 16461 205
rect 16481 205 16491 220
rect 16576 220 16616 230
rect 16576 205 16586 220
rect 16481 200 16586 205
rect 16606 205 16616 220
rect 16696 220 16736 230
rect 16696 205 16706 220
rect 16606 200 16706 205
rect 16726 205 16736 220
rect 16816 220 16856 230
rect 16816 205 16826 220
rect 16726 200 16826 205
rect 16846 205 16856 220
rect 16936 220 16976 230
rect 16936 205 16946 220
rect 16846 200 16946 205
rect 16966 205 16976 220
rect 17061 220 17101 230
rect 17061 205 17071 220
rect 16966 200 17071 205
rect 17091 205 17101 220
rect 17181 220 17221 230
rect 17181 205 17191 220
rect 17091 200 17191 205
rect 17211 205 17221 220
rect 17301 220 17341 230
rect 17301 205 17311 220
rect 17211 200 17311 205
rect 17331 205 17341 220
rect 17421 220 17461 230
rect 17421 205 17431 220
rect 17331 200 17431 205
rect 17451 205 17461 220
rect 17546 220 17586 230
rect 17546 205 17556 220
rect 17451 200 17556 205
rect 17576 205 17586 220
rect 17666 220 17706 230
rect 17666 205 17676 220
rect 17576 200 17676 205
rect 17696 205 17706 220
rect 17786 220 17826 230
rect 17786 205 17796 220
rect 17696 200 17796 205
rect 17816 205 17826 220
rect 17906 220 17946 230
rect 17906 205 17916 220
rect 17816 200 17916 205
rect 17936 205 17946 220
rect 18031 220 18071 230
rect 18031 205 18041 220
rect 17936 200 18041 205
rect 18061 205 18071 220
rect 18151 220 18191 230
rect 18151 205 18161 220
rect 18061 200 18161 205
rect 18181 205 18191 220
rect 18271 220 18311 230
rect 18271 205 18281 220
rect 18181 200 18281 205
rect 18301 205 18311 220
rect 18391 220 18431 230
rect 18391 205 18401 220
rect 18301 200 18401 205
rect 18421 205 18431 220
rect 18516 220 18556 230
rect 18516 205 18526 220
rect 18421 200 18526 205
rect 18546 205 18556 220
rect 18636 220 18676 230
rect 18636 205 18646 220
rect 18546 200 18646 205
rect 18666 205 18676 220
rect 18756 220 18796 230
rect 18756 205 18766 220
rect 18666 200 18766 205
rect 18786 205 18796 220
rect 18876 220 18916 230
rect 18876 205 18886 220
rect 18786 200 18886 205
rect 18906 205 18916 220
rect 19001 220 19041 230
rect 19001 205 19011 220
rect 18906 200 19011 205
rect 19031 205 19041 220
rect 19121 220 19161 230
rect 19121 205 19131 220
rect 19031 200 19131 205
rect 19151 205 19161 220
rect 19241 220 19281 230
rect 19241 205 19251 220
rect 19151 200 19251 205
rect 19271 205 19281 220
rect 19361 220 19401 230
rect 19361 205 19371 220
rect 19271 200 19371 205
rect 19391 205 19401 220
rect 19486 220 19526 230
rect 19486 205 19496 220
rect 19391 200 19496 205
rect 19516 205 19526 220
rect 19606 220 19646 230
rect 19606 205 19616 220
rect 19516 200 19616 205
rect 19636 205 19646 220
rect 19726 220 19766 230
rect 19726 205 19736 220
rect 19636 200 19736 205
rect 19756 205 19766 220
rect 19846 220 19886 230
rect 19846 205 19856 220
rect 19756 200 19856 205
rect 19876 205 19886 220
rect 19971 220 20011 230
rect 19971 205 19981 220
rect 19876 200 19981 205
rect 20001 205 20011 220
rect 20091 220 20131 230
rect 20091 205 20101 220
rect 20001 200 20101 205
rect 20121 205 20131 220
rect 20211 220 20251 230
rect 20211 205 20221 220
rect 20121 200 20221 205
rect 20241 205 20251 220
rect 20331 220 20371 230
rect 20331 205 20341 220
rect 20241 200 20341 205
rect 20361 205 20371 220
rect 20456 220 20496 230
rect 20456 205 20466 220
rect 20361 200 20466 205
rect 20486 205 20496 220
rect 20576 220 20616 230
rect 20576 205 20586 220
rect 20486 200 20586 205
rect 20606 205 20616 220
rect 20696 220 20736 230
rect 20696 205 20706 220
rect 20606 200 20706 205
rect 20726 205 20736 220
rect 20816 220 20856 230
rect 20816 205 20826 220
rect 20726 200 20826 205
rect 20846 205 20856 220
rect 20941 220 20981 230
rect 20941 205 20951 220
rect 20846 200 20951 205
rect 20971 205 20981 220
rect 21061 220 21101 230
rect 21061 205 21071 220
rect 20971 200 21071 205
rect 21091 200 21101 220
rect 5660 190 21101 200
rect 316 75 356 85
rect 316 55 326 75
rect 346 70 356 75
rect 431 75 471 85
rect 431 70 441 75
rect 346 55 441 70
rect 461 70 471 75
rect 551 75 591 85
rect 551 70 561 75
rect 461 55 561 70
rect 581 55 591 75
rect 316 45 356 55
rect 431 45 471 55
rect 551 45 591 55
rect 621 75 661 85
rect 621 55 631 75
rect 651 70 661 75
rect 736 75 776 85
rect 736 70 746 75
rect 651 55 746 70
rect 766 70 776 75
rect 856 75 906 85
rect 856 70 876 75
rect 766 55 876 70
rect 896 70 906 75
rect 981 75 1021 85
rect 981 70 991 75
rect 896 55 991 70
rect 1011 70 1021 75
rect 1101 75 1146 85
rect 1101 70 1116 75
rect 1011 55 1116 70
rect 1136 70 1146 75
rect 1221 75 1261 85
rect 1221 70 1231 75
rect 1136 55 1231 70
rect 1251 70 1261 75
rect 1341 75 1391 85
rect 1341 70 1361 75
rect 1251 55 1361 70
rect 1381 70 1391 75
rect 1466 75 1506 85
rect 1466 70 1476 75
rect 1381 55 1476 70
rect 1496 70 1506 75
rect 1586 75 1626 85
rect 1586 70 1596 75
rect 1496 55 1596 70
rect 1616 55 1626 75
rect 621 45 661 55
rect 736 45 776 55
rect 856 45 906 55
rect 981 45 1021 55
rect 1101 45 1146 55
rect 1221 45 1261 55
rect 1341 45 1391 55
rect 1466 45 1506 55
rect 1586 45 1626 55
rect 1656 75 1696 85
rect 1656 55 1666 75
rect 1686 70 1696 75
rect 1771 75 1811 85
rect 1771 70 1781 75
rect 1686 55 1781 70
rect 1801 70 1811 75
rect 1891 75 1941 85
rect 1891 70 1911 75
rect 1801 55 1911 70
rect 1931 70 1941 75
rect 2016 75 2056 85
rect 2016 70 2026 75
rect 1931 55 2026 70
rect 2046 70 2056 75
rect 2136 75 2181 85
rect 2136 70 2151 75
rect 2046 55 2151 70
rect 2171 70 2181 75
rect 2256 75 2296 85
rect 2256 70 2266 75
rect 2171 55 2266 70
rect 2286 70 2296 75
rect 2376 75 2426 85
rect 2376 70 2396 75
rect 2286 55 2396 70
rect 2416 70 2426 75
rect 2501 75 2541 85
rect 2501 70 2511 75
rect 2416 55 2511 70
rect 2531 70 2541 75
rect 2621 75 2666 85
rect 2621 70 2636 75
rect 2531 55 2636 70
rect 2656 70 2666 75
rect 2741 75 2781 85
rect 2741 70 2751 75
rect 2656 55 2751 70
rect 2771 70 2781 75
rect 2861 75 2911 85
rect 2861 70 2881 75
rect 2771 55 2881 70
rect 2901 70 2911 75
rect 2986 75 3026 85
rect 2986 70 2996 75
rect 2901 55 2996 70
rect 3016 70 3026 75
rect 3106 75 3151 85
rect 3106 70 3121 75
rect 3016 55 3121 70
rect 3141 70 3151 75
rect 3226 75 3266 85
rect 3226 70 3236 75
rect 3141 55 3236 70
rect 3256 70 3266 75
rect 3346 75 3396 85
rect 3346 70 3366 75
rect 3256 55 3366 70
rect 3386 70 3396 75
rect 3471 75 3511 85
rect 3471 70 3481 75
rect 3386 55 3481 70
rect 3501 70 3511 75
rect 3591 75 3636 85
rect 3591 70 3606 75
rect 3501 55 3606 70
rect 3626 70 3636 75
rect 3711 75 3751 85
rect 3711 70 3721 75
rect 3626 55 3721 70
rect 3741 70 3751 75
rect 3831 75 3881 85
rect 3831 70 3851 75
rect 3741 55 3851 70
rect 3871 70 3881 75
rect 3956 75 3996 85
rect 3956 70 3966 75
rect 3871 55 3966 70
rect 3986 70 3996 75
rect 4076 75 4121 85
rect 4076 70 4091 75
rect 3986 55 4091 70
rect 4111 70 4121 75
rect 4196 75 4236 85
rect 4196 70 4206 75
rect 4111 55 4206 70
rect 4226 70 4236 75
rect 4316 75 4366 85
rect 4316 70 4336 75
rect 4226 55 4336 70
rect 4356 70 4366 75
rect 4441 75 4481 85
rect 4441 70 4451 75
rect 4356 55 4451 70
rect 4471 70 4481 75
rect 4561 75 4606 85
rect 4561 70 4576 75
rect 4471 55 4576 70
rect 4596 70 4606 75
rect 4681 75 4721 85
rect 4681 70 4691 75
rect 4596 55 4691 70
rect 4711 70 4721 75
rect 4801 75 4851 85
rect 4801 70 4821 75
rect 4711 55 4821 70
rect 4841 70 4851 75
rect 4926 75 4966 85
rect 4926 70 4936 75
rect 4841 55 4936 70
rect 4956 70 4966 75
rect 5046 75 5091 85
rect 5046 70 5061 75
rect 4956 55 5061 70
rect 5081 70 5091 75
rect 5166 75 5206 85
rect 5166 70 5176 75
rect 5081 55 5176 70
rect 5196 70 5206 75
rect 5286 75 5336 85
rect 5286 70 5306 75
rect 5196 55 5306 70
rect 5326 70 5336 75
rect 5411 75 5451 85
rect 5411 70 5421 75
rect 5326 55 5421 70
rect 5441 70 5451 75
rect 5531 75 5571 85
rect 5531 70 5541 75
rect 5441 55 5541 70
rect 5561 55 5571 75
rect 1656 45 1696 55
rect 1771 45 1811 55
rect 1891 45 1941 55
rect 2016 45 2056 55
rect 2136 45 2181 55
rect 2256 45 2296 55
rect 2376 45 2426 55
rect 2501 45 2541 55
rect 2621 45 2666 55
rect 2741 45 2781 55
rect 2861 45 2911 55
rect 2986 45 3026 55
rect 3106 45 3151 55
rect 3226 45 3266 55
rect 3346 45 3396 55
rect 3471 45 3511 55
rect 3591 45 3636 55
rect 3711 45 3751 55
rect 3831 45 3881 55
rect 3956 45 3996 55
rect 4076 45 4121 55
rect 4196 45 4236 55
rect 4316 45 4366 55
rect 4441 45 4481 55
rect 4561 45 4606 55
rect 4681 45 4721 55
rect 4801 45 4851 55
rect 4926 45 4966 55
rect 5046 45 5091 55
rect 5166 45 5206 55
rect 5286 45 5336 55
rect 5411 45 5451 55
rect 5531 45 5571 55
rect 5601 75 5641 85
rect 5601 55 5611 75
rect 5631 70 5641 75
rect 5716 75 5756 85
rect 5716 70 5726 75
rect 5631 55 5726 70
rect 5746 70 5756 75
rect 5836 75 5886 85
rect 5836 70 5856 75
rect 5746 55 5856 70
rect 5876 70 5886 75
rect 5961 75 6001 85
rect 5961 70 5971 75
rect 5876 55 5971 70
rect 5991 70 6001 75
rect 6081 75 6126 85
rect 6081 70 6096 75
rect 5991 55 6096 70
rect 6116 70 6126 75
rect 6201 75 6241 85
rect 6201 70 6211 75
rect 6116 55 6211 70
rect 6231 70 6241 75
rect 6321 75 6371 85
rect 6321 70 6341 75
rect 6231 55 6341 70
rect 6361 70 6371 75
rect 6446 75 6486 85
rect 6446 70 6456 75
rect 6361 55 6456 70
rect 6476 70 6486 75
rect 6566 75 6611 85
rect 6566 70 6581 75
rect 6476 55 6581 70
rect 6601 70 6611 75
rect 6686 75 6726 85
rect 6686 70 6696 75
rect 6601 55 6696 70
rect 6716 70 6726 75
rect 6806 75 6856 85
rect 6806 70 6826 75
rect 6716 55 6826 70
rect 6846 70 6856 75
rect 6931 75 6971 85
rect 6931 70 6941 75
rect 6846 55 6941 70
rect 6961 70 6971 75
rect 7051 75 7096 85
rect 7051 70 7066 75
rect 6961 55 7066 70
rect 7086 70 7096 75
rect 7171 75 7211 85
rect 7171 70 7181 75
rect 7086 55 7181 70
rect 7201 70 7211 75
rect 7291 75 7336 85
rect 7291 70 7306 75
rect 7201 55 7306 70
rect 7326 70 7336 75
rect 7411 75 7451 85
rect 7411 70 7421 75
rect 7326 55 7421 70
rect 7441 70 7451 75
rect 7531 75 7576 85
rect 7531 70 7546 75
rect 7441 55 7546 70
rect 7566 70 7576 75
rect 7651 75 7691 85
rect 7651 70 7661 75
rect 7566 55 7661 70
rect 7681 70 7691 75
rect 7771 75 7821 85
rect 7771 70 7791 75
rect 7681 55 7791 70
rect 7811 70 7821 75
rect 7896 75 7936 85
rect 7896 70 7906 75
rect 7811 55 7906 70
rect 7926 70 7936 75
rect 8016 75 8061 85
rect 8016 70 8031 75
rect 7926 55 8031 70
rect 8051 70 8061 75
rect 8136 75 8176 85
rect 8136 70 8146 75
rect 8051 55 8146 70
rect 8166 70 8176 75
rect 8256 75 8306 85
rect 8256 70 8276 75
rect 8166 55 8276 70
rect 8296 70 8306 75
rect 8381 75 8421 85
rect 8381 70 8391 75
rect 8296 55 8391 70
rect 8411 70 8421 75
rect 8501 75 8546 85
rect 8501 70 8516 75
rect 8411 55 8516 70
rect 8536 70 8546 75
rect 8621 75 8661 85
rect 8621 70 8631 75
rect 8536 55 8631 70
rect 8651 70 8661 75
rect 8741 75 8791 85
rect 8741 70 8761 75
rect 8651 55 8761 70
rect 8781 70 8791 75
rect 8866 75 8906 85
rect 8866 70 8876 75
rect 8781 55 8876 70
rect 8896 70 8906 75
rect 8986 75 9031 85
rect 8986 70 9001 75
rect 8896 55 9001 70
rect 9021 70 9031 75
rect 9106 75 9146 85
rect 9106 70 9116 75
rect 9021 55 9116 70
rect 9136 70 9146 75
rect 9226 75 9276 85
rect 9226 70 9246 75
rect 9136 55 9246 70
rect 9266 70 9276 75
rect 9351 75 9391 85
rect 9351 70 9361 75
rect 9266 55 9361 70
rect 9381 70 9391 75
rect 9471 75 9521 85
rect 9471 70 9491 75
rect 9381 55 9491 70
rect 9511 70 9521 75
rect 9596 75 9636 85
rect 9596 70 9606 75
rect 9511 55 9606 70
rect 9626 70 9636 75
rect 9716 75 9766 85
rect 9716 70 9736 75
rect 9626 55 9736 70
rect 9756 70 9766 75
rect 9841 75 9881 85
rect 9841 70 9851 75
rect 9756 55 9851 70
rect 9871 70 9881 75
rect 9961 75 10006 85
rect 9961 70 9976 75
rect 9871 55 9976 70
rect 9996 70 10006 75
rect 10081 75 10121 85
rect 10081 70 10091 75
rect 9996 55 10091 70
rect 10111 70 10121 75
rect 10201 75 10251 85
rect 10201 70 10221 75
rect 10111 55 10221 70
rect 10241 70 10251 75
rect 10326 75 10366 85
rect 10326 70 10336 75
rect 10241 55 10336 70
rect 10356 70 10366 75
rect 10446 75 10491 85
rect 10446 70 10461 75
rect 10356 55 10461 70
rect 10481 70 10491 75
rect 10566 75 10606 85
rect 10566 70 10576 75
rect 10481 55 10576 70
rect 10596 70 10606 75
rect 10686 75 10736 85
rect 10686 70 10706 75
rect 10596 55 10706 70
rect 10726 70 10736 75
rect 10811 75 10851 85
rect 10811 70 10821 75
rect 10726 55 10821 70
rect 10841 70 10851 75
rect 10931 75 10976 85
rect 10931 70 10946 75
rect 10841 55 10946 70
rect 10966 70 10976 75
rect 11051 75 11091 85
rect 11051 70 11061 75
rect 10966 55 11061 70
rect 11081 70 11091 75
rect 11171 75 11221 85
rect 11171 70 11191 75
rect 11081 55 11191 70
rect 11211 70 11221 75
rect 11296 75 11336 85
rect 11296 70 11306 75
rect 11211 55 11306 70
rect 11326 70 11336 75
rect 11416 75 11461 85
rect 11416 70 11431 75
rect 11326 55 11431 70
rect 11451 70 11461 75
rect 11536 75 11576 85
rect 11536 70 11546 75
rect 11451 55 11546 70
rect 11566 70 11576 75
rect 11656 75 11706 85
rect 11656 70 11676 75
rect 11566 55 11676 70
rect 11696 70 11706 75
rect 11781 75 11821 85
rect 11781 70 11791 75
rect 11696 55 11791 70
rect 11811 70 11821 75
rect 11901 75 11946 85
rect 11901 70 11916 75
rect 11811 55 11916 70
rect 11936 70 11946 75
rect 12021 75 12061 85
rect 12021 70 12031 75
rect 11936 55 12031 70
rect 12051 70 12061 75
rect 12141 75 12191 85
rect 12141 70 12161 75
rect 12051 55 12161 70
rect 12181 70 12191 75
rect 12266 75 12306 85
rect 12266 70 12276 75
rect 12181 55 12276 70
rect 12296 70 12306 75
rect 12386 75 12431 85
rect 12386 70 12401 75
rect 12296 55 12401 70
rect 12421 70 12431 75
rect 12506 75 12546 85
rect 12506 70 12516 75
rect 12421 55 12516 70
rect 12536 70 12546 75
rect 12626 75 12676 85
rect 12626 70 12646 75
rect 12536 55 12646 70
rect 12666 70 12676 75
rect 12751 75 12791 85
rect 12751 70 12761 75
rect 12666 55 12761 70
rect 12781 70 12791 75
rect 12871 75 12916 85
rect 12871 70 12886 75
rect 12781 55 12886 70
rect 12906 70 12916 75
rect 12991 75 13031 85
rect 12991 70 13001 75
rect 12906 55 13001 70
rect 13021 70 13031 75
rect 13111 75 13161 85
rect 13111 70 13131 75
rect 13021 55 13131 70
rect 13151 70 13161 75
rect 13236 75 13276 85
rect 13236 70 13246 75
rect 13151 55 13246 70
rect 13266 70 13276 75
rect 13356 75 13401 85
rect 13356 70 13371 75
rect 13266 55 13371 70
rect 13391 70 13401 75
rect 13476 75 13516 85
rect 13476 70 13486 75
rect 13391 55 13486 70
rect 13506 70 13516 75
rect 13596 75 13646 85
rect 13596 70 13616 75
rect 13506 55 13616 70
rect 13636 70 13646 75
rect 13721 75 13761 85
rect 13721 70 13731 75
rect 13636 55 13731 70
rect 13751 70 13761 75
rect 13841 75 13886 85
rect 13841 70 13856 75
rect 13751 55 13856 70
rect 13876 70 13886 75
rect 13961 75 14001 85
rect 13961 70 13971 75
rect 13876 55 13971 70
rect 13991 70 14001 75
rect 14081 75 14131 85
rect 14081 70 14101 75
rect 13991 55 14101 70
rect 14121 70 14131 75
rect 14206 75 14246 85
rect 14206 70 14216 75
rect 14121 55 14216 70
rect 14236 70 14246 75
rect 14326 75 14371 85
rect 14326 70 14341 75
rect 14236 55 14341 70
rect 14361 70 14371 75
rect 14446 75 14486 85
rect 14446 70 14456 75
rect 14361 55 14456 70
rect 14476 70 14486 75
rect 14566 75 14616 85
rect 14566 70 14586 75
rect 14476 55 14586 70
rect 14606 70 14616 75
rect 14691 75 14731 85
rect 14691 70 14701 75
rect 14606 55 14701 70
rect 14721 70 14731 75
rect 14811 75 14856 85
rect 14811 70 14826 75
rect 14721 55 14826 70
rect 14846 70 14856 75
rect 14931 75 14971 85
rect 14931 70 14941 75
rect 14846 55 14941 70
rect 14961 70 14971 75
rect 15051 75 15101 85
rect 15051 70 15071 75
rect 14961 55 15071 70
rect 15091 70 15101 75
rect 15176 75 15216 85
rect 15176 70 15186 75
rect 15091 55 15186 70
rect 15206 70 15216 75
rect 15296 75 15341 85
rect 15296 70 15311 75
rect 15206 55 15311 70
rect 15331 70 15341 75
rect 15416 75 15456 85
rect 15416 70 15426 75
rect 15331 55 15426 70
rect 15446 70 15456 75
rect 15536 75 15586 85
rect 15536 70 15556 75
rect 15446 55 15556 70
rect 15576 70 15586 75
rect 15661 75 15701 85
rect 15661 70 15671 75
rect 15576 55 15671 70
rect 15691 70 15701 75
rect 15781 75 15826 85
rect 15781 70 15796 75
rect 15691 55 15796 70
rect 15816 70 15826 75
rect 15901 75 15941 85
rect 15901 70 15911 75
rect 15816 55 15911 70
rect 15931 70 15941 75
rect 16021 75 16071 85
rect 16021 70 16041 75
rect 15931 55 16041 70
rect 16061 70 16071 75
rect 16146 75 16186 85
rect 16146 70 16156 75
rect 16061 55 16156 70
rect 16176 70 16186 75
rect 16266 75 16311 85
rect 16266 70 16281 75
rect 16176 55 16281 70
rect 16301 70 16311 75
rect 16386 75 16426 85
rect 16386 70 16396 75
rect 16301 55 16396 70
rect 16416 70 16426 75
rect 16506 75 16556 85
rect 16506 70 16526 75
rect 16416 55 16526 70
rect 16546 70 16556 75
rect 16631 75 16671 85
rect 16631 70 16641 75
rect 16546 55 16641 70
rect 16661 70 16671 75
rect 16751 75 16796 85
rect 16751 70 16766 75
rect 16661 55 16766 70
rect 16786 70 16796 75
rect 16871 75 16911 85
rect 16871 70 16881 75
rect 16786 55 16881 70
rect 16901 70 16911 75
rect 16991 75 17041 85
rect 16991 70 17011 75
rect 16901 55 17011 70
rect 17031 70 17041 75
rect 17116 75 17156 85
rect 17116 70 17126 75
rect 17031 55 17126 70
rect 17146 70 17156 75
rect 17236 75 17281 85
rect 17236 70 17251 75
rect 17146 55 17251 70
rect 17271 70 17281 75
rect 17356 75 17396 85
rect 17356 70 17366 75
rect 17271 55 17366 70
rect 17386 70 17396 75
rect 17476 75 17526 85
rect 17476 70 17496 75
rect 17386 55 17496 70
rect 17516 70 17526 75
rect 17601 75 17641 85
rect 17601 70 17611 75
rect 17516 55 17611 70
rect 17631 70 17641 75
rect 17721 75 17766 85
rect 17721 70 17736 75
rect 17631 55 17736 70
rect 17756 70 17766 75
rect 17841 75 17881 85
rect 17841 70 17851 75
rect 17756 55 17851 70
rect 17871 70 17881 75
rect 17961 75 18011 85
rect 17961 70 17981 75
rect 17871 55 17981 70
rect 18001 70 18011 75
rect 18086 75 18126 85
rect 18086 70 18096 75
rect 18001 55 18096 70
rect 18116 70 18126 75
rect 18206 75 18251 85
rect 18206 70 18221 75
rect 18116 55 18221 70
rect 18241 70 18251 75
rect 18326 75 18366 85
rect 18326 70 18336 75
rect 18241 55 18336 70
rect 18356 70 18366 75
rect 18446 75 18496 85
rect 18446 70 18466 75
rect 18356 55 18466 70
rect 18486 70 18496 75
rect 18571 75 18611 85
rect 18571 70 18581 75
rect 18486 55 18581 70
rect 18601 70 18611 75
rect 18691 75 18736 85
rect 18691 70 18706 75
rect 18601 55 18706 70
rect 18726 70 18736 75
rect 18811 75 18851 85
rect 18811 70 18821 75
rect 18726 55 18821 70
rect 18841 70 18851 75
rect 18931 75 18981 85
rect 18931 70 18951 75
rect 18841 55 18951 70
rect 18971 70 18981 75
rect 19056 75 19096 85
rect 19056 70 19066 75
rect 18971 55 19066 70
rect 19086 70 19096 75
rect 19176 75 19221 85
rect 19176 70 19191 75
rect 19086 55 19191 70
rect 19211 70 19221 75
rect 19296 75 19336 85
rect 19296 70 19306 75
rect 19211 55 19306 70
rect 19326 70 19336 75
rect 19416 75 19466 85
rect 19416 70 19436 75
rect 19326 55 19436 70
rect 19456 70 19466 75
rect 19541 75 19581 85
rect 19541 70 19551 75
rect 19456 55 19551 70
rect 19571 70 19581 75
rect 19661 75 19706 85
rect 19661 70 19676 75
rect 19571 55 19676 70
rect 19696 70 19706 75
rect 19781 75 19821 85
rect 19781 70 19791 75
rect 19696 55 19791 70
rect 19811 70 19821 75
rect 19901 75 19951 85
rect 19901 70 19921 75
rect 19811 55 19921 70
rect 19941 70 19951 75
rect 20026 75 20066 85
rect 20026 70 20036 75
rect 19941 55 20036 70
rect 20056 70 20066 75
rect 20146 75 20191 85
rect 20146 70 20161 75
rect 20056 55 20161 70
rect 20181 70 20191 75
rect 20266 75 20306 85
rect 20266 70 20276 75
rect 20181 55 20276 70
rect 20296 70 20306 75
rect 20386 75 20436 85
rect 20386 70 20406 75
rect 20296 55 20406 70
rect 20426 70 20436 75
rect 20511 75 20551 85
rect 20511 70 20521 75
rect 20426 55 20521 70
rect 20541 70 20551 75
rect 20631 75 20676 85
rect 20631 70 20646 75
rect 20541 55 20646 70
rect 20666 70 20676 75
rect 20751 75 20791 85
rect 20751 70 20761 75
rect 20666 55 20761 70
rect 20781 70 20791 75
rect 20871 75 20921 85
rect 20871 70 20891 75
rect 20781 55 20891 70
rect 20911 70 20921 75
rect 20996 75 21036 85
rect 20996 70 21006 75
rect 20911 55 21006 70
rect 21026 70 21036 75
rect 21116 75 21156 85
rect 21116 70 21126 75
rect 21026 55 21126 70
rect 21146 55 21156 75
rect 5601 45 5641 55
rect 5716 45 5756 55
rect 5836 45 5886 55
rect 5961 45 6001 55
rect 6081 45 6126 55
rect 6201 45 6241 55
rect 6321 45 6371 55
rect 6446 45 6486 55
rect 6566 45 6611 55
rect 6686 45 6726 55
rect 6806 45 6856 55
rect 6931 45 6971 55
rect 7051 45 7096 55
rect 7171 45 7211 55
rect 7291 45 7336 55
rect 7411 45 7451 55
rect 7531 45 7576 55
rect 7651 45 7691 55
rect 7771 45 7821 55
rect 7896 45 7936 55
rect 8016 45 8061 55
rect 8136 45 8176 55
rect 8256 45 8306 55
rect 8381 45 8421 55
rect 8501 45 8546 55
rect 8621 45 8661 55
rect 8741 45 8791 55
rect 8866 45 8906 55
rect 8986 45 9031 55
rect 9106 45 9146 55
rect 9226 45 9276 55
rect 9351 45 9391 55
rect 9471 45 9521 55
rect 9596 45 9636 55
rect 9716 45 9766 55
rect 9841 45 9881 55
rect 9961 45 10006 55
rect 10081 45 10121 55
rect 10201 45 10251 55
rect 10326 45 10366 55
rect 10446 45 10491 55
rect 10566 45 10606 55
rect 10686 45 10736 55
rect 10811 45 10851 55
rect 10931 45 10976 55
rect 11051 45 11091 55
rect 11171 45 11221 55
rect 11296 45 11336 55
rect 11416 45 11461 55
rect 11536 45 11576 55
rect 11656 45 11706 55
rect 11781 45 11821 55
rect 11901 45 11946 55
rect 12021 45 12061 55
rect 12141 45 12191 55
rect 12266 45 12306 55
rect 12386 45 12431 55
rect 12506 45 12546 55
rect 12626 45 12676 55
rect 12751 45 12791 55
rect 12871 45 12916 55
rect 12991 45 13031 55
rect 13111 45 13161 55
rect 13236 45 13276 55
rect 13356 45 13401 55
rect 13476 45 13516 55
rect 13596 45 13646 55
rect 13721 45 13761 55
rect 13841 45 13886 55
rect 13961 45 14001 55
rect 14081 45 14131 55
rect 14206 45 14246 55
rect 14326 45 14371 55
rect 14446 45 14486 55
rect 14566 45 14616 55
rect 14691 45 14731 55
rect 14811 45 14856 55
rect 14931 45 14971 55
rect 15051 45 15101 55
rect 15176 45 15216 55
rect 15296 45 15341 55
rect 15416 45 15456 55
rect 15536 45 15586 55
rect 15661 45 15701 55
rect 15781 45 15826 55
rect 15901 45 15941 55
rect 16021 45 16071 55
rect 16146 45 16186 55
rect 16266 45 16311 55
rect 16386 45 16426 55
rect 16506 45 16556 55
rect 16631 45 16671 55
rect 16751 45 16796 55
rect 16871 45 16911 55
rect 16991 45 17041 55
rect 17116 45 17156 55
rect 17236 45 17281 55
rect 17356 45 17396 55
rect 17476 45 17526 55
rect 17601 45 17641 55
rect 17721 45 17766 55
rect 17841 45 17881 55
rect 17961 45 18011 55
rect 18086 45 18126 55
rect 18206 45 18251 55
rect 18326 45 18366 55
rect 18446 45 18496 55
rect 18571 45 18611 55
rect 18691 45 18736 55
rect 18811 45 18851 55
rect 18931 45 18981 55
rect 19056 45 19096 55
rect 19176 45 19221 55
rect 19296 45 19336 55
rect 19416 45 19466 55
rect 19541 45 19581 55
rect 19661 45 19706 55
rect 19781 45 19821 55
rect 19901 45 19951 55
rect 20026 45 20066 55
rect 20146 45 20191 55
rect 20266 45 20306 55
rect 20386 45 20436 55
rect 20511 45 20551 55
rect 20631 45 20676 55
rect 20751 45 20791 55
rect 20871 45 20921 55
rect 20996 45 21036 55
rect 21116 45 21156 55
rect 21150 15 21190 20
rect 21150 -15 21155 15
rect 21185 -15 21190 15
rect 21150 -20 21190 -15
rect 316 -45 356 -35
rect 316 -65 326 -45
rect 346 -50 356 -45
rect 436 -50 476 -40
rect 551 -50 591 -40
rect 346 -65 446 -50
rect 316 -75 356 -65
rect 436 -70 446 -65
rect 466 -65 561 -50
rect 466 -70 476 -65
rect 436 -80 476 -70
rect 551 -70 561 -65
rect 581 -70 591 -50
rect 551 -80 591 -70
rect 621 -45 661 -35
rect 866 -40 906 -35
rect 1106 -40 1146 -35
rect 1351 -40 1391 -35
rect 621 -65 631 -45
rect 651 -50 661 -45
rect 741 -50 781 -40
rect 856 -45 906 -40
rect 856 -50 876 -45
rect 651 -65 751 -50
rect 621 -75 661 -65
rect 741 -70 751 -65
rect 771 -65 876 -50
rect 896 -50 906 -45
rect 986 -50 1026 -40
rect 1101 -45 1146 -40
rect 1101 -50 1116 -45
rect 896 -65 996 -50
rect 771 -70 781 -65
rect 741 -80 781 -70
rect 856 -75 906 -65
rect 986 -70 996 -65
rect 1016 -65 1116 -50
rect 1136 -50 1146 -45
rect 1226 -50 1266 -40
rect 1341 -45 1391 -40
rect 1341 -50 1361 -45
rect 1136 -65 1236 -50
rect 1016 -70 1026 -65
rect 856 -80 896 -75
rect 986 -80 1026 -70
rect 1101 -75 1146 -65
rect 1226 -70 1236 -65
rect 1256 -65 1361 -50
rect 1381 -50 1391 -45
rect 1471 -50 1511 -40
rect 1586 -50 1626 -40
rect 1381 -65 1481 -50
rect 1256 -70 1266 -65
rect 1101 -80 1141 -75
rect 1226 -80 1266 -70
rect 1341 -75 1391 -65
rect 1471 -70 1481 -65
rect 1501 -65 1596 -50
rect 1501 -70 1511 -65
rect 1341 -80 1381 -75
rect 1471 -80 1511 -70
rect 1586 -70 1596 -65
rect 1616 -70 1626 -50
rect 1586 -80 1626 -70
rect 1656 -45 1696 -35
rect 1901 -40 1941 -35
rect 2141 -40 2181 -35
rect 2386 -40 2426 -35
rect 2626 -40 2666 -35
rect 2871 -40 2911 -35
rect 3111 -40 3151 -35
rect 3356 -40 3396 -35
rect 3596 -40 3636 -35
rect 3841 -40 3881 -35
rect 4081 -40 4121 -35
rect 4326 -40 4366 -35
rect 4566 -40 4606 -35
rect 4811 -40 4851 -35
rect 5051 -40 5091 -35
rect 5296 -40 5336 -35
rect 1656 -65 1666 -45
rect 1686 -50 1696 -45
rect 1776 -50 1816 -40
rect 1891 -45 1941 -40
rect 1891 -50 1911 -45
rect 1686 -65 1786 -50
rect 1656 -75 1696 -65
rect 1776 -70 1786 -65
rect 1806 -65 1911 -50
rect 1931 -50 1941 -45
rect 2021 -50 2061 -40
rect 2136 -45 2181 -40
rect 2136 -50 2151 -45
rect 1931 -65 2031 -50
rect 1806 -70 1816 -65
rect 1776 -80 1816 -70
rect 1891 -75 1941 -65
rect 2021 -70 2031 -65
rect 2051 -65 2151 -50
rect 2171 -50 2181 -45
rect 2261 -50 2301 -40
rect 2376 -45 2426 -40
rect 2376 -50 2396 -45
rect 2171 -65 2271 -50
rect 2051 -70 2061 -65
rect 1891 -80 1931 -75
rect 2021 -80 2061 -70
rect 2136 -75 2181 -65
rect 2261 -70 2271 -65
rect 2291 -65 2396 -50
rect 2416 -50 2426 -45
rect 2506 -50 2546 -40
rect 2621 -45 2666 -40
rect 2621 -50 2636 -45
rect 2416 -65 2516 -50
rect 2291 -70 2301 -65
rect 2136 -80 2176 -75
rect 2261 -80 2301 -70
rect 2376 -75 2426 -65
rect 2506 -70 2516 -65
rect 2536 -65 2636 -50
rect 2656 -50 2666 -45
rect 2746 -50 2786 -40
rect 2861 -45 2911 -40
rect 2861 -50 2881 -45
rect 2656 -65 2756 -50
rect 2536 -70 2546 -65
rect 2376 -80 2416 -75
rect 2506 -80 2546 -70
rect 2621 -75 2666 -65
rect 2746 -70 2756 -65
rect 2776 -65 2881 -50
rect 2901 -50 2911 -45
rect 2991 -50 3031 -40
rect 3106 -45 3151 -40
rect 3106 -50 3121 -45
rect 2901 -65 3001 -50
rect 2776 -70 2786 -65
rect 2621 -80 2661 -75
rect 2746 -80 2786 -70
rect 2861 -75 2911 -65
rect 2991 -70 3001 -65
rect 3021 -65 3121 -50
rect 3141 -50 3151 -45
rect 3231 -50 3271 -40
rect 3346 -45 3396 -40
rect 3346 -50 3366 -45
rect 3141 -65 3241 -50
rect 3021 -70 3031 -65
rect 2861 -80 2901 -75
rect 2991 -80 3031 -70
rect 3106 -75 3151 -65
rect 3231 -70 3241 -65
rect 3261 -65 3366 -50
rect 3386 -50 3396 -45
rect 3476 -50 3516 -40
rect 3591 -45 3636 -40
rect 3591 -50 3606 -45
rect 3386 -65 3486 -50
rect 3261 -70 3271 -65
rect 3106 -80 3146 -75
rect 3231 -80 3271 -70
rect 3346 -75 3396 -65
rect 3476 -70 3486 -65
rect 3506 -65 3606 -50
rect 3626 -50 3636 -45
rect 3716 -50 3756 -40
rect 3831 -45 3881 -40
rect 3831 -50 3851 -45
rect 3626 -65 3726 -50
rect 3506 -70 3516 -65
rect 3346 -80 3386 -75
rect 3476 -80 3516 -70
rect 3591 -75 3636 -65
rect 3716 -70 3726 -65
rect 3746 -65 3851 -50
rect 3871 -50 3881 -45
rect 3961 -50 4001 -40
rect 4076 -45 4121 -40
rect 4076 -50 4091 -45
rect 3871 -65 3971 -50
rect 3746 -70 3756 -65
rect 3591 -80 3626 -75
rect 3716 -80 3756 -70
rect 3831 -75 3881 -65
rect 3961 -70 3971 -65
rect 3991 -65 4091 -50
rect 4111 -50 4121 -45
rect 4201 -50 4241 -40
rect 4316 -45 4366 -40
rect 4316 -50 4336 -45
rect 4111 -65 4211 -50
rect 3991 -70 4001 -65
rect 3831 -80 3871 -75
rect 3961 -80 4001 -70
rect 4076 -75 4121 -65
rect 4201 -70 4211 -65
rect 4231 -65 4336 -50
rect 4356 -50 4366 -45
rect 4446 -50 4486 -40
rect 4561 -45 4606 -40
rect 4561 -50 4576 -45
rect 4356 -65 4456 -50
rect 4231 -70 4241 -65
rect 4076 -80 4116 -75
rect 4201 -80 4241 -70
rect 4316 -75 4366 -65
rect 4446 -70 4456 -65
rect 4476 -65 4576 -50
rect 4596 -50 4606 -45
rect 4686 -50 4726 -40
rect 4801 -45 4851 -40
rect 4801 -50 4821 -45
rect 4596 -65 4696 -50
rect 4476 -70 4486 -65
rect 4316 -80 4356 -75
rect 4446 -80 4486 -70
rect 4561 -75 4606 -65
rect 4686 -70 4696 -65
rect 4716 -65 4821 -50
rect 4841 -50 4851 -45
rect 4931 -50 4971 -40
rect 5046 -45 5091 -40
rect 5046 -50 5061 -45
rect 4841 -65 4941 -50
rect 4716 -70 4726 -65
rect 4561 -80 4601 -75
rect 4686 -80 4726 -70
rect 4801 -75 4851 -65
rect 4931 -70 4941 -65
rect 4961 -65 5061 -50
rect 5081 -50 5091 -45
rect 5171 -50 5211 -40
rect 5286 -45 5336 -40
rect 5286 -50 5306 -45
rect 5081 -65 5181 -50
rect 4961 -70 4971 -65
rect 4801 -80 4841 -75
rect 4931 -80 4971 -70
rect 5046 -75 5091 -65
rect 5171 -70 5181 -65
rect 5201 -65 5306 -50
rect 5326 -50 5336 -45
rect 5416 -50 5456 -40
rect 5531 -50 5571 -40
rect 5326 -65 5426 -50
rect 5201 -70 5211 -65
rect 5046 -80 5086 -75
rect 5171 -80 5211 -70
rect 5286 -75 5336 -65
rect 5416 -70 5426 -65
rect 5446 -65 5541 -50
rect 5446 -70 5456 -65
rect 5286 -80 5326 -75
rect 5416 -80 5456 -70
rect 5531 -70 5541 -65
rect 5561 -70 5571 -50
rect 5531 -80 5571 -70
rect 5601 -45 5641 -35
rect 5846 -40 5886 -35
rect 6086 -40 6126 -35
rect 6331 -40 6371 -35
rect 6571 -40 6611 -35
rect 6816 -40 6856 -35
rect 7056 -40 7096 -35
rect 7301 -40 7336 -35
rect 7536 -40 7576 -35
rect 7781 -40 7821 -35
rect 8021 -40 8061 -35
rect 8266 -40 8306 -35
rect 8506 -40 8546 -35
rect 8751 -40 8791 -35
rect 8991 -40 9031 -35
rect 9236 -40 9276 -35
rect 9481 -40 9521 -35
rect 9726 -40 9766 -35
rect 9966 -40 10006 -35
rect 10211 -40 10251 -35
rect 10451 -40 10491 -35
rect 10696 -40 10736 -35
rect 10936 -40 10976 -35
rect 11181 -40 11221 -35
rect 11421 -40 11461 -35
rect 11666 -40 11706 -35
rect 11906 -40 11946 -35
rect 12151 -40 12191 -35
rect 12391 -40 12431 -35
rect 12636 -40 12676 -35
rect 12876 -40 12916 -35
rect 13121 -40 13161 -35
rect 13361 -40 13401 -35
rect 13606 -40 13646 -35
rect 13846 -40 13886 -35
rect 14091 -40 14131 -35
rect 14331 -40 14371 -35
rect 14576 -40 14616 -35
rect 14816 -40 14856 -35
rect 15061 -40 15101 -35
rect 15301 -40 15341 -35
rect 15546 -40 15586 -35
rect 15786 -40 15826 -35
rect 16031 -40 16071 -35
rect 16271 -40 16311 -35
rect 16516 -40 16556 -35
rect 16756 -40 16796 -35
rect 17001 -40 17041 -35
rect 17241 -40 17281 -35
rect 17486 -40 17526 -35
rect 17726 -40 17766 -35
rect 17971 -40 18011 -35
rect 18211 -40 18251 -35
rect 18456 -40 18496 -35
rect 18696 -40 18736 -35
rect 18941 -40 18981 -35
rect 19181 -40 19221 -35
rect 19426 -40 19466 -35
rect 19666 -40 19706 -35
rect 19911 -40 19951 -35
rect 20151 -40 20191 -35
rect 20396 -40 20436 -35
rect 20636 -40 20676 -35
rect 20881 -40 20921 -35
rect 5601 -65 5611 -45
rect 5631 -50 5641 -45
rect 5721 -50 5761 -40
rect 5836 -45 5886 -40
rect 5836 -50 5856 -45
rect 5631 -65 5731 -50
rect 5601 -75 5641 -65
rect 5721 -70 5731 -65
rect 5751 -65 5856 -50
rect 5876 -50 5886 -45
rect 5966 -50 6006 -40
rect 6081 -45 6126 -40
rect 6081 -50 6096 -45
rect 5876 -65 5976 -50
rect 5751 -70 5761 -65
rect 5721 -80 5761 -70
rect 5836 -75 5886 -65
rect 5966 -70 5976 -65
rect 5996 -65 6096 -50
rect 6116 -50 6126 -45
rect 6206 -50 6246 -40
rect 6321 -45 6371 -40
rect 6321 -50 6341 -45
rect 6116 -65 6216 -50
rect 5996 -70 6006 -65
rect 5836 -80 5876 -75
rect 5966 -80 6006 -70
rect 6081 -75 6126 -65
rect 6206 -70 6216 -65
rect 6236 -65 6341 -50
rect 6361 -50 6371 -45
rect 6451 -50 6491 -40
rect 6566 -45 6611 -40
rect 6566 -50 6581 -45
rect 6361 -65 6461 -50
rect 6236 -70 6246 -65
rect 6081 -80 6121 -75
rect 6206 -80 6246 -70
rect 6321 -75 6371 -65
rect 6451 -70 6461 -65
rect 6481 -65 6581 -50
rect 6601 -50 6611 -45
rect 6691 -50 6731 -40
rect 6806 -45 6856 -40
rect 6806 -50 6826 -45
rect 6601 -65 6701 -50
rect 6481 -70 6491 -65
rect 6321 -80 6361 -75
rect 6451 -80 6491 -70
rect 6566 -75 6611 -65
rect 6691 -70 6701 -65
rect 6721 -65 6826 -50
rect 6846 -50 6856 -45
rect 6936 -50 6976 -40
rect 7051 -45 7096 -40
rect 7051 -50 7066 -45
rect 6846 -65 6946 -50
rect 6721 -70 6731 -65
rect 6566 -80 6606 -75
rect 6691 -80 6731 -70
rect 6806 -75 6856 -65
rect 6936 -70 6946 -65
rect 6966 -65 7066 -50
rect 7086 -50 7096 -45
rect 7176 -50 7216 -40
rect 7291 -45 7336 -40
rect 7291 -50 7306 -45
rect 7086 -65 7186 -50
rect 6966 -70 6976 -65
rect 6806 -80 6846 -75
rect 6936 -80 6976 -70
rect 7051 -75 7096 -65
rect 7176 -70 7186 -65
rect 7206 -65 7306 -50
rect 7326 -50 7336 -45
rect 7416 -50 7456 -40
rect 7531 -45 7576 -40
rect 7531 -50 7546 -45
rect 7326 -65 7426 -50
rect 7206 -70 7216 -65
rect 7051 -80 7091 -75
rect 7176 -80 7216 -70
rect 7291 -75 7336 -65
rect 7416 -70 7426 -65
rect 7446 -65 7546 -50
rect 7566 -50 7576 -45
rect 7656 -50 7696 -40
rect 7771 -45 7821 -40
rect 7771 -50 7791 -45
rect 7566 -65 7666 -50
rect 7446 -70 7456 -65
rect 7291 -80 7326 -75
rect 7416 -80 7456 -70
rect 7531 -75 7576 -65
rect 7656 -70 7666 -65
rect 7686 -65 7791 -50
rect 7811 -50 7821 -45
rect 7901 -50 7941 -40
rect 8016 -45 8061 -40
rect 8016 -50 8031 -45
rect 7811 -65 7911 -50
rect 7686 -70 7696 -65
rect 7531 -80 7566 -75
rect 7656 -80 7696 -70
rect 7771 -75 7821 -65
rect 7901 -70 7911 -65
rect 7931 -65 8031 -50
rect 8051 -50 8061 -45
rect 8141 -50 8181 -40
rect 8256 -45 8306 -40
rect 8256 -50 8276 -45
rect 8051 -65 8151 -50
rect 7931 -70 7941 -65
rect 7771 -80 7811 -75
rect 7901 -80 7941 -70
rect 8016 -75 8061 -65
rect 8141 -70 8151 -65
rect 8171 -65 8276 -50
rect 8296 -50 8306 -45
rect 8386 -50 8426 -40
rect 8501 -45 8546 -40
rect 8501 -50 8516 -45
rect 8296 -65 8396 -50
rect 8171 -70 8181 -65
rect 8016 -80 8056 -75
rect 8141 -80 8181 -70
rect 8256 -75 8306 -65
rect 8386 -70 8396 -65
rect 8416 -65 8516 -50
rect 8536 -50 8546 -45
rect 8626 -50 8666 -40
rect 8741 -45 8791 -40
rect 8741 -50 8761 -45
rect 8536 -65 8636 -50
rect 8416 -70 8426 -65
rect 8256 -80 8296 -75
rect 8386 -80 8426 -70
rect 8501 -75 8546 -65
rect 8626 -70 8636 -65
rect 8656 -65 8761 -50
rect 8781 -50 8791 -45
rect 8871 -50 8911 -40
rect 8986 -45 9031 -40
rect 8986 -50 9001 -45
rect 8781 -65 8881 -50
rect 8656 -70 8666 -65
rect 8501 -80 8541 -75
rect 8626 -80 8666 -70
rect 8741 -75 8791 -65
rect 8871 -70 8881 -65
rect 8901 -65 9001 -50
rect 9021 -50 9031 -45
rect 9111 -50 9151 -40
rect 9226 -45 9276 -40
rect 9226 -50 9246 -45
rect 9021 -65 9121 -50
rect 8901 -70 8911 -65
rect 8741 -80 8781 -75
rect 8871 -80 8911 -70
rect 8986 -75 9031 -65
rect 9111 -70 9121 -65
rect 9141 -65 9246 -50
rect 9266 -50 9276 -45
rect 9356 -50 9396 -40
rect 9471 -45 9521 -40
rect 9471 -50 9491 -45
rect 9266 -65 9366 -50
rect 9141 -70 9151 -65
rect 8986 -80 9026 -75
rect 9111 -80 9151 -70
rect 9226 -75 9276 -65
rect 9356 -70 9366 -65
rect 9386 -65 9491 -50
rect 9511 -50 9521 -45
rect 9601 -50 9641 -40
rect 9716 -45 9766 -40
rect 9716 -50 9736 -45
rect 9511 -65 9611 -50
rect 9386 -70 9396 -65
rect 9226 -80 9266 -75
rect 9356 -80 9396 -70
rect 9471 -75 9521 -65
rect 9601 -70 9611 -65
rect 9631 -65 9736 -50
rect 9756 -50 9766 -45
rect 9846 -50 9886 -40
rect 9961 -45 10006 -40
rect 9961 -50 9976 -45
rect 9756 -65 9856 -50
rect 9631 -70 9641 -65
rect 9471 -80 9511 -75
rect 9601 -80 9641 -70
rect 9716 -75 9766 -65
rect 9846 -70 9856 -65
rect 9876 -65 9976 -50
rect 9996 -50 10006 -45
rect 10086 -50 10126 -40
rect 10201 -45 10251 -40
rect 10201 -50 10221 -45
rect 9996 -65 10096 -50
rect 9876 -70 9886 -65
rect 9716 -80 9756 -75
rect 9846 -80 9886 -70
rect 9961 -75 10006 -65
rect 10086 -70 10096 -65
rect 10116 -65 10221 -50
rect 10241 -50 10251 -45
rect 10331 -50 10371 -40
rect 10446 -45 10491 -40
rect 10446 -50 10461 -45
rect 10241 -65 10341 -50
rect 10116 -70 10126 -65
rect 9961 -80 10001 -75
rect 10086 -80 10126 -70
rect 10201 -75 10251 -65
rect 10331 -70 10341 -65
rect 10361 -65 10461 -50
rect 10481 -50 10491 -45
rect 10571 -50 10611 -40
rect 10686 -45 10736 -40
rect 10686 -50 10706 -45
rect 10481 -65 10581 -50
rect 10361 -70 10371 -65
rect 10201 -80 10241 -75
rect 10331 -80 10371 -70
rect 10446 -75 10491 -65
rect 10571 -70 10581 -65
rect 10601 -65 10706 -50
rect 10726 -50 10736 -45
rect 10816 -50 10856 -40
rect 10931 -45 10976 -40
rect 10931 -50 10946 -45
rect 10726 -65 10826 -50
rect 10601 -70 10611 -65
rect 10446 -80 10486 -75
rect 10571 -80 10611 -70
rect 10686 -75 10736 -65
rect 10816 -70 10826 -65
rect 10846 -65 10946 -50
rect 10966 -50 10976 -45
rect 11056 -50 11096 -40
rect 11171 -45 11221 -40
rect 11171 -50 11191 -45
rect 10966 -65 11066 -50
rect 10846 -70 10856 -65
rect 10686 -80 10726 -75
rect 10816 -80 10856 -70
rect 10931 -75 10976 -65
rect 11056 -70 11066 -65
rect 11086 -65 11191 -50
rect 11211 -50 11221 -45
rect 11301 -50 11341 -40
rect 11416 -45 11461 -40
rect 11416 -50 11431 -45
rect 11211 -65 11311 -50
rect 11086 -70 11096 -65
rect 10931 -80 10971 -75
rect 11056 -80 11096 -70
rect 11171 -75 11221 -65
rect 11301 -70 11311 -65
rect 11331 -65 11431 -50
rect 11451 -50 11461 -45
rect 11541 -50 11581 -40
rect 11656 -45 11706 -40
rect 11656 -50 11676 -45
rect 11451 -65 11551 -50
rect 11331 -70 11341 -65
rect 11171 -80 11211 -75
rect 11301 -80 11341 -70
rect 11416 -75 11461 -65
rect 11541 -70 11551 -65
rect 11571 -65 11676 -50
rect 11696 -50 11706 -45
rect 11786 -50 11826 -40
rect 11901 -45 11946 -40
rect 11901 -50 11916 -45
rect 11696 -65 11796 -50
rect 11571 -70 11581 -65
rect 11416 -80 11451 -75
rect 11541 -80 11581 -70
rect 11656 -75 11706 -65
rect 11786 -70 11796 -65
rect 11816 -65 11916 -50
rect 11936 -50 11946 -45
rect 12026 -50 12066 -40
rect 12141 -45 12191 -40
rect 12141 -50 12161 -45
rect 11936 -65 12036 -50
rect 11816 -70 11826 -65
rect 11656 -80 11696 -75
rect 11786 -80 11826 -70
rect 11901 -75 11946 -65
rect 12026 -70 12036 -65
rect 12056 -65 12161 -50
rect 12181 -50 12191 -45
rect 12271 -50 12311 -40
rect 12386 -45 12431 -40
rect 12386 -50 12401 -45
rect 12181 -65 12281 -50
rect 12056 -70 12066 -65
rect 11901 -80 11941 -75
rect 12026 -80 12066 -70
rect 12141 -75 12191 -65
rect 12271 -70 12281 -65
rect 12301 -65 12401 -50
rect 12421 -50 12431 -45
rect 12511 -50 12551 -40
rect 12626 -45 12676 -40
rect 12626 -50 12646 -45
rect 12421 -65 12521 -50
rect 12301 -70 12311 -65
rect 12141 -80 12181 -75
rect 12271 -80 12311 -70
rect 12386 -75 12431 -65
rect 12511 -70 12521 -65
rect 12541 -65 12646 -50
rect 12666 -50 12676 -45
rect 12756 -50 12796 -40
rect 12871 -45 12916 -40
rect 12871 -50 12886 -45
rect 12666 -65 12766 -50
rect 12541 -70 12551 -65
rect 12386 -80 12426 -75
rect 12511 -80 12551 -70
rect 12626 -75 12676 -65
rect 12756 -70 12766 -65
rect 12786 -65 12886 -50
rect 12906 -50 12916 -45
rect 12996 -50 13036 -40
rect 13111 -45 13161 -40
rect 13111 -50 13131 -45
rect 12906 -65 13006 -50
rect 12786 -70 12796 -65
rect 12626 -80 12666 -75
rect 12756 -80 12796 -70
rect 12871 -75 12916 -65
rect 12996 -70 13006 -65
rect 13026 -65 13131 -50
rect 13151 -50 13161 -45
rect 13241 -50 13281 -40
rect 13356 -45 13401 -40
rect 13356 -50 13371 -45
rect 13151 -65 13251 -50
rect 13026 -70 13036 -65
rect 12871 -80 12911 -75
rect 12996 -80 13036 -70
rect 13111 -75 13161 -65
rect 13241 -70 13251 -65
rect 13271 -65 13371 -50
rect 13391 -50 13401 -45
rect 13481 -50 13521 -40
rect 13596 -45 13646 -40
rect 13596 -50 13616 -45
rect 13391 -65 13491 -50
rect 13271 -70 13281 -65
rect 13111 -80 13151 -75
rect 13241 -80 13281 -70
rect 13356 -75 13401 -65
rect 13481 -70 13491 -65
rect 13511 -65 13616 -50
rect 13636 -50 13646 -45
rect 13726 -50 13766 -40
rect 13841 -45 13886 -40
rect 13841 -50 13856 -45
rect 13636 -65 13736 -50
rect 13511 -70 13521 -65
rect 13356 -80 13396 -75
rect 13481 -80 13521 -70
rect 13596 -75 13646 -65
rect 13726 -70 13736 -65
rect 13756 -65 13856 -50
rect 13876 -50 13886 -45
rect 13966 -50 14006 -40
rect 14081 -45 14131 -40
rect 14081 -50 14101 -45
rect 13876 -65 13976 -50
rect 13756 -70 13766 -65
rect 13596 -80 13636 -75
rect 13726 -80 13766 -70
rect 13841 -75 13886 -65
rect 13966 -70 13976 -65
rect 13996 -65 14101 -50
rect 14121 -50 14131 -45
rect 14211 -50 14251 -40
rect 14326 -45 14371 -40
rect 14326 -50 14341 -45
rect 14121 -65 14221 -50
rect 13996 -70 14006 -65
rect 13841 -80 13881 -75
rect 13966 -80 14006 -70
rect 14081 -75 14131 -65
rect 14211 -70 14221 -65
rect 14241 -65 14341 -50
rect 14361 -50 14371 -45
rect 14451 -50 14491 -40
rect 14566 -45 14616 -40
rect 14566 -50 14586 -45
rect 14361 -65 14461 -50
rect 14241 -70 14251 -65
rect 14081 -80 14121 -75
rect 14211 -80 14251 -70
rect 14326 -75 14371 -65
rect 14451 -70 14461 -65
rect 14481 -65 14586 -50
rect 14606 -50 14616 -45
rect 14696 -50 14736 -40
rect 14811 -45 14856 -40
rect 14811 -50 14826 -45
rect 14606 -65 14706 -50
rect 14481 -70 14491 -65
rect 14326 -80 14366 -75
rect 14451 -80 14491 -70
rect 14566 -75 14616 -65
rect 14696 -70 14706 -65
rect 14726 -65 14826 -50
rect 14846 -50 14856 -45
rect 14936 -50 14976 -40
rect 15051 -45 15101 -40
rect 15051 -50 15071 -45
rect 14846 -65 14946 -50
rect 14726 -70 14736 -65
rect 14566 -80 14606 -75
rect 14696 -80 14736 -70
rect 14811 -75 14856 -65
rect 14936 -70 14946 -65
rect 14966 -65 15071 -50
rect 15091 -50 15101 -45
rect 15181 -50 15221 -40
rect 15296 -45 15341 -40
rect 15296 -50 15311 -45
rect 15091 -65 15191 -50
rect 14966 -70 14976 -65
rect 14811 -80 14851 -75
rect 14936 -80 14976 -70
rect 15051 -75 15101 -65
rect 15181 -70 15191 -65
rect 15211 -65 15311 -50
rect 15331 -50 15341 -45
rect 15421 -50 15461 -40
rect 15536 -45 15586 -40
rect 15536 -50 15556 -45
rect 15331 -65 15431 -50
rect 15211 -70 15221 -65
rect 15051 -80 15091 -75
rect 15181 -80 15221 -70
rect 15296 -75 15341 -65
rect 15421 -70 15431 -65
rect 15451 -65 15556 -50
rect 15576 -50 15586 -45
rect 15666 -50 15706 -40
rect 15781 -45 15826 -40
rect 15781 -50 15796 -45
rect 15576 -65 15676 -50
rect 15451 -70 15461 -65
rect 15296 -80 15331 -75
rect 15421 -80 15461 -70
rect 15536 -75 15586 -65
rect 15666 -70 15676 -65
rect 15696 -65 15796 -50
rect 15816 -50 15826 -45
rect 15906 -50 15946 -40
rect 16021 -45 16071 -40
rect 16021 -50 16041 -45
rect 15816 -65 15916 -50
rect 15696 -70 15706 -65
rect 15536 -80 15576 -75
rect 15666 -80 15706 -70
rect 15781 -75 15826 -65
rect 15906 -70 15916 -65
rect 15936 -65 16041 -50
rect 16061 -50 16071 -45
rect 16151 -50 16191 -40
rect 16266 -45 16311 -40
rect 16266 -50 16281 -45
rect 16061 -65 16161 -50
rect 15936 -70 15946 -65
rect 15781 -80 15821 -75
rect 15906 -80 15946 -70
rect 16021 -75 16071 -65
rect 16151 -70 16161 -65
rect 16181 -65 16281 -50
rect 16301 -50 16311 -45
rect 16391 -50 16431 -40
rect 16506 -45 16556 -40
rect 16506 -50 16526 -45
rect 16301 -65 16401 -50
rect 16181 -70 16191 -65
rect 16021 -80 16061 -75
rect 16151 -80 16191 -70
rect 16266 -75 16311 -65
rect 16391 -70 16401 -65
rect 16421 -65 16526 -50
rect 16546 -50 16556 -45
rect 16636 -50 16676 -40
rect 16751 -45 16796 -40
rect 16751 -50 16766 -45
rect 16546 -65 16646 -50
rect 16421 -70 16431 -65
rect 16266 -80 16306 -75
rect 16391 -80 16431 -70
rect 16506 -75 16556 -65
rect 16636 -70 16646 -65
rect 16666 -65 16766 -50
rect 16786 -50 16796 -45
rect 16876 -50 16916 -40
rect 16991 -45 17041 -40
rect 16991 -50 17011 -45
rect 16786 -65 16886 -50
rect 16666 -70 16676 -65
rect 16506 -80 16546 -75
rect 16636 -80 16676 -70
rect 16751 -75 16796 -65
rect 16876 -70 16886 -65
rect 16906 -65 17011 -50
rect 17031 -50 17041 -45
rect 17121 -50 17161 -40
rect 17236 -45 17281 -40
rect 17236 -50 17251 -45
rect 17031 -65 17131 -50
rect 16906 -70 16916 -65
rect 16751 -80 16791 -75
rect 16876 -80 16916 -70
rect 16991 -75 17041 -65
rect 17121 -70 17131 -65
rect 17151 -65 17251 -50
rect 17271 -50 17281 -45
rect 17361 -50 17401 -40
rect 17476 -45 17526 -40
rect 17476 -50 17496 -45
rect 17271 -65 17371 -50
rect 17151 -70 17161 -65
rect 16991 -80 17031 -75
rect 17121 -80 17161 -70
rect 17236 -75 17281 -65
rect 17361 -70 17371 -65
rect 17391 -65 17496 -50
rect 17516 -50 17526 -45
rect 17606 -50 17646 -40
rect 17721 -45 17766 -40
rect 17721 -50 17736 -45
rect 17516 -65 17616 -50
rect 17391 -70 17401 -65
rect 17236 -80 17276 -75
rect 17361 -80 17401 -70
rect 17476 -75 17526 -65
rect 17606 -70 17616 -65
rect 17636 -65 17736 -50
rect 17756 -50 17766 -45
rect 17846 -50 17886 -40
rect 17961 -45 18011 -40
rect 17961 -50 17981 -45
rect 17756 -65 17856 -50
rect 17636 -70 17646 -65
rect 17476 -80 17516 -75
rect 17606 -80 17646 -70
rect 17721 -75 17766 -65
rect 17846 -70 17856 -65
rect 17876 -65 17981 -50
rect 18001 -50 18011 -45
rect 18091 -50 18131 -40
rect 18206 -45 18251 -40
rect 18206 -50 18221 -45
rect 18001 -65 18101 -50
rect 17876 -70 17886 -65
rect 17721 -80 17761 -75
rect 17846 -80 17886 -70
rect 17961 -75 18011 -65
rect 18091 -70 18101 -65
rect 18121 -65 18221 -50
rect 18241 -50 18251 -45
rect 18331 -50 18371 -40
rect 18446 -45 18496 -40
rect 18446 -50 18466 -45
rect 18241 -65 18341 -50
rect 18121 -70 18131 -65
rect 17961 -80 18001 -75
rect 18091 -80 18131 -70
rect 18206 -75 18251 -65
rect 18331 -70 18341 -65
rect 18361 -65 18466 -50
rect 18486 -50 18496 -45
rect 18576 -50 18616 -40
rect 18691 -45 18736 -40
rect 18691 -50 18706 -45
rect 18486 -65 18586 -50
rect 18361 -70 18371 -65
rect 18206 -80 18246 -75
rect 18331 -80 18371 -70
rect 18446 -75 18496 -65
rect 18576 -70 18586 -65
rect 18606 -65 18706 -50
rect 18726 -50 18736 -45
rect 18816 -50 18856 -40
rect 18931 -45 18981 -40
rect 18931 -50 18951 -45
rect 18726 -65 18826 -50
rect 18606 -70 18616 -65
rect 18446 -80 18486 -75
rect 18576 -80 18616 -70
rect 18691 -75 18736 -65
rect 18816 -70 18826 -65
rect 18846 -65 18951 -50
rect 18971 -50 18981 -45
rect 19061 -50 19101 -40
rect 19176 -45 19221 -40
rect 19176 -50 19191 -45
rect 18971 -65 19071 -50
rect 18846 -70 18856 -65
rect 18691 -80 18731 -75
rect 18816 -80 18856 -70
rect 18931 -75 18981 -65
rect 19061 -70 19071 -65
rect 19091 -65 19191 -50
rect 19211 -50 19221 -45
rect 19301 -50 19341 -40
rect 19416 -45 19466 -40
rect 19416 -50 19436 -45
rect 19211 -65 19311 -50
rect 19091 -70 19101 -65
rect 18931 -80 18971 -75
rect 19061 -80 19101 -70
rect 19176 -75 19221 -65
rect 19301 -70 19311 -65
rect 19331 -65 19436 -50
rect 19456 -50 19466 -45
rect 19546 -50 19586 -40
rect 19661 -45 19706 -40
rect 19661 -50 19676 -45
rect 19456 -65 19556 -50
rect 19331 -70 19341 -65
rect 19176 -80 19211 -75
rect 19301 -80 19341 -70
rect 19416 -75 19466 -65
rect 19546 -70 19556 -65
rect 19576 -65 19676 -50
rect 19696 -50 19706 -45
rect 19786 -50 19826 -40
rect 19901 -45 19951 -40
rect 19901 -50 19921 -45
rect 19696 -65 19796 -50
rect 19576 -70 19586 -65
rect 19416 -80 19456 -75
rect 19546 -80 19586 -70
rect 19661 -75 19706 -65
rect 19786 -70 19796 -65
rect 19816 -65 19921 -50
rect 19941 -50 19951 -45
rect 20031 -50 20071 -40
rect 20146 -45 20191 -40
rect 20146 -50 20161 -45
rect 19941 -65 20041 -50
rect 19816 -70 19826 -65
rect 19661 -80 19701 -75
rect 19786 -80 19826 -70
rect 19901 -75 19951 -65
rect 20031 -70 20041 -65
rect 20061 -65 20161 -50
rect 20181 -50 20191 -45
rect 20271 -50 20311 -40
rect 20386 -45 20436 -40
rect 20386 -50 20406 -45
rect 20181 -65 20281 -50
rect 20061 -70 20071 -65
rect 19901 -80 19941 -75
rect 20031 -80 20071 -70
rect 20146 -75 20191 -65
rect 20271 -70 20281 -65
rect 20301 -65 20406 -50
rect 20426 -50 20436 -45
rect 20516 -50 20556 -40
rect 20631 -45 20676 -40
rect 20631 -50 20646 -45
rect 20426 -65 20526 -50
rect 20301 -70 20311 -65
rect 20146 -80 20186 -75
rect 20271 -80 20311 -70
rect 20386 -75 20436 -65
rect 20516 -70 20526 -65
rect 20546 -65 20646 -50
rect 20666 -50 20676 -45
rect 20756 -50 20796 -40
rect 20871 -45 20921 -40
rect 20871 -50 20891 -45
rect 20666 -65 20766 -50
rect 20546 -70 20556 -65
rect 20386 -80 20426 -75
rect 20516 -80 20556 -70
rect 20631 -75 20676 -65
rect 20756 -70 20766 -65
rect 20786 -65 20891 -50
rect 20911 -50 20921 -45
rect 21001 -50 21041 -40
rect 21116 -50 21156 -40
rect 20911 -65 21011 -50
rect 20786 -70 20796 -65
rect 20631 -80 20671 -75
rect 20756 -80 20796 -70
rect 20871 -75 20921 -65
rect 21001 -70 21011 -65
rect 21031 -65 21126 -50
rect 21031 -70 21041 -65
rect 20871 -80 20911 -75
rect 21001 -80 21041 -70
rect 21116 -70 21126 -65
rect 21146 -70 21156 -50
rect 21116 -80 21156 -70
rect 376 -120 416 -115
rect 496 -120 536 -115
rect 376 -125 536 -120
rect 376 -145 386 -125
rect 406 -135 506 -125
rect 406 -145 416 -135
rect 376 -150 416 -145
rect 496 -145 506 -135
rect 526 -145 536 -125
rect 680 -125 1571 -115
rect 1716 -120 1756 -115
rect 1836 -120 1876 -115
rect 1961 -120 2001 -115
rect 2081 -120 2121 -115
rect 2201 -120 2241 -115
rect 2321 -120 2361 -115
rect 2446 -120 2486 -115
rect 2566 -120 2606 -115
rect 2686 -120 2726 -115
rect 2806 -120 2846 -115
rect 2931 -120 2971 -115
rect 3051 -120 3091 -115
rect 3171 -120 3211 -115
rect 3291 -120 3331 -115
rect 3416 -120 3456 -115
rect 3536 -120 3576 -115
rect 3656 -120 3696 -115
rect 3776 -120 3816 -115
rect 3901 -120 3941 -115
rect 4021 -120 4061 -115
rect 4141 -120 4181 -115
rect 4261 -120 4301 -115
rect 4386 -120 4426 -115
rect 4506 -120 4546 -115
rect 4626 -120 4666 -115
rect 4746 -120 4786 -115
rect 4871 -120 4911 -115
rect 4991 -120 5031 -115
rect 5111 -120 5151 -115
rect 5231 -120 5271 -115
rect 5356 -120 5396 -115
rect 5476 -120 5516 -115
rect 5661 -120 5701 -115
rect 5781 -120 5821 -115
rect 5906 -120 5946 -115
rect 6026 -120 6066 -115
rect 6146 -120 6186 -115
rect 6266 -120 6306 -115
rect 6391 -120 6431 -115
rect 6511 -120 6551 -115
rect 6631 -120 6671 -115
rect 6751 -120 6791 -115
rect 6876 -120 6916 -115
rect 6996 -120 7036 -115
rect 7116 -120 7156 -115
rect 7236 -120 7276 -115
rect 7356 -120 7396 -115
rect 7476 -120 7516 -115
rect 7596 -120 7636 -115
rect 7716 -120 7756 -115
rect 7841 -120 7881 -115
rect 7961 -120 8001 -115
rect 8081 -120 8121 -115
rect 8201 -120 8241 -115
rect 8326 -120 8366 -115
rect 8446 -120 8486 -115
rect 8566 -120 8606 -115
rect 8686 -120 8726 -115
rect 8811 -120 8851 -115
rect 8931 -120 8971 -115
rect 9051 -120 9091 -115
rect 9171 -120 9211 -115
rect 9296 -120 9336 -115
rect 9416 -120 9456 -115
rect 9541 -120 9581 -115
rect 9661 -120 9701 -115
rect 9786 -120 9826 -115
rect 9906 -120 9946 -115
rect 10026 -120 10066 -115
rect 10146 -120 10186 -115
rect 10271 -120 10311 -115
rect 10391 -120 10431 -115
rect 10511 -120 10551 -115
rect 10631 -120 10671 -115
rect 10756 -120 10796 -115
rect 10876 -120 10916 -115
rect 10996 -120 11036 -115
rect 11116 -120 11156 -115
rect 11241 -120 11281 -115
rect 11361 -120 11401 -115
rect 11481 -120 11521 -115
rect 11601 -120 11641 -115
rect 11726 -120 11766 -115
rect 11846 -120 11886 -115
rect 11966 -120 12006 -115
rect 12086 -120 12126 -115
rect 12211 -120 12251 -115
rect 12331 -120 12371 -115
rect 12451 -120 12491 -115
rect 12571 -120 12611 -115
rect 12696 -120 12736 -115
rect 12816 -120 12856 -115
rect 12936 -120 12976 -115
rect 13056 -120 13096 -115
rect 13181 -120 13221 -115
rect 13301 -120 13341 -115
rect 13421 -120 13461 -115
rect 13541 -120 13581 -115
rect 13666 -120 13706 -115
rect 13786 -120 13826 -115
rect 13906 -120 13946 -115
rect 14026 -120 14066 -115
rect 14151 -120 14191 -115
rect 14271 -120 14311 -115
rect 14391 -120 14431 -115
rect 14511 -120 14551 -115
rect 14636 -120 14676 -115
rect 14756 -120 14796 -115
rect 14876 -120 14916 -115
rect 14996 -120 15036 -115
rect 15121 -120 15161 -115
rect 15241 -120 15281 -115
rect 15361 -120 15401 -115
rect 15481 -120 15521 -115
rect 15606 -120 15646 -115
rect 15726 -120 15766 -115
rect 15846 -120 15886 -115
rect 15966 -120 16006 -115
rect 16091 -120 16131 -115
rect 16211 -120 16251 -115
rect 16331 -120 16371 -115
rect 16451 -120 16491 -115
rect 16576 -120 16616 -115
rect 16696 -120 16736 -115
rect 16816 -120 16856 -115
rect 16936 -120 16976 -115
rect 17061 -120 17101 -115
rect 17181 -120 17221 -115
rect 17301 -120 17341 -115
rect 17421 -120 17461 -115
rect 17546 -120 17586 -115
rect 17666 -120 17706 -115
rect 17786 -120 17826 -115
rect 17906 -120 17946 -115
rect 18031 -120 18071 -115
rect 18151 -120 18191 -115
rect 18271 -120 18311 -115
rect 18391 -120 18431 -115
rect 18516 -120 18556 -115
rect 18636 -120 18676 -115
rect 18756 -120 18796 -115
rect 18876 -120 18916 -115
rect 19001 -120 19041 -115
rect 19121 -120 19161 -115
rect 19241 -120 19281 -115
rect 19361 -120 19401 -115
rect 19486 -120 19526 -115
rect 19606 -120 19646 -115
rect 19726 -120 19766 -115
rect 19846 -120 19886 -115
rect 19971 -120 20011 -115
rect 20091 -120 20131 -115
rect 20211 -120 20251 -115
rect 20331 -120 20371 -115
rect 20456 -120 20496 -115
rect 20576 -120 20616 -115
rect 20696 -120 20736 -115
rect 20816 -120 20856 -115
rect 20941 -120 20981 -115
rect 21061 -120 21101 -115
rect 680 -145 691 -125
rect 711 -145 811 -125
rect 831 -145 936 -125
rect 956 -145 1056 -125
rect 1076 -145 1176 -125
rect 1196 -145 1296 -125
rect 1316 -145 1421 -125
rect 1441 -145 1541 -125
rect 1561 -145 1571 -125
rect 1715 -125 5516 -120
rect 1715 -140 1726 -125
rect 496 -150 536 -145
rect 681 -150 721 -145
rect 801 -150 841 -145
rect 926 -150 966 -145
rect 1046 -150 1086 -145
rect 1166 -150 1206 -145
rect 1286 -150 1326 -145
rect 1411 -150 1451 -145
rect 1531 -150 1571 -145
rect 1716 -145 1726 -140
rect 1746 -140 1846 -125
rect 1746 -145 1756 -140
rect 1716 -150 1756 -145
rect 1836 -145 1846 -140
rect 1866 -140 1971 -125
rect 1866 -145 1876 -140
rect 1836 -150 1876 -145
rect 1961 -145 1971 -140
rect 1991 -140 2091 -125
rect 1991 -145 2001 -140
rect 1961 -150 2001 -145
rect 2081 -145 2091 -140
rect 2111 -140 2211 -125
rect 2111 -145 2121 -140
rect 2081 -150 2121 -145
rect 2201 -145 2211 -140
rect 2231 -140 2331 -125
rect 2231 -145 2241 -140
rect 2201 -150 2241 -145
rect 2321 -145 2331 -140
rect 2351 -140 2456 -125
rect 2351 -145 2361 -140
rect 2321 -150 2361 -145
rect 2446 -145 2456 -140
rect 2476 -140 2576 -125
rect 2476 -145 2486 -140
rect 2446 -150 2486 -145
rect 2566 -145 2576 -140
rect 2596 -140 2696 -125
rect 2596 -145 2606 -140
rect 2566 -150 2606 -145
rect 2686 -145 2696 -140
rect 2716 -140 2816 -125
rect 2716 -145 2726 -140
rect 2686 -150 2726 -145
rect 2806 -145 2816 -140
rect 2836 -140 2941 -125
rect 2836 -145 2846 -140
rect 2806 -150 2846 -145
rect 2931 -145 2941 -140
rect 2961 -140 3061 -125
rect 2961 -145 2971 -140
rect 2931 -150 2971 -145
rect 3051 -145 3061 -140
rect 3081 -140 3181 -125
rect 3081 -145 3091 -140
rect 3051 -150 3091 -145
rect 3171 -145 3181 -140
rect 3201 -140 3301 -125
rect 3201 -145 3211 -140
rect 3171 -150 3211 -145
rect 3291 -145 3301 -140
rect 3321 -140 3426 -125
rect 3321 -145 3331 -140
rect 3291 -150 3331 -145
rect 3416 -145 3426 -140
rect 3446 -140 3546 -125
rect 3446 -145 3456 -140
rect 3416 -150 3456 -145
rect 3536 -145 3546 -140
rect 3566 -140 3666 -125
rect 3566 -145 3576 -140
rect 3536 -150 3576 -145
rect 3656 -145 3666 -140
rect 3686 -140 3786 -125
rect 3686 -145 3696 -140
rect 3656 -150 3696 -145
rect 3776 -145 3786 -140
rect 3806 -140 3911 -125
rect 3806 -145 3816 -140
rect 3776 -150 3816 -145
rect 3901 -145 3911 -140
rect 3931 -140 4031 -125
rect 3931 -145 3941 -140
rect 3901 -150 3941 -145
rect 4021 -145 4031 -140
rect 4051 -140 4151 -125
rect 4051 -145 4061 -140
rect 4021 -150 4061 -145
rect 4141 -145 4151 -140
rect 4171 -140 4271 -125
rect 4171 -145 4181 -140
rect 4141 -150 4181 -145
rect 4261 -145 4271 -140
rect 4291 -140 4396 -125
rect 4291 -145 4301 -140
rect 4261 -150 4301 -145
rect 4386 -145 4396 -140
rect 4416 -140 4516 -125
rect 4416 -145 4426 -140
rect 4386 -150 4426 -145
rect 4506 -145 4516 -140
rect 4536 -140 4636 -125
rect 4536 -145 4546 -140
rect 4506 -150 4546 -145
rect 4626 -145 4636 -140
rect 4656 -140 4756 -125
rect 4656 -145 4666 -140
rect 4626 -150 4666 -145
rect 4746 -145 4756 -140
rect 4776 -140 4881 -125
rect 4776 -145 4786 -140
rect 4746 -150 4786 -145
rect 4871 -145 4881 -140
rect 4901 -140 5001 -125
rect 4901 -145 4911 -140
rect 4871 -150 4911 -145
rect 4991 -145 5001 -140
rect 5021 -140 5121 -125
rect 5021 -145 5031 -140
rect 4991 -150 5031 -145
rect 5111 -145 5121 -140
rect 5141 -140 5241 -125
rect 5141 -145 5151 -140
rect 5111 -150 5151 -145
rect 5231 -145 5241 -140
rect 5261 -140 5366 -125
rect 5261 -145 5271 -140
rect 5231 -150 5271 -145
rect 5356 -145 5366 -140
rect 5386 -140 5486 -125
rect 5386 -145 5396 -140
rect 5356 -150 5396 -145
rect 5476 -145 5486 -140
rect 5506 -145 5516 -125
rect 5660 -125 6401 -120
rect 5660 -140 5671 -125
rect 5476 -150 5516 -145
rect 5661 -145 5671 -140
rect 5691 -140 5791 -125
rect 5691 -145 5701 -140
rect 5661 -150 5701 -145
rect 5781 -145 5791 -140
rect 5811 -140 5916 -125
rect 5811 -145 5821 -140
rect 5781 -150 5821 -145
rect 5906 -145 5916 -140
rect 5936 -140 6036 -125
rect 5936 -145 5946 -140
rect 5906 -150 5946 -145
rect 6026 -145 6036 -140
rect 6056 -140 6156 -125
rect 6056 -145 6066 -140
rect 6026 -150 6066 -145
rect 6146 -145 6156 -140
rect 6176 -140 6276 -125
rect 6176 -145 6186 -140
rect 6146 -150 6186 -145
rect 6266 -145 6276 -140
rect 6296 -140 6401 -125
rect 6421 -125 9551 -120
rect 6421 -140 6521 -125
rect 6296 -145 6306 -140
rect 6391 -145 6430 -140
rect 6511 -145 6521 -140
rect 6541 -140 6641 -125
rect 6541 -145 6551 -140
rect 6266 -150 6306 -145
rect 6511 -150 6551 -145
rect 6631 -145 6641 -140
rect 6661 -140 6761 -125
rect 6661 -145 6671 -140
rect 6631 -150 6671 -145
rect 6751 -145 6761 -140
rect 6781 -140 6886 -125
rect 6781 -145 6791 -140
rect 6751 -150 6791 -145
rect 6876 -145 6886 -140
rect 6906 -140 7006 -125
rect 6906 -145 6916 -140
rect 6876 -150 6916 -145
rect 6996 -145 7006 -140
rect 7026 -140 7126 -125
rect 7026 -145 7036 -140
rect 6996 -150 7036 -145
rect 7116 -145 7126 -140
rect 7146 -140 7246 -125
rect 7146 -145 7156 -140
rect 7116 -150 7156 -145
rect 7236 -145 7246 -140
rect 7266 -140 7366 -125
rect 7266 -145 7276 -140
rect 7236 -150 7276 -145
rect 7356 -145 7366 -140
rect 7386 -140 7486 -125
rect 7386 -145 7396 -140
rect 7356 -150 7396 -145
rect 7476 -145 7486 -140
rect 7506 -140 7606 -125
rect 7506 -145 7516 -140
rect 7476 -150 7516 -145
rect 7596 -145 7606 -140
rect 7626 -140 7726 -125
rect 7626 -145 7636 -140
rect 7596 -150 7636 -145
rect 7716 -145 7726 -140
rect 7746 -140 7851 -125
rect 7746 -145 7756 -140
rect 7716 -150 7756 -145
rect 7841 -145 7851 -140
rect 7871 -140 7971 -125
rect 7871 -145 7881 -140
rect 7841 -150 7881 -145
rect 7961 -145 7971 -140
rect 7991 -140 8091 -125
rect 7991 -145 8001 -140
rect 7961 -150 8001 -145
rect 8081 -145 8091 -140
rect 8111 -140 8211 -125
rect 8111 -145 8121 -140
rect 8081 -150 8121 -145
rect 8201 -145 8211 -140
rect 8231 -140 8336 -125
rect 8231 -145 8241 -140
rect 8201 -150 8241 -145
rect 8326 -145 8336 -140
rect 8356 -140 8456 -125
rect 8356 -145 8366 -140
rect 8326 -150 8366 -145
rect 8446 -145 8456 -140
rect 8476 -140 8576 -125
rect 8476 -145 8486 -140
rect 8446 -150 8486 -145
rect 8566 -145 8576 -140
rect 8596 -140 8696 -125
rect 8596 -145 8606 -140
rect 8566 -150 8606 -145
rect 8686 -145 8696 -140
rect 8716 -140 8821 -125
rect 8716 -145 8726 -140
rect 8686 -150 8726 -145
rect 8811 -145 8821 -140
rect 8841 -140 8941 -125
rect 8841 -145 8851 -140
rect 8811 -150 8851 -145
rect 8931 -145 8941 -140
rect 8961 -140 9061 -125
rect 8961 -145 8971 -140
rect 8931 -150 8971 -145
rect 9051 -145 9061 -140
rect 9081 -140 9181 -125
rect 9081 -145 9091 -140
rect 9051 -150 9091 -145
rect 9171 -145 9181 -140
rect 9201 -140 9306 -125
rect 9201 -145 9211 -140
rect 9171 -150 9211 -145
rect 9296 -145 9306 -140
rect 9326 -140 9426 -125
rect 9326 -145 9336 -140
rect 9296 -150 9336 -145
rect 9416 -145 9426 -140
rect 9446 -140 9551 -125
rect 9571 -125 21101 -120
rect 9571 -140 9671 -125
rect 9446 -145 9456 -140
rect 9541 -145 9580 -140
rect 9661 -145 9671 -140
rect 9691 -140 9796 -125
rect 9691 -145 9701 -140
rect 9416 -150 9456 -145
rect 9661 -150 9701 -145
rect 9786 -145 9796 -140
rect 9816 -140 9916 -125
rect 9816 -145 9826 -140
rect 9786 -150 9826 -145
rect 9906 -145 9916 -140
rect 9936 -140 10036 -125
rect 9936 -145 9946 -140
rect 9906 -150 9946 -145
rect 10026 -145 10036 -140
rect 10056 -140 10156 -125
rect 10056 -145 10066 -140
rect 10026 -150 10066 -145
rect 10146 -145 10156 -140
rect 10176 -140 10281 -125
rect 10176 -145 10186 -140
rect 10146 -150 10186 -145
rect 10271 -145 10281 -140
rect 10301 -140 10401 -125
rect 10301 -145 10311 -140
rect 10271 -150 10311 -145
rect 10391 -145 10401 -140
rect 10421 -140 10521 -125
rect 10421 -145 10431 -140
rect 10391 -150 10431 -145
rect 10511 -145 10521 -140
rect 10541 -140 10641 -125
rect 10541 -145 10551 -140
rect 10511 -150 10551 -145
rect 10631 -145 10641 -140
rect 10661 -140 10766 -125
rect 10661 -145 10671 -140
rect 10631 -150 10671 -145
rect 10756 -145 10766 -140
rect 10786 -140 10886 -125
rect 10786 -145 10796 -140
rect 10756 -150 10796 -145
rect 10876 -145 10886 -140
rect 10906 -140 11006 -125
rect 10906 -145 10916 -140
rect 10876 -150 10916 -145
rect 10996 -145 11006 -140
rect 11026 -140 11126 -125
rect 11026 -145 11036 -140
rect 10996 -150 11036 -145
rect 11116 -145 11126 -140
rect 11146 -140 11251 -125
rect 11146 -145 11156 -140
rect 11116 -150 11156 -145
rect 11241 -145 11251 -140
rect 11271 -140 11371 -125
rect 11271 -145 11281 -140
rect 11241 -150 11281 -145
rect 11361 -145 11371 -140
rect 11391 -140 11491 -125
rect 11391 -145 11401 -140
rect 11361 -150 11401 -145
rect 11481 -145 11491 -140
rect 11511 -140 11611 -125
rect 11511 -145 11521 -140
rect 11481 -150 11521 -145
rect 11601 -145 11611 -140
rect 11631 -140 11736 -125
rect 11631 -145 11641 -140
rect 11601 -150 11641 -145
rect 11726 -145 11736 -140
rect 11756 -140 11856 -125
rect 11756 -145 11766 -140
rect 11726 -150 11766 -145
rect 11846 -145 11856 -140
rect 11876 -140 11976 -125
rect 11876 -145 11886 -140
rect 11846 -150 11886 -145
rect 11966 -145 11976 -140
rect 11996 -140 12096 -125
rect 11996 -145 12006 -140
rect 11966 -150 12006 -145
rect 12086 -145 12096 -140
rect 12116 -140 12221 -125
rect 12116 -145 12126 -140
rect 12086 -150 12126 -145
rect 12211 -145 12221 -140
rect 12241 -140 12341 -125
rect 12241 -145 12251 -140
rect 12211 -150 12251 -145
rect 12331 -145 12341 -140
rect 12361 -140 12461 -125
rect 12361 -145 12371 -140
rect 12331 -150 12371 -145
rect 12451 -145 12461 -140
rect 12481 -140 12581 -125
rect 12481 -145 12491 -140
rect 12451 -150 12491 -145
rect 12571 -145 12581 -140
rect 12601 -140 12706 -125
rect 12601 -145 12611 -140
rect 12571 -150 12611 -145
rect 12696 -145 12706 -140
rect 12726 -140 12826 -125
rect 12726 -145 12736 -140
rect 12696 -150 12736 -145
rect 12816 -145 12826 -140
rect 12846 -140 12946 -125
rect 12846 -145 12856 -140
rect 12816 -150 12856 -145
rect 12936 -145 12946 -140
rect 12966 -140 13066 -125
rect 12966 -145 12976 -140
rect 12936 -150 12976 -145
rect 13056 -145 13066 -140
rect 13086 -140 13191 -125
rect 13086 -145 13096 -140
rect 13056 -150 13096 -145
rect 13181 -145 13191 -140
rect 13211 -140 13311 -125
rect 13211 -145 13221 -140
rect 13181 -150 13221 -145
rect 13301 -145 13311 -140
rect 13331 -140 13431 -125
rect 13331 -145 13341 -140
rect 13301 -150 13341 -145
rect 13421 -145 13431 -140
rect 13451 -140 13551 -125
rect 13451 -145 13461 -140
rect 13421 -150 13461 -145
rect 13541 -145 13551 -140
rect 13571 -140 13676 -125
rect 13571 -145 13581 -140
rect 13541 -150 13581 -145
rect 13666 -145 13676 -140
rect 13696 -140 13796 -125
rect 13696 -145 13706 -140
rect 13666 -150 13706 -145
rect 13786 -145 13796 -140
rect 13816 -140 13916 -125
rect 13816 -145 13826 -140
rect 13786 -150 13826 -145
rect 13906 -145 13916 -140
rect 13936 -140 14036 -125
rect 13936 -145 13946 -140
rect 13906 -150 13946 -145
rect 14026 -145 14036 -140
rect 14056 -140 14161 -125
rect 14056 -145 14066 -140
rect 14026 -150 14066 -145
rect 14151 -145 14161 -140
rect 14181 -140 14281 -125
rect 14181 -145 14191 -140
rect 14151 -150 14191 -145
rect 14271 -145 14281 -140
rect 14301 -140 14401 -125
rect 14301 -145 14311 -140
rect 14271 -150 14311 -145
rect 14391 -145 14401 -140
rect 14421 -140 14521 -125
rect 14421 -145 14431 -140
rect 14391 -150 14431 -145
rect 14511 -145 14521 -140
rect 14541 -140 14646 -125
rect 14541 -145 14551 -140
rect 14511 -150 14551 -145
rect 14636 -145 14646 -140
rect 14666 -140 14766 -125
rect 14666 -145 14676 -140
rect 14636 -150 14676 -145
rect 14756 -145 14766 -140
rect 14786 -140 14886 -125
rect 14786 -145 14796 -140
rect 14756 -150 14796 -145
rect 14876 -145 14886 -140
rect 14906 -140 15006 -125
rect 14906 -145 14916 -140
rect 14876 -150 14916 -145
rect 14996 -145 15006 -140
rect 15026 -140 15131 -125
rect 15026 -145 15036 -140
rect 14996 -150 15036 -145
rect 15121 -145 15131 -140
rect 15151 -140 15251 -125
rect 15151 -145 15161 -140
rect 15121 -150 15161 -145
rect 15241 -145 15251 -140
rect 15271 -140 15371 -125
rect 15271 -145 15281 -140
rect 15241 -150 15281 -145
rect 15361 -145 15371 -140
rect 15391 -140 15491 -125
rect 15391 -145 15401 -140
rect 15361 -150 15401 -145
rect 15481 -145 15491 -140
rect 15511 -140 15616 -125
rect 15511 -145 15521 -140
rect 15481 -150 15521 -145
rect 15606 -145 15616 -140
rect 15636 -140 15736 -125
rect 15636 -145 15646 -140
rect 15606 -150 15646 -145
rect 15726 -145 15736 -140
rect 15756 -140 15856 -125
rect 15756 -145 15766 -140
rect 15726 -150 15766 -145
rect 15846 -145 15856 -140
rect 15876 -140 15976 -125
rect 15876 -145 15886 -140
rect 15846 -150 15886 -145
rect 15966 -145 15976 -140
rect 15996 -140 16101 -125
rect 15996 -145 16006 -140
rect 15966 -150 16006 -145
rect 16091 -145 16101 -140
rect 16121 -140 16221 -125
rect 16121 -145 16131 -140
rect 16091 -150 16131 -145
rect 16211 -145 16221 -140
rect 16241 -140 16341 -125
rect 16241 -145 16251 -140
rect 16211 -150 16251 -145
rect 16331 -145 16341 -140
rect 16361 -140 16461 -125
rect 16361 -145 16371 -140
rect 16331 -150 16371 -145
rect 16451 -145 16461 -140
rect 16481 -140 16586 -125
rect 16481 -145 16491 -140
rect 16451 -150 16491 -145
rect 16576 -145 16586 -140
rect 16606 -140 16706 -125
rect 16606 -145 16616 -140
rect 16576 -150 16616 -145
rect 16696 -145 16706 -140
rect 16726 -140 16826 -125
rect 16726 -145 16736 -140
rect 16696 -150 16736 -145
rect 16816 -145 16826 -140
rect 16846 -140 16946 -125
rect 16846 -145 16856 -140
rect 16816 -150 16856 -145
rect 16936 -145 16946 -140
rect 16966 -140 17071 -125
rect 16966 -145 16976 -140
rect 16936 -150 16976 -145
rect 17061 -145 17071 -140
rect 17091 -140 17191 -125
rect 17091 -145 17101 -140
rect 17061 -150 17101 -145
rect 17181 -145 17191 -140
rect 17211 -140 17311 -125
rect 17211 -145 17221 -140
rect 17181 -150 17221 -145
rect 17301 -145 17311 -140
rect 17331 -140 17431 -125
rect 17331 -145 17341 -140
rect 17301 -150 17341 -145
rect 17421 -145 17431 -140
rect 17451 -140 17556 -125
rect 17451 -145 17461 -140
rect 17421 -150 17461 -145
rect 17546 -145 17556 -140
rect 17576 -140 17676 -125
rect 17576 -145 17586 -140
rect 17546 -150 17586 -145
rect 17666 -145 17676 -140
rect 17696 -140 17796 -125
rect 17696 -145 17706 -140
rect 17666 -150 17706 -145
rect 17786 -145 17796 -140
rect 17816 -140 17916 -125
rect 17816 -145 17826 -140
rect 17786 -150 17826 -145
rect 17906 -145 17916 -140
rect 17936 -140 18041 -125
rect 17936 -145 17946 -140
rect 17906 -150 17946 -145
rect 18031 -145 18041 -140
rect 18061 -140 18161 -125
rect 18061 -145 18071 -140
rect 18031 -150 18071 -145
rect 18151 -145 18161 -140
rect 18181 -140 18281 -125
rect 18181 -145 18191 -140
rect 18151 -150 18191 -145
rect 18271 -145 18281 -140
rect 18301 -140 18401 -125
rect 18301 -145 18311 -140
rect 18271 -150 18311 -145
rect 18391 -145 18401 -140
rect 18421 -140 18526 -125
rect 18421 -145 18431 -140
rect 18391 -150 18431 -145
rect 18516 -145 18526 -140
rect 18546 -140 18646 -125
rect 18546 -145 18556 -140
rect 18516 -150 18556 -145
rect 18636 -145 18646 -140
rect 18666 -140 18766 -125
rect 18666 -145 18676 -140
rect 18636 -150 18676 -145
rect 18756 -145 18766 -140
rect 18786 -140 18886 -125
rect 18786 -145 18796 -140
rect 18756 -150 18796 -145
rect 18876 -145 18886 -140
rect 18906 -140 19011 -125
rect 18906 -145 18916 -140
rect 18876 -150 18916 -145
rect 19001 -145 19011 -140
rect 19031 -140 19131 -125
rect 19031 -145 19041 -140
rect 19001 -150 19041 -145
rect 19121 -145 19131 -140
rect 19151 -140 19251 -125
rect 19151 -145 19161 -140
rect 19121 -150 19161 -145
rect 19241 -145 19251 -140
rect 19271 -140 19371 -125
rect 19271 -145 19281 -140
rect 19241 -150 19281 -145
rect 19361 -145 19371 -140
rect 19391 -140 19496 -125
rect 19391 -145 19401 -140
rect 19361 -150 19401 -145
rect 19486 -145 19496 -140
rect 19516 -140 19616 -125
rect 19516 -145 19526 -140
rect 19486 -150 19526 -145
rect 19606 -145 19616 -140
rect 19636 -140 19736 -125
rect 19636 -145 19646 -140
rect 19606 -150 19646 -145
rect 19726 -145 19736 -140
rect 19756 -140 19856 -125
rect 19756 -145 19766 -140
rect 19726 -150 19766 -145
rect 19846 -145 19856 -140
rect 19876 -140 19981 -125
rect 19876 -145 19886 -140
rect 19846 -150 19886 -145
rect 19971 -145 19981 -140
rect 20001 -140 20101 -125
rect 20001 -145 20011 -140
rect 19971 -150 20011 -145
rect 20091 -145 20101 -140
rect 20121 -140 20221 -125
rect 20121 -145 20131 -140
rect 20091 -150 20131 -145
rect 20211 -145 20221 -140
rect 20241 -140 20341 -125
rect 20241 -145 20251 -140
rect 20211 -150 20251 -145
rect 20331 -145 20341 -140
rect 20361 -140 20466 -125
rect 20361 -145 20371 -140
rect 20331 -150 20371 -145
rect 20456 -145 20466 -140
rect 20486 -140 20586 -125
rect 20486 -145 20496 -140
rect 20456 -150 20496 -145
rect 20576 -145 20586 -140
rect 20606 -140 20706 -125
rect 20606 -145 20616 -140
rect 20576 -150 20616 -145
rect 20696 -145 20706 -140
rect 20726 -140 20826 -125
rect 20726 -145 20736 -140
rect 20696 -150 20736 -145
rect 20816 -145 20826 -140
rect 20846 -140 20951 -125
rect 20846 -145 20856 -140
rect 20816 -150 20856 -145
rect 20941 -145 20951 -140
rect 20971 -140 21071 -125
rect 20971 -145 20981 -140
rect 20941 -150 20981 -145
rect 21061 -145 21071 -140
rect 21091 -145 21101 -125
rect 21061 -150 21101 -145
rect 181 -165 221 -160
rect -425 -190 -355 -180
rect -425 -240 -415 -190
rect -365 -240 -355 -190
rect 181 -195 186 -165
rect 216 -195 221 -165
rect 181 -200 221 -195
rect 426 -165 466 -160
rect 426 -195 431 -165
rect 461 -195 466 -165
rect 426 -200 466 -195
rect 731 -165 771 -160
rect 731 -195 736 -165
rect 766 -195 771 -165
rect 731 -200 771 -195
rect 976 -165 1016 -160
rect 976 -195 981 -165
rect 1011 -195 1016 -165
rect 976 -200 1016 -195
rect 1216 -165 1256 -160
rect 1216 -195 1221 -165
rect 1251 -195 1256 -165
rect 1216 -200 1256 -195
rect 1461 -165 1501 -160
rect 1461 -195 1466 -165
rect 1496 -195 1501 -165
rect 1766 -165 1806 -160
rect 1461 -200 1501 -195
rect 1625 -200 1685 -190
rect 1766 -195 1771 -165
rect 1801 -195 1806 -165
rect 1766 -200 1806 -195
rect 2011 -165 2051 -160
rect 2011 -195 2016 -165
rect 2046 -195 2051 -165
rect 2011 -200 2051 -195
rect 2251 -165 2291 -160
rect 2251 -195 2256 -165
rect 2286 -195 2291 -165
rect 2251 -200 2291 -195
rect 2496 -165 2536 -160
rect 2496 -195 2501 -165
rect 2531 -195 2536 -165
rect 2496 -200 2536 -195
rect 2736 -165 2776 -160
rect 2736 -195 2741 -165
rect 2771 -195 2776 -165
rect 2736 -200 2776 -195
rect 2981 -165 3021 -160
rect 2981 -195 2986 -165
rect 3016 -195 3021 -165
rect 2981 -200 3021 -195
rect 3221 -165 3261 -160
rect 3221 -195 3226 -165
rect 3256 -195 3261 -165
rect 3221 -200 3261 -195
rect 3466 -165 3506 -160
rect 3466 -195 3471 -165
rect 3501 -195 3506 -165
rect 3466 -200 3506 -195
rect 3706 -165 3746 -160
rect 3706 -195 3711 -165
rect 3741 -195 3746 -165
rect 3706 -200 3746 -195
rect 3951 -165 3991 -160
rect 3951 -195 3956 -165
rect 3986 -195 3991 -165
rect 4191 -165 4231 -160
rect 3951 -200 3991 -195
rect 4050 -195 4110 -185
rect 1625 -240 1635 -200
rect 1675 -240 1685 -200
rect 4050 -235 4060 -195
rect 4100 -235 4110 -195
rect 4191 -195 4196 -165
rect 4226 -195 4231 -165
rect 4191 -200 4231 -195
rect 4436 -165 4476 -160
rect 4436 -195 4441 -165
rect 4471 -195 4476 -165
rect 4436 -200 4476 -195
rect 4676 -165 4716 -160
rect 4676 -195 4681 -165
rect 4711 -195 4716 -165
rect 4676 -200 4716 -195
rect 4921 -165 4961 -160
rect 4921 -195 4926 -165
rect 4956 -195 4961 -165
rect 4921 -200 4961 -195
rect 5161 -165 5201 -160
rect 5161 -195 5166 -165
rect 5196 -195 5201 -165
rect 5161 -200 5201 -195
rect 5406 -165 5446 -160
rect 5406 -195 5411 -165
rect 5441 -195 5446 -165
rect 5406 -200 5446 -195
rect 5711 -165 5751 -160
rect 5711 -195 5716 -165
rect 5746 -195 5751 -165
rect 5711 -200 5751 -195
rect 5956 -165 5996 -160
rect 5956 -195 5961 -165
rect 5991 -195 5996 -165
rect 5956 -200 5996 -195
rect 6196 -165 6236 -160
rect 6196 -195 6201 -165
rect 6231 -195 6236 -165
rect 6196 -200 6236 -195
rect 6681 -165 6721 -160
rect 6681 -195 6686 -165
rect 6716 -195 6721 -165
rect 6681 -200 6721 -195
rect 6926 -165 6966 -160
rect 6926 -195 6931 -165
rect 6961 -195 6966 -165
rect 6926 -200 6966 -195
rect 7166 -165 7206 -160
rect 7166 -195 7171 -165
rect 7201 -195 7206 -165
rect 7166 -200 7206 -195
rect 7406 -165 7446 -160
rect 7406 -195 7411 -165
rect 7441 -195 7446 -165
rect 7406 -200 7446 -195
rect 7646 -165 7686 -160
rect 7646 -195 7651 -165
rect 7681 -195 7686 -165
rect 7646 -200 7686 -195
rect 8131 -165 8171 -160
rect 8131 -195 8136 -165
rect 8166 -195 8171 -165
rect 8131 -200 8171 -195
rect 8376 -165 8416 -160
rect 8376 -195 8381 -165
rect 8411 -195 8416 -165
rect 8376 -200 8416 -195
rect 8616 -165 8656 -160
rect 8616 -195 8621 -165
rect 8651 -195 8656 -165
rect 8616 -200 8656 -195
rect 8861 -165 8901 -160
rect 8861 -195 8866 -165
rect 8896 -195 8901 -165
rect 8861 -200 8901 -195
rect 9101 -165 9141 -160
rect 9101 -195 9106 -165
rect 9136 -195 9141 -165
rect 9101 -200 9141 -195
rect 9346 -165 9386 -160
rect 9346 -195 9351 -165
rect 9381 -195 9386 -165
rect 9346 -200 9386 -195
rect 9836 -165 9876 -160
rect 9836 -195 9841 -165
rect 9871 -195 9876 -165
rect 9836 -200 9876 -195
rect 10076 -165 10116 -160
rect 10076 -195 10081 -165
rect 10111 -195 10116 -165
rect 10076 -200 10116 -195
rect 10321 -165 10361 -160
rect 10321 -195 10326 -165
rect 10356 -195 10361 -165
rect 10321 -200 10361 -195
rect 10561 -165 10601 -160
rect 10561 -195 10566 -165
rect 10596 -195 10601 -165
rect 10561 -200 10601 -195
rect 10806 -165 10846 -160
rect 10806 -195 10811 -165
rect 10841 -195 10846 -165
rect 10806 -200 10846 -195
rect 11046 -165 11086 -160
rect 11046 -195 11051 -165
rect 11081 -195 11086 -165
rect 11046 -200 11086 -195
rect 11291 -165 11331 -160
rect 11291 -195 11296 -165
rect 11326 -195 11331 -165
rect 11291 -200 11331 -195
rect 11531 -165 11571 -160
rect 11531 -195 11536 -165
rect 11566 -195 11571 -165
rect 11531 -200 11571 -195
rect 11776 -165 11816 -160
rect 11776 -195 11781 -165
rect 11811 -195 11816 -165
rect 11776 -200 11816 -195
rect 12261 -165 12301 -160
rect 12261 -195 12266 -165
rect 12296 -195 12301 -165
rect 12261 -200 12301 -195
rect 12501 -165 12541 -160
rect 12501 -195 12506 -165
rect 12536 -195 12541 -165
rect 12501 -200 12541 -195
rect 12746 -165 12786 -160
rect 12746 -195 12751 -165
rect 12781 -195 12786 -165
rect 12746 -200 12786 -195
rect 12986 -165 13026 -160
rect 12986 -195 12991 -165
rect 13021 -195 13026 -165
rect 12986 -200 13026 -195
rect 13231 -165 13271 -160
rect 13231 -195 13236 -165
rect 13266 -195 13271 -165
rect 13231 -200 13271 -195
rect 13471 -165 13511 -160
rect 13471 -195 13476 -165
rect 13506 -195 13511 -165
rect 13471 -200 13511 -195
rect 13716 -165 13756 -160
rect 13716 -195 13721 -165
rect 13751 -195 13756 -165
rect 13716 -200 13756 -195
rect 14201 -165 14241 -160
rect 14201 -195 14206 -165
rect 14236 -195 14241 -165
rect 14201 -200 14241 -195
rect 14441 -165 14481 -160
rect 14441 -195 14446 -165
rect 14476 -195 14481 -165
rect 14441 -200 14481 -195
rect 14686 -165 14726 -160
rect 14686 -195 14691 -165
rect 14721 -195 14726 -165
rect 14686 -200 14726 -195
rect 14926 -165 14966 -160
rect 14926 -195 14931 -165
rect 14961 -195 14966 -165
rect 14926 -200 14966 -195
rect 15171 -165 15211 -160
rect 15171 -195 15176 -165
rect 15206 -195 15211 -165
rect 15171 -200 15211 -195
rect 15411 -165 15451 -160
rect 15411 -195 15416 -165
rect 15446 -195 15451 -165
rect 15411 -200 15451 -195
rect 15656 -165 15696 -160
rect 15656 -195 15661 -165
rect 15691 -195 15696 -165
rect 15656 -200 15696 -195
rect 16141 -165 16181 -160
rect 16141 -195 16146 -165
rect 16176 -195 16181 -165
rect 16141 -200 16181 -195
rect 16381 -165 16421 -160
rect 16381 -195 16386 -165
rect 16416 -195 16421 -165
rect 16381 -200 16421 -195
rect 16626 -165 16666 -160
rect 16626 -195 16631 -165
rect 16661 -195 16666 -165
rect 16626 -200 16666 -195
rect 16866 -165 16906 -160
rect 16866 -195 16871 -165
rect 16901 -195 16906 -165
rect 16866 -200 16906 -195
rect 17111 -165 17151 -160
rect 17111 -195 17116 -165
rect 17146 -195 17151 -165
rect 17111 -200 17151 -195
rect 17351 -165 17391 -160
rect 17351 -195 17356 -165
rect 17386 -195 17391 -165
rect 17351 -200 17391 -195
rect 17596 -165 17636 -160
rect 17596 -195 17601 -165
rect 17631 -195 17636 -165
rect 17596 -200 17636 -195
rect 17836 -165 17876 -160
rect 17836 -195 17841 -165
rect 17871 -195 17876 -165
rect 17836 -200 17876 -195
rect 18081 -165 18121 -160
rect 18081 -195 18086 -165
rect 18116 -195 18121 -165
rect 18081 -200 18121 -195
rect 18321 -165 18361 -160
rect 18321 -195 18326 -165
rect 18356 -195 18361 -165
rect 18321 -200 18361 -195
rect 18566 -165 18606 -160
rect 18566 -195 18571 -165
rect 18601 -195 18606 -165
rect 18566 -200 18606 -195
rect 18806 -165 18846 -160
rect 18806 -195 18811 -165
rect 18841 -195 18846 -165
rect 18806 -200 18846 -195
rect 19051 -165 19091 -160
rect 19051 -195 19056 -165
rect 19086 -195 19091 -165
rect 19051 -200 19091 -195
rect 19291 -165 19331 -160
rect 19291 -195 19296 -165
rect 19326 -195 19331 -165
rect 19291 -200 19331 -195
rect 19536 -165 19576 -160
rect 19536 -195 19541 -165
rect 19571 -195 19576 -165
rect 19536 -200 19576 -195
rect 19776 -165 19816 -160
rect 19776 -195 19781 -165
rect 19811 -195 19816 -165
rect 19776 -200 19816 -195
rect 20021 -165 20061 -160
rect 20021 -195 20026 -165
rect 20056 -195 20061 -165
rect 20021 -200 20061 -195
rect 20261 -165 20301 -160
rect 20261 -195 20266 -165
rect 20296 -195 20301 -165
rect 20261 -200 20301 -195
rect 20506 -165 20546 -160
rect 20506 -195 20511 -165
rect 20541 -195 20546 -165
rect 20506 -200 20546 -195
rect 20746 -165 20786 -160
rect 20746 -195 20751 -165
rect 20781 -195 20786 -165
rect 20746 -200 20786 -195
rect 20991 -165 21031 -160
rect 20991 -195 20996 -165
rect 21026 -195 21031 -165
rect 20991 -200 21031 -195
rect 9560 -210 9620 -200
rect 17695 -210 17755 -200
rect -425 -250 -355 -240
rect 85 -245 125 -240
rect 85 -275 90 -245
rect 120 -275 125 -245
rect 85 -280 125 -275
rect 325 -245 365 -240
rect 325 -275 330 -245
rect 360 -275 365 -245
rect 325 -280 365 -275
rect 565 -245 605 -240
rect 565 -275 570 -245
rect 600 -275 605 -245
rect 565 -280 605 -275
rect 805 -245 845 -240
rect 805 -275 810 -245
rect 840 -275 845 -245
rect 805 -280 845 -275
rect 1045 -245 1085 -240
rect 1045 -275 1050 -245
rect 1080 -275 1085 -245
rect 1045 -280 1085 -275
rect 1285 -245 1325 -240
rect 1285 -275 1290 -245
rect 1320 -275 1325 -245
rect 1285 -280 1325 -275
rect 1525 -245 1565 -240
rect 1525 -275 1530 -245
rect 1560 -275 1565 -245
rect 1625 -250 1685 -240
rect 1765 -245 1805 -240
rect 1525 -280 1565 -275
rect 1765 -275 1770 -245
rect 1800 -275 1805 -245
rect 1765 -280 1805 -275
rect 2005 -245 2045 -240
rect 2005 -275 2010 -245
rect 2040 -275 2045 -245
rect 2005 -280 2045 -275
rect 2245 -245 2285 -240
rect 2245 -275 2250 -245
rect 2280 -275 2285 -245
rect 2245 -280 2285 -275
rect 2485 -245 2525 -240
rect 2485 -275 2490 -245
rect 2520 -275 2525 -245
rect 2485 -280 2525 -275
rect 2725 -245 2765 -240
rect 2725 -275 2730 -245
rect 2760 -275 2765 -245
rect 2725 -280 2765 -275
rect 2965 -245 3005 -240
rect 2965 -275 2970 -245
rect 3000 -275 3005 -245
rect 2965 -280 3005 -275
rect 3205 -245 3245 -240
rect 3205 -275 3210 -245
rect 3240 -275 3245 -245
rect 3205 -280 3245 -275
rect 3445 -245 3485 -240
rect 3445 -275 3450 -245
rect 3480 -275 3485 -245
rect 3445 -280 3485 -275
rect 3685 -245 3725 -240
rect 3685 -275 3690 -245
rect 3720 -275 3725 -245
rect 3685 -280 3725 -275
rect 3925 -245 3965 -240
rect 4050 -245 4110 -235
rect 6445 -220 6505 -210
rect 4165 -245 4205 -240
rect 3925 -275 3930 -245
rect 3960 -275 3965 -245
rect 3925 -280 3965 -275
rect 4165 -275 4170 -245
rect 4200 -275 4205 -245
rect 4165 -280 4205 -275
rect 4405 -245 4445 -240
rect 4405 -275 4410 -245
rect 4440 -275 4445 -245
rect 4405 -280 4445 -275
rect 4645 -245 4685 -240
rect 4645 -275 4650 -245
rect 4680 -275 4685 -245
rect 4645 -280 4685 -275
rect 4885 -245 4925 -240
rect 4885 -275 4890 -245
rect 4920 -275 4925 -245
rect 4885 -280 4925 -275
rect 5125 -245 5165 -240
rect 5125 -275 5130 -245
rect 5160 -275 5165 -245
rect 5125 -280 5165 -275
rect 5365 -245 5405 -240
rect 5365 -275 5370 -245
rect 5400 -275 5405 -245
rect 5365 -280 5405 -275
rect 5605 -245 5645 -240
rect 5605 -275 5610 -245
rect 5640 -275 5645 -245
rect 5605 -280 5645 -275
rect 5845 -245 5885 -240
rect 5845 -275 5850 -245
rect 5880 -275 5885 -245
rect 5845 -280 5885 -275
rect 6085 -245 6125 -240
rect 6085 -275 6090 -245
rect 6120 -275 6125 -245
rect 6085 -280 6125 -275
rect 6325 -245 6365 -240
rect 6325 -275 6330 -245
rect 6360 -275 6365 -245
rect 6445 -260 6455 -220
rect 6495 -260 6505 -220
rect 7870 -220 7930 -210
rect 6445 -270 6505 -260
rect 6565 -245 6605 -240
rect 6325 -280 6365 -275
rect 6565 -275 6570 -245
rect 6600 -275 6605 -245
rect 6565 -280 6605 -275
rect 6805 -245 6845 -240
rect 6805 -275 6810 -245
rect 6840 -275 6845 -245
rect 6805 -280 6845 -275
rect 7045 -245 7085 -240
rect 7045 -275 7050 -245
rect 7080 -275 7085 -245
rect 7045 -280 7085 -275
rect 7285 -245 7325 -240
rect 7285 -275 7290 -245
rect 7320 -275 7325 -245
rect 7285 -280 7325 -275
rect 7525 -245 7565 -240
rect 7525 -275 7530 -245
rect 7560 -275 7565 -245
rect 7525 -280 7565 -275
rect 7765 -245 7805 -240
rect 7765 -275 7770 -245
rect 7800 -275 7805 -245
rect 7870 -260 7880 -220
rect 7920 -260 7930 -220
rect 7870 -270 7930 -260
rect 8005 -245 8045 -240
rect 7765 -280 7805 -275
rect 8005 -275 8010 -245
rect 8040 -275 8045 -245
rect 8005 -280 8045 -275
rect 8245 -245 8285 -240
rect 8245 -275 8250 -245
rect 8280 -275 8285 -245
rect 8245 -280 8285 -275
rect 8485 -245 8525 -240
rect 8485 -275 8490 -245
rect 8520 -275 8525 -245
rect 8485 -280 8525 -275
rect 8725 -245 8765 -240
rect 8725 -275 8730 -245
rect 8760 -275 8765 -245
rect 8725 -280 8765 -275
rect 8965 -245 9005 -240
rect 8965 -275 8970 -245
rect 9000 -275 9005 -245
rect 8965 -280 9005 -275
rect 9205 -245 9245 -240
rect 9205 -275 9210 -245
rect 9240 -275 9245 -245
rect 9205 -280 9245 -275
rect 9445 -245 9485 -240
rect 9445 -275 9450 -245
rect 9480 -275 9485 -245
rect 9560 -250 9570 -210
rect 9610 -250 9620 -210
rect 11940 -220 12000 -210
rect 9560 -260 9620 -250
rect 9685 -245 9725 -240
rect 9445 -280 9485 -275
rect 9685 -275 9690 -245
rect 9720 -275 9725 -245
rect 9685 -280 9725 -275
rect 9925 -245 9965 -240
rect 9925 -275 9930 -245
rect 9960 -275 9965 -245
rect 9925 -280 9965 -275
rect 10165 -245 10205 -240
rect 10165 -275 10170 -245
rect 10200 -275 10205 -245
rect 10165 -280 10205 -275
rect 10405 -245 10445 -240
rect 10405 -275 10410 -245
rect 10440 -275 10445 -245
rect 10405 -280 10445 -275
rect 10645 -245 10685 -240
rect 10645 -275 10650 -245
rect 10680 -275 10685 -245
rect 10645 -280 10685 -275
rect 10885 -245 10925 -240
rect 10885 -275 10890 -245
rect 10920 -275 10925 -245
rect 10885 -280 10925 -275
rect 11125 -245 11165 -240
rect 11125 -275 11130 -245
rect 11160 -275 11165 -245
rect 11125 -280 11165 -275
rect 11365 -245 11405 -240
rect 11365 -275 11370 -245
rect 11400 -275 11405 -245
rect 11365 -280 11405 -275
rect 11605 -245 11645 -240
rect 11605 -275 11610 -245
rect 11640 -275 11645 -245
rect 11605 -280 11645 -275
rect 11845 -245 11885 -240
rect 11845 -275 11850 -245
rect 11880 -275 11885 -245
rect 11940 -260 11950 -220
rect 11990 -260 12000 -220
rect 13860 -220 13920 -210
rect 11940 -270 12000 -260
rect 12085 -245 12125 -240
rect 11845 -280 11885 -275
rect 12085 -275 12090 -245
rect 12120 -275 12125 -245
rect 12085 -280 12125 -275
rect 12325 -245 12365 -240
rect 12325 -275 12330 -245
rect 12360 -275 12365 -245
rect 12325 -280 12365 -275
rect 12565 -245 12605 -240
rect 12565 -275 12570 -245
rect 12600 -275 12605 -245
rect 12565 -280 12605 -275
rect 12805 -245 12845 -240
rect 12805 -275 12810 -245
rect 12840 -275 12845 -245
rect 12805 -280 12845 -275
rect 13045 -245 13085 -240
rect 13045 -275 13050 -245
rect 13080 -275 13085 -245
rect 13045 -280 13085 -275
rect 13285 -245 13325 -240
rect 13285 -275 13290 -245
rect 13320 -275 13325 -245
rect 13285 -280 13325 -275
rect 13525 -245 13565 -240
rect 13525 -275 13530 -245
rect 13560 -275 13565 -245
rect 13525 -280 13565 -275
rect 13765 -245 13805 -240
rect 13765 -275 13770 -245
rect 13800 -275 13805 -245
rect 13860 -260 13870 -220
rect 13910 -260 13920 -220
rect 15805 -220 15865 -210
rect 13860 -270 13920 -260
rect 14005 -245 14045 -240
rect 13765 -280 13805 -275
rect 14005 -275 14010 -245
rect 14040 -275 14045 -245
rect 14005 -280 14045 -275
rect 14245 -245 14285 -240
rect 14245 -275 14250 -245
rect 14280 -275 14285 -245
rect 14245 -280 14285 -275
rect 14485 -245 14525 -240
rect 14485 -275 14490 -245
rect 14520 -275 14525 -245
rect 14485 -280 14525 -275
rect 14725 -245 14765 -240
rect 14725 -275 14730 -245
rect 14760 -275 14765 -245
rect 14725 -280 14765 -275
rect 14965 -245 15005 -240
rect 14965 -275 14970 -245
rect 15000 -275 15005 -245
rect 14965 -280 15005 -275
rect 15205 -245 15245 -240
rect 15205 -275 15210 -245
rect 15240 -275 15245 -245
rect 15205 -280 15245 -275
rect 15445 -245 15485 -240
rect 15445 -275 15450 -245
rect 15480 -275 15485 -245
rect 15445 -280 15485 -275
rect 15685 -245 15725 -240
rect 15685 -275 15690 -245
rect 15720 -275 15725 -245
rect 15805 -260 15815 -220
rect 15855 -260 15865 -220
rect 15805 -270 15865 -260
rect 15925 -245 15965 -240
rect 15685 -280 15725 -275
rect 15925 -275 15930 -245
rect 15960 -275 15965 -245
rect 15925 -280 15965 -275
rect 16165 -245 16205 -240
rect 16165 -275 16170 -245
rect 16200 -275 16205 -245
rect 16165 -280 16205 -275
rect 16405 -245 16445 -240
rect 16405 -275 16410 -245
rect 16440 -275 16445 -245
rect 16405 -280 16445 -275
rect 16645 -245 16685 -240
rect 16645 -275 16650 -245
rect 16680 -275 16685 -245
rect 16645 -280 16685 -275
rect 16885 -245 16925 -240
rect 16885 -275 16890 -245
rect 16920 -275 16925 -245
rect 16885 -280 16925 -275
rect 17125 -245 17165 -240
rect 17125 -275 17130 -245
rect 17160 -275 17165 -245
rect 17125 -280 17165 -275
rect 17365 -245 17405 -240
rect 17365 -275 17370 -245
rect 17400 -275 17405 -245
rect 17365 -280 17405 -275
rect 17605 -245 17645 -240
rect 17605 -275 17610 -245
rect 17640 -275 17645 -245
rect 17695 -250 17705 -210
rect 17745 -250 17755 -210
rect 19635 -210 19695 -200
rect 17695 -260 17755 -250
rect 17845 -245 17885 -240
rect 17605 -280 17645 -275
rect 17845 -275 17850 -245
rect 17880 -275 17885 -245
rect 17845 -280 17885 -275
rect 18085 -245 18125 -240
rect 18085 -275 18090 -245
rect 18120 -275 18125 -245
rect 18085 -280 18125 -275
rect 18325 -245 18365 -240
rect 18325 -275 18330 -245
rect 18360 -275 18365 -245
rect 18325 -280 18365 -275
rect 18565 -245 18605 -240
rect 18565 -275 18570 -245
rect 18600 -275 18605 -245
rect 18565 -280 18605 -275
rect 18805 -245 18845 -240
rect 18805 -275 18810 -245
rect 18840 -275 18845 -245
rect 18805 -280 18845 -275
rect 19045 -245 19085 -240
rect 19045 -275 19050 -245
rect 19080 -275 19085 -245
rect 19045 -280 19085 -275
rect 19285 -245 19325 -240
rect 19285 -275 19290 -245
rect 19320 -275 19325 -245
rect 19285 -280 19325 -275
rect 19525 -245 19565 -240
rect 19525 -275 19530 -245
rect 19560 -275 19565 -245
rect 19635 -250 19645 -210
rect 19685 -250 19695 -210
rect 19635 -260 19695 -250
rect 19765 -245 19805 -240
rect 19525 -280 19565 -275
rect 19765 -275 19770 -245
rect 19800 -275 19805 -245
rect 19765 -280 19805 -275
rect 20005 -245 20045 -240
rect 20005 -275 20010 -245
rect 20040 -275 20045 -245
rect 20005 -280 20045 -275
rect 20245 -245 20285 -240
rect 20245 -275 20250 -245
rect 20280 -275 20285 -245
rect 20245 -280 20285 -275
rect 20485 -245 20525 -240
rect 20485 -275 20490 -245
rect 20520 -275 20525 -245
rect 20485 -280 20525 -275
rect 20725 -245 20765 -240
rect 20725 -275 20730 -245
rect 20760 -275 20765 -245
rect 20725 -280 20765 -275
rect 20965 -245 21005 -240
rect 20965 -275 20970 -245
rect 21000 -275 21005 -245
rect 20965 -280 21005 -275
rect 21205 -245 21245 -240
rect 21205 -275 21210 -245
rect 21240 -275 21245 -245
rect 21205 -280 21245 -275
rect 21445 -245 21485 -240
rect 21445 -275 21450 -245
rect 21480 -275 21485 -245
rect 21445 -280 21485 -275
rect 21685 -245 21725 -240
rect 21685 -275 21690 -245
rect 21720 -275 21725 -245
rect 21685 -280 21725 -275
rect 21925 -245 21965 -240
rect 21925 -275 21930 -245
rect 21960 -275 21965 -245
rect 21925 -280 21965 -275
rect 22165 -245 22205 -240
rect 22165 -275 22170 -245
rect 22200 -275 22205 -245
rect 22165 -280 22205 -275
rect 22405 -245 22445 -240
rect 22405 -275 22410 -245
rect 22440 -275 22445 -245
rect 22405 -280 22445 -275
rect 22645 -245 22685 -240
rect 22645 -275 22650 -245
rect 22680 -275 22685 -245
rect 22645 -280 22685 -275
rect 22885 -245 22925 -240
rect 22885 -275 22890 -245
rect 22920 -275 22925 -245
rect 22885 -280 22925 -275
rect 23125 -245 23165 -240
rect 23125 -275 23130 -245
rect 23160 -275 23165 -245
rect 23125 -280 23165 -275
rect 23365 -245 23405 -240
rect 23365 -275 23370 -245
rect 23400 -275 23405 -245
rect 23365 -280 23405 -275
rect 23605 -245 23645 -240
rect 23605 -275 23610 -245
rect 23640 -275 23645 -245
rect 23605 -280 23645 -275
rect 23845 -245 23885 -240
rect 23845 -275 23850 -245
rect 23880 -275 23885 -245
rect 23845 -280 23885 -275
rect 24085 -245 24125 -240
rect 24085 -275 24090 -245
rect 24120 -275 24125 -245
rect 24085 -280 24125 -275
rect 24325 -245 24365 -240
rect 24325 -275 24330 -245
rect 24360 -275 24365 -245
rect 24325 -280 24365 -275
rect 24565 -245 24605 -240
rect 24565 -275 24570 -245
rect 24600 -275 24605 -245
rect 24565 -280 24605 -275
rect 24805 -245 24845 -240
rect 24805 -275 24810 -245
rect 24840 -275 24845 -245
rect 24805 -280 24845 -275
rect 25045 -245 25085 -240
rect 25045 -275 25050 -245
rect 25080 -275 25085 -245
rect 25045 -280 25085 -275
rect 25285 -245 25325 -240
rect 25285 -275 25290 -245
rect 25320 -275 25325 -245
rect 25285 -280 25325 -275
rect 25525 -245 25565 -240
rect 25525 -275 25530 -245
rect 25560 -275 25565 -245
rect 25525 -280 25565 -275
rect 25765 -245 25805 -240
rect 25765 -275 25770 -245
rect 25800 -275 25805 -245
rect 25765 -280 25805 -275
rect 26005 -245 26045 -240
rect 26005 -275 26010 -245
rect 26040 -275 26045 -245
rect 26005 -280 26045 -275
rect 26245 -245 26285 -240
rect 26245 -275 26250 -245
rect 26280 -275 26285 -245
rect 26245 -280 26285 -275
rect 26485 -245 26525 -240
rect 26485 -275 26490 -245
rect 26520 -275 26525 -245
rect 26485 -280 26525 -275
rect 26725 -245 26765 -240
rect 26725 -275 26730 -245
rect 26760 -275 26765 -245
rect 26725 -280 26765 -275
rect 26965 -245 27005 -240
rect 26965 -275 26970 -245
rect 27000 -275 27005 -245
rect 26965 -280 27005 -275
rect 27205 -245 27245 -240
rect 27205 -275 27210 -245
rect 27240 -275 27245 -245
rect 27205 -280 27245 -275
rect 27445 -245 27485 -240
rect 27445 -275 27450 -245
rect 27480 -275 27485 -245
rect 27445 -280 27485 -275
rect 27685 -245 27725 -240
rect 27685 -275 27690 -245
rect 27720 -275 27725 -245
rect 27685 -280 27725 -275
rect 27925 -245 27965 -240
rect 27925 -275 27930 -245
rect 27960 -275 27965 -245
rect 27925 -280 27965 -275
rect 28165 -245 28205 -240
rect 28165 -275 28170 -245
rect 28200 -275 28205 -245
rect 28165 -280 28205 -275
rect 28405 -245 28445 -240
rect 28405 -275 28410 -245
rect 28440 -275 28445 -245
rect 28405 -280 28445 -275
rect 28645 -245 28685 -240
rect 28645 -275 28650 -245
rect 28680 -275 28685 -245
rect 28645 -280 28685 -275
rect 28885 -245 28925 -240
rect 28885 -275 28890 -245
rect 28920 -275 28925 -245
rect 28885 -280 28925 -275
rect 29125 -245 29165 -240
rect 29125 -275 29130 -245
rect 29160 -275 29165 -245
rect 29125 -280 29165 -275
rect 29365 -245 29405 -240
rect 29365 -275 29370 -245
rect 29400 -275 29405 -245
rect 29365 -280 29405 -275
rect 29605 -245 29645 -240
rect 29605 -275 29610 -245
rect 29640 -275 29645 -245
rect 29605 -280 29645 -275
rect 29845 -245 29885 -240
rect 29845 -275 29850 -245
rect 29880 -275 29885 -245
rect 29845 -280 29885 -275
rect 30085 -245 30125 -240
rect 30085 -275 30090 -245
rect 30120 -275 30125 -245
rect 30085 -280 30125 -275
rect 30325 -245 30365 -240
rect 30325 -275 30330 -245
rect 30360 -275 30365 -245
rect 30325 -280 30365 -275
rect 30565 -245 30605 -240
rect 30565 -275 30570 -245
rect 30600 -275 30605 -245
rect 30565 -280 30605 -275
rect 15 -295 55 -290
rect 15 -315 25 -295
rect 45 -305 55 -295
rect 135 -295 175 -290
rect 135 -305 145 -295
rect 45 -315 145 -305
rect 165 -305 175 -295
rect 255 -295 295 -290
rect 255 -305 265 -295
rect 165 -315 265 -305
rect 285 -305 295 -295
rect 375 -295 415 -290
rect 375 -305 385 -295
rect 285 -315 385 -305
rect 405 -305 415 -295
rect 495 -295 535 -290
rect 495 -305 505 -295
rect 405 -315 505 -305
rect 525 -305 535 -295
rect 615 -295 655 -290
rect 615 -305 625 -295
rect 525 -315 625 -305
rect 645 -305 655 -295
rect 735 -295 775 -290
rect 735 -305 745 -295
rect 645 -315 745 -305
rect 765 -305 775 -295
rect 855 -295 895 -290
rect 855 -305 865 -295
rect 765 -315 865 -305
rect 885 -305 895 -295
rect 975 -295 1015 -290
rect 975 -305 985 -295
rect 885 -315 985 -305
rect 1005 -305 1015 -295
rect 1095 -295 1135 -290
rect 1095 -305 1105 -295
rect 1005 -315 1105 -305
rect 1125 -305 1135 -295
rect 1215 -295 1255 -290
rect 1215 -305 1225 -295
rect 1125 -315 1225 -305
rect 1245 -305 1255 -295
rect 1335 -295 1375 -290
rect 1335 -305 1345 -295
rect 1245 -315 1345 -305
rect 1365 -305 1375 -295
rect 1455 -295 1495 -290
rect 1455 -305 1465 -295
rect 1365 -315 1465 -305
rect 1485 -305 1495 -295
rect 1575 -295 1615 -290
rect 1575 -305 1585 -295
rect 1485 -315 1585 -305
rect 1605 -305 1615 -295
rect 1695 -295 1735 -290
rect 1695 -305 1705 -295
rect 1605 -315 1705 -305
rect 1725 -305 1735 -295
rect 1815 -295 1855 -290
rect 1815 -305 1825 -295
rect 1725 -315 1825 -305
rect 1845 -305 1855 -295
rect 1935 -295 1975 -290
rect 1935 -305 1945 -295
rect 1845 -315 1945 -305
rect 1965 -305 1975 -295
rect 2055 -295 2095 -290
rect 2055 -305 2065 -295
rect 1965 -315 2065 -305
rect 2085 -305 2095 -295
rect 2175 -295 2215 -290
rect 2175 -305 2185 -295
rect 2085 -315 2185 -305
rect 2205 -305 2215 -295
rect 2295 -295 2335 -290
rect 2295 -305 2305 -295
rect 2205 -315 2305 -305
rect 2325 -305 2335 -295
rect 2415 -295 2455 -290
rect 2415 -305 2425 -295
rect 2325 -315 2425 -305
rect 2445 -305 2455 -295
rect 2535 -295 2575 -290
rect 2535 -305 2545 -295
rect 2445 -315 2545 -305
rect 2565 -305 2575 -295
rect 2655 -295 2695 -290
rect 2655 -305 2665 -295
rect 2565 -315 2665 -305
rect 2685 -305 2695 -295
rect 2775 -295 2815 -290
rect 2775 -305 2785 -295
rect 2685 -315 2785 -305
rect 2805 -305 2815 -295
rect 2895 -295 2935 -290
rect 2895 -305 2905 -295
rect 2805 -315 2905 -305
rect 2925 -305 2935 -295
rect 3015 -295 3055 -290
rect 3015 -305 3025 -295
rect 2925 -315 3025 -305
rect 3045 -305 3055 -295
rect 3135 -295 3175 -290
rect 3135 -305 3145 -295
rect 3045 -315 3145 -305
rect 3165 -305 3175 -295
rect 3255 -295 3295 -290
rect 3255 -305 3265 -295
rect 3165 -315 3265 -305
rect 3285 -305 3295 -295
rect 3375 -295 3415 -290
rect 3375 -305 3385 -295
rect 3285 -315 3385 -305
rect 3405 -305 3415 -295
rect 3495 -295 3535 -290
rect 3495 -305 3505 -295
rect 3405 -315 3505 -305
rect 3525 -305 3535 -295
rect 3615 -295 3655 -290
rect 3615 -305 3625 -295
rect 3525 -315 3625 -305
rect 3645 -305 3655 -295
rect 3735 -295 3775 -290
rect 3735 -305 3745 -295
rect 3645 -315 3745 -305
rect 3765 -305 3775 -295
rect 3855 -295 3895 -290
rect 3855 -305 3865 -295
rect 3765 -315 3865 -305
rect 3885 -305 3895 -295
rect 3975 -295 4015 -290
rect 3975 -305 3985 -295
rect 3885 -315 3985 -305
rect 4005 -305 4015 -295
rect 4095 -295 4135 -290
rect 4095 -305 4105 -295
rect 4005 -315 4105 -305
rect 4125 -305 4135 -295
rect 4215 -295 4255 -290
rect 4215 -305 4225 -295
rect 4125 -315 4225 -305
rect 4245 -305 4255 -295
rect 4335 -295 4375 -290
rect 4335 -305 4345 -295
rect 4245 -315 4345 -305
rect 4365 -305 4375 -295
rect 4455 -295 4495 -290
rect 4455 -305 4465 -295
rect 4365 -315 4465 -305
rect 4485 -305 4495 -295
rect 4575 -295 4615 -290
rect 4575 -305 4585 -295
rect 4485 -315 4585 -305
rect 4605 -305 4615 -295
rect 4695 -295 4735 -290
rect 4695 -305 4705 -295
rect 4605 -315 4705 -305
rect 4725 -305 4735 -295
rect 4815 -295 4855 -290
rect 4815 -305 4825 -295
rect 4725 -315 4825 -305
rect 4845 -305 4855 -295
rect 4935 -295 4975 -290
rect 4935 -305 4945 -295
rect 4845 -315 4945 -305
rect 4965 -305 4975 -295
rect 5055 -295 5095 -290
rect 5055 -305 5065 -295
rect 4965 -315 5065 -305
rect 5085 -305 5095 -295
rect 5175 -295 5215 -290
rect 5175 -305 5185 -295
rect 5085 -315 5185 -305
rect 5205 -305 5215 -295
rect 5295 -295 5335 -290
rect 5295 -305 5305 -295
rect 5205 -315 5305 -305
rect 5325 -305 5335 -295
rect 5415 -295 5455 -290
rect 5415 -305 5425 -295
rect 5325 -315 5425 -305
rect 5445 -305 5455 -295
rect 5535 -295 5575 -290
rect 5535 -305 5545 -295
rect 5445 -315 5545 -305
rect 5565 -305 5575 -295
rect 5655 -295 5695 -290
rect 5655 -305 5665 -295
rect 5565 -315 5665 -305
rect 5685 -305 5695 -295
rect 5775 -295 5815 -290
rect 5775 -305 5785 -295
rect 5685 -315 5785 -305
rect 5805 -305 5815 -295
rect 5895 -295 5935 -290
rect 5895 -305 5905 -295
rect 5805 -315 5905 -305
rect 5925 -305 5935 -295
rect 6015 -295 6055 -290
rect 6015 -305 6025 -295
rect 5925 -315 6025 -305
rect 6045 -305 6055 -295
rect 6135 -295 6175 -290
rect 6135 -305 6145 -295
rect 6045 -315 6145 -305
rect 6165 -305 6175 -295
rect 6255 -295 6295 -290
rect 6255 -305 6265 -295
rect 6165 -315 6265 -305
rect 6285 -305 6295 -295
rect 6375 -295 6415 -290
rect 6375 -305 6385 -295
rect 6285 -315 6385 -305
rect 6405 -305 6415 -295
rect 6495 -295 6535 -290
rect 6495 -305 6505 -295
rect 6405 -315 6505 -305
rect 6525 -305 6535 -295
rect 6615 -295 6655 -290
rect 6615 -305 6625 -295
rect 6525 -315 6625 -305
rect 6645 -305 6655 -295
rect 6735 -295 6775 -290
rect 6735 -305 6745 -295
rect 6645 -315 6745 -305
rect 6765 -305 6775 -295
rect 6855 -295 6895 -290
rect 6855 -305 6865 -295
rect 6765 -315 6865 -305
rect 6885 -305 6895 -295
rect 6975 -295 7015 -290
rect 6975 -305 6985 -295
rect 6885 -315 6985 -305
rect 7005 -305 7015 -295
rect 7095 -295 7135 -290
rect 7095 -305 7105 -295
rect 7005 -315 7105 -305
rect 7125 -305 7135 -295
rect 7215 -295 7255 -290
rect 7215 -305 7225 -295
rect 7125 -315 7225 -305
rect 7245 -305 7255 -295
rect 7335 -295 7375 -290
rect 7335 -305 7345 -295
rect 7245 -315 7345 -305
rect 7365 -305 7375 -295
rect 7455 -295 7495 -290
rect 7455 -305 7465 -295
rect 7365 -315 7465 -305
rect 7485 -305 7495 -295
rect 7575 -295 7615 -290
rect 7575 -305 7585 -295
rect 7485 -315 7585 -305
rect 7605 -305 7615 -295
rect 7695 -295 7735 -290
rect 7695 -305 7705 -295
rect 7605 -315 7705 -305
rect 7725 -305 7735 -295
rect 7815 -295 7855 -290
rect 7815 -305 7825 -295
rect 7725 -315 7825 -305
rect 7845 -305 7855 -295
rect 7935 -295 7975 -290
rect 7935 -305 7945 -295
rect 7845 -315 7945 -305
rect 7965 -305 7975 -295
rect 8055 -295 8095 -290
rect 8055 -305 8065 -295
rect 7965 -315 8065 -305
rect 8085 -305 8095 -295
rect 8175 -295 8215 -290
rect 8175 -305 8185 -295
rect 8085 -315 8185 -305
rect 8205 -305 8215 -295
rect 8295 -295 8335 -290
rect 8295 -305 8305 -295
rect 8205 -315 8305 -305
rect 8325 -305 8335 -295
rect 8415 -295 8455 -290
rect 8415 -305 8425 -295
rect 8325 -315 8425 -305
rect 8445 -305 8455 -295
rect 8535 -295 8575 -290
rect 8535 -305 8545 -295
rect 8445 -315 8545 -305
rect 8565 -305 8575 -295
rect 8655 -295 8695 -290
rect 8655 -305 8665 -295
rect 8565 -315 8665 -305
rect 8685 -305 8695 -295
rect 8775 -295 8815 -290
rect 8775 -305 8785 -295
rect 8685 -315 8785 -305
rect 8805 -305 8815 -295
rect 8895 -295 8935 -290
rect 8895 -305 8905 -295
rect 8805 -315 8905 -305
rect 8925 -305 8935 -295
rect 9015 -295 9055 -290
rect 9015 -305 9025 -295
rect 8925 -315 9025 -305
rect 9045 -305 9055 -295
rect 9135 -295 9175 -290
rect 9135 -305 9145 -295
rect 9045 -315 9145 -305
rect 9165 -305 9175 -295
rect 9255 -295 9295 -290
rect 9255 -305 9265 -295
rect 9165 -315 9265 -305
rect 9285 -305 9295 -295
rect 9375 -295 9415 -290
rect 9375 -305 9385 -295
rect 9285 -315 9385 -305
rect 9405 -305 9415 -295
rect 9495 -295 9535 -290
rect 9495 -305 9505 -295
rect 9405 -315 9505 -305
rect 9525 -305 9535 -295
rect 9615 -295 9655 -290
rect 9615 -305 9625 -295
rect 9525 -315 9625 -305
rect 9645 -305 9655 -295
rect 9735 -295 9775 -290
rect 9735 -305 9745 -295
rect 9645 -315 9745 -305
rect 9765 -305 9775 -295
rect 9855 -295 9895 -290
rect 9855 -305 9865 -295
rect 9765 -315 9865 -305
rect 9885 -305 9895 -295
rect 9975 -295 10015 -290
rect 9975 -305 9985 -295
rect 9885 -315 9985 -305
rect 10005 -305 10015 -295
rect 10095 -295 10135 -290
rect 10095 -305 10105 -295
rect 10005 -315 10105 -305
rect 10125 -305 10135 -295
rect 10215 -295 10255 -290
rect 10215 -305 10225 -295
rect 10125 -315 10225 -305
rect 10245 -305 10255 -295
rect 10335 -295 10375 -290
rect 10335 -305 10345 -295
rect 10245 -315 10345 -305
rect 10365 -305 10375 -295
rect 10455 -295 10495 -290
rect 10455 -305 10465 -295
rect 10365 -315 10465 -305
rect 10485 -305 10495 -295
rect 10575 -295 10615 -290
rect 10575 -305 10585 -295
rect 10485 -315 10585 -305
rect 10605 -305 10615 -295
rect 10695 -295 10735 -290
rect 10695 -305 10705 -295
rect 10605 -315 10705 -305
rect 10725 -305 10735 -295
rect 10815 -295 10855 -290
rect 10815 -305 10825 -295
rect 10725 -315 10825 -305
rect 10845 -305 10855 -295
rect 10935 -295 10975 -290
rect 10935 -305 10945 -295
rect 10845 -315 10945 -305
rect 10965 -305 10975 -295
rect 11055 -295 11095 -290
rect 11055 -305 11065 -295
rect 10965 -315 11065 -305
rect 11085 -305 11095 -295
rect 11175 -295 11215 -290
rect 11175 -305 11185 -295
rect 11085 -315 11185 -305
rect 11205 -305 11215 -295
rect 11295 -295 11335 -290
rect 11295 -305 11305 -295
rect 11205 -315 11305 -305
rect 11325 -305 11335 -295
rect 11415 -295 11455 -290
rect 11415 -305 11425 -295
rect 11325 -315 11425 -305
rect 11445 -305 11455 -295
rect 11535 -295 11575 -290
rect 11535 -305 11545 -295
rect 11445 -315 11545 -305
rect 11565 -305 11575 -295
rect 11655 -295 11695 -290
rect 11655 -305 11665 -295
rect 11565 -315 11665 -305
rect 11685 -305 11695 -295
rect 11775 -295 11815 -290
rect 11775 -305 11785 -295
rect 11685 -315 11785 -305
rect 11805 -305 11815 -295
rect 11895 -295 11935 -290
rect 11895 -305 11905 -295
rect 11805 -315 11905 -305
rect 11925 -305 11935 -295
rect 12015 -295 12055 -290
rect 12015 -305 12025 -295
rect 11925 -315 12025 -305
rect 12045 -305 12055 -295
rect 12135 -295 12175 -290
rect 12135 -305 12145 -295
rect 12045 -315 12145 -305
rect 12165 -305 12175 -295
rect 12255 -295 12295 -290
rect 12255 -305 12265 -295
rect 12165 -315 12265 -305
rect 12285 -305 12295 -295
rect 12375 -295 12415 -290
rect 12375 -305 12385 -295
rect 12285 -315 12385 -305
rect 12405 -305 12415 -295
rect 12495 -295 12535 -290
rect 12495 -305 12505 -295
rect 12405 -315 12505 -305
rect 12525 -305 12535 -295
rect 12615 -295 12655 -290
rect 12615 -305 12625 -295
rect 12525 -315 12625 -305
rect 12645 -305 12655 -295
rect 12735 -295 12775 -290
rect 12735 -305 12745 -295
rect 12645 -315 12745 -305
rect 12765 -305 12775 -295
rect 12855 -295 12895 -290
rect 12855 -305 12865 -295
rect 12765 -315 12865 -305
rect 12885 -305 12895 -295
rect 12975 -295 13015 -290
rect 12975 -305 12985 -295
rect 12885 -315 12985 -305
rect 13005 -305 13015 -295
rect 13095 -295 13135 -290
rect 13095 -305 13105 -295
rect 13005 -315 13105 -305
rect 13125 -305 13135 -295
rect 13215 -295 13255 -290
rect 13215 -305 13225 -295
rect 13125 -315 13225 -305
rect 13245 -305 13255 -295
rect 13335 -295 13375 -290
rect 13335 -305 13345 -295
rect 13245 -315 13345 -305
rect 13365 -305 13375 -295
rect 13455 -295 13495 -290
rect 13455 -305 13465 -295
rect 13365 -315 13465 -305
rect 13485 -305 13495 -295
rect 13575 -295 13615 -290
rect 13575 -305 13585 -295
rect 13485 -315 13585 -305
rect 13605 -305 13615 -295
rect 13695 -295 13735 -290
rect 13695 -305 13705 -295
rect 13605 -315 13705 -305
rect 13725 -305 13735 -295
rect 13815 -295 13855 -290
rect 13815 -305 13825 -295
rect 13725 -315 13825 -305
rect 13845 -305 13855 -295
rect 13935 -295 13975 -290
rect 13935 -305 13945 -295
rect 13845 -315 13945 -305
rect 13965 -305 13975 -295
rect 14055 -295 14095 -290
rect 14055 -305 14065 -295
rect 13965 -315 14065 -305
rect 14085 -305 14095 -295
rect 14175 -295 14215 -290
rect 14175 -305 14185 -295
rect 14085 -315 14185 -305
rect 14205 -305 14215 -295
rect 14295 -295 14335 -290
rect 14295 -305 14305 -295
rect 14205 -315 14305 -305
rect 14325 -305 14335 -295
rect 14415 -295 14455 -290
rect 14415 -305 14425 -295
rect 14325 -315 14425 -305
rect 14445 -305 14455 -295
rect 14535 -295 14575 -290
rect 14535 -305 14545 -295
rect 14445 -315 14545 -305
rect 14565 -305 14575 -295
rect 14655 -295 14695 -290
rect 14655 -305 14665 -295
rect 14565 -315 14665 -305
rect 14685 -305 14695 -295
rect 14775 -295 14815 -290
rect 14775 -305 14785 -295
rect 14685 -315 14785 -305
rect 14805 -305 14815 -295
rect 14895 -295 14935 -290
rect 14895 -305 14905 -295
rect 14805 -315 14905 -305
rect 14925 -305 14935 -295
rect 15015 -295 15055 -290
rect 15015 -305 15025 -295
rect 14925 -315 15025 -305
rect 15045 -305 15055 -295
rect 15135 -295 15175 -290
rect 15135 -305 15145 -295
rect 15045 -315 15145 -305
rect 15165 -305 15175 -295
rect 15255 -295 15295 -290
rect 15255 -305 15265 -295
rect 15165 -315 15265 -305
rect 15285 -305 15295 -295
rect 15375 -295 15415 -290
rect 15375 -305 15385 -295
rect 15285 -315 15385 -305
rect 15405 -305 15415 -295
rect 15495 -295 15535 -290
rect 15495 -305 15505 -295
rect 15405 -315 15505 -305
rect 15525 -305 15535 -295
rect 15615 -295 15655 -290
rect 15615 -305 15625 -295
rect 15525 -315 15625 -305
rect 15645 -305 15655 -295
rect 15735 -295 15775 -290
rect 15735 -305 15745 -295
rect 15645 -315 15745 -305
rect 15765 -305 15775 -295
rect 15855 -295 15895 -290
rect 15855 -305 15865 -295
rect 15765 -315 15865 -305
rect 15885 -305 15895 -295
rect 15975 -295 16015 -290
rect 15975 -305 15985 -295
rect 15885 -315 15985 -305
rect 16005 -305 16015 -295
rect 16095 -295 16135 -290
rect 16095 -305 16105 -295
rect 16005 -315 16105 -305
rect 16125 -305 16135 -295
rect 16215 -295 16255 -290
rect 16215 -305 16225 -295
rect 16125 -315 16225 -305
rect 16245 -305 16255 -295
rect 16335 -295 16375 -290
rect 16335 -305 16345 -295
rect 16245 -315 16345 -305
rect 16365 -305 16375 -295
rect 16455 -295 16495 -290
rect 16455 -305 16465 -295
rect 16365 -315 16465 -305
rect 16485 -305 16495 -295
rect 16575 -295 16615 -290
rect 16575 -305 16585 -295
rect 16485 -315 16585 -305
rect 16605 -305 16615 -295
rect 16695 -295 16735 -290
rect 16695 -305 16705 -295
rect 16605 -315 16705 -305
rect 16725 -305 16735 -295
rect 16815 -295 16855 -290
rect 16815 -305 16825 -295
rect 16725 -315 16825 -305
rect 16845 -305 16855 -295
rect 16935 -295 16975 -290
rect 16935 -305 16945 -295
rect 16845 -315 16945 -305
rect 16965 -305 16975 -295
rect 17055 -295 17095 -290
rect 17055 -305 17065 -295
rect 16965 -315 17065 -305
rect 17085 -305 17095 -295
rect 17175 -295 17215 -290
rect 17175 -305 17185 -295
rect 17085 -315 17185 -305
rect 17205 -305 17215 -295
rect 17295 -295 17335 -290
rect 17295 -305 17305 -295
rect 17205 -315 17305 -305
rect 17325 -305 17335 -295
rect 17415 -295 17455 -290
rect 17415 -305 17425 -295
rect 17325 -315 17425 -305
rect 17445 -305 17455 -295
rect 17535 -295 17575 -290
rect 17535 -305 17545 -295
rect 17445 -315 17545 -305
rect 17565 -305 17575 -295
rect 17655 -295 17695 -290
rect 17655 -305 17665 -295
rect 17565 -315 17665 -305
rect 17685 -305 17695 -295
rect 17775 -295 17815 -290
rect 17775 -305 17785 -295
rect 17685 -315 17785 -305
rect 17805 -305 17815 -295
rect 17895 -295 17935 -290
rect 17895 -305 17905 -295
rect 17805 -315 17905 -305
rect 17925 -305 17935 -295
rect 18015 -295 18055 -290
rect 18015 -305 18025 -295
rect 17925 -315 18025 -305
rect 18045 -305 18055 -295
rect 18135 -295 18175 -290
rect 18135 -305 18145 -295
rect 18045 -315 18145 -305
rect 18165 -305 18175 -295
rect 18255 -295 18295 -290
rect 18255 -305 18265 -295
rect 18165 -315 18265 -305
rect 18285 -305 18295 -295
rect 18375 -295 18415 -290
rect 18375 -305 18385 -295
rect 18285 -315 18385 -305
rect 18405 -305 18415 -295
rect 18495 -295 18535 -290
rect 18495 -305 18505 -295
rect 18405 -315 18505 -305
rect 18525 -305 18535 -295
rect 18615 -295 18655 -290
rect 18615 -305 18625 -295
rect 18525 -315 18625 -305
rect 18645 -305 18655 -295
rect 18735 -295 18775 -290
rect 18735 -305 18745 -295
rect 18645 -315 18745 -305
rect 18765 -305 18775 -295
rect 18855 -295 18895 -290
rect 18855 -305 18865 -295
rect 18765 -315 18865 -305
rect 18885 -305 18895 -295
rect 18975 -295 19015 -290
rect 18975 -305 18985 -295
rect 18885 -315 18985 -305
rect 19005 -305 19015 -295
rect 19095 -295 19135 -290
rect 19095 -305 19105 -295
rect 19005 -315 19105 -305
rect 19125 -305 19135 -295
rect 19215 -295 19255 -290
rect 19215 -305 19225 -295
rect 19125 -315 19225 -305
rect 19245 -305 19255 -295
rect 19335 -295 19375 -290
rect 19335 -305 19345 -295
rect 19245 -315 19345 -305
rect 19365 -305 19375 -295
rect 19455 -295 19495 -290
rect 19455 -305 19465 -295
rect 19365 -315 19465 -305
rect 19485 -305 19495 -295
rect 19575 -295 19615 -290
rect 19575 -305 19585 -295
rect 19485 -315 19585 -305
rect 19605 -305 19615 -295
rect 19695 -295 19735 -290
rect 19695 -305 19705 -295
rect 19605 -315 19705 -305
rect 19725 -305 19735 -295
rect 19815 -295 19855 -290
rect 19815 -305 19825 -295
rect 19725 -315 19825 -305
rect 19845 -305 19855 -295
rect 19935 -295 19975 -290
rect 19935 -305 19945 -295
rect 19845 -315 19945 -305
rect 19965 -305 19975 -295
rect 20055 -295 20095 -290
rect 20055 -305 20065 -295
rect 19965 -315 20065 -305
rect 20085 -305 20095 -295
rect 20175 -295 20215 -290
rect 20175 -305 20185 -295
rect 20085 -315 20185 -305
rect 20205 -305 20215 -295
rect 20295 -295 20335 -290
rect 20295 -305 20305 -295
rect 20205 -315 20305 -305
rect 20325 -305 20335 -295
rect 20415 -295 20455 -290
rect 20415 -305 20425 -295
rect 20325 -315 20425 -305
rect 20445 -305 20455 -295
rect 20535 -295 20575 -290
rect 20535 -305 20545 -295
rect 20445 -315 20545 -305
rect 20565 -305 20575 -295
rect 20655 -295 20695 -290
rect 20655 -305 20665 -295
rect 20565 -315 20665 -305
rect 20685 -305 20695 -295
rect 20775 -295 20815 -290
rect 20775 -305 20785 -295
rect 20685 -315 20785 -305
rect 20805 -305 20815 -295
rect 20895 -295 20935 -290
rect 20895 -305 20905 -295
rect 20805 -315 20905 -305
rect 20925 -305 20935 -295
rect 21015 -295 21055 -290
rect 21015 -305 21025 -295
rect 20925 -315 21025 -305
rect 21045 -305 21055 -295
rect 21135 -295 21175 -290
rect 21135 -305 21145 -295
rect 21045 -315 21145 -305
rect 21165 -305 21175 -295
rect 21255 -295 21295 -290
rect 21255 -305 21265 -295
rect 21165 -315 21265 -305
rect 21285 -305 21295 -295
rect 21375 -295 21415 -290
rect 21375 -305 21385 -295
rect 21285 -315 21385 -305
rect 21405 -305 21415 -295
rect 21495 -295 21535 -290
rect 21495 -305 21505 -295
rect 21405 -315 21505 -305
rect 21525 -305 21535 -295
rect 21615 -295 21655 -290
rect 21615 -305 21625 -295
rect 21525 -315 21625 -305
rect 21645 -305 21655 -295
rect 21735 -295 21775 -290
rect 21735 -305 21745 -295
rect 21645 -315 21745 -305
rect 21765 -305 21775 -295
rect 21855 -295 21895 -290
rect 21855 -305 21865 -295
rect 21765 -315 21865 -305
rect 21885 -305 21895 -295
rect 21975 -295 22015 -290
rect 21975 -305 21985 -295
rect 21885 -315 21985 -305
rect 22005 -305 22015 -295
rect 22095 -295 22135 -290
rect 22095 -305 22105 -295
rect 22005 -315 22105 -305
rect 22125 -305 22135 -295
rect 22215 -295 22255 -290
rect 22215 -305 22225 -295
rect 22125 -315 22225 -305
rect 22245 -305 22255 -295
rect 22335 -295 22375 -290
rect 22335 -305 22345 -295
rect 22245 -315 22345 -305
rect 22365 -305 22375 -295
rect 22455 -295 22495 -290
rect 22455 -305 22465 -295
rect 22365 -315 22465 -305
rect 22485 -305 22495 -295
rect 22575 -295 22615 -290
rect 22575 -305 22585 -295
rect 22485 -315 22585 -305
rect 22605 -305 22615 -295
rect 22695 -295 22735 -290
rect 22695 -305 22705 -295
rect 22605 -315 22705 -305
rect 22725 -305 22735 -295
rect 22815 -295 22855 -290
rect 22815 -305 22825 -295
rect 22725 -315 22825 -305
rect 22845 -305 22855 -295
rect 22935 -295 22975 -290
rect 22935 -305 22945 -295
rect 22845 -315 22945 -305
rect 22965 -305 22975 -295
rect 23055 -295 23095 -290
rect 23055 -305 23065 -295
rect 22965 -315 23065 -305
rect 23085 -305 23095 -295
rect 23175 -295 23215 -290
rect 23175 -305 23185 -295
rect 23085 -315 23185 -305
rect 23205 -305 23215 -295
rect 23295 -295 23335 -290
rect 23295 -305 23305 -295
rect 23205 -315 23305 -305
rect 23325 -305 23335 -295
rect 23415 -295 23455 -290
rect 23415 -305 23425 -295
rect 23325 -315 23425 -305
rect 23445 -305 23455 -295
rect 23535 -295 23575 -290
rect 23535 -305 23545 -295
rect 23445 -315 23545 -305
rect 23565 -305 23575 -295
rect 23655 -295 23695 -290
rect 23655 -305 23665 -295
rect 23565 -315 23665 -305
rect 23685 -305 23695 -295
rect 23775 -295 23815 -290
rect 23775 -305 23785 -295
rect 23685 -315 23785 -305
rect 23805 -305 23815 -295
rect 23895 -295 23935 -290
rect 23895 -305 23905 -295
rect 23805 -315 23905 -305
rect 23925 -305 23935 -295
rect 24015 -295 24055 -290
rect 24015 -305 24025 -295
rect 23925 -315 24025 -305
rect 24045 -305 24055 -295
rect 24135 -295 24175 -290
rect 24135 -305 24145 -295
rect 24045 -315 24145 -305
rect 24165 -305 24175 -295
rect 24255 -295 24295 -290
rect 24255 -305 24265 -295
rect 24165 -315 24265 -305
rect 24285 -305 24295 -295
rect 24375 -295 24415 -290
rect 24375 -305 24385 -295
rect 24285 -315 24385 -305
rect 24405 -305 24415 -295
rect 24495 -295 24535 -290
rect 24495 -305 24505 -295
rect 24405 -315 24505 -305
rect 24525 -305 24535 -295
rect 24615 -295 24655 -290
rect 24615 -305 24625 -295
rect 24525 -315 24625 -305
rect 24645 -305 24655 -295
rect 24735 -295 24775 -290
rect 24735 -305 24745 -295
rect 24645 -315 24745 -305
rect 24765 -305 24775 -295
rect 24855 -295 24895 -290
rect 24855 -305 24865 -295
rect 24765 -315 24865 -305
rect 24885 -305 24895 -295
rect 24975 -295 25015 -290
rect 24975 -305 24985 -295
rect 24885 -315 24985 -305
rect 25005 -305 25015 -295
rect 25095 -295 25135 -290
rect 25095 -305 25105 -295
rect 25005 -315 25105 -305
rect 25125 -305 25135 -295
rect 25215 -295 25255 -290
rect 25215 -305 25225 -295
rect 25125 -315 25225 -305
rect 25245 -305 25255 -295
rect 25335 -295 25375 -290
rect 25335 -305 25345 -295
rect 25245 -315 25345 -305
rect 25365 -305 25375 -295
rect 25455 -295 25495 -290
rect 25455 -305 25465 -295
rect 25365 -315 25465 -305
rect 25485 -305 25495 -295
rect 25575 -295 25615 -290
rect 25575 -305 25585 -295
rect 25485 -315 25585 -305
rect 25605 -305 25615 -295
rect 25695 -295 25735 -290
rect 25695 -305 25705 -295
rect 25605 -315 25705 -305
rect 25725 -305 25735 -295
rect 25815 -295 25855 -290
rect 25815 -305 25825 -295
rect 25725 -315 25825 -305
rect 25845 -305 25855 -295
rect 25935 -295 25975 -290
rect 25935 -305 25945 -295
rect 25845 -315 25945 -305
rect 25965 -305 25975 -295
rect 26055 -295 26095 -290
rect 26055 -305 26065 -295
rect 25965 -315 26065 -305
rect 26085 -305 26095 -295
rect 26175 -295 26215 -290
rect 26175 -305 26185 -295
rect 26085 -315 26185 -305
rect 26205 -305 26215 -295
rect 26295 -295 26335 -290
rect 26295 -305 26305 -295
rect 26205 -315 26305 -305
rect 26325 -305 26335 -295
rect 26415 -295 26455 -290
rect 26415 -305 26425 -295
rect 26325 -315 26425 -305
rect 26445 -305 26455 -295
rect 26535 -295 26575 -290
rect 26535 -305 26545 -295
rect 26445 -315 26545 -305
rect 26565 -305 26575 -295
rect 26655 -295 26695 -290
rect 26655 -305 26665 -295
rect 26565 -315 26665 -305
rect 26685 -305 26695 -295
rect 26775 -295 26815 -290
rect 26775 -305 26785 -295
rect 26685 -315 26785 -305
rect 26805 -305 26815 -295
rect 26895 -295 26935 -290
rect 26895 -305 26905 -295
rect 26805 -315 26905 -305
rect 26925 -305 26935 -295
rect 27015 -295 27055 -290
rect 27015 -305 27025 -295
rect 26925 -315 27025 -305
rect 27045 -305 27055 -295
rect 27135 -295 27175 -290
rect 27135 -305 27145 -295
rect 27045 -315 27145 -305
rect 27165 -305 27175 -295
rect 27255 -295 27295 -290
rect 27255 -305 27265 -295
rect 27165 -315 27265 -305
rect 27285 -305 27295 -295
rect 27375 -295 27415 -290
rect 27375 -305 27385 -295
rect 27285 -315 27385 -305
rect 27405 -305 27415 -295
rect 27495 -295 27535 -290
rect 27495 -305 27505 -295
rect 27405 -315 27505 -305
rect 27525 -305 27535 -295
rect 27615 -295 27655 -290
rect 27615 -305 27625 -295
rect 27525 -315 27625 -305
rect 27645 -305 27655 -295
rect 27735 -295 27775 -290
rect 27735 -305 27745 -295
rect 27645 -315 27745 -305
rect 27765 -305 27775 -295
rect 27855 -295 27895 -290
rect 27855 -305 27865 -295
rect 27765 -315 27865 -305
rect 27885 -305 27895 -295
rect 27975 -295 28015 -290
rect 27975 -305 27985 -295
rect 27885 -315 27985 -305
rect 28005 -305 28015 -295
rect 28095 -295 28135 -290
rect 28095 -305 28105 -295
rect 28005 -315 28105 -305
rect 28125 -305 28135 -295
rect 28215 -295 28255 -290
rect 28215 -305 28225 -295
rect 28125 -315 28225 -305
rect 28245 -305 28255 -295
rect 28335 -295 28375 -290
rect 28335 -305 28345 -295
rect 28245 -315 28345 -305
rect 28365 -305 28375 -295
rect 28455 -295 28495 -290
rect 28455 -305 28465 -295
rect 28365 -315 28465 -305
rect 28485 -305 28495 -295
rect 28575 -295 28615 -290
rect 28575 -305 28585 -295
rect 28485 -315 28585 -305
rect 28605 -305 28615 -295
rect 28695 -295 28735 -290
rect 28695 -305 28705 -295
rect 28605 -315 28705 -305
rect 28725 -305 28735 -295
rect 28815 -295 28855 -290
rect 28815 -305 28825 -295
rect 28725 -315 28825 -305
rect 28845 -305 28855 -295
rect 28935 -295 28975 -290
rect 28935 -305 28945 -295
rect 28845 -315 28945 -305
rect 28965 -305 28975 -295
rect 29055 -295 29095 -290
rect 29055 -305 29065 -295
rect 28965 -315 29065 -305
rect 29085 -305 29095 -295
rect 29175 -295 29215 -290
rect 29175 -305 29185 -295
rect 29085 -315 29185 -305
rect 29205 -305 29215 -295
rect 29295 -295 29335 -290
rect 29295 -305 29305 -295
rect 29205 -315 29305 -305
rect 29325 -305 29335 -295
rect 29415 -295 29455 -290
rect 29415 -305 29425 -295
rect 29325 -315 29425 -305
rect 29445 -305 29455 -295
rect 29535 -295 29575 -290
rect 29535 -305 29545 -295
rect 29445 -315 29545 -305
rect 29565 -305 29575 -295
rect 29655 -295 29695 -290
rect 29655 -305 29665 -295
rect 29565 -315 29665 -305
rect 29685 -305 29695 -295
rect 29775 -295 29815 -290
rect 29775 -305 29785 -295
rect 29685 -315 29785 -305
rect 29805 -305 29815 -295
rect 29895 -295 29935 -290
rect 29895 -305 29905 -295
rect 29805 -315 29905 -305
rect 29925 -305 29935 -295
rect 30015 -295 30055 -290
rect 30015 -305 30025 -295
rect 29925 -315 30025 -305
rect 30045 -305 30055 -295
rect 30135 -295 30175 -290
rect 30135 -305 30145 -295
rect 30045 -315 30145 -305
rect 30165 -305 30175 -295
rect 30255 -295 30295 -290
rect 30255 -305 30265 -295
rect 30165 -315 30265 -305
rect 30285 -305 30295 -295
rect 30375 -295 30415 -290
rect 30375 -305 30385 -295
rect 30285 -315 30385 -305
rect 30405 -305 30415 -295
rect 30495 -295 30535 -290
rect 30495 -305 30505 -295
rect 30405 -315 30505 -305
rect 30525 -305 30535 -295
rect 30615 -295 30655 -290
rect 30615 -305 30625 -295
rect 30525 -315 30625 -305
rect 30645 -315 30655 -295
rect 15 -320 30655 -315
rect 15 -325 55 -320
rect 135 -325 175 -320
rect 255 -325 295 -320
rect 375 -325 415 -320
rect 495 -325 535 -320
rect 615 -325 655 -320
rect 735 -325 775 -320
rect 855 -325 895 -320
rect 975 -325 1015 -320
rect 1095 -325 1135 -320
rect 1215 -325 1255 -320
rect 1335 -325 1375 -320
rect 1455 -325 1495 -320
rect 1575 -325 1615 -320
rect 1695 -325 1735 -320
rect 1815 -325 1855 -320
rect 1935 -325 1975 -320
rect 2055 -325 2095 -320
rect 2175 -325 2215 -320
rect 2295 -325 2335 -320
rect 2415 -325 2455 -320
rect 2535 -325 2575 -320
rect 2655 -325 2695 -320
rect 2775 -325 2815 -320
rect 2895 -325 2935 -320
rect 3015 -325 3055 -320
rect 3135 -325 3175 -320
rect 3255 -325 3295 -320
rect 3375 -325 3415 -320
rect 3495 -325 3535 -320
rect 3615 -325 3655 -320
rect 3735 -325 3775 -320
rect 3855 -325 3895 -320
rect 3975 -325 4015 -320
rect 4095 -325 4135 -320
rect 4215 -325 4255 -320
rect 4335 -325 4375 -320
rect 4455 -325 4495 -320
rect 4575 -325 4615 -320
rect 4695 -325 4735 -320
rect 4815 -325 4855 -320
rect 4935 -325 4975 -320
rect 5055 -325 5095 -320
rect 5175 -325 5215 -320
rect 5295 -325 5335 -320
rect 5415 -325 5455 -320
rect 5535 -325 5575 -320
rect 5655 -325 5695 -320
rect 5775 -325 5815 -320
rect 5895 -325 5935 -320
rect 6015 -325 6055 -320
rect 6135 -325 6175 -320
rect 6255 -325 6295 -320
rect 6375 -325 6415 -320
rect 6495 -325 6535 -320
rect 6615 -325 6655 -320
rect 6735 -325 6775 -320
rect 6855 -325 6895 -320
rect 6975 -325 7015 -320
rect 7095 -325 7135 -320
rect 7215 -325 7255 -320
rect 7335 -325 7375 -320
rect 7455 -325 7495 -320
rect 7575 -325 7615 -320
rect 7695 -325 7735 -320
rect 7815 -325 7855 -320
rect 7935 -325 7975 -320
rect 8055 -325 8095 -320
rect 8175 -325 8215 -320
rect 8295 -325 8335 -320
rect 8415 -325 8455 -320
rect 8535 -325 8575 -320
rect 8655 -325 8695 -320
rect 8775 -325 8815 -320
rect 8895 -325 8935 -320
rect 9015 -325 9055 -320
rect 9135 -325 9175 -320
rect 9255 -325 9295 -320
rect 9375 -325 9415 -320
rect 9495 -325 9535 -320
rect 9615 -325 9655 -320
rect 9735 -325 9775 -320
rect 9855 -325 9895 -320
rect 9975 -325 10015 -320
rect 10095 -325 10135 -320
rect 10215 -325 10255 -320
rect 10335 -325 10375 -320
rect 10455 -325 10495 -320
rect 10575 -325 10615 -320
rect 10695 -325 10735 -320
rect 10815 -325 10855 -320
rect 10935 -325 10975 -320
rect 11055 -325 11095 -320
rect 11175 -325 11215 -320
rect 11295 -325 11335 -320
rect 11415 -325 11455 -320
rect 11535 -325 11575 -320
rect 11655 -325 11695 -320
rect 11775 -325 11815 -320
rect 11895 -325 11935 -320
rect 12015 -325 12055 -320
rect 12135 -325 12175 -320
rect 12255 -325 12295 -320
rect 12375 -325 12415 -320
rect 12495 -325 12535 -320
rect 12615 -325 12655 -320
rect 12735 -325 12775 -320
rect 12855 -325 12895 -320
rect 12975 -325 13015 -320
rect 13095 -325 13135 -320
rect 13215 -325 13255 -320
rect 13335 -325 13375 -320
rect 13455 -325 13495 -320
rect 13575 -325 13615 -320
rect 13695 -325 13735 -320
rect 13815 -325 13855 -320
rect 13935 -325 13975 -320
rect 14055 -325 14095 -320
rect 14175 -325 14215 -320
rect 14295 -325 14335 -320
rect 14415 -325 14455 -320
rect 14535 -325 14575 -320
rect 14655 -325 14695 -320
rect 14775 -325 14815 -320
rect 14895 -325 14935 -320
rect 15015 -325 15055 -320
rect 15135 -325 15175 -320
rect 15255 -325 15295 -320
rect 15375 -325 15415 -320
rect 15495 -325 15535 -320
rect 15615 -325 15655 -320
rect 15735 -325 15775 -320
rect 15855 -325 15895 -320
rect 15975 -325 16015 -320
rect 16095 -325 16135 -320
rect 16215 -325 16255 -320
rect 16335 -325 16375 -320
rect 16455 -325 16495 -320
rect 16575 -325 16615 -320
rect 16695 -325 16735 -320
rect 16815 -325 16855 -320
rect 16935 -325 16975 -320
rect 17055 -325 17095 -320
rect 17175 -325 17215 -320
rect 17295 -325 17335 -320
rect 17415 -325 17455 -320
rect 17535 -325 17575 -320
rect 17655 -325 17695 -320
rect 17775 -325 17815 -320
rect 17895 -325 17935 -320
rect 18015 -325 18055 -320
rect 18135 -325 18175 -320
rect 18255 -325 18295 -320
rect 18375 -325 18415 -320
rect 18495 -325 18535 -320
rect 18615 -325 18655 -320
rect 18735 -325 18775 -320
rect 18855 -325 18895 -320
rect 18975 -325 19015 -320
rect 19095 -325 19135 -320
rect 19215 -325 19255 -320
rect 19335 -325 19375 -320
rect 19455 -325 19495 -320
rect 19575 -325 19615 -320
rect 19695 -325 19735 -320
rect 19815 -325 19855 -320
rect 19935 -325 19975 -320
rect 20055 -325 20095 -320
rect 20175 -325 20215 -320
rect 20295 -325 20335 -320
rect 20415 -325 20455 -320
rect 20535 -325 20575 -320
rect 20655 -325 20695 -320
rect 20775 -325 20815 -320
rect 20895 -325 20935 -320
rect 21015 -325 21055 -320
rect 21135 -325 21175 -320
rect 21255 -325 21295 -320
rect 21375 -325 21415 -320
rect 21495 -325 21535 -320
rect 21615 -325 21655 -320
rect 21735 -325 21775 -320
rect 21855 -325 21895 -320
rect 21975 -325 22015 -320
rect 22095 -325 22135 -320
rect 22215 -325 22255 -320
rect 22335 -325 22375 -320
rect 22455 -325 22495 -320
rect 22575 -325 22615 -320
rect 22695 -325 22735 -320
rect 22815 -325 22855 -320
rect 22935 -325 22975 -320
rect 23055 -325 23095 -320
rect 23175 -325 23215 -320
rect 23295 -325 23335 -320
rect 23415 -325 23455 -320
rect 23535 -325 23575 -320
rect 23655 -325 23695 -320
rect 23775 -325 23815 -320
rect 23895 -325 23935 -320
rect 24015 -325 24055 -320
rect 24135 -325 24175 -320
rect 24255 -325 24295 -320
rect 24375 -325 24415 -320
rect 24495 -325 24535 -320
rect 24615 -325 24655 -320
rect 24735 -325 24775 -320
rect 24855 -325 24895 -320
rect 24975 -325 25015 -320
rect 25095 -325 25135 -320
rect 25215 -325 25255 -320
rect 25335 -325 25375 -320
rect 25455 -325 25495 -320
rect 25575 -325 25615 -320
rect 25695 -325 25735 -320
rect 25815 -325 25855 -320
rect 25935 -325 25975 -320
rect 26055 -325 26095 -320
rect 26175 -325 26215 -320
rect 26295 -325 26335 -320
rect 26415 -325 26455 -320
rect 26535 -325 26575 -320
rect 26655 -325 26695 -320
rect 26775 -325 26815 -320
rect 26895 -325 26935 -320
rect 27015 -325 27055 -320
rect 27135 -325 27175 -320
rect 27255 -325 27295 -320
rect 27375 -325 27415 -320
rect 27495 -325 27535 -320
rect 27615 -325 27655 -320
rect 27735 -325 27775 -320
rect 27855 -325 27895 -320
rect 27975 -325 28015 -320
rect 28095 -325 28135 -320
rect 28215 -325 28255 -320
rect 28335 -325 28375 -320
rect 28455 -325 28495 -320
rect 28575 -325 28615 -320
rect 28695 -325 28735 -320
rect 28815 -325 28855 -320
rect 28935 -325 28975 -320
rect 29055 -325 29095 -320
rect 29175 -325 29215 -320
rect 29295 -325 29335 -320
rect 29415 -325 29455 -320
rect 29535 -325 29575 -320
rect 29655 -325 29695 -320
rect 29775 -325 29815 -320
rect 29895 -325 29935 -320
rect 30015 -325 30055 -320
rect 30135 -325 30175 -320
rect 30255 -325 30295 -320
rect 30375 -325 30415 -320
rect 30495 -325 30535 -320
rect 30615 -325 30655 -320
rect -40 -420 0 -410
rect -40 -440 -30 -420
rect -10 -425 0 -420
rect 75 -420 115 -410
rect 200 -415 240 -410
rect 75 -425 85 -420
rect -10 -440 85 -425
rect 105 -425 115 -420
rect 195 -420 240 -415
rect 195 -425 210 -420
rect 105 -440 210 -425
rect 230 -425 240 -420
rect 315 -420 355 -410
rect 440 -415 480 -410
rect 315 -425 325 -420
rect 230 -440 325 -425
rect 345 -425 355 -420
rect 435 -420 480 -415
rect 435 -425 450 -420
rect 345 -440 450 -425
rect 470 -425 480 -420
rect 555 -420 595 -410
rect 680 -415 720 -410
rect 555 -425 565 -420
rect 470 -440 565 -425
rect 585 -425 595 -420
rect 675 -420 720 -415
rect 675 -425 690 -420
rect 585 -440 690 -425
rect 710 -425 720 -420
rect 795 -420 835 -410
rect 920 -415 960 -410
rect 795 -425 805 -420
rect 710 -440 805 -425
rect 825 -425 835 -420
rect 915 -420 960 -415
rect 915 -425 930 -420
rect 825 -440 930 -425
rect 950 -425 960 -420
rect 1035 -420 1075 -410
rect 1160 -415 1200 -410
rect 1035 -425 1045 -420
rect 950 -440 1045 -425
rect 1065 -425 1075 -420
rect 1155 -420 1200 -415
rect 1155 -425 1170 -420
rect 1065 -440 1170 -425
rect 1190 -425 1200 -420
rect 1275 -420 1315 -410
rect 1400 -415 1440 -410
rect 1275 -425 1285 -420
rect 1190 -440 1285 -425
rect 1305 -425 1315 -420
rect 1395 -420 1440 -415
rect 1395 -425 1410 -420
rect 1305 -440 1410 -425
rect 1430 -425 1440 -420
rect 1515 -420 1555 -410
rect 1640 -415 1680 -410
rect 1515 -425 1525 -420
rect 1430 -440 1525 -425
rect 1545 -425 1555 -420
rect 1635 -420 1680 -415
rect 1635 -425 1650 -420
rect 1545 -440 1650 -425
rect 1670 -425 1680 -420
rect 1755 -420 1795 -410
rect 1880 -415 1920 -410
rect 1755 -425 1765 -420
rect 1670 -440 1765 -425
rect 1785 -425 1795 -420
rect 1875 -420 1920 -415
rect 1875 -425 1890 -420
rect 1785 -440 1890 -425
rect 1910 -425 1920 -420
rect 1995 -420 2035 -410
rect 2120 -415 2160 -410
rect 1995 -425 2005 -420
rect 1910 -440 2005 -425
rect 2025 -425 2035 -420
rect 2115 -420 2160 -415
rect 2115 -425 2130 -420
rect 2025 -440 2130 -425
rect 2150 -425 2160 -420
rect 2235 -420 2275 -410
rect 2360 -415 2400 -410
rect 2235 -425 2245 -420
rect 2150 -440 2245 -425
rect 2265 -425 2275 -420
rect 2355 -420 2400 -415
rect 2355 -425 2370 -420
rect 2265 -440 2370 -425
rect 2390 -425 2400 -420
rect 2475 -420 2515 -410
rect 2600 -415 2640 -410
rect 2475 -425 2485 -420
rect 2390 -440 2485 -425
rect 2505 -425 2515 -420
rect 2595 -420 2640 -415
rect 2595 -425 2610 -420
rect 2505 -440 2610 -425
rect 2630 -425 2640 -420
rect 2715 -420 2755 -410
rect 2840 -415 2880 -410
rect 2715 -425 2725 -420
rect 2630 -440 2725 -425
rect 2745 -425 2755 -420
rect 2835 -420 2880 -415
rect 2835 -425 2850 -420
rect 2745 -440 2850 -425
rect 2870 -425 2880 -420
rect 2955 -420 2995 -410
rect 3080 -415 3120 -410
rect 2955 -425 2965 -420
rect 2870 -440 2965 -425
rect 2985 -425 2995 -420
rect 3075 -420 3120 -415
rect 3075 -425 3090 -420
rect 2985 -440 3090 -425
rect 3110 -425 3120 -420
rect 3195 -420 3235 -410
rect 3320 -415 3360 -410
rect 3195 -425 3205 -420
rect 3110 -440 3205 -425
rect 3225 -425 3235 -420
rect 3315 -420 3360 -415
rect 3315 -425 3330 -420
rect 3225 -440 3330 -425
rect 3350 -425 3360 -420
rect 3435 -420 3475 -410
rect 3560 -415 3600 -410
rect 3435 -425 3445 -420
rect 3350 -440 3445 -425
rect 3465 -425 3475 -420
rect 3555 -420 3600 -415
rect 3555 -425 3570 -420
rect 3465 -440 3570 -425
rect 3590 -425 3600 -420
rect 3675 -420 3715 -410
rect 3800 -415 3840 -410
rect 3675 -425 3685 -420
rect 3590 -440 3685 -425
rect 3705 -425 3715 -420
rect 3795 -420 3840 -415
rect 3795 -425 3810 -420
rect 3705 -440 3810 -425
rect 3830 -425 3840 -420
rect 3915 -420 3955 -410
rect 4040 -415 4080 -410
rect 3915 -425 3925 -420
rect 3830 -440 3925 -425
rect 3945 -425 3955 -420
rect 4035 -420 4080 -415
rect 4035 -425 4050 -420
rect 3945 -440 4050 -425
rect 4070 -425 4080 -420
rect 4155 -420 4195 -410
rect 4280 -415 4320 -410
rect 4155 -425 4165 -420
rect 4070 -440 4165 -425
rect 4185 -425 4195 -420
rect 4275 -420 4320 -415
rect 4275 -425 4290 -420
rect 4185 -440 4290 -425
rect 4310 -425 4320 -420
rect 4395 -420 4435 -410
rect 4520 -415 4560 -410
rect 4395 -425 4405 -420
rect 4310 -440 4405 -425
rect 4425 -425 4435 -420
rect 4515 -420 4560 -415
rect 4515 -425 4530 -420
rect 4425 -440 4530 -425
rect 4550 -425 4560 -420
rect 4635 -420 4675 -410
rect 4760 -415 4800 -410
rect 4635 -425 4645 -420
rect 4550 -440 4645 -425
rect 4665 -425 4675 -420
rect 4755 -420 4800 -415
rect 4755 -425 4770 -420
rect 4665 -440 4770 -425
rect 4790 -425 4800 -420
rect 4875 -420 4915 -410
rect 5000 -415 5040 -410
rect 4875 -425 4885 -420
rect 4790 -440 4885 -425
rect 4905 -425 4915 -420
rect 4995 -420 5040 -415
rect 4995 -425 5010 -420
rect 4905 -440 5010 -425
rect 5030 -425 5040 -420
rect 5115 -420 5155 -410
rect 5240 -415 5280 -410
rect 5115 -425 5125 -420
rect 5030 -440 5125 -425
rect 5145 -425 5155 -420
rect 5235 -420 5280 -415
rect 5235 -425 5250 -420
rect 5145 -440 5250 -425
rect 5270 -425 5280 -420
rect 5355 -420 5395 -410
rect 5480 -415 5520 -410
rect 5355 -425 5365 -420
rect 5270 -440 5365 -425
rect 5385 -425 5395 -420
rect 5475 -420 5520 -415
rect 5475 -425 5490 -420
rect 5385 -440 5490 -425
rect 5510 -425 5520 -420
rect 5595 -420 5635 -410
rect 5720 -415 5760 -410
rect 5595 -425 5605 -420
rect 5510 -440 5605 -425
rect 5625 -425 5635 -420
rect 5715 -420 5760 -415
rect 5715 -425 5730 -420
rect 5625 -440 5730 -425
rect 5750 -425 5760 -420
rect 5835 -420 5875 -410
rect 5960 -415 6000 -410
rect 5835 -425 5845 -420
rect 5750 -440 5845 -425
rect 5865 -425 5875 -420
rect 5955 -420 6000 -415
rect 5955 -425 5970 -420
rect 5865 -440 5970 -425
rect 5990 -425 6000 -420
rect 6075 -420 6115 -410
rect 6200 -415 6240 -410
rect 6075 -425 6085 -420
rect 5990 -440 6085 -425
rect 6105 -425 6115 -420
rect 6195 -420 6240 -415
rect 6195 -425 6210 -420
rect 6105 -440 6210 -425
rect 6230 -425 6240 -420
rect 6315 -420 6355 -410
rect 6440 -415 6480 -410
rect 6315 -425 6325 -420
rect 6230 -440 6325 -425
rect 6345 -425 6355 -420
rect 6435 -420 6480 -415
rect 6435 -425 6450 -420
rect 6345 -440 6450 -425
rect 6470 -425 6480 -420
rect 6555 -420 6595 -410
rect 6680 -415 6720 -410
rect 6555 -425 6565 -420
rect 6470 -440 6565 -425
rect 6585 -425 6595 -420
rect 6675 -420 6720 -415
rect 6675 -425 6690 -420
rect 6585 -440 6690 -425
rect 6710 -425 6720 -420
rect 6795 -420 6835 -410
rect 6920 -415 6960 -410
rect 6795 -425 6805 -420
rect 6710 -440 6805 -425
rect 6825 -425 6835 -420
rect 6915 -420 6960 -415
rect 6915 -425 6930 -420
rect 6825 -440 6930 -425
rect 6950 -425 6960 -420
rect 7035 -420 7075 -410
rect 7160 -415 7200 -410
rect 7035 -425 7045 -420
rect 6950 -440 7045 -425
rect 7065 -425 7075 -420
rect 7155 -420 7200 -415
rect 7155 -425 7170 -420
rect 7065 -440 7170 -425
rect 7190 -425 7200 -420
rect 7275 -420 7315 -410
rect 7400 -415 7440 -410
rect 7275 -425 7285 -420
rect 7190 -440 7285 -425
rect 7305 -425 7315 -420
rect 7395 -420 7440 -415
rect 7395 -425 7410 -420
rect 7305 -440 7410 -425
rect 7430 -425 7440 -420
rect 7515 -420 7555 -410
rect 7640 -415 7680 -410
rect 7515 -425 7525 -420
rect 7430 -440 7525 -425
rect 7545 -425 7555 -420
rect 7635 -420 7680 -415
rect 7635 -425 7650 -420
rect 7545 -440 7650 -425
rect 7670 -425 7680 -420
rect 7755 -420 7795 -410
rect 7880 -415 7920 -410
rect 7755 -425 7765 -420
rect 7670 -440 7765 -425
rect 7785 -425 7795 -420
rect 7875 -420 7920 -415
rect 7875 -425 7890 -420
rect 7785 -440 7890 -425
rect 7910 -425 7920 -420
rect 7995 -420 8035 -410
rect 8120 -415 8160 -410
rect 7995 -425 8005 -420
rect 7910 -440 8005 -425
rect 8025 -425 8035 -420
rect 8115 -420 8160 -415
rect 8115 -425 8130 -420
rect 8025 -440 8130 -425
rect 8150 -425 8160 -420
rect 8235 -420 8275 -410
rect 8360 -415 8400 -410
rect 8235 -425 8245 -420
rect 8150 -440 8245 -425
rect 8265 -425 8275 -420
rect 8355 -420 8400 -415
rect 8355 -425 8370 -420
rect 8265 -440 8370 -425
rect 8390 -425 8400 -420
rect 8475 -420 8515 -410
rect 8600 -415 8640 -410
rect 8475 -425 8485 -420
rect 8390 -440 8485 -425
rect 8505 -425 8515 -420
rect 8595 -420 8640 -415
rect 8595 -425 8610 -420
rect 8505 -440 8610 -425
rect 8630 -425 8640 -420
rect 8715 -420 8755 -410
rect 8840 -415 8880 -410
rect 8715 -425 8725 -420
rect 8630 -440 8725 -425
rect 8745 -425 8755 -420
rect 8835 -420 8880 -415
rect 8835 -425 8850 -420
rect 8745 -440 8850 -425
rect 8870 -425 8880 -420
rect 8955 -420 8995 -410
rect 9080 -415 9120 -410
rect 8955 -425 8965 -420
rect 8870 -440 8965 -425
rect 8985 -425 8995 -420
rect 9075 -420 9120 -415
rect 9075 -425 9090 -420
rect 8985 -440 9090 -425
rect 9110 -425 9120 -420
rect 9195 -420 9235 -410
rect 9320 -415 9360 -410
rect 9195 -425 9205 -420
rect 9110 -440 9205 -425
rect 9225 -425 9235 -420
rect 9315 -420 9360 -415
rect 9315 -425 9330 -420
rect 9225 -440 9330 -425
rect 9350 -425 9360 -420
rect 9435 -420 9475 -410
rect 9560 -415 9600 -410
rect 9435 -425 9445 -420
rect 9350 -440 9445 -425
rect 9465 -425 9475 -420
rect 9555 -420 9600 -415
rect 9555 -425 9570 -420
rect 9465 -440 9570 -425
rect 9590 -425 9600 -420
rect 9675 -420 9715 -410
rect 9800 -415 9840 -410
rect 9675 -425 9685 -420
rect 9590 -440 9685 -425
rect 9705 -425 9715 -420
rect 9795 -420 9840 -415
rect 9795 -425 9810 -420
rect 9705 -440 9810 -425
rect 9830 -425 9840 -420
rect 9915 -420 9955 -410
rect 10040 -415 10080 -410
rect 9915 -425 9925 -420
rect 9830 -440 9925 -425
rect 9945 -425 9955 -420
rect 10035 -420 10080 -415
rect 10035 -425 10050 -420
rect 9945 -440 10050 -425
rect 10070 -425 10080 -420
rect 10155 -420 10195 -410
rect 10280 -415 10320 -410
rect 10155 -425 10165 -420
rect 10070 -440 10165 -425
rect 10185 -425 10195 -420
rect 10275 -420 10320 -415
rect 10275 -425 10290 -420
rect 10185 -440 10290 -425
rect 10310 -425 10320 -420
rect 10395 -420 10435 -410
rect 10520 -415 10560 -410
rect 10395 -425 10405 -420
rect 10310 -440 10405 -425
rect 10425 -425 10435 -420
rect 10515 -420 10560 -415
rect 10515 -425 10530 -420
rect 10425 -440 10530 -425
rect 10550 -425 10560 -420
rect 10635 -420 10675 -410
rect 10760 -415 10800 -410
rect 10635 -425 10645 -420
rect 10550 -440 10645 -425
rect 10665 -425 10675 -420
rect 10755 -420 10800 -415
rect 10755 -425 10770 -420
rect 10665 -440 10770 -425
rect 10790 -425 10800 -420
rect 10875 -420 10915 -410
rect 11000 -415 11040 -410
rect 10875 -425 10885 -420
rect 10790 -440 10885 -425
rect 10905 -425 10915 -420
rect 10995 -420 11040 -415
rect 10995 -425 11010 -420
rect 10905 -440 11010 -425
rect 11030 -425 11040 -420
rect 11115 -420 11155 -410
rect 11240 -415 11280 -410
rect 11115 -425 11125 -420
rect 11030 -440 11125 -425
rect 11145 -425 11155 -420
rect 11235 -420 11280 -415
rect 11235 -425 11250 -420
rect 11145 -440 11250 -425
rect 11270 -425 11280 -420
rect 11355 -420 11395 -410
rect 11480 -415 11520 -410
rect 11355 -425 11365 -420
rect 11270 -440 11365 -425
rect 11385 -425 11395 -420
rect 11475 -420 11520 -415
rect 11475 -425 11490 -420
rect 11385 -440 11490 -425
rect 11510 -425 11520 -420
rect 11595 -420 11635 -410
rect 11720 -415 11760 -410
rect 11595 -425 11605 -420
rect 11510 -440 11605 -425
rect 11625 -425 11635 -420
rect 11715 -420 11760 -415
rect 11715 -425 11730 -420
rect 11625 -440 11730 -425
rect 11750 -425 11760 -420
rect 11835 -420 11875 -410
rect 11960 -415 12000 -410
rect 11835 -425 11845 -420
rect 11750 -440 11845 -425
rect 11865 -425 11875 -420
rect 11955 -420 12000 -415
rect 11955 -425 11970 -420
rect 11865 -440 11970 -425
rect 11990 -425 12000 -420
rect 12075 -420 12115 -410
rect 12200 -415 12240 -410
rect 12075 -425 12085 -420
rect 11990 -440 12085 -425
rect 12105 -425 12115 -420
rect 12195 -420 12240 -415
rect 12195 -425 12210 -420
rect 12105 -440 12210 -425
rect 12230 -425 12240 -420
rect 12315 -420 12355 -410
rect 12440 -415 12480 -410
rect 12315 -425 12325 -420
rect 12230 -440 12325 -425
rect 12345 -425 12355 -420
rect 12435 -420 12480 -415
rect 12435 -425 12450 -420
rect 12345 -440 12450 -425
rect 12470 -425 12480 -420
rect 12555 -420 12595 -410
rect 12680 -415 12720 -410
rect 12555 -425 12565 -420
rect 12470 -440 12565 -425
rect 12585 -425 12595 -420
rect 12675 -420 12720 -415
rect 12675 -425 12690 -420
rect 12585 -440 12690 -425
rect 12710 -425 12720 -420
rect 12795 -420 12835 -410
rect 12920 -415 12960 -410
rect 12795 -425 12805 -420
rect 12710 -440 12805 -425
rect 12825 -425 12835 -420
rect 12915 -420 12960 -415
rect 12915 -425 12930 -420
rect 12825 -440 12930 -425
rect 12950 -425 12960 -420
rect 13035 -420 13075 -410
rect 13160 -415 13200 -410
rect 13035 -425 13045 -420
rect 12950 -440 13045 -425
rect 13065 -425 13075 -420
rect 13155 -420 13200 -415
rect 13155 -425 13170 -420
rect 13065 -440 13170 -425
rect 13190 -425 13200 -420
rect 13275 -420 13315 -410
rect 13400 -415 13440 -410
rect 13275 -425 13285 -420
rect 13190 -440 13285 -425
rect 13305 -425 13315 -420
rect 13395 -420 13440 -415
rect 13395 -425 13410 -420
rect 13305 -440 13410 -425
rect 13430 -425 13440 -420
rect 13515 -420 13555 -410
rect 13640 -415 13680 -410
rect 13515 -425 13525 -420
rect 13430 -440 13525 -425
rect 13545 -425 13555 -420
rect 13635 -420 13680 -415
rect 13635 -425 13650 -420
rect 13545 -440 13650 -425
rect 13670 -425 13680 -420
rect 13755 -420 13795 -410
rect 13880 -415 13920 -410
rect 13755 -425 13765 -420
rect 13670 -440 13765 -425
rect 13785 -425 13795 -420
rect 13875 -420 13920 -415
rect 13875 -425 13890 -420
rect 13785 -440 13890 -425
rect 13910 -425 13920 -420
rect 13995 -420 14035 -410
rect 14120 -415 14160 -410
rect 13995 -425 14005 -420
rect 13910 -440 14005 -425
rect 14025 -425 14035 -420
rect 14115 -420 14160 -415
rect 14115 -425 14130 -420
rect 14025 -440 14130 -425
rect 14150 -425 14160 -420
rect 14235 -420 14275 -410
rect 14360 -415 14400 -410
rect 14235 -425 14245 -420
rect 14150 -440 14245 -425
rect 14265 -425 14275 -420
rect 14355 -420 14400 -415
rect 14355 -425 14370 -420
rect 14265 -440 14370 -425
rect 14390 -425 14400 -420
rect 14475 -420 14515 -410
rect 14600 -415 14640 -410
rect 14475 -425 14485 -420
rect 14390 -440 14485 -425
rect 14505 -425 14515 -420
rect 14595 -420 14640 -415
rect 14595 -425 14610 -420
rect 14505 -440 14610 -425
rect 14630 -425 14640 -420
rect 14715 -420 14755 -410
rect 14840 -415 14880 -410
rect 14715 -425 14725 -420
rect 14630 -440 14725 -425
rect 14745 -425 14755 -420
rect 14835 -420 14880 -415
rect 14835 -425 14850 -420
rect 14745 -440 14850 -425
rect 14870 -425 14880 -420
rect 14955 -420 14995 -410
rect 15080 -415 15120 -410
rect 14955 -425 14965 -420
rect 14870 -440 14965 -425
rect 14985 -425 14995 -420
rect 15075 -420 15120 -415
rect 15075 -425 15090 -420
rect 14985 -440 15090 -425
rect 15110 -425 15120 -420
rect 15195 -420 15235 -410
rect 15320 -415 15360 -410
rect 15195 -425 15205 -420
rect 15110 -440 15205 -425
rect 15225 -425 15235 -420
rect 15315 -420 15360 -415
rect 15315 -425 15330 -420
rect 15225 -440 15330 -425
rect 15350 -425 15360 -420
rect 15435 -420 15475 -410
rect 15560 -415 15600 -410
rect 15435 -425 15445 -420
rect 15350 -440 15445 -425
rect 15465 -425 15475 -420
rect 15555 -420 15600 -415
rect 15555 -425 15570 -420
rect 15465 -440 15570 -425
rect 15590 -425 15600 -420
rect 15675 -420 15715 -410
rect 15800 -415 15840 -410
rect 15675 -425 15685 -420
rect 15590 -440 15685 -425
rect 15705 -425 15715 -420
rect 15795 -420 15840 -415
rect 15795 -425 15810 -420
rect 15705 -440 15810 -425
rect 15830 -425 15840 -420
rect 15915 -420 15955 -410
rect 16040 -415 16080 -410
rect 15915 -425 15925 -420
rect 15830 -440 15925 -425
rect 15945 -425 15955 -420
rect 16035 -420 16080 -415
rect 16035 -425 16050 -420
rect 15945 -440 16050 -425
rect 16070 -425 16080 -420
rect 16155 -420 16195 -410
rect 16280 -415 16320 -410
rect 16155 -425 16165 -420
rect 16070 -440 16165 -425
rect 16185 -425 16195 -420
rect 16275 -420 16320 -415
rect 16275 -425 16290 -420
rect 16185 -440 16290 -425
rect 16310 -425 16320 -420
rect 16395 -420 16435 -410
rect 16520 -415 16560 -410
rect 16395 -425 16405 -420
rect 16310 -440 16405 -425
rect 16425 -425 16435 -420
rect 16515 -420 16560 -415
rect 16515 -425 16530 -420
rect 16425 -440 16530 -425
rect 16550 -425 16560 -420
rect 16635 -420 16675 -410
rect 16760 -415 16800 -410
rect 16635 -425 16645 -420
rect 16550 -440 16645 -425
rect 16665 -425 16675 -420
rect 16755 -420 16800 -415
rect 16755 -425 16770 -420
rect 16665 -440 16770 -425
rect 16790 -425 16800 -420
rect 16875 -420 16915 -410
rect 17000 -415 17040 -410
rect 16875 -425 16885 -420
rect 16790 -440 16885 -425
rect 16905 -425 16915 -420
rect 16995 -420 17040 -415
rect 16995 -425 17010 -420
rect 16905 -440 17010 -425
rect 17030 -425 17040 -420
rect 17115 -420 17155 -410
rect 17240 -415 17280 -410
rect 17115 -425 17125 -420
rect 17030 -440 17125 -425
rect 17145 -425 17155 -420
rect 17235 -420 17280 -415
rect 17235 -425 17250 -420
rect 17145 -440 17250 -425
rect 17270 -425 17280 -420
rect 17355 -420 17395 -410
rect 17480 -415 17520 -410
rect 17355 -425 17365 -420
rect 17270 -440 17365 -425
rect 17385 -425 17395 -420
rect 17475 -420 17520 -415
rect 17475 -425 17490 -420
rect 17385 -440 17490 -425
rect 17510 -425 17520 -420
rect 17595 -420 17635 -410
rect 17720 -415 17760 -410
rect 17595 -425 17605 -420
rect 17510 -440 17605 -425
rect 17625 -425 17635 -420
rect 17715 -420 17760 -415
rect 17715 -425 17730 -420
rect 17625 -440 17730 -425
rect 17750 -425 17760 -420
rect 17835 -420 17875 -410
rect 17960 -415 18000 -410
rect 17835 -425 17845 -420
rect 17750 -440 17845 -425
rect 17865 -425 17875 -420
rect 17955 -420 18000 -415
rect 17955 -425 17970 -420
rect 17865 -440 17970 -425
rect 17990 -425 18000 -420
rect 18075 -420 18115 -410
rect 18200 -415 18240 -410
rect 18075 -425 18085 -420
rect 17990 -440 18085 -425
rect 18105 -425 18115 -420
rect 18195 -420 18240 -415
rect 18195 -425 18210 -420
rect 18105 -440 18210 -425
rect 18230 -425 18240 -420
rect 18315 -420 18355 -410
rect 18440 -415 18480 -410
rect 18315 -425 18325 -420
rect 18230 -440 18325 -425
rect 18345 -425 18355 -420
rect 18435 -420 18480 -415
rect 18435 -425 18450 -420
rect 18345 -440 18450 -425
rect 18470 -425 18480 -420
rect 18555 -420 18595 -410
rect 18680 -415 18720 -410
rect 18555 -425 18565 -420
rect 18470 -440 18565 -425
rect 18585 -425 18595 -420
rect 18675 -420 18720 -415
rect 18675 -425 18690 -420
rect 18585 -440 18690 -425
rect 18710 -425 18720 -420
rect 18795 -420 18835 -410
rect 18920 -415 18960 -410
rect 18795 -425 18805 -420
rect 18710 -440 18805 -425
rect 18825 -425 18835 -420
rect 18915 -420 18960 -415
rect 18915 -425 18930 -420
rect 18825 -440 18930 -425
rect 18950 -425 18960 -420
rect 19035 -420 19075 -410
rect 19160 -415 19200 -410
rect 19035 -425 19045 -420
rect 18950 -440 19045 -425
rect 19065 -425 19075 -420
rect 19155 -420 19200 -415
rect 19155 -425 19170 -420
rect 19065 -440 19170 -425
rect 19190 -425 19200 -420
rect 19275 -420 19315 -410
rect 19400 -415 19440 -410
rect 19275 -425 19285 -420
rect 19190 -440 19285 -425
rect 19305 -425 19315 -420
rect 19395 -420 19440 -415
rect 19395 -425 19410 -420
rect 19305 -440 19410 -425
rect 19430 -425 19440 -420
rect 19515 -420 19555 -410
rect 19640 -415 19680 -410
rect 19515 -425 19525 -420
rect 19430 -440 19525 -425
rect 19545 -425 19555 -420
rect 19635 -420 19680 -415
rect 19635 -425 19650 -420
rect 19545 -440 19650 -425
rect 19670 -425 19680 -420
rect 19755 -420 19795 -410
rect 19880 -415 19920 -410
rect 19755 -425 19765 -420
rect 19670 -440 19765 -425
rect 19785 -425 19795 -420
rect 19875 -420 19920 -415
rect 19875 -425 19890 -420
rect 19785 -440 19890 -425
rect 19910 -425 19920 -420
rect 19995 -420 20035 -410
rect 20120 -415 20160 -410
rect 19995 -425 20005 -420
rect 19910 -440 20005 -425
rect 20025 -425 20035 -420
rect 20115 -420 20160 -415
rect 20115 -425 20130 -420
rect 20025 -440 20130 -425
rect 20150 -425 20160 -420
rect 20235 -420 20275 -410
rect 20360 -415 20400 -410
rect 20235 -425 20245 -420
rect 20150 -440 20245 -425
rect 20265 -425 20275 -420
rect 20355 -420 20400 -415
rect 20355 -425 20370 -420
rect 20265 -440 20370 -425
rect 20390 -425 20400 -420
rect 20475 -420 20515 -410
rect 20600 -415 20640 -410
rect 20475 -425 20485 -420
rect 20390 -440 20485 -425
rect 20505 -425 20515 -420
rect 20595 -420 20640 -415
rect 20595 -425 20610 -420
rect 20505 -440 20610 -425
rect 20630 -425 20640 -420
rect 20715 -420 20755 -410
rect 20840 -415 20880 -410
rect 20715 -425 20725 -420
rect 20630 -440 20725 -425
rect 20745 -425 20755 -420
rect 20835 -420 20880 -415
rect 20835 -425 20850 -420
rect 20745 -440 20850 -425
rect 20870 -425 20880 -420
rect 20955 -420 20995 -410
rect 21080 -415 21120 -410
rect 20955 -425 20965 -420
rect 20870 -440 20965 -425
rect 20985 -425 20995 -420
rect 21075 -420 21120 -415
rect 21075 -425 21090 -420
rect 20985 -440 21090 -425
rect 21110 -425 21120 -420
rect 21195 -420 21235 -410
rect 21320 -415 21360 -410
rect 21195 -425 21205 -420
rect 21110 -440 21205 -425
rect 21225 -425 21235 -420
rect 21315 -420 21360 -415
rect 21315 -425 21330 -420
rect 21225 -440 21330 -425
rect 21350 -425 21360 -420
rect 21435 -420 21475 -410
rect 21560 -415 21600 -410
rect 21435 -425 21445 -420
rect 21350 -440 21445 -425
rect 21465 -425 21475 -420
rect 21555 -420 21600 -415
rect 21555 -425 21570 -420
rect 21465 -440 21570 -425
rect 21590 -425 21600 -420
rect 21675 -420 21715 -410
rect 21800 -415 21840 -410
rect 21675 -425 21685 -420
rect 21590 -440 21685 -425
rect 21705 -425 21715 -420
rect 21795 -420 21840 -415
rect 21795 -425 21810 -420
rect 21705 -440 21810 -425
rect 21830 -425 21840 -420
rect 21915 -420 21955 -410
rect 22040 -415 22080 -410
rect 21915 -425 21925 -420
rect 21830 -440 21925 -425
rect 21945 -425 21955 -420
rect 22035 -420 22080 -415
rect 22035 -425 22050 -420
rect 21945 -440 22050 -425
rect 22070 -425 22080 -420
rect 22155 -420 22195 -410
rect 22280 -415 22320 -410
rect 22155 -425 22165 -420
rect 22070 -440 22165 -425
rect 22185 -425 22195 -420
rect 22275 -420 22320 -415
rect 22275 -425 22290 -420
rect 22185 -440 22290 -425
rect 22310 -425 22320 -420
rect 22395 -420 22435 -410
rect 22520 -415 22560 -410
rect 22395 -425 22405 -420
rect 22310 -440 22405 -425
rect 22425 -425 22435 -420
rect 22515 -420 22560 -415
rect 22515 -425 22530 -420
rect 22425 -440 22530 -425
rect 22550 -425 22560 -420
rect 22635 -420 22675 -410
rect 22760 -415 22800 -410
rect 22635 -425 22645 -420
rect 22550 -440 22645 -425
rect 22665 -425 22675 -420
rect 22755 -420 22800 -415
rect 22755 -425 22770 -420
rect 22665 -440 22770 -425
rect 22790 -425 22800 -420
rect 22875 -420 22915 -410
rect 23000 -415 23040 -410
rect 22875 -425 22885 -420
rect 22790 -440 22885 -425
rect 22905 -425 22915 -420
rect 22995 -420 23040 -415
rect 22995 -425 23010 -420
rect 22905 -440 23010 -425
rect 23030 -425 23040 -420
rect 23115 -420 23155 -410
rect 23240 -415 23280 -410
rect 23115 -425 23125 -420
rect 23030 -440 23125 -425
rect 23145 -425 23155 -420
rect 23235 -420 23280 -415
rect 23235 -425 23250 -420
rect 23145 -440 23250 -425
rect 23270 -425 23280 -420
rect 23355 -420 23395 -410
rect 23480 -415 23520 -410
rect 23355 -425 23365 -420
rect 23270 -440 23365 -425
rect 23385 -425 23395 -420
rect 23475 -420 23520 -415
rect 23475 -425 23490 -420
rect 23385 -440 23490 -425
rect 23510 -425 23520 -420
rect 23595 -420 23635 -410
rect 23720 -415 23760 -410
rect 23595 -425 23605 -420
rect 23510 -440 23605 -425
rect 23625 -425 23635 -420
rect 23715 -420 23760 -415
rect 23715 -425 23730 -420
rect 23625 -440 23730 -425
rect 23750 -425 23760 -420
rect 23835 -420 23875 -410
rect 23960 -415 24000 -410
rect 23835 -425 23845 -420
rect 23750 -440 23845 -425
rect 23865 -425 23875 -420
rect 23955 -420 24000 -415
rect 23955 -425 23970 -420
rect 23865 -440 23970 -425
rect 23990 -425 24000 -420
rect 24075 -420 24115 -410
rect 24200 -415 24240 -410
rect 24075 -425 24085 -420
rect 23990 -440 24085 -425
rect 24105 -425 24115 -420
rect 24195 -420 24240 -415
rect 24195 -425 24210 -420
rect 24105 -440 24210 -425
rect 24230 -425 24240 -420
rect 24315 -420 24355 -410
rect 24440 -415 24480 -410
rect 24315 -425 24325 -420
rect 24230 -440 24325 -425
rect 24345 -425 24355 -420
rect 24435 -420 24480 -415
rect 24435 -425 24450 -420
rect 24345 -440 24450 -425
rect 24470 -425 24480 -420
rect 24555 -420 24595 -410
rect 24680 -415 24720 -410
rect 24555 -425 24565 -420
rect 24470 -440 24565 -425
rect 24585 -425 24595 -420
rect 24675 -420 24720 -415
rect 24675 -425 24690 -420
rect 24585 -440 24690 -425
rect 24710 -425 24720 -420
rect 24795 -420 24835 -410
rect 24920 -415 24960 -410
rect 24795 -425 24805 -420
rect 24710 -440 24805 -425
rect 24825 -425 24835 -420
rect 24915 -420 24960 -415
rect 24915 -425 24930 -420
rect 24825 -440 24930 -425
rect 24950 -425 24960 -420
rect 25035 -420 25075 -410
rect 25160 -415 25200 -410
rect 25035 -425 25045 -420
rect 24950 -440 25045 -425
rect 25065 -425 25075 -420
rect 25155 -420 25200 -415
rect 25155 -425 25170 -420
rect 25065 -440 25170 -425
rect 25190 -425 25200 -420
rect 25275 -420 25315 -410
rect 25400 -415 25440 -410
rect 25275 -425 25285 -420
rect 25190 -440 25285 -425
rect 25305 -425 25315 -420
rect 25395 -420 25440 -415
rect 25395 -425 25410 -420
rect 25305 -440 25410 -425
rect 25430 -425 25440 -420
rect 25515 -420 25555 -410
rect 25640 -415 25680 -410
rect 25515 -425 25525 -420
rect 25430 -440 25525 -425
rect 25545 -425 25555 -420
rect 25635 -420 25680 -415
rect 25635 -425 25650 -420
rect 25545 -440 25650 -425
rect 25670 -425 25680 -420
rect 25755 -420 25795 -410
rect 25880 -415 25920 -410
rect 25755 -425 25765 -420
rect 25670 -440 25765 -425
rect 25785 -425 25795 -420
rect 25875 -420 25920 -415
rect 25875 -425 25890 -420
rect 25785 -440 25890 -425
rect 25910 -425 25920 -420
rect 25995 -420 26035 -410
rect 26120 -415 26160 -410
rect 25995 -425 26005 -420
rect 25910 -440 26005 -425
rect 26025 -425 26035 -420
rect 26115 -420 26160 -415
rect 26115 -425 26130 -420
rect 26025 -440 26130 -425
rect 26150 -425 26160 -420
rect 26235 -420 26275 -410
rect 26360 -415 26400 -410
rect 26235 -425 26245 -420
rect 26150 -440 26245 -425
rect 26265 -425 26275 -420
rect 26355 -420 26400 -415
rect 26355 -425 26370 -420
rect 26265 -440 26370 -425
rect 26390 -425 26400 -420
rect 26475 -420 26515 -410
rect 26600 -415 26640 -410
rect 26475 -425 26485 -420
rect 26390 -440 26485 -425
rect 26505 -425 26515 -420
rect 26595 -420 26640 -415
rect 26595 -425 26610 -420
rect 26505 -440 26610 -425
rect 26630 -425 26640 -420
rect 26715 -420 26755 -410
rect 26840 -415 26880 -410
rect 26715 -425 26725 -420
rect 26630 -440 26725 -425
rect 26745 -425 26755 -420
rect 26835 -420 26880 -415
rect 26835 -425 26850 -420
rect 26745 -440 26850 -425
rect 26870 -425 26880 -420
rect 26955 -420 26995 -410
rect 27080 -415 27120 -410
rect 26955 -425 26965 -420
rect 26870 -440 26965 -425
rect 26985 -425 26995 -420
rect 27075 -420 27120 -415
rect 27075 -425 27090 -420
rect 26985 -440 27090 -425
rect 27110 -425 27120 -420
rect 27195 -420 27235 -410
rect 27320 -415 27360 -410
rect 27195 -425 27205 -420
rect 27110 -440 27205 -425
rect 27225 -425 27235 -420
rect 27315 -420 27360 -415
rect 27315 -425 27330 -420
rect 27225 -440 27330 -425
rect 27350 -425 27360 -420
rect 27435 -420 27475 -410
rect 27560 -415 27600 -410
rect 27435 -425 27445 -420
rect 27350 -440 27445 -425
rect 27465 -425 27475 -420
rect 27555 -420 27600 -415
rect 27555 -425 27570 -420
rect 27465 -440 27570 -425
rect 27590 -425 27600 -420
rect 27675 -420 27715 -410
rect 27800 -415 27840 -410
rect 27675 -425 27685 -420
rect 27590 -440 27685 -425
rect 27705 -425 27715 -420
rect 27795 -420 27840 -415
rect 27795 -425 27810 -420
rect 27705 -440 27810 -425
rect 27830 -425 27840 -420
rect 27915 -420 27955 -410
rect 28040 -415 28080 -410
rect 27915 -425 27925 -420
rect 27830 -440 27925 -425
rect 27945 -425 27955 -420
rect 28035 -420 28080 -415
rect 28035 -425 28050 -420
rect 27945 -440 28050 -425
rect 28070 -425 28080 -420
rect 28155 -420 28195 -410
rect 28280 -415 28320 -410
rect 28155 -425 28165 -420
rect 28070 -440 28165 -425
rect 28185 -425 28195 -420
rect 28275 -420 28320 -415
rect 28275 -425 28290 -420
rect 28185 -440 28290 -425
rect 28310 -425 28320 -420
rect 28395 -420 28435 -410
rect 28520 -415 28560 -410
rect 28395 -425 28405 -420
rect 28310 -440 28405 -425
rect 28425 -425 28435 -420
rect 28515 -420 28560 -415
rect 28515 -425 28530 -420
rect 28425 -440 28530 -425
rect 28550 -425 28560 -420
rect 28635 -420 28675 -410
rect 28760 -415 28800 -410
rect 28635 -425 28645 -420
rect 28550 -440 28645 -425
rect 28665 -425 28675 -420
rect 28755 -420 28800 -415
rect 28755 -425 28770 -420
rect 28665 -440 28770 -425
rect 28790 -425 28800 -420
rect 28875 -420 28915 -410
rect 29000 -415 29040 -410
rect 28875 -425 28885 -420
rect 28790 -440 28885 -425
rect 28905 -425 28915 -420
rect 28995 -420 29040 -415
rect 28995 -425 29010 -420
rect 28905 -440 29010 -425
rect 29030 -425 29040 -420
rect 29115 -420 29155 -410
rect 29240 -415 29280 -410
rect 29115 -425 29125 -420
rect 29030 -440 29125 -425
rect 29145 -425 29155 -420
rect 29235 -420 29280 -415
rect 29235 -425 29250 -420
rect 29145 -440 29250 -425
rect 29270 -425 29280 -420
rect 29355 -420 29395 -410
rect 29480 -415 29520 -410
rect 29355 -425 29365 -420
rect 29270 -440 29365 -425
rect 29385 -425 29395 -420
rect 29475 -420 29520 -415
rect 29475 -425 29490 -420
rect 29385 -440 29490 -425
rect 29510 -425 29520 -420
rect 29595 -420 29635 -410
rect 29720 -415 29760 -410
rect 29595 -425 29605 -420
rect 29510 -440 29605 -425
rect 29625 -425 29635 -420
rect 29715 -420 29760 -415
rect 29715 -425 29730 -420
rect 29625 -440 29730 -425
rect 29750 -425 29760 -420
rect 29835 -420 29875 -410
rect 29960 -415 30000 -410
rect 29835 -425 29845 -420
rect 29750 -440 29845 -425
rect 29865 -425 29875 -420
rect 29955 -420 30000 -415
rect 29955 -425 29970 -420
rect 29865 -440 29970 -425
rect 29990 -425 30000 -420
rect 30075 -420 30115 -410
rect 30200 -415 30240 -410
rect 30075 -425 30085 -420
rect 29990 -440 30085 -425
rect 30105 -425 30115 -420
rect 30195 -420 30240 -415
rect 30195 -425 30210 -420
rect 30105 -440 30210 -425
rect 30230 -425 30240 -420
rect 30315 -420 30355 -410
rect 30440 -415 30480 -410
rect 30315 -425 30325 -420
rect 30230 -440 30325 -425
rect 30345 -425 30355 -420
rect 30435 -420 30480 -415
rect 30435 -425 30450 -420
rect 30345 -440 30450 -425
rect 30470 -425 30480 -420
rect 30555 -420 30595 -410
rect 30555 -425 30565 -420
rect 30470 -440 30565 -425
rect 30585 -425 30595 -420
rect 30675 -425 30715 -415
rect 30585 -440 30685 -425
rect -40 -450 0 -440
rect 75 -450 115 -440
rect 195 -450 240 -440
rect 315 -450 355 -440
rect 435 -450 480 -440
rect 555 -450 595 -440
rect 675 -450 720 -440
rect 795 -450 835 -440
rect 915 -450 960 -440
rect 1035 -450 1075 -440
rect 1155 -450 1200 -440
rect 1275 -450 1315 -440
rect 1395 -450 1440 -440
rect 1515 -450 1555 -440
rect 1635 -450 1680 -440
rect 1755 -450 1795 -440
rect 1875 -450 1920 -440
rect 1995 -450 2035 -440
rect 2115 -450 2160 -440
rect 2235 -450 2275 -440
rect 2355 -450 2400 -440
rect 2475 -450 2515 -440
rect 2595 -450 2640 -440
rect 2715 -450 2755 -440
rect 2835 -450 2880 -440
rect 2955 -450 2995 -440
rect 3075 -450 3120 -440
rect 3195 -450 3235 -440
rect 3315 -450 3360 -440
rect 3435 -450 3475 -440
rect 3555 -450 3600 -440
rect 3675 -450 3715 -440
rect 3795 -450 3840 -440
rect 3915 -450 3955 -440
rect 4035 -450 4080 -440
rect 4155 -450 4195 -440
rect 4275 -450 4320 -440
rect 4395 -450 4435 -440
rect 4515 -450 4560 -440
rect 4635 -450 4675 -440
rect 4755 -450 4800 -440
rect 4875 -450 4915 -440
rect 4995 -450 5040 -440
rect 5115 -450 5155 -440
rect 5235 -450 5280 -440
rect 5355 -450 5395 -440
rect 5475 -450 5520 -440
rect 5595 -450 5635 -440
rect 5715 -450 5760 -440
rect 5835 -450 5875 -440
rect 5955 -450 6000 -440
rect 6075 -450 6115 -440
rect 6195 -450 6240 -440
rect 6315 -450 6355 -440
rect 6435 -450 6480 -440
rect 6555 -450 6595 -440
rect 6675 -450 6720 -440
rect 6795 -450 6835 -440
rect 6915 -450 6960 -440
rect 7035 -450 7075 -440
rect 7155 -450 7200 -440
rect 7275 -450 7315 -440
rect 7395 -450 7440 -440
rect 7515 -450 7555 -440
rect 7635 -450 7680 -440
rect 7755 -450 7795 -440
rect 7875 -450 7920 -440
rect 7995 -450 8035 -440
rect 8115 -450 8160 -440
rect 8235 -450 8275 -440
rect 8355 -450 8400 -440
rect 8475 -450 8515 -440
rect 8595 -450 8640 -440
rect 8715 -450 8755 -440
rect 8835 -450 8880 -440
rect 8955 -450 8995 -440
rect 9075 -450 9120 -440
rect 9195 -450 9235 -440
rect 9315 -450 9360 -440
rect 9435 -450 9475 -440
rect 9555 -450 9600 -440
rect 9675 -450 9715 -440
rect 9795 -450 9840 -440
rect 9915 -450 9955 -440
rect 10035 -450 10080 -440
rect 10155 -450 10195 -440
rect 10275 -450 10320 -440
rect 10395 -450 10435 -440
rect 10515 -450 10560 -440
rect 10635 -450 10675 -440
rect 10755 -450 10800 -440
rect 10875 -450 10915 -440
rect 10995 -450 11040 -440
rect 11115 -450 11155 -440
rect 11235 -450 11280 -440
rect 11355 -450 11395 -440
rect 11475 -450 11520 -440
rect 11595 -450 11635 -440
rect 11715 -450 11760 -440
rect 11835 -450 11875 -440
rect 11955 -450 12000 -440
rect 12075 -450 12115 -440
rect 12195 -450 12240 -440
rect 12315 -450 12355 -440
rect 12435 -450 12480 -440
rect 12555 -450 12595 -440
rect 12675 -450 12720 -440
rect 12795 -450 12835 -440
rect 12915 -450 12960 -440
rect 13035 -450 13075 -440
rect 13155 -450 13200 -440
rect 13275 -450 13315 -440
rect 13395 -450 13440 -440
rect 13515 -450 13555 -440
rect 13635 -450 13680 -440
rect 13755 -450 13795 -440
rect 13875 -450 13920 -440
rect 13995 -450 14035 -440
rect 14115 -450 14160 -440
rect 14235 -450 14275 -440
rect 14355 -450 14400 -440
rect 14475 -450 14515 -440
rect 14595 -450 14640 -440
rect 14715 -450 14755 -440
rect 14835 -450 14880 -440
rect 14955 -450 14995 -440
rect 15075 -450 15120 -440
rect 15195 -450 15235 -440
rect 15315 -450 15360 -440
rect 15435 -450 15475 -440
rect 15555 -450 15600 -440
rect 15675 -450 15715 -440
rect 15795 -450 15840 -440
rect 15915 -450 15955 -440
rect 16035 -450 16080 -440
rect 16155 -450 16195 -440
rect 16275 -450 16320 -440
rect 16395 -450 16435 -440
rect 16515 -450 16560 -440
rect 16635 -450 16675 -440
rect 16755 -450 16800 -440
rect 16875 -450 16915 -440
rect 16995 -450 17040 -440
rect 17115 -450 17155 -440
rect 17235 -450 17280 -440
rect 17355 -450 17395 -440
rect 17475 -450 17520 -440
rect 17595 -450 17635 -440
rect 17715 -450 17760 -440
rect 17835 -450 17875 -440
rect 17955 -450 18000 -440
rect 18075 -450 18115 -440
rect 18195 -450 18240 -440
rect 18315 -450 18355 -440
rect 18435 -450 18480 -440
rect 18555 -450 18595 -440
rect 18675 -450 18720 -440
rect 18795 -450 18835 -440
rect 18915 -450 18960 -440
rect 19035 -450 19075 -440
rect 19155 -450 19200 -440
rect 19275 -450 19315 -440
rect 19395 -450 19440 -440
rect 19515 -450 19555 -440
rect 19635 -450 19680 -440
rect 19755 -450 19795 -440
rect 19875 -450 19920 -440
rect 19995 -450 20035 -440
rect 20115 -450 20160 -440
rect 20235 -450 20275 -440
rect 20355 -450 20400 -440
rect 20475 -450 20515 -440
rect 20595 -450 20640 -440
rect 20715 -450 20755 -440
rect 20835 -450 20880 -440
rect 20955 -450 20995 -440
rect 21075 -450 21120 -440
rect 21195 -450 21235 -440
rect 21315 -450 21360 -440
rect 21435 -450 21475 -440
rect 21555 -450 21600 -440
rect 21675 -450 21715 -440
rect 21795 -450 21840 -440
rect 21915 -450 21955 -440
rect 22035 -450 22080 -440
rect 22155 -450 22195 -440
rect 22275 -450 22320 -440
rect 22395 -450 22435 -440
rect 22515 -450 22560 -440
rect 22635 -450 22675 -440
rect 22755 -450 22800 -440
rect 22875 -450 22915 -440
rect 22995 -450 23040 -440
rect 23115 -450 23155 -440
rect 23235 -450 23280 -440
rect 23355 -450 23395 -440
rect 23475 -450 23520 -440
rect 23595 -450 23635 -440
rect 23715 -450 23760 -440
rect 23835 -450 23875 -440
rect 23955 -450 24000 -440
rect 24075 -450 24115 -440
rect 24195 -450 24240 -440
rect 24315 -450 24355 -440
rect 24435 -450 24480 -440
rect 24555 -450 24595 -440
rect 24675 -450 24720 -440
rect 24795 -450 24835 -440
rect 24915 -450 24960 -440
rect 25035 -450 25075 -440
rect 25155 -450 25200 -440
rect 25275 -450 25315 -440
rect 25395 -450 25440 -440
rect 25515 -450 25555 -440
rect 25635 -450 25680 -440
rect 25755 -450 25795 -440
rect 25875 -450 25920 -440
rect 25995 -450 26035 -440
rect 26115 -450 26160 -440
rect 26235 -450 26275 -440
rect 26355 -450 26400 -440
rect 26475 -450 26515 -440
rect 26595 -450 26640 -440
rect 26715 -450 26755 -440
rect 26835 -450 26880 -440
rect 26955 -450 26995 -440
rect 27075 -450 27120 -440
rect 27195 -450 27235 -440
rect 27315 -450 27360 -440
rect 27435 -450 27475 -440
rect 27555 -450 27600 -440
rect 27675 -450 27715 -440
rect 27795 -450 27840 -440
rect 27915 -450 27955 -440
rect 28035 -450 28080 -440
rect 28155 -450 28195 -440
rect 28275 -450 28320 -440
rect 28395 -450 28435 -440
rect 28515 -450 28560 -440
rect 28635 -450 28675 -440
rect 28755 -450 28800 -440
rect 28875 -450 28915 -440
rect 28995 -450 29040 -440
rect 29115 -450 29155 -440
rect 29235 -450 29280 -440
rect 29355 -450 29395 -440
rect 29475 -450 29520 -440
rect 29595 -450 29635 -440
rect 29715 -450 29760 -440
rect 29835 -450 29875 -440
rect 29955 -450 30000 -440
rect 30075 -450 30115 -440
rect 30195 -450 30240 -440
rect 30315 -450 30355 -440
rect 30435 -450 30480 -440
rect 30555 -450 30595 -440
rect 30675 -445 30685 -440
rect 30705 -445 30715 -425
rect 195 -455 235 -450
rect 435 -455 475 -450
rect 675 -455 715 -450
rect 915 -455 955 -450
rect 1155 -455 1195 -450
rect 1395 -455 1435 -450
rect 1635 -455 1675 -450
rect 1875 -455 1915 -450
rect 2115 -455 2155 -450
rect 2355 -455 2395 -450
rect 2595 -455 2635 -450
rect 2835 -455 2875 -450
rect 3075 -455 3115 -450
rect 3315 -455 3355 -450
rect 3555 -455 3595 -450
rect 3795 -455 3835 -450
rect 4035 -455 4075 -450
rect 4275 -455 4315 -450
rect 4515 -455 4555 -450
rect 4755 -455 4795 -450
rect 4995 -455 5035 -450
rect 5235 -455 5275 -450
rect 5475 -455 5515 -450
rect 5715 -455 5755 -450
rect 5955 -455 5995 -450
rect 6195 -455 6235 -450
rect 6435 -455 6475 -450
rect 6675 -455 6715 -450
rect 6915 -455 6955 -450
rect 7155 -455 7195 -450
rect 7395 -455 7435 -450
rect 7635 -455 7675 -450
rect 7875 -455 7915 -450
rect 8115 -455 8155 -450
rect 8355 -455 8395 -450
rect 8595 -455 8635 -450
rect 8835 -455 8875 -450
rect 9075 -455 9115 -450
rect 9315 -455 9355 -450
rect 9555 -455 9595 -450
rect 9795 -455 9835 -450
rect 10035 -455 10075 -450
rect 10275 -455 10315 -450
rect 10515 -455 10555 -450
rect 10755 -455 10795 -450
rect 10995 -455 11035 -450
rect 11235 -455 11275 -450
rect 11475 -455 11515 -450
rect 11715 -455 11755 -450
rect 11955 -455 11995 -450
rect 12195 -455 12235 -450
rect 12435 -455 12475 -450
rect 12675 -455 12715 -450
rect 12915 -455 12955 -450
rect 13155 -455 13195 -450
rect 13395 -455 13435 -450
rect 13635 -455 13675 -450
rect 13875 -455 13915 -450
rect 14115 -455 14155 -450
rect 14355 -455 14395 -450
rect 14595 -455 14635 -450
rect 14835 -455 14875 -450
rect 15075 -455 15115 -450
rect 15315 -455 15355 -450
rect 15555 -455 15595 -450
rect 15795 -455 15835 -450
rect 16035 -455 16075 -450
rect 16275 -455 16315 -450
rect 16515 -455 16555 -450
rect 16755 -455 16795 -450
rect 16995 -455 17035 -450
rect 17235 -455 17275 -450
rect 17475 -455 17515 -450
rect 17715 -455 17755 -450
rect 17955 -455 17995 -450
rect 18195 -455 18235 -450
rect 18435 -455 18475 -450
rect 18675 -455 18715 -450
rect 18915 -455 18955 -450
rect 19155 -455 19195 -450
rect 19395 -455 19435 -450
rect 19635 -455 19675 -450
rect 19875 -455 19915 -450
rect 20115 -455 20155 -450
rect 20355 -455 20395 -450
rect 20595 -455 20635 -450
rect 20835 -455 20875 -450
rect 21075 -455 21115 -450
rect 21315 -455 21355 -450
rect 21555 -455 21595 -450
rect 21795 -455 21835 -450
rect 22035 -455 22075 -450
rect 22275 -455 22315 -450
rect 22515 -455 22555 -450
rect 22755 -455 22795 -450
rect 22995 -455 23035 -450
rect 23235 -455 23275 -450
rect 23475 -455 23515 -450
rect 23715 -455 23755 -450
rect 23955 -455 23995 -450
rect 24195 -455 24235 -450
rect 24435 -455 24475 -450
rect 24675 -455 24715 -450
rect 24915 -455 24955 -450
rect 25155 -455 25195 -450
rect 25395 -455 25435 -450
rect 25635 -455 25675 -450
rect 25875 -455 25915 -450
rect 26115 -455 26155 -450
rect 26355 -455 26395 -450
rect 26595 -455 26635 -450
rect 26835 -455 26875 -450
rect 27075 -455 27115 -450
rect 27315 -455 27355 -450
rect 27555 -455 27595 -450
rect 27795 -455 27835 -450
rect 28035 -455 28075 -450
rect 28275 -455 28315 -450
rect 28515 -455 28555 -450
rect 28755 -455 28795 -450
rect 28995 -455 29035 -450
rect 29235 -455 29275 -450
rect 29475 -455 29515 -450
rect 29715 -455 29755 -450
rect 29955 -455 29995 -450
rect 30195 -455 30235 -450
rect 30435 -455 30475 -450
rect 30675 -455 30715 -445
rect 30730 -480 30770 -475
rect 30730 -510 30735 -480
rect 30765 -510 30770 -480
rect 30730 -515 30770 -510
rect -40 -545 0 -535
rect 80 -545 120 -535
rect 195 -545 240 -535
rect 320 -545 360 -535
rect 435 -545 480 -535
rect 560 -545 600 -535
rect 675 -545 720 -535
rect 800 -545 840 -535
rect 915 -545 960 -535
rect 1040 -545 1080 -535
rect 1155 -545 1200 -535
rect 1280 -545 1320 -535
rect 1395 -545 1440 -535
rect 1520 -545 1560 -535
rect 1635 -545 1680 -535
rect 1760 -545 1800 -535
rect 1875 -545 1920 -535
rect 2000 -545 2040 -535
rect 2115 -545 2160 -535
rect 2240 -545 2280 -535
rect 2355 -545 2400 -535
rect 2480 -545 2520 -535
rect 2595 -545 2640 -535
rect 2720 -545 2760 -535
rect 2835 -545 2880 -535
rect 2960 -545 3000 -535
rect 3075 -545 3120 -535
rect 3200 -545 3240 -535
rect 3315 -545 3360 -535
rect 3440 -545 3480 -535
rect 3555 -545 3600 -535
rect 3680 -545 3720 -535
rect 3795 -545 3840 -535
rect 3920 -545 3960 -535
rect 4035 -545 4080 -535
rect 4160 -545 4200 -535
rect 4275 -545 4320 -535
rect 4400 -545 4440 -535
rect 4515 -545 4560 -535
rect 4640 -545 4680 -535
rect 4755 -545 4800 -535
rect 4880 -545 4920 -535
rect 4995 -545 5040 -535
rect 5120 -545 5160 -535
rect 5235 -545 5280 -535
rect 5360 -545 5400 -535
rect 5475 -545 5520 -535
rect 5600 -545 5640 -535
rect 5715 -545 5760 -535
rect 5840 -545 5880 -535
rect 5955 -545 6000 -535
rect 6080 -545 6120 -535
rect 6195 -545 6240 -535
rect 6320 -545 6360 -535
rect 6435 -545 6480 -535
rect 6560 -545 6600 -535
rect 6675 -545 6720 -535
rect 6800 -545 6840 -535
rect 6915 -545 6960 -535
rect 7040 -545 7080 -535
rect 7155 -545 7200 -535
rect 7280 -545 7320 -535
rect 7395 -545 7440 -535
rect 7520 -545 7560 -535
rect 7635 -545 7680 -535
rect 7760 -545 7800 -535
rect 7875 -545 7920 -535
rect 8000 -545 8040 -535
rect 8115 -545 8160 -535
rect 8240 -545 8280 -535
rect 8355 -545 8400 -535
rect 8480 -545 8520 -535
rect 8595 -545 8640 -535
rect 8720 -545 8760 -535
rect 8835 -545 8880 -535
rect 8960 -545 9000 -535
rect 9075 -545 9120 -535
rect 9200 -545 9240 -535
rect 9315 -545 9360 -535
rect 9440 -545 9480 -535
rect 9555 -545 9600 -535
rect 9680 -545 9720 -535
rect 9795 -545 9840 -535
rect 9920 -545 9960 -535
rect 10035 -545 10080 -535
rect 10160 -545 10200 -535
rect 10275 -545 10320 -535
rect 10400 -545 10440 -535
rect 10515 -545 10560 -535
rect 10640 -545 10680 -535
rect 10755 -545 10800 -535
rect 10880 -545 10920 -535
rect 10995 -545 11040 -535
rect 11120 -545 11160 -535
rect 11235 -545 11280 -535
rect 11360 -545 11400 -535
rect 11475 -545 11520 -535
rect 11600 -545 11640 -535
rect 11715 -545 11760 -535
rect 11840 -545 11880 -535
rect 11955 -545 12000 -535
rect 12080 -545 12120 -535
rect 12195 -545 12240 -535
rect 12320 -545 12360 -535
rect 12435 -545 12480 -535
rect 12560 -545 12600 -535
rect 12675 -545 12720 -535
rect 12800 -545 12840 -535
rect 12915 -545 12960 -535
rect 13040 -545 13080 -535
rect 13155 -545 13200 -535
rect 13280 -545 13320 -535
rect 13395 -545 13440 -535
rect 13520 -545 13560 -535
rect 13635 -545 13680 -535
rect 13760 -545 13800 -535
rect 13875 -545 13920 -535
rect 14000 -545 14040 -535
rect 14115 -545 14160 -535
rect 14240 -545 14280 -535
rect 14355 -545 14400 -535
rect 14480 -545 14520 -535
rect 14595 -545 14640 -535
rect 14720 -545 14760 -535
rect 14835 -545 14880 -535
rect 14960 -545 15000 -535
rect 15075 -545 15120 -535
rect 15200 -545 15240 -535
rect 15315 -545 15360 -535
rect 15440 -545 15480 -535
rect 15555 -545 15600 -535
rect 15680 -545 15720 -535
rect 15795 -545 15840 -535
rect 15920 -545 15960 -535
rect 16035 -545 16080 -535
rect 16160 -545 16200 -535
rect 16275 -545 16320 -535
rect 16400 -545 16440 -535
rect 16515 -545 16560 -535
rect 16640 -545 16680 -535
rect 16755 -545 16800 -535
rect 16880 -545 16920 -535
rect 16995 -545 17040 -535
rect 17120 -545 17160 -535
rect 17235 -545 17280 -535
rect 17360 -545 17400 -535
rect 17475 -545 17520 -535
rect 17600 -545 17640 -535
rect 17715 -545 17760 -535
rect 17840 -545 17880 -535
rect 17955 -545 18000 -535
rect 18080 -545 18120 -535
rect 18195 -545 18240 -535
rect 18320 -545 18360 -535
rect 18435 -545 18480 -535
rect 18560 -545 18600 -535
rect 18675 -545 18720 -535
rect 18800 -545 18840 -535
rect 18915 -545 18960 -535
rect 19040 -545 19080 -535
rect 19155 -545 19200 -535
rect 19280 -545 19320 -535
rect 19395 -545 19440 -535
rect 19520 -545 19560 -535
rect 19635 -545 19680 -535
rect 19760 -545 19800 -535
rect 19875 -545 19920 -535
rect 20000 -545 20040 -535
rect 20115 -545 20160 -535
rect 20240 -545 20280 -535
rect 20355 -545 20400 -535
rect 20480 -545 20520 -535
rect 20595 -545 20640 -535
rect 20720 -545 20760 -535
rect 20835 -545 20880 -535
rect 20960 -545 21000 -535
rect 21075 -545 21120 -535
rect 21200 -545 21240 -535
rect 21315 -545 21360 -535
rect 21440 -545 21480 -535
rect 21555 -545 21600 -535
rect 21680 -545 21720 -535
rect 21795 -545 21840 -535
rect 21920 -545 21960 -535
rect 22035 -545 22080 -535
rect 22160 -545 22200 -535
rect 22275 -545 22320 -535
rect 22400 -545 22440 -535
rect 22515 -545 22560 -535
rect 22640 -545 22680 -535
rect 22755 -545 22800 -535
rect 22880 -545 22920 -535
rect 22995 -545 23040 -535
rect 23120 -545 23160 -535
rect 23235 -545 23280 -535
rect 23360 -545 23400 -535
rect 23475 -545 23520 -535
rect 23600 -545 23640 -535
rect 23715 -545 23760 -535
rect 23840 -545 23880 -535
rect 23955 -545 24000 -535
rect 24080 -545 24120 -535
rect 24195 -545 24240 -535
rect 24320 -545 24360 -535
rect 24435 -545 24480 -535
rect 24560 -545 24600 -535
rect 24675 -545 24720 -535
rect 24800 -545 24840 -535
rect 24915 -545 24960 -535
rect 25040 -545 25080 -535
rect 25155 -545 25200 -535
rect 25280 -545 25320 -535
rect 25395 -545 25440 -535
rect 25520 -545 25560 -535
rect 25635 -545 25680 -535
rect 25760 -545 25800 -535
rect 25875 -545 25920 -535
rect 26000 -545 26040 -535
rect 26115 -545 26160 -535
rect 26240 -545 26280 -535
rect 26355 -545 26400 -535
rect 26480 -545 26520 -535
rect 26595 -545 26640 -535
rect 26720 -545 26760 -535
rect 26835 -545 26880 -535
rect 26960 -545 27000 -535
rect 27075 -545 27120 -535
rect 27200 -545 27240 -535
rect 27315 -545 27360 -535
rect 27440 -545 27480 -535
rect 27555 -545 27600 -535
rect 27680 -545 27720 -535
rect 27795 -545 27840 -535
rect 27920 -545 27960 -535
rect 28035 -545 28080 -535
rect 28160 -545 28200 -535
rect 28275 -545 28320 -535
rect 28400 -545 28440 -535
rect 28515 -545 28560 -535
rect 28640 -545 28680 -535
rect 28755 -545 28800 -535
rect 28880 -545 28920 -535
rect 28995 -545 29040 -535
rect 29120 -545 29160 -535
rect 29235 -545 29280 -535
rect 29360 -545 29400 -535
rect 29475 -545 29520 -535
rect 29600 -545 29640 -535
rect 29715 -545 29760 -535
rect 29840 -545 29880 -535
rect 29955 -545 30000 -535
rect 30080 -545 30120 -535
rect 30195 -545 30240 -535
rect 30320 -545 30360 -535
rect 30435 -545 30480 -535
rect 30560 -545 30600 -535
rect 30675 -545 30715 -535
rect -40 -565 -30 -545
rect -10 -560 90 -545
rect -10 -565 0 -560
rect -40 -575 0 -565
rect 80 -565 90 -560
rect 110 -560 210 -545
rect 110 -565 120 -560
rect 80 -575 120 -565
rect 195 -565 210 -560
rect 230 -560 330 -545
rect 230 -565 240 -560
rect 195 -575 240 -565
rect 320 -565 330 -560
rect 350 -560 450 -545
rect 350 -565 360 -560
rect 320 -575 360 -565
rect 435 -565 450 -560
rect 470 -560 570 -545
rect 470 -565 480 -560
rect 435 -575 480 -565
rect 560 -565 570 -560
rect 590 -560 690 -545
rect 590 -565 600 -560
rect 560 -575 600 -565
rect 675 -565 690 -560
rect 710 -560 810 -545
rect 710 -565 720 -560
rect 675 -575 720 -565
rect 800 -565 810 -560
rect 830 -560 930 -545
rect 830 -565 840 -560
rect 800 -575 840 -565
rect 915 -565 930 -560
rect 950 -560 1050 -545
rect 950 -565 960 -560
rect 915 -575 960 -565
rect 1040 -565 1050 -560
rect 1070 -560 1170 -545
rect 1070 -565 1080 -560
rect 1040 -575 1080 -565
rect 1155 -565 1170 -560
rect 1190 -560 1290 -545
rect 1190 -565 1200 -560
rect 1155 -575 1200 -565
rect 1280 -565 1290 -560
rect 1310 -560 1410 -545
rect 1310 -565 1320 -560
rect 1280 -575 1320 -565
rect 1395 -565 1410 -560
rect 1430 -560 1530 -545
rect 1430 -565 1440 -560
rect 1395 -575 1440 -565
rect 1520 -565 1530 -560
rect 1550 -560 1650 -545
rect 1550 -565 1560 -560
rect 1520 -575 1560 -565
rect 1635 -565 1650 -560
rect 1670 -560 1770 -545
rect 1670 -565 1680 -560
rect 1635 -575 1680 -565
rect 1760 -565 1770 -560
rect 1790 -560 1890 -545
rect 1790 -565 1800 -560
rect 1760 -575 1800 -565
rect 1875 -565 1890 -560
rect 1910 -560 2010 -545
rect 1910 -565 1920 -560
rect 1875 -575 1920 -565
rect 2000 -565 2010 -560
rect 2030 -560 2130 -545
rect 2030 -565 2040 -560
rect 2000 -575 2040 -565
rect 2115 -565 2130 -560
rect 2150 -560 2250 -545
rect 2150 -565 2160 -560
rect 2115 -575 2160 -565
rect 2240 -565 2250 -560
rect 2270 -560 2370 -545
rect 2270 -565 2280 -560
rect 2240 -575 2280 -565
rect 2355 -565 2370 -560
rect 2390 -560 2490 -545
rect 2390 -565 2400 -560
rect 2355 -575 2400 -565
rect 2480 -565 2490 -560
rect 2510 -560 2610 -545
rect 2510 -565 2520 -560
rect 2480 -575 2520 -565
rect 2595 -565 2610 -560
rect 2630 -560 2730 -545
rect 2630 -565 2640 -560
rect 2595 -575 2640 -565
rect 2720 -565 2730 -560
rect 2750 -560 2850 -545
rect 2750 -565 2760 -560
rect 2720 -575 2760 -565
rect 2835 -565 2850 -560
rect 2870 -560 2970 -545
rect 2870 -565 2880 -560
rect 2835 -575 2880 -565
rect 2960 -565 2970 -560
rect 2990 -560 3090 -545
rect 2990 -565 3000 -560
rect 2960 -575 3000 -565
rect 3075 -565 3090 -560
rect 3110 -560 3210 -545
rect 3110 -565 3120 -560
rect 3075 -575 3120 -565
rect 3200 -565 3210 -560
rect 3230 -560 3330 -545
rect 3230 -565 3240 -560
rect 3200 -575 3240 -565
rect 3315 -565 3330 -560
rect 3350 -560 3450 -545
rect 3350 -565 3360 -560
rect 3315 -575 3360 -565
rect 3440 -565 3450 -560
rect 3470 -560 3570 -545
rect 3470 -565 3480 -560
rect 3440 -575 3480 -565
rect 3555 -565 3570 -560
rect 3590 -560 3690 -545
rect 3590 -565 3600 -560
rect 3555 -575 3600 -565
rect 3680 -565 3690 -560
rect 3710 -560 3810 -545
rect 3710 -565 3720 -560
rect 3680 -575 3720 -565
rect 3795 -565 3810 -560
rect 3830 -560 3930 -545
rect 3830 -565 3840 -560
rect 3795 -575 3840 -565
rect 3920 -565 3930 -560
rect 3950 -560 4050 -545
rect 3950 -565 3960 -560
rect 3920 -575 3960 -565
rect 4035 -565 4050 -560
rect 4070 -560 4170 -545
rect 4070 -565 4080 -560
rect 4035 -575 4080 -565
rect 4160 -565 4170 -560
rect 4190 -560 4290 -545
rect 4190 -565 4200 -560
rect 4160 -575 4200 -565
rect 4275 -565 4290 -560
rect 4310 -560 4410 -545
rect 4310 -565 4320 -560
rect 4275 -575 4320 -565
rect 4400 -565 4410 -560
rect 4430 -560 4530 -545
rect 4430 -565 4440 -560
rect 4400 -575 4440 -565
rect 4515 -565 4530 -560
rect 4550 -560 4650 -545
rect 4550 -565 4560 -560
rect 4515 -575 4560 -565
rect 4640 -565 4650 -560
rect 4670 -560 4770 -545
rect 4670 -565 4680 -560
rect 4640 -575 4680 -565
rect 4755 -565 4770 -560
rect 4790 -560 4890 -545
rect 4790 -565 4800 -560
rect 4755 -575 4800 -565
rect 4880 -565 4890 -560
rect 4910 -560 5010 -545
rect 4910 -565 4920 -560
rect 4880 -575 4920 -565
rect 4995 -565 5010 -560
rect 5030 -560 5130 -545
rect 5030 -565 5040 -560
rect 4995 -575 5040 -565
rect 5120 -565 5130 -560
rect 5150 -560 5250 -545
rect 5150 -565 5160 -560
rect 5120 -575 5160 -565
rect 5235 -565 5250 -560
rect 5270 -560 5370 -545
rect 5270 -565 5280 -560
rect 5235 -575 5280 -565
rect 5360 -565 5370 -560
rect 5390 -560 5490 -545
rect 5390 -565 5400 -560
rect 5360 -575 5400 -565
rect 5475 -565 5490 -560
rect 5510 -560 5610 -545
rect 5510 -565 5520 -560
rect 5475 -575 5520 -565
rect 5600 -565 5610 -560
rect 5630 -560 5730 -545
rect 5630 -565 5640 -560
rect 5600 -575 5640 -565
rect 5715 -565 5730 -560
rect 5750 -560 5850 -545
rect 5750 -565 5760 -560
rect 5715 -575 5760 -565
rect 5840 -565 5850 -560
rect 5870 -560 5970 -545
rect 5870 -565 5880 -560
rect 5840 -575 5880 -565
rect 5955 -565 5970 -560
rect 5990 -560 6090 -545
rect 5990 -565 6000 -560
rect 5955 -575 6000 -565
rect 6080 -565 6090 -560
rect 6110 -560 6210 -545
rect 6110 -565 6120 -560
rect 6080 -575 6120 -565
rect 6195 -565 6210 -560
rect 6230 -560 6330 -545
rect 6230 -565 6240 -560
rect 6195 -575 6240 -565
rect 6320 -565 6330 -560
rect 6350 -560 6450 -545
rect 6350 -565 6360 -560
rect 6320 -575 6360 -565
rect 6435 -565 6450 -560
rect 6470 -560 6570 -545
rect 6470 -565 6480 -560
rect 6435 -575 6480 -565
rect 6560 -565 6570 -560
rect 6590 -560 6690 -545
rect 6590 -565 6600 -560
rect 6560 -575 6600 -565
rect 6675 -565 6690 -560
rect 6710 -560 6810 -545
rect 6710 -565 6720 -560
rect 6675 -575 6720 -565
rect 6800 -565 6810 -560
rect 6830 -560 6930 -545
rect 6830 -565 6840 -560
rect 6800 -575 6840 -565
rect 6915 -565 6930 -560
rect 6950 -560 7050 -545
rect 6950 -565 6960 -560
rect 6915 -575 6960 -565
rect 7040 -565 7050 -560
rect 7070 -560 7170 -545
rect 7070 -565 7080 -560
rect 7040 -575 7080 -565
rect 7155 -565 7170 -560
rect 7190 -560 7290 -545
rect 7190 -565 7200 -560
rect 7155 -575 7200 -565
rect 7280 -565 7290 -560
rect 7310 -560 7410 -545
rect 7310 -565 7320 -560
rect 7280 -575 7320 -565
rect 7395 -565 7410 -560
rect 7430 -560 7530 -545
rect 7430 -565 7440 -560
rect 7395 -575 7440 -565
rect 7520 -565 7530 -560
rect 7550 -560 7650 -545
rect 7550 -565 7560 -560
rect 7520 -575 7560 -565
rect 7635 -565 7650 -560
rect 7670 -560 7770 -545
rect 7670 -565 7680 -560
rect 7635 -575 7680 -565
rect 7760 -565 7770 -560
rect 7790 -560 7890 -545
rect 7790 -565 7800 -560
rect 7760 -575 7800 -565
rect 7875 -565 7890 -560
rect 7910 -560 8010 -545
rect 7910 -565 7920 -560
rect 7875 -575 7920 -565
rect 8000 -565 8010 -560
rect 8030 -560 8130 -545
rect 8030 -565 8040 -560
rect 8000 -575 8040 -565
rect 8115 -565 8130 -560
rect 8150 -560 8250 -545
rect 8150 -565 8160 -560
rect 8115 -575 8160 -565
rect 8240 -565 8250 -560
rect 8270 -560 8370 -545
rect 8270 -565 8280 -560
rect 8240 -575 8280 -565
rect 8355 -565 8370 -560
rect 8390 -560 8490 -545
rect 8390 -565 8400 -560
rect 8355 -575 8400 -565
rect 8480 -565 8490 -560
rect 8510 -560 8610 -545
rect 8510 -565 8520 -560
rect 8480 -575 8520 -565
rect 8595 -565 8610 -560
rect 8630 -560 8730 -545
rect 8630 -565 8640 -560
rect 8595 -575 8640 -565
rect 8720 -565 8730 -560
rect 8750 -560 8850 -545
rect 8750 -565 8760 -560
rect 8720 -575 8760 -565
rect 8835 -565 8850 -560
rect 8870 -560 8970 -545
rect 8870 -565 8880 -560
rect 8835 -575 8880 -565
rect 8960 -565 8970 -560
rect 8990 -560 9090 -545
rect 8990 -565 9000 -560
rect 8960 -575 9000 -565
rect 9075 -565 9090 -560
rect 9110 -560 9210 -545
rect 9110 -565 9120 -560
rect 9075 -575 9120 -565
rect 9200 -565 9210 -560
rect 9230 -560 9330 -545
rect 9230 -565 9240 -560
rect 9200 -575 9240 -565
rect 9315 -565 9330 -560
rect 9350 -560 9450 -545
rect 9350 -565 9360 -560
rect 9315 -575 9360 -565
rect 9440 -565 9450 -560
rect 9470 -560 9570 -545
rect 9470 -565 9480 -560
rect 9440 -575 9480 -565
rect 9555 -565 9570 -560
rect 9590 -560 9690 -545
rect 9590 -565 9600 -560
rect 9555 -575 9600 -565
rect 9680 -565 9690 -560
rect 9710 -560 9810 -545
rect 9710 -565 9720 -560
rect 9680 -575 9720 -565
rect 9795 -565 9810 -560
rect 9830 -560 9930 -545
rect 9830 -565 9840 -560
rect 9795 -575 9840 -565
rect 9920 -565 9930 -560
rect 9950 -560 10050 -545
rect 9950 -565 9960 -560
rect 9920 -575 9960 -565
rect 10035 -565 10050 -560
rect 10070 -560 10170 -545
rect 10070 -565 10080 -560
rect 10035 -575 10080 -565
rect 10160 -565 10170 -560
rect 10190 -560 10290 -545
rect 10190 -565 10200 -560
rect 10160 -575 10200 -565
rect 10275 -565 10290 -560
rect 10310 -560 10410 -545
rect 10310 -565 10320 -560
rect 10275 -575 10320 -565
rect 10400 -565 10410 -560
rect 10430 -560 10530 -545
rect 10430 -565 10440 -560
rect 10400 -575 10440 -565
rect 10515 -565 10530 -560
rect 10550 -560 10650 -545
rect 10550 -565 10560 -560
rect 10515 -575 10560 -565
rect 10640 -565 10650 -560
rect 10670 -560 10770 -545
rect 10670 -565 10680 -560
rect 10640 -575 10680 -565
rect 10755 -565 10770 -560
rect 10790 -560 10890 -545
rect 10790 -565 10800 -560
rect 10755 -575 10800 -565
rect 10880 -565 10890 -560
rect 10910 -560 11010 -545
rect 10910 -565 10920 -560
rect 10880 -575 10920 -565
rect 10995 -565 11010 -560
rect 11030 -560 11130 -545
rect 11030 -565 11040 -560
rect 10995 -575 11040 -565
rect 11120 -565 11130 -560
rect 11150 -560 11250 -545
rect 11150 -565 11160 -560
rect 11120 -575 11160 -565
rect 11235 -565 11250 -560
rect 11270 -560 11370 -545
rect 11270 -565 11280 -560
rect 11235 -575 11280 -565
rect 11360 -565 11370 -560
rect 11390 -560 11490 -545
rect 11390 -565 11400 -560
rect 11360 -575 11400 -565
rect 11475 -565 11490 -560
rect 11510 -560 11610 -545
rect 11510 -565 11520 -560
rect 11475 -575 11520 -565
rect 11600 -565 11610 -560
rect 11630 -560 11730 -545
rect 11630 -565 11640 -560
rect 11600 -575 11640 -565
rect 11715 -565 11730 -560
rect 11750 -560 11850 -545
rect 11750 -565 11760 -560
rect 11715 -575 11760 -565
rect 11840 -565 11850 -560
rect 11870 -560 11970 -545
rect 11870 -565 11880 -560
rect 11840 -575 11880 -565
rect 11955 -565 11970 -560
rect 11990 -560 12090 -545
rect 11990 -565 12000 -560
rect 11955 -575 12000 -565
rect 12080 -565 12090 -560
rect 12110 -560 12210 -545
rect 12110 -565 12120 -560
rect 12080 -575 12120 -565
rect 12195 -565 12210 -560
rect 12230 -560 12330 -545
rect 12230 -565 12240 -560
rect 12195 -575 12240 -565
rect 12320 -565 12330 -560
rect 12350 -560 12450 -545
rect 12350 -565 12360 -560
rect 12320 -575 12360 -565
rect 12435 -565 12450 -560
rect 12470 -560 12570 -545
rect 12470 -565 12480 -560
rect 12435 -575 12480 -565
rect 12560 -565 12570 -560
rect 12590 -560 12690 -545
rect 12590 -565 12600 -560
rect 12560 -575 12600 -565
rect 12675 -565 12690 -560
rect 12710 -560 12810 -545
rect 12710 -565 12720 -560
rect 12675 -575 12720 -565
rect 12800 -565 12810 -560
rect 12830 -560 12930 -545
rect 12830 -565 12840 -560
rect 12800 -575 12840 -565
rect 12915 -565 12930 -560
rect 12950 -560 13050 -545
rect 12950 -565 12960 -560
rect 12915 -575 12960 -565
rect 13040 -565 13050 -560
rect 13070 -560 13170 -545
rect 13070 -565 13080 -560
rect 13040 -575 13080 -565
rect 13155 -565 13170 -560
rect 13190 -560 13290 -545
rect 13190 -565 13200 -560
rect 13155 -575 13200 -565
rect 13280 -565 13290 -560
rect 13310 -560 13410 -545
rect 13310 -565 13320 -560
rect 13280 -575 13320 -565
rect 13395 -565 13410 -560
rect 13430 -560 13530 -545
rect 13430 -565 13440 -560
rect 13395 -575 13440 -565
rect 13520 -565 13530 -560
rect 13550 -560 13650 -545
rect 13550 -565 13560 -560
rect 13520 -575 13560 -565
rect 13635 -565 13650 -560
rect 13670 -560 13770 -545
rect 13670 -565 13680 -560
rect 13635 -575 13680 -565
rect 13760 -565 13770 -560
rect 13790 -560 13890 -545
rect 13790 -565 13800 -560
rect 13760 -575 13800 -565
rect 13875 -565 13890 -560
rect 13910 -560 14010 -545
rect 13910 -565 13920 -560
rect 13875 -575 13920 -565
rect 14000 -565 14010 -560
rect 14030 -560 14130 -545
rect 14030 -565 14040 -560
rect 14000 -575 14040 -565
rect 14115 -565 14130 -560
rect 14150 -560 14250 -545
rect 14150 -565 14160 -560
rect 14115 -575 14160 -565
rect 14240 -565 14250 -560
rect 14270 -560 14370 -545
rect 14270 -565 14280 -560
rect 14240 -575 14280 -565
rect 14355 -565 14370 -560
rect 14390 -560 14490 -545
rect 14390 -565 14400 -560
rect 14355 -575 14400 -565
rect 14480 -565 14490 -560
rect 14510 -560 14610 -545
rect 14510 -565 14520 -560
rect 14480 -575 14520 -565
rect 14595 -565 14610 -560
rect 14630 -560 14730 -545
rect 14630 -565 14640 -560
rect 14595 -575 14640 -565
rect 14720 -565 14730 -560
rect 14750 -560 14850 -545
rect 14750 -565 14760 -560
rect 14720 -575 14760 -565
rect 14835 -565 14850 -560
rect 14870 -560 14970 -545
rect 14870 -565 14880 -560
rect 14835 -575 14880 -565
rect 14960 -565 14970 -560
rect 14990 -560 15090 -545
rect 14990 -565 15000 -560
rect 14960 -575 15000 -565
rect 15075 -565 15090 -560
rect 15110 -560 15210 -545
rect 15110 -565 15120 -560
rect 15075 -575 15120 -565
rect 15200 -565 15210 -560
rect 15230 -560 15330 -545
rect 15230 -565 15240 -560
rect 15200 -575 15240 -565
rect 15315 -565 15330 -560
rect 15350 -560 15450 -545
rect 15350 -565 15360 -560
rect 15315 -575 15360 -565
rect 15440 -565 15450 -560
rect 15470 -560 15570 -545
rect 15470 -565 15480 -560
rect 15440 -575 15480 -565
rect 15555 -565 15570 -560
rect 15590 -560 15690 -545
rect 15590 -565 15600 -560
rect 15555 -575 15600 -565
rect 15680 -565 15690 -560
rect 15710 -560 15810 -545
rect 15710 -565 15720 -560
rect 15680 -575 15720 -565
rect 15795 -565 15810 -560
rect 15830 -560 15930 -545
rect 15830 -565 15840 -560
rect 15795 -575 15840 -565
rect 15920 -565 15930 -560
rect 15950 -560 16050 -545
rect 15950 -565 15960 -560
rect 15920 -575 15960 -565
rect 16035 -565 16050 -560
rect 16070 -560 16170 -545
rect 16070 -565 16080 -560
rect 16035 -575 16080 -565
rect 16160 -565 16170 -560
rect 16190 -560 16290 -545
rect 16190 -565 16200 -560
rect 16160 -575 16200 -565
rect 16275 -565 16290 -560
rect 16310 -560 16410 -545
rect 16310 -565 16320 -560
rect 16275 -575 16320 -565
rect 16400 -565 16410 -560
rect 16430 -560 16530 -545
rect 16430 -565 16440 -560
rect 16400 -575 16440 -565
rect 16515 -565 16530 -560
rect 16550 -560 16650 -545
rect 16550 -565 16560 -560
rect 16515 -575 16560 -565
rect 16640 -565 16650 -560
rect 16670 -560 16770 -545
rect 16670 -565 16680 -560
rect 16640 -575 16680 -565
rect 16755 -565 16770 -560
rect 16790 -560 16890 -545
rect 16790 -565 16800 -560
rect 16755 -575 16800 -565
rect 16880 -565 16890 -560
rect 16910 -560 17010 -545
rect 16910 -565 16920 -560
rect 16880 -575 16920 -565
rect 16995 -565 17010 -560
rect 17030 -560 17130 -545
rect 17030 -565 17040 -560
rect 16995 -575 17040 -565
rect 17120 -565 17130 -560
rect 17150 -560 17250 -545
rect 17150 -565 17160 -560
rect 17120 -575 17160 -565
rect 17235 -565 17250 -560
rect 17270 -560 17370 -545
rect 17270 -565 17280 -560
rect 17235 -575 17280 -565
rect 17360 -565 17370 -560
rect 17390 -560 17490 -545
rect 17390 -565 17400 -560
rect 17360 -575 17400 -565
rect 17475 -565 17490 -560
rect 17510 -560 17610 -545
rect 17510 -565 17520 -560
rect 17475 -575 17520 -565
rect 17600 -565 17610 -560
rect 17630 -560 17730 -545
rect 17630 -565 17640 -560
rect 17600 -575 17640 -565
rect 17715 -565 17730 -560
rect 17750 -560 17850 -545
rect 17750 -565 17760 -560
rect 17715 -575 17760 -565
rect 17840 -565 17850 -560
rect 17870 -560 17970 -545
rect 17870 -565 17880 -560
rect 17840 -575 17880 -565
rect 17955 -565 17970 -560
rect 17990 -560 18090 -545
rect 17990 -565 18000 -560
rect 17955 -575 18000 -565
rect 18080 -565 18090 -560
rect 18110 -560 18210 -545
rect 18110 -565 18120 -560
rect 18080 -575 18120 -565
rect 18195 -565 18210 -560
rect 18230 -560 18330 -545
rect 18230 -565 18240 -560
rect 18195 -575 18240 -565
rect 18320 -565 18330 -560
rect 18350 -560 18450 -545
rect 18350 -565 18360 -560
rect 18320 -575 18360 -565
rect 18435 -565 18450 -560
rect 18470 -560 18570 -545
rect 18470 -565 18480 -560
rect 18435 -575 18480 -565
rect 18560 -565 18570 -560
rect 18590 -560 18690 -545
rect 18590 -565 18600 -560
rect 18560 -575 18600 -565
rect 18675 -565 18690 -560
rect 18710 -560 18810 -545
rect 18710 -565 18720 -560
rect 18675 -575 18720 -565
rect 18800 -565 18810 -560
rect 18830 -560 18930 -545
rect 18830 -565 18840 -560
rect 18800 -575 18840 -565
rect 18915 -565 18930 -560
rect 18950 -560 19050 -545
rect 18950 -565 18960 -560
rect 18915 -575 18960 -565
rect 19040 -565 19050 -560
rect 19070 -560 19170 -545
rect 19070 -565 19080 -560
rect 19040 -575 19080 -565
rect 19155 -565 19170 -560
rect 19190 -560 19290 -545
rect 19190 -565 19200 -560
rect 19155 -575 19200 -565
rect 19280 -565 19290 -560
rect 19310 -560 19410 -545
rect 19310 -565 19320 -560
rect 19280 -575 19320 -565
rect 19395 -565 19410 -560
rect 19430 -560 19530 -545
rect 19430 -565 19440 -560
rect 19395 -575 19440 -565
rect 19520 -565 19530 -560
rect 19550 -560 19650 -545
rect 19550 -565 19560 -560
rect 19520 -575 19560 -565
rect 19635 -565 19650 -560
rect 19670 -560 19770 -545
rect 19670 -565 19680 -560
rect 19635 -575 19680 -565
rect 19760 -565 19770 -560
rect 19790 -560 19890 -545
rect 19790 -565 19800 -560
rect 19760 -575 19800 -565
rect 19875 -565 19890 -560
rect 19910 -560 20010 -545
rect 19910 -565 19920 -560
rect 19875 -575 19920 -565
rect 20000 -565 20010 -560
rect 20030 -560 20130 -545
rect 20030 -565 20040 -560
rect 20000 -575 20040 -565
rect 20115 -565 20130 -560
rect 20150 -560 20250 -545
rect 20150 -565 20160 -560
rect 20115 -575 20160 -565
rect 20240 -565 20250 -560
rect 20270 -560 20370 -545
rect 20270 -565 20280 -560
rect 20240 -575 20280 -565
rect 20355 -565 20370 -560
rect 20390 -560 20490 -545
rect 20390 -565 20400 -560
rect 20355 -575 20400 -565
rect 20480 -565 20490 -560
rect 20510 -560 20610 -545
rect 20510 -565 20520 -560
rect 20480 -575 20520 -565
rect 20595 -565 20610 -560
rect 20630 -560 20730 -545
rect 20630 -565 20640 -560
rect 20595 -575 20640 -565
rect 20720 -565 20730 -560
rect 20750 -560 20850 -545
rect 20750 -565 20760 -560
rect 20720 -575 20760 -565
rect 20835 -565 20850 -560
rect 20870 -560 20970 -545
rect 20870 -565 20880 -560
rect 20835 -575 20880 -565
rect 20960 -565 20970 -560
rect 20990 -560 21090 -545
rect 20990 -565 21000 -560
rect 20960 -575 21000 -565
rect 21075 -565 21090 -560
rect 21110 -560 21210 -545
rect 21110 -565 21120 -560
rect 21075 -575 21120 -565
rect 21200 -565 21210 -560
rect 21230 -560 21330 -545
rect 21230 -565 21240 -560
rect 21200 -575 21240 -565
rect 21315 -565 21330 -560
rect 21350 -560 21450 -545
rect 21350 -565 21360 -560
rect 21315 -575 21360 -565
rect 21440 -565 21450 -560
rect 21470 -560 21570 -545
rect 21470 -565 21480 -560
rect 21440 -575 21480 -565
rect 21555 -565 21570 -560
rect 21590 -560 21690 -545
rect 21590 -565 21600 -560
rect 21555 -575 21600 -565
rect 21680 -565 21690 -560
rect 21710 -560 21810 -545
rect 21710 -565 21720 -560
rect 21680 -575 21720 -565
rect 21795 -565 21810 -560
rect 21830 -560 21930 -545
rect 21830 -565 21840 -560
rect 21795 -575 21840 -565
rect 21920 -565 21930 -560
rect 21950 -560 22050 -545
rect 21950 -565 21960 -560
rect 21920 -575 21960 -565
rect 22035 -565 22050 -560
rect 22070 -560 22170 -545
rect 22070 -565 22080 -560
rect 22035 -575 22080 -565
rect 22160 -565 22170 -560
rect 22190 -560 22290 -545
rect 22190 -565 22200 -560
rect 22160 -575 22200 -565
rect 22275 -565 22290 -560
rect 22310 -560 22410 -545
rect 22310 -565 22320 -560
rect 22275 -575 22320 -565
rect 22400 -565 22410 -560
rect 22430 -560 22530 -545
rect 22430 -565 22440 -560
rect 22400 -575 22440 -565
rect 22515 -565 22530 -560
rect 22550 -560 22650 -545
rect 22550 -565 22560 -560
rect 22515 -575 22560 -565
rect 22640 -565 22650 -560
rect 22670 -560 22770 -545
rect 22670 -565 22680 -560
rect 22640 -575 22680 -565
rect 22755 -565 22770 -560
rect 22790 -560 22890 -545
rect 22790 -565 22800 -560
rect 22755 -575 22800 -565
rect 22880 -565 22890 -560
rect 22910 -560 23010 -545
rect 22910 -565 22920 -560
rect 22880 -575 22920 -565
rect 22995 -565 23010 -560
rect 23030 -560 23130 -545
rect 23030 -565 23040 -560
rect 22995 -575 23040 -565
rect 23120 -565 23130 -560
rect 23150 -560 23250 -545
rect 23150 -565 23160 -560
rect 23120 -575 23160 -565
rect 23235 -565 23250 -560
rect 23270 -560 23370 -545
rect 23270 -565 23280 -560
rect 23235 -575 23280 -565
rect 23360 -565 23370 -560
rect 23390 -560 23490 -545
rect 23390 -565 23400 -560
rect 23360 -575 23400 -565
rect 23475 -565 23490 -560
rect 23510 -560 23610 -545
rect 23510 -565 23520 -560
rect 23475 -575 23520 -565
rect 23600 -565 23610 -560
rect 23630 -560 23730 -545
rect 23630 -565 23640 -560
rect 23600 -575 23640 -565
rect 23715 -565 23730 -560
rect 23750 -560 23850 -545
rect 23750 -565 23760 -560
rect 23715 -575 23760 -565
rect 23840 -565 23850 -560
rect 23870 -560 23970 -545
rect 23870 -565 23880 -560
rect 23840 -575 23880 -565
rect 23955 -565 23970 -560
rect 23990 -560 24090 -545
rect 23990 -565 24000 -560
rect 23955 -575 24000 -565
rect 24080 -565 24090 -560
rect 24110 -560 24210 -545
rect 24110 -565 24120 -560
rect 24080 -575 24120 -565
rect 24195 -565 24210 -560
rect 24230 -560 24330 -545
rect 24230 -565 24240 -560
rect 24195 -575 24240 -565
rect 24320 -565 24330 -560
rect 24350 -560 24450 -545
rect 24350 -565 24360 -560
rect 24320 -575 24360 -565
rect 24435 -565 24450 -560
rect 24470 -560 24570 -545
rect 24470 -565 24480 -560
rect 24435 -575 24480 -565
rect 24560 -565 24570 -560
rect 24590 -560 24690 -545
rect 24590 -565 24600 -560
rect 24560 -575 24600 -565
rect 24675 -565 24690 -560
rect 24710 -560 24810 -545
rect 24710 -565 24720 -560
rect 24675 -575 24720 -565
rect 24800 -565 24810 -560
rect 24830 -560 24930 -545
rect 24830 -565 24840 -560
rect 24800 -575 24840 -565
rect 24915 -565 24930 -560
rect 24950 -560 25050 -545
rect 24950 -565 24960 -560
rect 24915 -575 24960 -565
rect 25040 -565 25050 -560
rect 25070 -560 25170 -545
rect 25070 -565 25080 -560
rect 25040 -575 25080 -565
rect 25155 -565 25170 -560
rect 25190 -560 25290 -545
rect 25190 -565 25200 -560
rect 25155 -575 25200 -565
rect 25280 -565 25290 -560
rect 25310 -560 25410 -545
rect 25310 -565 25320 -560
rect 25280 -575 25320 -565
rect 25395 -565 25410 -560
rect 25430 -560 25530 -545
rect 25430 -565 25440 -560
rect 25395 -575 25440 -565
rect 25520 -565 25530 -560
rect 25550 -560 25650 -545
rect 25550 -565 25560 -560
rect 25520 -575 25560 -565
rect 25635 -565 25650 -560
rect 25670 -560 25770 -545
rect 25670 -565 25680 -560
rect 25635 -575 25680 -565
rect 25760 -565 25770 -560
rect 25790 -560 25890 -545
rect 25790 -565 25800 -560
rect 25760 -575 25800 -565
rect 25875 -565 25890 -560
rect 25910 -560 26010 -545
rect 25910 -565 25920 -560
rect 25875 -575 25920 -565
rect 26000 -565 26010 -560
rect 26030 -560 26130 -545
rect 26030 -565 26040 -560
rect 26000 -575 26040 -565
rect 26115 -565 26130 -560
rect 26150 -560 26250 -545
rect 26150 -565 26160 -560
rect 26115 -575 26160 -565
rect 26240 -565 26250 -560
rect 26270 -560 26370 -545
rect 26270 -565 26280 -560
rect 26240 -575 26280 -565
rect 26355 -565 26370 -560
rect 26390 -560 26490 -545
rect 26390 -565 26400 -560
rect 26355 -575 26400 -565
rect 26480 -565 26490 -560
rect 26510 -560 26610 -545
rect 26510 -565 26520 -560
rect 26480 -575 26520 -565
rect 26595 -565 26610 -560
rect 26630 -560 26730 -545
rect 26630 -565 26640 -560
rect 26595 -575 26640 -565
rect 26720 -565 26730 -560
rect 26750 -560 26850 -545
rect 26750 -565 26760 -560
rect 26720 -575 26760 -565
rect 26835 -565 26850 -560
rect 26870 -560 26970 -545
rect 26870 -565 26880 -560
rect 26835 -575 26880 -565
rect 26960 -565 26970 -560
rect 26990 -560 27090 -545
rect 26990 -565 27000 -560
rect 26960 -575 27000 -565
rect 27075 -565 27090 -560
rect 27110 -560 27210 -545
rect 27110 -565 27120 -560
rect 27075 -575 27120 -565
rect 27200 -565 27210 -560
rect 27230 -560 27330 -545
rect 27230 -565 27240 -560
rect 27200 -575 27240 -565
rect 27315 -565 27330 -560
rect 27350 -560 27450 -545
rect 27350 -565 27360 -560
rect 27315 -575 27360 -565
rect 27440 -565 27450 -560
rect 27470 -560 27570 -545
rect 27470 -565 27480 -560
rect 27440 -575 27480 -565
rect 27555 -565 27570 -560
rect 27590 -560 27690 -545
rect 27590 -565 27600 -560
rect 27555 -575 27600 -565
rect 27680 -565 27690 -560
rect 27710 -560 27810 -545
rect 27710 -565 27720 -560
rect 27680 -575 27720 -565
rect 27795 -565 27810 -560
rect 27830 -560 27930 -545
rect 27830 -565 27840 -560
rect 27795 -575 27840 -565
rect 27920 -565 27930 -560
rect 27950 -560 28050 -545
rect 27950 -565 27960 -560
rect 27920 -575 27960 -565
rect 28035 -565 28050 -560
rect 28070 -560 28170 -545
rect 28070 -565 28080 -560
rect 28035 -575 28080 -565
rect 28160 -565 28170 -560
rect 28190 -560 28290 -545
rect 28190 -565 28200 -560
rect 28160 -575 28200 -565
rect 28275 -565 28290 -560
rect 28310 -560 28410 -545
rect 28310 -565 28320 -560
rect 28275 -575 28320 -565
rect 28400 -565 28410 -560
rect 28430 -560 28530 -545
rect 28430 -565 28440 -560
rect 28400 -575 28440 -565
rect 28515 -565 28530 -560
rect 28550 -560 28650 -545
rect 28550 -565 28560 -560
rect 28515 -575 28560 -565
rect 28640 -565 28650 -560
rect 28670 -560 28770 -545
rect 28670 -565 28680 -560
rect 28640 -575 28680 -565
rect 28755 -565 28770 -560
rect 28790 -560 28890 -545
rect 28790 -565 28800 -560
rect 28755 -575 28800 -565
rect 28880 -565 28890 -560
rect 28910 -560 29010 -545
rect 28910 -565 28920 -560
rect 28880 -575 28920 -565
rect 28995 -565 29010 -560
rect 29030 -560 29130 -545
rect 29030 -565 29040 -560
rect 28995 -575 29040 -565
rect 29120 -565 29130 -560
rect 29150 -560 29250 -545
rect 29150 -565 29160 -560
rect 29120 -575 29160 -565
rect 29235 -565 29250 -560
rect 29270 -560 29370 -545
rect 29270 -565 29280 -560
rect 29235 -575 29280 -565
rect 29360 -565 29370 -560
rect 29390 -560 29490 -545
rect 29390 -565 29400 -560
rect 29360 -575 29400 -565
rect 29475 -565 29490 -560
rect 29510 -560 29610 -545
rect 29510 -565 29520 -560
rect 29475 -575 29520 -565
rect 29600 -565 29610 -560
rect 29630 -560 29730 -545
rect 29630 -565 29640 -560
rect 29600 -575 29640 -565
rect 29715 -565 29730 -560
rect 29750 -560 29850 -545
rect 29750 -565 29760 -560
rect 29715 -575 29760 -565
rect 29840 -565 29850 -560
rect 29870 -560 29970 -545
rect 29870 -565 29880 -560
rect 29840 -575 29880 -565
rect 29955 -565 29970 -560
rect 29990 -560 30090 -545
rect 29990 -565 30000 -560
rect 29955 -575 30000 -565
rect 30080 -565 30090 -560
rect 30110 -560 30210 -545
rect 30110 -565 30120 -560
rect 30080 -575 30120 -565
rect 30195 -565 30210 -560
rect 30230 -560 30330 -545
rect 30230 -565 30240 -560
rect 30195 -575 30240 -565
rect 30320 -565 30330 -560
rect 30350 -560 30450 -545
rect 30350 -565 30360 -560
rect 30320 -575 30360 -565
rect 30435 -565 30450 -560
rect 30470 -560 30570 -545
rect 30470 -565 30480 -560
rect 30435 -575 30480 -565
rect 30560 -565 30570 -560
rect 30590 -560 30685 -545
rect 30590 -565 30600 -560
rect 30560 -575 30600 -565
rect 30675 -565 30685 -560
rect 30705 -565 30715 -545
rect 30675 -575 30715 -565
rect 15 -785 30655 -775
rect 15 -805 25 -785
rect 45 -790 145 -785
rect 45 -805 55 -790
rect 15 -815 55 -805
rect 135 -805 145 -790
rect 165 -790 265 -785
rect 165 -805 175 -790
rect 135 -815 175 -805
rect 255 -805 265 -790
rect 285 -790 385 -785
rect 285 -805 295 -790
rect 255 -815 295 -805
rect 375 -805 385 -790
rect 405 -790 505 -785
rect 405 -805 415 -790
rect 375 -815 415 -805
rect 495 -805 505 -790
rect 525 -790 625 -785
rect 525 -805 535 -790
rect 495 -815 535 -805
rect 615 -805 625 -790
rect 645 -790 745 -785
rect 645 -805 655 -790
rect 615 -815 655 -805
rect 735 -805 745 -790
rect 765 -790 865 -785
rect 765 -805 775 -790
rect 735 -815 775 -805
rect 855 -805 865 -790
rect 885 -790 985 -785
rect 885 -805 895 -790
rect 855 -815 895 -805
rect 975 -805 985 -790
rect 1005 -790 1105 -785
rect 1005 -805 1015 -790
rect 975 -815 1015 -805
rect 1095 -805 1105 -790
rect 1125 -790 1225 -785
rect 1125 -805 1135 -790
rect 1095 -815 1135 -805
rect 1215 -805 1225 -790
rect 1245 -790 1345 -785
rect 1245 -805 1255 -790
rect 1215 -815 1255 -805
rect 1335 -805 1345 -790
rect 1365 -790 1465 -785
rect 1365 -805 1375 -790
rect 1335 -815 1375 -805
rect 1455 -805 1465 -790
rect 1485 -790 1585 -785
rect 1485 -805 1495 -790
rect 1455 -815 1495 -805
rect 1575 -805 1585 -790
rect 1605 -790 1705 -785
rect 1605 -805 1615 -790
rect 1575 -815 1615 -805
rect 1695 -805 1705 -790
rect 1725 -790 1825 -785
rect 1725 -805 1735 -790
rect 1695 -815 1735 -805
rect 1815 -805 1825 -790
rect 1845 -790 1945 -785
rect 1845 -805 1855 -790
rect 1815 -815 1855 -805
rect 1935 -805 1945 -790
rect 1965 -790 2065 -785
rect 1965 -805 1975 -790
rect 1935 -815 1975 -805
rect 2055 -805 2065 -790
rect 2085 -790 2185 -785
rect 2085 -805 2095 -790
rect 2055 -815 2095 -805
rect 2175 -805 2185 -790
rect 2205 -790 2305 -785
rect 2205 -805 2215 -790
rect 2175 -815 2215 -805
rect 2295 -805 2305 -790
rect 2325 -790 2425 -785
rect 2325 -805 2335 -790
rect 2295 -815 2335 -805
rect 2415 -805 2425 -790
rect 2445 -790 2545 -785
rect 2445 -805 2455 -790
rect 2415 -815 2455 -805
rect 2535 -805 2545 -790
rect 2565 -790 2665 -785
rect 2565 -805 2575 -790
rect 2535 -815 2575 -805
rect 2655 -805 2665 -790
rect 2685 -790 2785 -785
rect 2685 -805 2695 -790
rect 2655 -815 2695 -805
rect 2775 -805 2785 -790
rect 2805 -790 2905 -785
rect 2805 -805 2815 -790
rect 2775 -815 2815 -805
rect 2895 -805 2905 -790
rect 2925 -790 3025 -785
rect 2925 -805 2935 -790
rect 2895 -815 2935 -805
rect 3015 -805 3025 -790
rect 3045 -790 3145 -785
rect 3045 -805 3055 -790
rect 3015 -815 3055 -805
rect 3135 -805 3145 -790
rect 3165 -790 3265 -785
rect 3165 -805 3175 -790
rect 3135 -815 3175 -805
rect 3255 -805 3265 -790
rect 3285 -790 3385 -785
rect 3285 -805 3295 -790
rect 3255 -815 3295 -805
rect 3375 -805 3385 -790
rect 3405 -790 3505 -785
rect 3405 -805 3415 -790
rect 3375 -815 3415 -805
rect 3495 -805 3505 -790
rect 3525 -790 3625 -785
rect 3525 -805 3535 -790
rect 3495 -815 3535 -805
rect 3615 -805 3625 -790
rect 3645 -790 3745 -785
rect 3645 -805 3655 -790
rect 3615 -815 3655 -805
rect 3735 -805 3745 -790
rect 3765 -790 3865 -785
rect 3765 -805 3775 -790
rect 3735 -815 3775 -805
rect 3855 -805 3865 -790
rect 3885 -790 3985 -785
rect 3885 -805 3895 -790
rect 3855 -815 3895 -805
rect 3975 -805 3985 -790
rect 4005 -790 4105 -785
rect 4005 -805 4015 -790
rect 3975 -815 4015 -805
rect 4095 -805 4105 -790
rect 4125 -790 4225 -785
rect 4125 -805 4135 -790
rect 4095 -815 4135 -805
rect 4215 -805 4225 -790
rect 4245 -790 4345 -785
rect 4245 -805 4255 -790
rect 4215 -815 4255 -805
rect 4335 -805 4345 -790
rect 4365 -790 4465 -785
rect 4365 -805 4375 -790
rect 4335 -815 4375 -805
rect 4455 -805 4465 -790
rect 4485 -790 4585 -785
rect 4485 -805 4495 -790
rect 4455 -815 4495 -805
rect 4575 -805 4585 -790
rect 4605 -790 4705 -785
rect 4605 -805 4615 -790
rect 4575 -815 4615 -805
rect 4695 -805 4705 -790
rect 4725 -790 4825 -785
rect 4725 -805 4735 -790
rect 4695 -815 4735 -805
rect 4815 -805 4825 -790
rect 4845 -790 4945 -785
rect 4845 -805 4855 -790
rect 4815 -815 4855 -805
rect 4935 -805 4945 -790
rect 4965 -790 5065 -785
rect 4965 -805 4975 -790
rect 4935 -815 4975 -805
rect 5055 -805 5065 -790
rect 5085 -790 5185 -785
rect 5085 -805 5095 -790
rect 5055 -815 5095 -805
rect 5175 -805 5185 -790
rect 5205 -790 5305 -785
rect 5205 -805 5215 -790
rect 5175 -815 5215 -805
rect 5295 -805 5305 -790
rect 5325 -790 5425 -785
rect 5325 -805 5335 -790
rect 5295 -815 5335 -805
rect 5415 -805 5425 -790
rect 5445 -790 5545 -785
rect 5445 -805 5455 -790
rect 5415 -815 5455 -805
rect 5535 -805 5545 -790
rect 5565 -790 5665 -785
rect 5565 -805 5575 -790
rect 5535 -815 5575 -805
rect 5655 -805 5665 -790
rect 5685 -790 5785 -785
rect 5685 -805 5695 -790
rect 5655 -815 5695 -805
rect 5775 -805 5785 -790
rect 5805 -790 5905 -785
rect 5805 -805 5815 -790
rect 5775 -815 5815 -805
rect 5895 -805 5905 -790
rect 5925 -790 6025 -785
rect 5925 -805 5935 -790
rect 5895 -815 5935 -805
rect 6015 -805 6025 -790
rect 6045 -790 6145 -785
rect 6045 -805 6055 -790
rect 6015 -815 6055 -805
rect 6135 -805 6145 -790
rect 6165 -790 6265 -785
rect 6165 -805 6175 -790
rect 6135 -815 6175 -805
rect 6255 -805 6265 -790
rect 6285 -790 6385 -785
rect 6285 -805 6295 -790
rect 6255 -815 6295 -805
rect 6375 -805 6385 -790
rect 6405 -790 6505 -785
rect 6405 -805 6415 -790
rect 6375 -815 6415 -805
rect 6495 -805 6505 -790
rect 6525 -790 6625 -785
rect 6525 -805 6535 -790
rect 6495 -815 6535 -805
rect 6615 -805 6625 -790
rect 6645 -790 6745 -785
rect 6645 -805 6655 -790
rect 6615 -815 6655 -805
rect 6735 -805 6745 -790
rect 6765 -790 6865 -785
rect 6765 -805 6775 -790
rect 6735 -815 6775 -805
rect 6855 -805 6865 -790
rect 6885 -790 6985 -785
rect 6885 -805 6895 -790
rect 6855 -815 6895 -805
rect 6975 -805 6985 -790
rect 7005 -790 7105 -785
rect 7005 -805 7015 -790
rect 6975 -815 7015 -805
rect 7095 -805 7105 -790
rect 7125 -790 7225 -785
rect 7125 -805 7135 -790
rect 7095 -815 7135 -805
rect 7215 -805 7225 -790
rect 7245 -790 7345 -785
rect 7245 -805 7255 -790
rect 7215 -815 7255 -805
rect 7335 -805 7345 -790
rect 7365 -790 7465 -785
rect 7365 -805 7375 -790
rect 7335 -815 7375 -805
rect 7455 -805 7465 -790
rect 7485 -790 7585 -785
rect 7485 -805 7495 -790
rect 7455 -815 7495 -805
rect 7575 -805 7585 -790
rect 7605 -790 7705 -785
rect 7605 -805 7615 -790
rect 7575 -815 7615 -805
rect 7695 -805 7705 -790
rect 7725 -790 7825 -785
rect 7725 -805 7735 -790
rect 7695 -815 7735 -805
rect 7815 -805 7825 -790
rect 7845 -790 7945 -785
rect 7845 -805 7855 -790
rect 7815 -815 7855 -805
rect 7935 -805 7945 -790
rect 7965 -790 8065 -785
rect 7965 -805 7975 -790
rect 7935 -815 7975 -805
rect 8055 -805 8065 -790
rect 8085 -790 8185 -785
rect 8085 -805 8095 -790
rect 8055 -815 8095 -805
rect 8175 -805 8185 -790
rect 8205 -790 8305 -785
rect 8205 -805 8215 -790
rect 8175 -815 8215 -805
rect 8295 -805 8305 -790
rect 8325 -790 8425 -785
rect 8325 -805 8335 -790
rect 8295 -815 8335 -805
rect 8415 -805 8425 -790
rect 8445 -790 8545 -785
rect 8445 -805 8455 -790
rect 8415 -815 8455 -805
rect 8535 -805 8545 -790
rect 8565 -790 8665 -785
rect 8565 -805 8575 -790
rect 8535 -815 8575 -805
rect 8655 -805 8665 -790
rect 8685 -790 8785 -785
rect 8685 -805 8695 -790
rect 8655 -815 8695 -805
rect 8775 -805 8785 -790
rect 8805 -790 8905 -785
rect 8805 -805 8815 -790
rect 8775 -815 8815 -805
rect 8895 -805 8905 -790
rect 8925 -790 9025 -785
rect 8925 -805 8935 -790
rect 8895 -815 8935 -805
rect 9015 -805 9025 -790
rect 9045 -790 9145 -785
rect 9045 -805 9055 -790
rect 9015 -815 9055 -805
rect 9135 -805 9145 -790
rect 9165 -790 9265 -785
rect 9165 -805 9175 -790
rect 9135 -815 9175 -805
rect 9255 -805 9265 -790
rect 9285 -790 9385 -785
rect 9285 -805 9295 -790
rect 9255 -815 9295 -805
rect 9375 -805 9385 -790
rect 9405 -790 9505 -785
rect 9405 -805 9415 -790
rect 9375 -815 9415 -805
rect 9495 -805 9505 -790
rect 9525 -790 9625 -785
rect 9525 -805 9535 -790
rect 9495 -815 9535 -805
rect 9615 -805 9625 -790
rect 9645 -790 9745 -785
rect 9645 -805 9655 -790
rect 9615 -815 9655 -805
rect 9735 -805 9745 -790
rect 9765 -790 9865 -785
rect 9765 -805 9775 -790
rect 9735 -815 9775 -805
rect 9855 -805 9865 -790
rect 9885 -790 9985 -785
rect 9885 -805 9895 -790
rect 9855 -815 9895 -805
rect 9975 -805 9985 -790
rect 10005 -790 10105 -785
rect 10005 -805 10015 -790
rect 9975 -815 10015 -805
rect 10095 -805 10105 -790
rect 10125 -790 10225 -785
rect 10125 -805 10135 -790
rect 10095 -815 10135 -805
rect 10215 -805 10225 -790
rect 10245 -790 10345 -785
rect 10245 -805 10255 -790
rect 10215 -815 10255 -805
rect 10335 -805 10345 -790
rect 10365 -790 10465 -785
rect 10365 -805 10375 -790
rect 10335 -815 10375 -805
rect 10455 -805 10465 -790
rect 10485 -790 10585 -785
rect 10485 -805 10495 -790
rect 10455 -815 10495 -805
rect 10575 -805 10585 -790
rect 10605 -790 10705 -785
rect 10605 -805 10615 -790
rect 10575 -815 10615 -805
rect 10695 -805 10705 -790
rect 10725 -790 10825 -785
rect 10725 -805 10735 -790
rect 10695 -815 10735 -805
rect 10815 -805 10825 -790
rect 10845 -790 10945 -785
rect 10845 -805 10855 -790
rect 10815 -815 10855 -805
rect 10935 -805 10945 -790
rect 10965 -790 11065 -785
rect 10965 -805 10975 -790
rect 10935 -815 10975 -805
rect 11055 -805 11065 -790
rect 11085 -790 11185 -785
rect 11085 -805 11095 -790
rect 11055 -815 11095 -805
rect 11175 -805 11185 -790
rect 11205 -790 11305 -785
rect 11205 -805 11215 -790
rect 11175 -815 11215 -805
rect 11295 -805 11305 -790
rect 11325 -790 11425 -785
rect 11325 -805 11335 -790
rect 11295 -815 11335 -805
rect 11415 -805 11425 -790
rect 11445 -790 11545 -785
rect 11445 -805 11455 -790
rect 11415 -815 11455 -805
rect 11535 -805 11545 -790
rect 11565 -790 11665 -785
rect 11565 -805 11575 -790
rect 11535 -815 11575 -805
rect 11655 -805 11665 -790
rect 11685 -790 11785 -785
rect 11685 -805 11695 -790
rect 11655 -815 11695 -805
rect 11775 -805 11785 -790
rect 11805 -790 11905 -785
rect 11805 -805 11815 -790
rect 11775 -815 11815 -805
rect 11895 -805 11905 -790
rect 11925 -790 12025 -785
rect 11925 -805 11935 -790
rect 11895 -815 11935 -805
rect 12015 -805 12025 -790
rect 12045 -790 12145 -785
rect 12045 -805 12055 -790
rect 12015 -815 12055 -805
rect 12135 -805 12145 -790
rect 12165 -790 12265 -785
rect 12165 -805 12175 -790
rect 12135 -815 12175 -805
rect 12255 -805 12265 -790
rect 12285 -790 12385 -785
rect 12285 -805 12295 -790
rect 12255 -815 12295 -805
rect 12375 -805 12385 -790
rect 12405 -790 12505 -785
rect 12405 -805 12415 -790
rect 12375 -815 12415 -805
rect 12495 -805 12505 -790
rect 12525 -790 12625 -785
rect 12525 -805 12535 -790
rect 12495 -815 12535 -805
rect 12615 -805 12625 -790
rect 12645 -790 12745 -785
rect 12645 -805 12655 -790
rect 12615 -815 12655 -805
rect 12735 -805 12745 -790
rect 12765 -790 12865 -785
rect 12765 -805 12775 -790
rect 12735 -815 12775 -805
rect 12855 -805 12865 -790
rect 12885 -790 12985 -785
rect 12885 -805 12895 -790
rect 12855 -815 12895 -805
rect 12975 -805 12985 -790
rect 13005 -790 13105 -785
rect 13005 -805 13015 -790
rect 12975 -815 13015 -805
rect 13095 -805 13105 -790
rect 13125 -790 13225 -785
rect 13125 -805 13135 -790
rect 13095 -815 13135 -805
rect 13215 -805 13225 -790
rect 13245 -790 13345 -785
rect 13245 -805 13255 -790
rect 13215 -815 13255 -805
rect 13335 -805 13345 -790
rect 13365 -790 13465 -785
rect 13365 -805 13375 -790
rect 13335 -815 13375 -805
rect 13455 -805 13465 -790
rect 13485 -790 13585 -785
rect 13485 -805 13495 -790
rect 13455 -815 13495 -805
rect 13575 -805 13585 -790
rect 13605 -790 13705 -785
rect 13605 -805 13615 -790
rect 13575 -815 13615 -805
rect 13695 -805 13705 -790
rect 13725 -790 13825 -785
rect 13725 -805 13735 -790
rect 13695 -815 13735 -805
rect 13815 -805 13825 -790
rect 13845 -790 13945 -785
rect 13845 -805 13855 -790
rect 13815 -815 13855 -805
rect 13935 -805 13945 -790
rect 13965 -790 14065 -785
rect 13965 -805 13975 -790
rect 13935 -815 13975 -805
rect 14055 -805 14065 -790
rect 14085 -790 14185 -785
rect 14085 -805 14095 -790
rect 14055 -815 14095 -805
rect 14175 -805 14185 -790
rect 14205 -790 14305 -785
rect 14205 -805 14215 -790
rect 14175 -815 14215 -805
rect 14295 -805 14305 -790
rect 14325 -790 14425 -785
rect 14325 -805 14335 -790
rect 14295 -815 14335 -805
rect 14415 -805 14425 -790
rect 14445 -790 14545 -785
rect 14445 -805 14455 -790
rect 14415 -815 14455 -805
rect 14535 -805 14545 -790
rect 14565 -790 14665 -785
rect 14565 -805 14575 -790
rect 14535 -815 14575 -805
rect 14655 -805 14665 -790
rect 14685 -790 14785 -785
rect 14685 -805 14695 -790
rect 14655 -815 14695 -805
rect 14775 -805 14785 -790
rect 14805 -790 14905 -785
rect 14805 -805 14815 -790
rect 14775 -815 14815 -805
rect 14895 -805 14905 -790
rect 14925 -790 15025 -785
rect 14925 -805 14935 -790
rect 14895 -815 14935 -805
rect 15015 -805 15025 -790
rect 15045 -790 15145 -785
rect 15045 -805 15055 -790
rect 15015 -815 15055 -805
rect 15135 -805 15145 -790
rect 15165 -790 15265 -785
rect 15165 -805 15175 -790
rect 15135 -815 15175 -805
rect 15255 -805 15265 -790
rect 15285 -790 15385 -785
rect 15285 -805 15295 -790
rect 15255 -815 15295 -805
rect 15375 -805 15385 -790
rect 15405 -790 15505 -785
rect 15405 -805 15415 -790
rect 15375 -815 15415 -805
rect 15495 -805 15505 -790
rect 15525 -790 15625 -785
rect 15525 -805 15535 -790
rect 15495 -815 15535 -805
rect 15615 -805 15625 -790
rect 15645 -790 15745 -785
rect 15645 -805 15655 -790
rect 15615 -815 15655 -805
rect 15735 -805 15745 -790
rect 15765 -790 15865 -785
rect 15765 -805 15775 -790
rect 15735 -815 15775 -805
rect 15855 -805 15865 -790
rect 15885 -790 15985 -785
rect 15885 -805 15895 -790
rect 15855 -815 15895 -805
rect 15975 -805 15985 -790
rect 16005 -790 16105 -785
rect 16005 -805 16015 -790
rect 15975 -815 16015 -805
rect 16095 -805 16105 -790
rect 16125 -790 16225 -785
rect 16125 -805 16135 -790
rect 16095 -815 16135 -805
rect 16215 -805 16225 -790
rect 16245 -790 16345 -785
rect 16245 -805 16255 -790
rect 16215 -815 16255 -805
rect 16335 -805 16345 -790
rect 16365 -790 16465 -785
rect 16365 -805 16375 -790
rect 16335 -815 16375 -805
rect 16455 -805 16465 -790
rect 16485 -790 16585 -785
rect 16485 -805 16495 -790
rect 16455 -815 16495 -805
rect 16575 -805 16585 -790
rect 16605 -790 16705 -785
rect 16605 -805 16615 -790
rect 16575 -815 16615 -805
rect 16695 -805 16705 -790
rect 16725 -790 16825 -785
rect 16725 -805 16735 -790
rect 16695 -815 16735 -805
rect 16815 -805 16825 -790
rect 16845 -790 16945 -785
rect 16845 -805 16855 -790
rect 16815 -815 16855 -805
rect 16935 -805 16945 -790
rect 16965 -790 17065 -785
rect 16965 -805 16975 -790
rect 16935 -815 16975 -805
rect 17055 -805 17065 -790
rect 17085 -790 17185 -785
rect 17085 -805 17095 -790
rect 17055 -815 17095 -805
rect 17175 -805 17185 -790
rect 17205 -790 17305 -785
rect 17205 -805 17215 -790
rect 17175 -815 17215 -805
rect 17295 -805 17305 -790
rect 17325 -790 17425 -785
rect 17325 -805 17335 -790
rect 17295 -815 17335 -805
rect 17415 -805 17425 -790
rect 17445 -790 17545 -785
rect 17445 -805 17455 -790
rect 17415 -815 17455 -805
rect 17535 -805 17545 -790
rect 17565 -790 17665 -785
rect 17565 -805 17575 -790
rect 17535 -815 17575 -805
rect 17655 -805 17665 -790
rect 17685 -790 17785 -785
rect 17685 -805 17695 -790
rect 17655 -815 17695 -805
rect 17775 -805 17785 -790
rect 17805 -790 17905 -785
rect 17805 -805 17815 -790
rect 17775 -815 17815 -805
rect 17895 -805 17905 -790
rect 17925 -790 18025 -785
rect 17925 -805 17935 -790
rect 17895 -815 17935 -805
rect 18015 -805 18025 -790
rect 18045 -790 18145 -785
rect 18045 -805 18055 -790
rect 18015 -815 18055 -805
rect 18135 -805 18145 -790
rect 18165 -790 18265 -785
rect 18165 -805 18175 -790
rect 18135 -815 18175 -805
rect 18255 -805 18265 -790
rect 18285 -790 18385 -785
rect 18285 -805 18295 -790
rect 18255 -815 18295 -805
rect 18375 -805 18385 -790
rect 18405 -790 18505 -785
rect 18405 -805 18415 -790
rect 18375 -815 18415 -805
rect 18495 -805 18505 -790
rect 18525 -790 18625 -785
rect 18525 -805 18535 -790
rect 18495 -815 18535 -805
rect 18615 -805 18625 -790
rect 18645 -790 18745 -785
rect 18645 -805 18655 -790
rect 18615 -815 18655 -805
rect 18735 -805 18745 -790
rect 18765 -790 18865 -785
rect 18765 -805 18775 -790
rect 18735 -815 18775 -805
rect 18855 -805 18865 -790
rect 18885 -790 18985 -785
rect 18885 -805 18895 -790
rect 18855 -815 18895 -805
rect 18975 -805 18985 -790
rect 19005 -790 19105 -785
rect 19005 -805 19015 -790
rect 18975 -815 19015 -805
rect 19095 -805 19105 -790
rect 19125 -790 19225 -785
rect 19125 -805 19135 -790
rect 19095 -815 19135 -805
rect 19215 -805 19225 -790
rect 19245 -790 19345 -785
rect 19245 -805 19255 -790
rect 19215 -815 19255 -805
rect 19335 -805 19345 -790
rect 19365 -790 19465 -785
rect 19365 -805 19375 -790
rect 19335 -815 19375 -805
rect 19455 -805 19465 -790
rect 19485 -790 19585 -785
rect 19485 -805 19495 -790
rect 19455 -815 19495 -805
rect 19575 -805 19585 -790
rect 19605 -790 19705 -785
rect 19605 -805 19615 -790
rect 19575 -815 19615 -805
rect 19695 -805 19705 -790
rect 19725 -790 19825 -785
rect 19725 -805 19735 -790
rect 19695 -815 19735 -805
rect 19815 -805 19825 -790
rect 19845 -790 19945 -785
rect 19845 -805 19855 -790
rect 19815 -815 19855 -805
rect 19935 -805 19945 -790
rect 19965 -790 20065 -785
rect 19965 -805 19975 -790
rect 19935 -815 19975 -805
rect 20055 -805 20065 -790
rect 20085 -790 20185 -785
rect 20085 -805 20095 -790
rect 20055 -815 20095 -805
rect 20175 -805 20185 -790
rect 20205 -790 20305 -785
rect 20205 -805 20215 -790
rect 20175 -815 20215 -805
rect 20295 -805 20305 -790
rect 20325 -790 20425 -785
rect 20325 -805 20335 -790
rect 20295 -815 20335 -805
rect 20415 -805 20425 -790
rect 20445 -790 20545 -785
rect 20445 -805 20455 -790
rect 20415 -815 20455 -805
rect 20535 -805 20545 -790
rect 20565 -790 20665 -785
rect 20565 -805 20575 -790
rect 20535 -815 20575 -805
rect 20655 -805 20665 -790
rect 20685 -790 20785 -785
rect 20685 -805 20695 -790
rect 20655 -815 20695 -805
rect 20775 -805 20785 -790
rect 20805 -790 20905 -785
rect 20805 -805 20815 -790
rect 20775 -815 20815 -805
rect 20895 -805 20905 -790
rect 20925 -790 21025 -785
rect 20925 -805 20935 -790
rect 20895 -815 20935 -805
rect 21015 -805 21025 -790
rect 21045 -790 21145 -785
rect 21045 -805 21055 -790
rect 21015 -815 21055 -805
rect 21135 -805 21145 -790
rect 21165 -790 21265 -785
rect 21165 -805 21175 -790
rect 21135 -815 21175 -805
rect 21255 -805 21265 -790
rect 21285 -790 21385 -785
rect 21285 -805 21295 -790
rect 21255 -815 21295 -805
rect 21375 -805 21385 -790
rect 21405 -790 21505 -785
rect 21405 -805 21415 -790
rect 21375 -815 21415 -805
rect 21495 -805 21505 -790
rect 21525 -790 21625 -785
rect 21525 -805 21535 -790
rect 21495 -815 21535 -805
rect 21615 -805 21625 -790
rect 21645 -790 21745 -785
rect 21645 -805 21655 -790
rect 21615 -815 21655 -805
rect 21735 -805 21745 -790
rect 21765 -790 21865 -785
rect 21765 -805 21775 -790
rect 21735 -815 21775 -805
rect 21855 -805 21865 -790
rect 21885 -790 21985 -785
rect 21885 -805 21895 -790
rect 21855 -815 21895 -805
rect 21975 -805 21985 -790
rect 22005 -790 22105 -785
rect 22005 -805 22015 -790
rect 21975 -815 22015 -805
rect 22095 -805 22105 -790
rect 22125 -790 22225 -785
rect 22125 -805 22135 -790
rect 22095 -815 22135 -805
rect 22215 -805 22225 -790
rect 22245 -790 22345 -785
rect 22245 -805 22255 -790
rect 22215 -815 22255 -805
rect 22335 -805 22345 -790
rect 22365 -790 22465 -785
rect 22365 -805 22375 -790
rect 22335 -815 22375 -805
rect 22455 -805 22465 -790
rect 22485 -790 22585 -785
rect 22485 -805 22495 -790
rect 22455 -815 22495 -805
rect 22575 -805 22585 -790
rect 22605 -790 22705 -785
rect 22605 -805 22615 -790
rect 22575 -815 22615 -805
rect 22695 -805 22705 -790
rect 22725 -790 22825 -785
rect 22725 -805 22735 -790
rect 22695 -815 22735 -805
rect 22815 -805 22825 -790
rect 22845 -790 22945 -785
rect 22845 -805 22855 -790
rect 22815 -815 22855 -805
rect 22935 -805 22945 -790
rect 22965 -790 23065 -785
rect 22965 -805 22975 -790
rect 22935 -815 22975 -805
rect 23055 -805 23065 -790
rect 23085 -790 23185 -785
rect 23085 -805 23095 -790
rect 23055 -815 23095 -805
rect 23175 -805 23185 -790
rect 23205 -790 23305 -785
rect 23205 -805 23215 -790
rect 23175 -815 23215 -805
rect 23295 -805 23305 -790
rect 23325 -790 23425 -785
rect 23325 -805 23335 -790
rect 23295 -815 23335 -805
rect 23415 -805 23425 -790
rect 23445 -790 23545 -785
rect 23445 -805 23455 -790
rect 23415 -815 23455 -805
rect 23535 -805 23545 -790
rect 23565 -790 23665 -785
rect 23565 -805 23575 -790
rect 23535 -815 23575 -805
rect 23655 -805 23665 -790
rect 23685 -790 23785 -785
rect 23685 -805 23695 -790
rect 23655 -815 23695 -805
rect 23775 -805 23785 -790
rect 23805 -790 23905 -785
rect 23805 -805 23815 -790
rect 23775 -815 23815 -805
rect 23895 -805 23905 -790
rect 23925 -790 24025 -785
rect 23925 -805 23935 -790
rect 23895 -815 23935 -805
rect 24015 -805 24025 -790
rect 24045 -790 24145 -785
rect 24045 -805 24055 -790
rect 24015 -815 24055 -805
rect 24135 -805 24145 -790
rect 24165 -790 24265 -785
rect 24165 -805 24175 -790
rect 24135 -815 24175 -805
rect 24255 -805 24265 -790
rect 24285 -790 24385 -785
rect 24285 -805 24295 -790
rect 24255 -815 24295 -805
rect 24375 -805 24385 -790
rect 24405 -790 24505 -785
rect 24405 -805 24415 -790
rect 24375 -815 24415 -805
rect 24495 -805 24505 -790
rect 24525 -790 24625 -785
rect 24525 -805 24535 -790
rect 24495 -815 24535 -805
rect 24615 -805 24625 -790
rect 24645 -790 24745 -785
rect 24645 -805 24655 -790
rect 24615 -815 24655 -805
rect 24735 -805 24745 -790
rect 24765 -790 24865 -785
rect 24765 -805 24775 -790
rect 24735 -815 24775 -805
rect 24855 -805 24865 -790
rect 24885 -790 24985 -785
rect 24885 -805 24895 -790
rect 24855 -815 24895 -805
rect 24975 -805 24985 -790
rect 25005 -790 25105 -785
rect 25005 -805 25015 -790
rect 24975 -815 25015 -805
rect 25095 -805 25105 -790
rect 25125 -790 25225 -785
rect 25125 -805 25135 -790
rect 25095 -815 25135 -805
rect 25215 -805 25225 -790
rect 25245 -790 25345 -785
rect 25245 -805 25255 -790
rect 25215 -815 25255 -805
rect 25335 -805 25345 -790
rect 25365 -790 25465 -785
rect 25365 -805 25375 -790
rect 25335 -815 25375 -805
rect 25455 -805 25465 -790
rect 25485 -790 25585 -785
rect 25485 -805 25495 -790
rect 25455 -815 25495 -805
rect 25575 -805 25585 -790
rect 25605 -790 25705 -785
rect 25605 -805 25615 -790
rect 25575 -815 25615 -805
rect 25695 -805 25705 -790
rect 25725 -790 25825 -785
rect 25725 -805 25735 -790
rect 25695 -815 25735 -805
rect 25815 -805 25825 -790
rect 25845 -790 25945 -785
rect 25845 -805 25855 -790
rect 25815 -815 25855 -805
rect 25935 -805 25945 -790
rect 25965 -790 26065 -785
rect 25965 -805 25975 -790
rect 25935 -815 25975 -805
rect 26055 -805 26065 -790
rect 26085 -790 26185 -785
rect 26085 -805 26095 -790
rect 26055 -815 26095 -805
rect 26175 -805 26185 -790
rect 26205 -790 26305 -785
rect 26205 -805 26215 -790
rect 26175 -815 26215 -805
rect 26295 -805 26305 -790
rect 26325 -790 26425 -785
rect 26325 -805 26335 -790
rect 26295 -815 26335 -805
rect 26415 -805 26425 -790
rect 26445 -790 26545 -785
rect 26445 -805 26455 -790
rect 26415 -815 26455 -805
rect 26535 -805 26545 -790
rect 26565 -790 26665 -785
rect 26565 -805 26575 -790
rect 26535 -815 26575 -805
rect 26655 -805 26665 -790
rect 26685 -790 26785 -785
rect 26685 -805 26695 -790
rect 26655 -815 26695 -805
rect 26775 -805 26785 -790
rect 26805 -790 26905 -785
rect 26805 -805 26815 -790
rect 26775 -815 26815 -805
rect 26895 -805 26905 -790
rect 26925 -790 27025 -785
rect 26925 -805 26935 -790
rect 26895 -815 26935 -805
rect 27015 -805 27025 -790
rect 27045 -790 27145 -785
rect 27045 -805 27055 -790
rect 27015 -815 27055 -805
rect 27135 -805 27145 -790
rect 27165 -790 27265 -785
rect 27165 -805 27175 -790
rect 27135 -815 27175 -805
rect 27255 -805 27265 -790
rect 27285 -790 27385 -785
rect 27285 -805 27295 -790
rect 27255 -815 27295 -805
rect 27375 -805 27385 -790
rect 27405 -790 27505 -785
rect 27405 -805 27415 -790
rect 27375 -815 27415 -805
rect 27495 -805 27505 -790
rect 27525 -790 27625 -785
rect 27525 -805 27535 -790
rect 27495 -815 27535 -805
rect 27615 -805 27625 -790
rect 27645 -790 27745 -785
rect 27645 -805 27655 -790
rect 27615 -815 27655 -805
rect 27735 -805 27745 -790
rect 27765 -790 27865 -785
rect 27765 -805 27775 -790
rect 27735 -815 27775 -805
rect 27855 -805 27865 -790
rect 27885 -790 27985 -785
rect 27885 -805 27895 -790
rect 27855 -815 27895 -805
rect 27975 -805 27985 -790
rect 28005 -790 28105 -785
rect 28005 -805 28015 -790
rect 27975 -815 28015 -805
rect 28095 -805 28105 -790
rect 28125 -790 28225 -785
rect 28125 -805 28135 -790
rect 28095 -815 28135 -805
rect 28215 -805 28225 -790
rect 28245 -790 28345 -785
rect 28245 -805 28255 -790
rect 28215 -815 28255 -805
rect 28335 -805 28345 -790
rect 28365 -790 28465 -785
rect 28365 -805 28375 -790
rect 28335 -815 28375 -805
rect 28455 -805 28465 -790
rect 28485 -790 28585 -785
rect 28485 -805 28495 -790
rect 28455 -815 28495 -805
rect 28575 -805 28585 -790
rect 28605 -790 28705 -785
rect 28605 -805 28615 -790
rect 28575 -815 28615 -805
rect 28695 -805 28705 -790
rect 28725 -790 28825 -785
rect 28725 -805 28735 -790
rect 28695 -815 28735 -805
rect 28815 -805 28825 -790
rect 28845 -790 28945 -785
rect 28845 -805 28855 -790
rect 28815 -815 28855 -805
rect 28935 -805 28945 -790
rect 28965 -790 29065 -785
rect 28965 -805 28975 -790
rect 28935 -815 28975 -805
rect 29055 -805 29065 -790
rect 29085 -790 29185 -785
rect 29085 -805 29095 -790
rect 29055 -815 29095 -805
rect 29175 -805 29185 -790
rect 29205 -790 29305 -785
rect 29205 -805 29215 -790
rect 29175 -815 29215 -805
rect 29295 -805 29305 -790
rect 29325 -790 29425 -785
rect 29325 -805 29335 -790
rect 29295 -815 29335 -805
rect 29415 -805 29425 -790
rect 29445 -790 29545 -785
rect 29445 -805 29455 -790
rect 29415 -815 29455 -805
rect 29535 -805 29545 -790
rect 29565 -790 29665 -785
rect 29565 -805 29575 -790
rect 29535 -815 29575 -805
rect 29655 -805 29665 -790
rect 29685 -790 29785 -785
rect 29685 -805 29695 -790
rect 29655 -815 29695 -805
rect 29775 -805 29785 -790
rect 29805 -790 29905 -785
rect 29805 -805 29815 -790
rect 29775 -815 29815 -805
rect 29895 -805 29905 -790
rect 29925 -790 30025 -785
rect 29925 -805 29935 -790
rect 29895 -815 29935 -805
rect 30015 -805 30025 -790
rect 30045 -790 30145 -785
rect 30045 -805 30055 -790
rect 30015 -815 30055 -805
rect 30135 -805 30145 -790
rect 30165 -790 30265 -785
rect 30165 -805 30175 -790
rect 30135 -815 30175 -805
rect 30255 -805 30265 -790
rect 30285 -790 30385 -785
rect 30285 -805 30295 -790
rect 30255 -815 30295 -805
rect 30375 -805 30385 -790
rect 30405 -790 30505 -785
rect 30405 -805 30415 -790
rect 30375 -815 30415 -805
rect 30495 -805 30505 -790
rect 30525 -790 30625 -785
rect 30525 -805 30535 -790
rect 30495 -815 30535 -805
rect 30615 -805 30625 -790
rect 30645 -805 30655 -785
rect 30615 -815 30655 -805
rect 80 -820 120 -815
rect 80 -850 85 -820
rect 115 -850 120 -820
rect 80 -855 120 -850
rect 320 -820 360 -815
rect 320 -850 325 -820
rect 355 -850 360 -820
rect 320 -855 360 -850
rect 560 -820 600 -815
rect 560 -850 565 -820
rect 595 -850 600 -820
rect 1040 -820 1080 -815
rect 560 -855 600 -850
rect 790 -835 845 -825
rect 790 -870 800 -835
rect 835 -870 845 -835
rect 1040 -850 1045 -820
rect 1075 -850 1080 -820
rect 1040 -855 1080 -850
rect 1280 -820 1320 -815
rect 1280 -850 1285 -820
rect 1315 -850 1320 -820
rect 1280 -855 1320 -850
rect 1520 -820 1560 -815
rect 1520 -850 1525 -820
rect 1555 -850 1560 -820
rect 1520 -855 1560 -850
rect 1760 -820 1800 -815
rect 1760 -850 1765 -820
rect 1795 -850 1800 -820
rect 1760 -855 1800 -850
rect 2000 -820 2040 -815
rect 2000 -850 2005 -820
rect 2035 -850 2040 -820
rect 2000 -855 2040 -850
rect 2240 -820 2280 -815
rect 2240 -850 2245 -820
rect 2275 -850 2280 -820
rect 2240 -855 2280 -850
rect 2480 -820 2520 -815
rect 2480 -850 2485 -820
rect 2515 -850 2520 -820
rect 2480 -855 2520 -850
rect 2720 -820 2760 -815
rect 2720 -850 2725 -820
rect 2755 -850 2760 -820
rect 3200 -820 3240 -815
rect 2720 -855 2760 -850
rect 2950 -835 3005 -825
rect 790 -880 845 -870
rect 2950 -870 2960 -835
rect 2995 -870 3005 -835
rect 3200 -850 3205 -820
rect 3235 -850 3240 -820
rect 3200 -855 3240 -850
rect 3440 -820 3480 -815
rect 3440 -850 3445 -820
rect 3475 -850 3480 -820
rect 3440 -855 3480 -850
rect 3680 -820 3720 -815
rect 3680 -850 3685 -820
rect 3715 -850 3720 -820
rect 3680 -855 3720 -850
rect 3920 -820 3960 -815
rect 3920 -850 3925 -820
rect 3955 -850 3960 -820
rect 3920 -855 3960 -850
rect 4160 -820 4200 -815
rect 4160 -850 4165 -820
rect 4195 -850 4200 -820
rect 4160 -855 4200 -850
rect 4400 -820 4440 -815
rect 4400 -850 4405 -820
rect 4435 -850 4440 -820
rect 4400 -855 4440 -850
rect 4640 -820 4680 -815
rect 4640 -850 4645 -820
rect 4675 -850 4680 -820
rect 4640 -855 4680 -850
rect 4880 -820 4920 -815
rect 4880 -850 4885 -820
rect 4915 -850 4920 -820
rect 5360 -820 5400 -815
rect 4880 -855 4920 -850
rect 5110 -835 5165 -825
rect 2950 -880 3005 -870
rect 5110 -870 5120 -835
rect 5155 -870 5165 -835
rect 5360 -850 5365 -820
rect 5395 -850 5400 -820
rect 5360 -855 5400 -850
rect 5600 -820 5640 -815
rect 5600 -850 5605 -820
rect 5635 -850 5640 -820
rect 5600 -855 5640 -850
rect 5840 -820 5880 -815
rect 5840 -850 5845 -820
rect 5875 -850 5880 -820
rect 5840 -855 5880 -850
rect 6080 -820 6120 -815
rect 6080 -850 6085 -820
rect 6115 -850 6120 -820
rect 6080 -855 6120 -850
rect 6320 -820 6360 -815
rect 6320 -850 6325 -820
rect 6355 -850 6360 -820
rect 6320 -855 6360 -850
rect 6560 -820 6600 -815
rect 6560 -850 6565 -820
rect 6595 -850 6600 -820
rect 6560 -855 6600 -850
rect 6800 -820 6840 -815
rect 6800 -850 6805 -820
rect 6835 -850 6840 -820
rect 6800 -855 6840 -850
rect 7040 -820 7080 -815
rect 7040 -850 7045 -820
rect 7075 -850 7080 -820
rect 7520 -820 7560 -815
rect 7040 -855 7080 -850
rect 7270 -835 7325 -825
rect 5110 -880 5165 -870
rect 7270 -870 7280 -835
rect 7315 -870 7325 -835
rect 7520 -850 7525 -820
rect 7555 -850 7560 -820
rect 7520 -855 7560 -850
rect 7760 -820 7800 -815
rect 7760 -850 7765 -820
rect 7795 -850 7800 -820
rect 7760 -855 7800 -850
rect 8000 -820 8040 -815
rect 8000 -850 8005 -820
rect 8035 -850 8040 -820
rect 8000 -855 8040 -850
rect 8240 -820 8280 -815
rect 8240 -850 8245 -820
rect 8275 -850 8280 -820
rect 8240 -855 8280 -850
rect 8480 -820 8520 -815
rect 8480 -850 8485 -820
rect 8515 -850 8520 -820
rect 8480 -855 8520 -850
rect 8720 -820 8760 -815
rect 8720 -850 8725 -820
rect 8755 -850 8760 -820
rect 8720 -855 8760 -850
rect 8960 -820 9000 -815
rect 8960 -850 8965 -820
rect 8995 -850 9000 -820
rect 8960 -855 9000 -850
rect 9200 -820 9240 -815
rect 9200 -850 9205 -820
rect 9235 -850 9240 -820
rect 9680 -820 9720 -815
rect 9200 -855 9240 -850
rect 9430 -835 9485 -825
rect 7270 -880 7325 -870
rect 9430 -870 9440 -835
rect 9475 -870 9485 -835
rect 9680 -850 9685 -820
rect 9715 -850 9720 -820
rect 9680 -855 9720 -850
rect 9920 -820 9960 -815
rect 9920 -850 9925 -820
rect 9955 -850 9960 -820
rect 9920 -855 9960 -850
rect 10160 -820 10200 -815
rect 10160 -850 10165 -820
rect 10195 -850 10200 -820
rect 10160 -855 10200 -850
rect 10400 -820 10440 -815
rect 10400 -850 10405 -820
rect 10435 -850 10440 -820
rect 10400 -855 10440 -850
rect 10640 -820 10680 -815
rect 10640 -850 10645 -820
rect 10675 -850 10680 -820
rect 10640 -855 10680 -850
rect 10880 -820 10920 -815
rect 10880 -850 10885 -820
rect 10915 -850 10920 -820
rect 10880 -855 10920 -850
rect 11120 -820 11160 -815
rect 11120 -850 11125 -820
rect 11155 -850 11160 -820
rect 11120 -855 11160 -850
rect 11360 -820 11400 -815
rect 11360 -850 11365 -820
rect 11395 -850 11400 -820
rect 11840 -820 11880 -815
rect 11360 -855 11400 -850
rect 11590 -835 11645 -825
rect 9430 -880 9485 -870
rect 11590 -870 11600 -835
rect 11635 -870 11645 -835
rect 11840 -850 11845 -820
rect 11875 -850 11880 -820
rect 11840 -855 11880 -850
rect 12080 -820 12120 -815
rect 12080 -850 12085 -820
rect 12115 -850 12120 -820
rect 12080 -855 12120 -850
rect 12320 -820 12360 -815
rect 12320 -850 12325 -820
rect 12355 -850 12360 -820
rect 12320 -855 12360 -850
rect 12560 -820 12600 -815
rect 12560 -850 12565 -820
rect 12595 -850 12600 -820
rect 12560 -855 12600 -850
rect 12800 -820 12840 -815
rect 12800 -850 12805 -820
rect 12835 -850 12840 -820
rect 12800 -855 12840 -850
rect 13040 -820 13080 -815
rect 13040 -850 13045 -820
rect 13075 -850 13080 -820
rect 13040 -855 13080 -850
rect 13280 -820 13320 -815
rect 13280 -850 13285 -820
rect 13315 -850 13320 -820
rect 13280 -855 13320 -850
rect 13520 -820 13560 -815
rect 13520 -850 13525 -820
rect 13555 -850 13560 -820
rect 14000 -820 14040 -815
rect 13520 -855 13560 -850
rect 13750 -835 13805 -825
rect 11590 -880 11645 -870
rect 13750 -870 13760 -835
rect 13795 -870 13805 -835
rect 14000 -850 14005 -820
rect 14035 -850 14040 -820
rect 14000 -855 14040 -850
rect 14240 -820 14280 -815
rect 14240 -850 14245 -820
rect 14275 -850 14280 -820
rect 14240 -855 14280 -850
rect 14480 -820 14520 -815
rect 14480 -850 14485 -820
rect 14515 -850 14520 -820
rect 14480 -855 14520 -850
rect 14720 -820 14760 -815
rect 14720 -850 14725 -820
rect 14755 -850 14760 -820
rect 14720 -855 14760 -850
rect 14960 -820 15000 -815
rect 14960 -850 14965 -820
rect 14995 -850 15000 -820
rect 14960 -855 15000 -850
rect 15200 -820 15240 -815
rect 15200 -850 15205 -820
rect 15235 -850 15240 -820
rect 15200 -855 15240 -850
rect 15440 -820 15480 -815
rect 15440 -850 15445 -820
rect 15475 -850 15480 -820
rect 15440 -855 15480 -850
rect 15680 -820 15720 -815
rect 15680 -850 15685 -820
rect 15715 -850 15720 -820
rect 16160 -820 16200 -815
rect 15680 -855 15720 -850
rect 15910 -835 15965 -825
rect 13750 -880 13805 -870
rect 15910 -870 15920 -835
rect 15955 -870 15965 -835
rect 16160 -850 16165 -820
rect 16195 -850 16200 -820
rect 16160 -855 16200 -850
rect 16400 -820 16440 -815
rect 16400 -850 16405 -820
rect 16435 -850 16440 -820
rect 16400 -855 16440 -850
rect 16640 -820 16680 -815
rect 16640 -850 16645 -820
rect 16675 -850 16680 -820
rect 16640 -855 16680 -850
rect 16880 -820 16920 -815
rect 16880 -850 16885 -820
rect 16915 -850 16920 -820
rect 16880 -855 16920 -850
rect 17120 -820 17160 -815
rect 17120 -850 17125 -820
rect 17155 -850 17160 -820
rect 17120 -855 17160 -850
rect 17360 -820 17400 -815
rect 17360 -850 17365 -820
rect 17395 -850 17400 -820
rect 17360 -855 17400 -850
rect 17600 -820 17640 -815
rect 17600 -850 17605 -820
rect 17635 -850 17640 -820
rect 17600 -855 17640 -850
rect 17840 -820 17880 -815
rect 17840 -850 17845 -820
rect 17875 -850 17880 -820
rect 18320 -820 18360 -815
rect 17840 -855 17880 -850
rect 18070 -835 18125 -825
rect 15910 -880 15965 -870
rect 18070 -870 18080 -835
rect 18115 -870 18125 -835
rect 18320 -850 18325 -820
rect 18355 -850 18360 -820
rect 18320 -855 18360 -850
rect 18560 -820 18600 -815
rect 18560 -850 18565 -820
rect 18595 -850 18600 -820
rect 18560 -855 18600 -850
rect 18800 -820 18840 -815
rect 18800 -850 18805 -820
rect 18835 -850 18840 -820
rect 18800 -855 18840 -850
rect 19040 -820 19080 -815
rect 19040 -850 19045 -820
rect 19075 -850 19080 -820
rect 19040 -855 19080 -850
rect 19280 -820 19320 -815
rect 19280 -850 19285 -820
rect 19315 -850 19320 -820
rect 19280 -855 19320 -850
rect 19520 -820 19560 -815
rect 19520 -850 19525 -820
rect 19555 -850 19560 -820
rect 19520 -855 19560 -850
rect 19760 -820 19800 -815
rect 19760 -850 19765 -820
rect 19795 -850 19800 -820
rect 19760 -855 19800 -850
rect 20000 -820 20040 -815
rect 20000 -850 20005 -820
rect 20035 -850 20040 -820
rect 20480 -820 20520 -815
rect 20000 -855 20040 -850
rect 20230 -835 20285 -825
rect 18070 -880 18125 -870
rect 20230 -870 20240 -835
rect 20275 -870 20285 -835
rect 20480 -850 20485 -820
rect 20515 -850 20520 -820
rect 20480 -855 20520 -850
rect 20720 -820 20760 -815
rect 20720 -850 20725 -820
rect 20755 -850 20760 -820
rect 20720 -855 20760 -850
rect 20960 -820 21000 -815
rect 20960 -850 20965 -820
rect 20995 -850 21000 -820
rect 20960 -855 21000 -850
rect 21200 -820 21240 -815
rect 21200 -850 21205 -820
rect 21235 -850 21240 -820
rect 21200 -855 21240 -850
rect 21440 -820 21480 -815
rect 21440 -850 21445 -820
rect 21475 -850 21480 -820
rect 21440 -855 21480 -850
rect 21680 -820 21720 -815
rect 21680 -850 21685 -820
rect 21715 -850 21720 -820
rect 21680 -855 21720 -850
rect 21920 -820 21960 -815
rect 21920 -850 21925 -820
rect 21955 -850 21960 -820
rect 21920 -855 21960 -850
rect 22160 -820 22200 -815
rect 22160 -850 22165 -820
rect 22195 -850 22200 -820
rect 22640 -820 22680 -815
rect 22160 -855 22200 -850
rect 22390 -835 22445 -825
rect 20230 -880 20285 -870
rect 22390 -870 22400 -835
rect 22435 -870 22445 -835
rect 22640 -850 22645 -820
rect 22675 -850 22680 -820
rect 22640 -855 22680 -850
rect 22880 -820 22920 -815
rect 22880 -850 22885 -820
rect 22915 -850 22920 -820
rect 22880 -855 22920 -850
rect 23120 -820 23160 -815
rect 23120 -850 23125 -820
rect 23155 -850 23160 -820
rect 23120 -855 23160 -850
rect 23360 -820 23400 -815
rect 23360 -850 23365 -820
rect 23395 -850 23400 -820
rect 23360 -855 23400 -850
rect 23600 -820 23640 -815
rect 23600 -850 23605 -820
rect 23635 -850 23640 -820
rect 23600 -855 23640 -850
rect 23840 -820 23880 -815
rect 23840 -850 23845 -820
rect 23875 -850 23880 -820
rect 23840 -855 23880 -850
rect 24080 -820 24120 -815
rect 24080 -850 24085 -820
rect 24115 -850 24120 -820
rect 24560 -820 24600 -815
rect 24080 -855 24120 -850
rect 24310 -835 24365 -825
rect 22390 -880 22445 -870
rect 24310 -870 24320 -835
rect 24355 -870 24365 -835
rect 24560 -850 24565 -820
rect 24595 -850 24600 -820
rect 24560 -855 24600 -850
rect 24800 -820 24840 -815
rect 24800 -850 24805 -820
rect 24835 -850 24840 -820
rect 24800 -855 24840 -850
rect 25040 -820 25080 -815
rect 25040 -850 25045 -820
rect 25075 -850 25080 -820
rect 25040 -855 25080 -850
rect 25280 -820 25320 -815
rect 25280 -850 25285 -820
rect 25315 -850 25320 -820
rect 25280 -855 25320 -850
rect 25520 -820 25560 -815
rect 25520 -850 25525 -820
rect 25555 -850 25560 -820
rect 25520 -855 25560 -850
rect 25760 -820 25800 -815
rect 25760 -850 25765 -820
rect 25795 -850 25800 -820
rect 25760 -855 25800 -850
rect 26000 -820 26040 -815
rect 26000 -850 26005 -820
rect 26035 -850 26040 -820
rect 26480 -820 26520 -815
rect 26000 -855 26040 -850
rect 26230 -835 26285 -825
rect 24310 -880 24365 -870
rect 26230 -870 26240 -835
rect 26275 -870 26285 -835
rect 26480 -850 26485 -820
rect 26515 -850 26520 -820
rect 26480 -855 26520 -850
rect 26720 -820 26760 -815
rect 26720 -850 26725 -820
rect 26755 -850 26760 -820
rect 26720 -855 26760 -850
rect 26960 -820 27000 -815
rect 26960 -850 26965 -820
rect 26995 -850 27000 -820
rect 26960 -855 27000 -850
rect 27200 -820 27240 -815
rect 27200 -850 27205 -820
rect 27235 -850 27240 -820
rect 27200 -855 27240 -850
rect 27440 -820 27480 -815
rect 27440 -850 27445 -820
rect 27475 -850 27480 -820
rect 27440 -855 27480 -850
rect 27680 -820 27720 -815
rect 27680 -850 27685 -820
rect 27715 -850 27720 -820
rect 27680 -855 27720 -850
rect 27920 -820 27960 -815
rect 27920 -850 27925 -820
rect 27955 -850 27960 -820
rect 28400 -820 28440 -815
rect 27920 -855 27960 -850
rect 28150 -835 28205 -825
rect 26230 -880 26285 -870
rect 28150 -870 28160 -835
rect 28195 -870 28205 -835
rect 28400 -850 28405 -820
rect 28435 -850 28440 -820
rect 28400 -855 28440 -850
rect 28640 -820 28680 -815
rect 28640 -850 28645 -820
rect 28675 -850 28680 -820
rect 28640 -855 28680 -850
rect 28880 -820 28920 -815
rect 28880 -850 28885 -820
rect 28915 -850 28920 -820
rect 28880 -855 28920 -850
rect 29120 -820 29160 -815
rect 29120 -850 29125 -820
rect 29155 -850 29160 -820
rect 29120 -855 29160 -850
rect 29360 -820 29400 -815
rect 29360 -850 29365 -820
rect 29395 -850 29400 -820
rect 29360 -855 29400 -850
rect 29600 -820 29640 -815
rect 29600 -850 29605 -820
rect 29635 -850 29640 -820
rect 30080 -820 30120 -815
rect 29600 -855 29640 -850
rect 29830 -835 29885 -825
rect 28150 -880 28205 -870
rect 29830 -870 29840 -835
rect 29875 -870 29885 -835
rect 30080 -850 30085 -820
rect 30115 -850 30120 -820
rect 30080 -855 30120 -850
rect 30320 -820 30360 -815
rect 30320 -850 30325 -820
rect 30355 -850 30360 -820
rect 30320 -855 30360 -850
rect 30560 -820 30600 -815
rect 30560 -850 30565 -820
rect 30595 -850 30600 -820
rect 30560 -855 30600 -850
rect 29830 -880 29885 -870
<< via1 >>
rect 195 240 230 275
rect 2265 270 2300 305
rect 4205 270 4240 305
rect 6455 270 6490 305
rect 9360 270 9395 305
rect 11305 270 11340 305
rect 13000 270 13035 305
rect 15185 270 15220 305
rect 17365 270 17400 305
rect 19550 270 19585 305
rect 20760 270 20795 305
rect 436 260 466 265
rect 436 240 441 260
rect 441 240 461 260
rect 461 240 466 260
rect 436 235 466 240
rect 741 260 771 265
rect 741 240 746 260
rect 746 240 766 260
rect 766 240 771 260
rect 741 235 771 240
rect 986 260 1016 265
rect 986 240 991 260
rect 991 240 1011 260
rect 1011 240 1016 260
rect 986 235 1016 240
rect 1226 260 1256 265
rect 1226 240 1231 260
rect 1231 240 1251 260
rect 1251 240 1256 260
rect 1226 235 1256 240
rect 1471 260 1501 265
rect 1471 240 1476 260
rect 1476 240 1496 260
rect 1496 240 1501 260
rect 1471 235 1501 240
rect 1776 260 1806 265
rect 1776 240 1781 260
rect 1781 240 1801 260
rect 1801 240 1806 260
rect 1776 235 1806 240
rect 2021 260 2051 265
rect 2021 240 2026 260
rect 2026 240 2046 260
rect 2046 240 2051 260
rect 2021 235 2051 240
rect 2506 260 2536 265
rect 2506 240 2511 260
rect 2511 240 2531 260
rect 2531 240 2536 260
rect 2506 235 2536 240
rect 2746 260 2776 265
rect 2746 240 2751 260
rect 2751 240 2771 260
rect 2771 240 2776 260
rect 2746 235 2776 240
rect 2991 260 3021 265
rect 2991 240 2996 260
rect 2996 240 3016 260
rect 3016 240 3021 260
rect 2991 235 3021 240
rect 3231 260 3261 265
rect 3231 240 3236 260
rect 3236 240 3256 260
rect 3256 240 3261 260
rect 3231 235 3261 240
rect 3476 260 3506 265
rect 3476 240 3481 260
rect 3481 240 3501 260
rect 3501 240 3506 260
rect 3476 235 3506 240
rect 3716 260 3746 265
rect 3716 240 3721 260
rect 3721 240 3741 260
rect 3741 240 3746 260
rect 3716 235 3746 240
rect 3961 260 3991 265
rect 3961 240 3966 260
rect 3966 240 3986 260
rect 3986 240 3991 260
rect 3961 235 3991 240
rect 4446 260 4476 265
rect 4446 240 4451 260
rect 4451 240 4471 260
rect 4471 240 4476 260
rect 4446 235 4476 240
rect 4686 260 4716 265
rect 4686 240 4691 260
rect 4691 240 4711 260
rect 4711 240 4716 260
rect 4686 235 4716 240
rect 4931 260 4961 265
rect 4931 240 4936 260
rect 4936 240 4956 260
rect 4956 240 4961 260
rect 4931 235 4961 240
rect 5171 260 5201 265
rect 5171 240 5176 260
rect 5176 240 5196 260
rect 5196 240 5201 260
rect 5171 235 5201 240
rect 5416 260 5446 265
rect 5416 240 5421 260
rect 5421 240 5441 260
rect 5441 240 5446 260
rect 5416 235 5446 240
rect 5721 260 5751 265
rect 5721 240 5726 260
rect 5726 240 5746 260
rect 5746 240 5751 260
rect 5721 235 5751 240
rect 5966 260 5996 265
rect 5966 240 5971 260
rect 5971 240 5991 260
rect 5991 240 5996 260
rect 5966 235 5996 240
rect 6206 260 6236 265
rect 6206 240 6211 260
rect 6211 240 6231 260
rect 6231 240 6236 260
rect 6206 235 6236 240
rect 6691 260 6721 265
rect 6691 240 6696 260
rect 6696 240 6716 260
rect 6716 240 6721 260
rect 6691 235 6721 240
rect 6936 260 6966 265
rect 6936 240 6941 260
rect 6941 240 6961 260
rect 6961 240 6966 260
rect 6936 235 6966 240
rect 7176 260 7206 265
rect 7176 240 7181 260
rect 7181 240 7201 260
rect 7201 240 7206 260
rect 7176 235 7206 240
rect 7416 260 7446 265
rect 7416 240 7421 260
rect 7421 240 7441 260
rect 7441 240 7446 260
rect 7416 235 7446 240
rect 7656 260 7686 265
rect 7656 240 7661 260
rect 7661 240 7681 260
rect 7681 240 7686 260
rect 7656 235 7686 240
rect 7901 260 7931 265
rect 7901 240 7906 260
rect 7906 240 7926 260
rect 7926 240 7931 260
rect 7901 235 7931 240
rect 8141 260 8171 265
rect 8141 240 8146 260
rect 8146 240 8166 260
rect 8166 240 8171 260
rect 8141 235 8171 240
rect 8386 260 8416 265
rect 8386 240 8391 260
rect 8391 240 8411 260
rect 8411 240 8416 260
rect 8386 235 8416 240
rect 8626 260 8656 265
rect 8626 240 8631 260
rect 8631 240 8651 260
rect 8651 240 8656 260
rect 8626 235 8656 240
rect 8871 260 8901 265
rect 8871 240 8876 260
rect 8876 240 8896 260
rect 8896 240 8901 260
rect 8871 235 8901 240
rect 9111 260 9141 265
rect 9111 240 9116 260
rect 9116 240 9136 260
rect 9136 240 9141 260
rect 9111 235 9141 240
rect 9601 260 9631 265
rect 9601 240 9606 260
rect 9606 240 9626 260
rect 9626 240 9631 260
rect 9601 235 9631 240
rect 9846 260 9876 265
rect 9846 240 9851 260
rect 9851 240 9871 260
rect 9871 240 9876 260
rect 9846 235 9876 240
rect 10086 260 10116 265
rect 10086 240 10091 260
rect 10091 240 10111 260
rect 10111 240 10116 260
rect 10086 235 10116 240
rect 10331 260 10361 265
rect 10331 240 10336 260
rect 10336 240 10356 260
rect 10356 240 10361 260
rect 10331 235 10361 240
rect 10571 260 10601 265
rect 10571 240 10576 260
rect 10576 240 10596 260
rect 10596 240 10601 260
rect 10571 235 10601 240
rect 10816 260 10846 265
rect 10816 240 10821 260
rect 10821 240 10841 260
rect 10841 240 10846 260
rect 10816 235 10846 240
rect 11056 260 11086 265
rect 11056 240 11061 260
rect 11061 240 11081 260
rect 11081 240 11086 260
rect 11056 235 11086 240
rect 11541 260 11571 265
rect 11541 240 11546 260
rect 11546 240 11566 260
rect 11566 240 11571 260
rect 11541 235 11571 240
rect 11786 260 11816 265
rect 11786 240 11791 260
rect 11791 240 11811 260
rect 11811 240 11816 260
rect 11786 235 11816 240
rect 12026 260 12056 265
rect 12026 240 12031 260
rect 12031 240 12051 260
rect 12051 240 12056 260
rect 12026 235 12056 240
rect 12271 260 12301 265
rect 12271 240 12276 260
rect 12276 240 12296 260
rect 12296 240 12301 260
rect 12271 235 12301 240
rect 12511 260 12541 265
rect 12511 240 12516 260
rect 12516 240 12536 260
rect 12536 240 12541 260
rect 12511 235 12541 240
rect 12756 260 12786 265
rect 12756 240 12761 260
rect 12761 240 12781 260
rect 12781 240 12786 260
rect 12756 235 12786 240
rect 13241 260 13271 265
rect 13241 240 13246 260
rect 13246 240 13266 260
rect 13266 240 13271 260
rect 13241 235 13271 240
rect 13481 260 13511 265
rect 13481 240 13486 260
rect 13486 240 13506 260
rect 13506 240 13511 260
rect 13481 235 13511 240
rect 13726 260 13756 265
rect 13726 240 13731 260
rect 13731 240 13751 260
rect 13751 240 13756 260
rect 13726 235 13756 240
rect 13966 260 13996 265
rect 13966 240 13971 260
rect 13971 240 13991 260
rect 13991 240 13996 260
rect 13966 235 13996 240
rect 14211 260 14241 265
rect 14211 240 14216 260
rect 14216 240 14236 260
rect 14236 240 14241 260
rect 14211 235 14241 240
rect 14451 260 14481 265
rect 14451 240 14456 260
rect 14456 240 14476 260
rect 14476 240 14481 260
rect 14451 235 14481 240
rect 14696 260 14726 265
rect 14696 240 14701 260
rect 14701 240 14721 260
rect 14721 240 14726 260
rect 14696 235 14726 240
rect 14936 260 14966 265
rect 14936 240 14941 260
rect 14941 240 14961 260
rect 14961 240 14966 260
rect 14936 235 14966 240
rect 15421 260 15451 265
rect 15421 240 15426 260
rect 15426 240 15446 260
rect 15446 240 15451 260
rect 15421 235 15451 240
rect 15666 260 15696 265
rect 15666 240 15671 260
rect 15671 240 15691 260
rect 15691 240 15696 260
rect 15666 235 15696 240
rect 15906 260 15936 265
rect 15906 240 15911 260
rect 15911 240 15931 260
rect 15931 240 15936 260
rect 15906 235 15936 240
rect 16151 260 16181 265
rect 16151 240 16156 260
rect 16156 240 16176 260
rect 16176 240 16181 260
rect 16151 235 16181 240
rect 16391 260 16421 265
rect 16391 240 16396 260
rect 16396 240 16416 260
rect 16416 240 16421 260
rect 16391 235 16421 240
rect 16636 260 16666 265
rect 16636 240 16641 260
rect 16641 240 16661 260
rect 16661 240 16666 260
rect 16636 235 16666 240
rect 16876 260 16906 265
rect 16876 240 16881 260
rect 16881 240 16901 260
rect 16901 240 16906 260
rect 16876 235 16906 240
rect 17121 260 17151 265
rect 17121 240 17126 260
rect 17126 240 17146 260
rect 17146 240 17151 260
rect 17121 235 17151 240
rect 17606 260 17636 265
rect 17606 240 17611 260
rect 17611 240 17631 260
rect 17631 240 17636 260
rect 17606 235 17636 240
rect 17846 260 17876 265
rect 17846 240 17851 260
rect 17851 240 17871 260
rect 17871 240 17876 260
rect 17846 235 17876 240
rect 18091 260 18121 265
rect 18091 240 18096 260
rect 18096 240 18116 260
rect 18116 240 18121 260
rect 18091 235 18121 240
rect 18331 260 18361 265
rect 18331 240 18336 260
rect 18336 240 18356 260
rect 18356 240 18361 260
rect 18331 235 18361 240
rect 18576 260 18606 265
rect 18576 240 18581 260
rect 18581 240 18601 260
rect 18601 240 18606 260
rect 18576 235 18606 240
rect 18816 260 18846 265
rect 18816 240 18821 260
rect 18821 240 18841 260
rect 18841 240 18846 260
rect 18816 235 18846 240
rect 19061 260 19091 265
rect 19061 240 19066 260
rect 19066 240 19086 260
rect 19086 240 19091 260
rect 19061 235 19091 240
rect 19301 260 19331 265
rect 19301 240 19306 260
rect 19306 240 19326 260
rect 19326 240 19331 260
rect 19301 235 19331 240
rect 19786 260 19816 265
rect 19786 240 19791 260
rect 19791 240 19811 260
rect 19811 240 19816 260
rect 19786 235 19816 240
rect 20031 260 20061 265
rect 20031 240 20036 260
rect 20036 240 20056 260
rect 20056 240 20061 260
rect 20031 235 20061 240
rect 20271 260 20301 265
rect 20271 240 20276 260
rect 20276 240 20296 260
rect 20296 240 20301 260
rect 20271 235 20301 240
rect 20516 260 20546 265
rect 20516 240 20521 260
rect 20521 240 20541 260
rect 20541 240 20546 260
rect 20516 235 20546 240
rect 21001 260 21031 265
rect 21001 240 21006 260
rect 21006 240 21026 260
rect 21026 240 21031 260
rect 21001 235 21031 240
rect 21155 10 21185 15
rect 21155 -10 21160 10
rect 21160 -10 21180 10
rect 21180 -10 21185 10
rect 21155 -15 21185 -10
rect -415 -240 -365 -190
rect 186 -170 216 -165
rect 186 -190 191 -170
rect 191 -190 211 -170
rect 211 -190 216 -170
rect 186 -195 216 -190
rect 431 -170 461 -165
rect 431 -190 436 -170
rect 436 -190 456 -170
rect 456 -190 461 -170
rect 431 -195 461 -190
rect 736 -170 766 -165
rect 736 -190 741 -170
rect 741 -190 761 -170
rect 761 -190 766 -170
rect 736 -195 766 -190
rect 981 -170 1011 -165
rect 981 -190 986 -170
rect 986 -190 1006 -170
rect 1006 -190 1011 -170
rect 981 -195 1011 -190
rect 1221 -170 1251 -165
rect 1221 -190 1226 -170
rect 1226 -190 1246 -170
rect 1246 -190 1251 -170
rect 1221 -195 1251 -190
rect 1466 -170 1496 -165
rect 1466 -190 1471 -170
rect 1471 -190 1491 -170
rect 1491 -190 1496 -170
rect 1466 -195 1496 -190
rect 1771 -170 1801 -165
rect 1771 -190 1776 -170
rect 1776 -190 1796 -170
rect 1796 -190 1801 -170
rect 1771 -195 1801 -190
rect 2016 -170 2046 -165
rect 2016 -190 2021 -170
rect 2021 -190 2041 -170
rect 2041 -190 2046 -170
rect 2016 -195 2046 -190
rect 2256 -170 2286 -165
rect 2256 -190 2261 -170
rect 2261 -190 2281 -170
rect 2281 -190 2286 -170
rect 2256 -195 2286 -190
rect 2501 -170 2531 -165
rect 2501 -190 2506 -170
rect 2506 -190 2526 -170
rect 2526 -190 2531 -170
rect 2501 -195 2531 -190
rect 2741 -170 2771 -165
rect 2741 -190 2746 -170
rect 2746 -190 2766 -170
rect 2766 -190 2771 -170
rect 2741 -195 2771 -190
rect 2986 -170 3016 -165
rect 2986 -190 2991 -170
rect 2991 -190 3011 -170
rect 3011 -190 3016 -170
rect 2986 -195 3016 -190
rect 3226 -170 3256 -165
rect 3226 -190 3231 -170
rect 3231 -190 3251 -170
rect 3251 -190 3256 -170
rect 3226 -195 3256 -190
rect 3471 -170 3501 -165
rect 3471 -190 3476 -170
rect 3476 -190 3496 -170
rect 3496 -190 3501 -170
rect 3471 -195 3501 -190
rect 3711 -170 3741 -165
rect 3711 -190 3716 -170
rect 3716 -190 3736 -170
rect 3736 -190 3741 -170
rect 3711 -195 3741 -190
rect 3956 -170 3986 -165
rect 3956 -190 3961 -170
rect 3961 -190 3981 -170
rect 3981 -190 3986 -170
rect 3956 -195 3986 -190
rect 1635 -240 1675 -200
rect 4060 -235 4100 -195
rect 4196 -170 4226 -165
rect 4196 -190 4201 -170
rect 4201 -190 4221 -170
rect 4221 -190 4226 -170
rect 4196 -195 4226 -190
rect 4441 -170 4471 -165
rect 4441 -190 4446 -170
rect 4446 -190 4466 -170
rect 4466 -190 4471 -170
rect 4441 -195 4471 -190
rect 4681 -170 4711 -165
rect 4681 -190 4686 -170
rect 4686 -190 4706 -170
rect 4706 -190 4711 -170
rect 4681 -195 4711 -190
rect 4926 -170 4956 -165
rect 4926 -190 4931 -170
rect 4931 -190 4951 -170
rect 4951 -190 4956 -170
rect 4926 -195 4956 -190
rect 5166 -170 5196 -165
rect 5166 -190 5171 -170
rect 5171 -190 5191 -170
rect 5191 -190 5196 -170
rect 5166 -195 5196 -190
rect 5411 -170 5441 -165
rect 5411 -190 5416 -170
rect 5416 -190 5436 -170
rect 5436 -190 5441 -170
rect 5411 -195 5441 -190
rect 5716 -170 5746 -165
rect 5716 -190 5721 -170
rect 5721 -190 5741 -170
rect 5741 -190 5746 -170
rect 5716 -195 5746 -190
rect 5961 -170 5991 -165
rect 5961 -190 5966 -170
rect 5966 -190 5986 -170
rect 5986 -190 5991 -170
rect 5961 -195 5991 -190
rect 6201 -170 6231 -165
rect 6201 -190 6206 -170
rect 6206 -190 6226 -170
rect 6226 -190 6231 -170
rect 6201 -195 6231 -190
rect 6686 -170 6716 -165
rect 6686 -190 6691 -170
rect 6691 -190 6711 -170
rect 6711 -190 6716 -170
rect 6686 -195 6716 -190
rect 6931 -170 6961 -165
rect 6931 -190 6936 -170
rect 6936 -190 6956 -170
rect 6956 -190 6961 -170
rect 6931 -195 6961 -190
rect 7171 -170 7201 -165
rect 7171 -190 7176 -170
rect 7176 -190 7196 -170
rect 7196 -190 7201 -170
rect 7171 -195 7201 -190
rect 7411 -170 7441 -165
rect 7411 -190 7416 -170
rect 7416 -190 7436 -170
rect 7436 -190 7441 -170
rect 7411 -195 7441 -190
rect 7651 -170 7681 -165
rect 7651 -190 7656 -170
rect 7656 -190 7676 -170
rect 7676 -190 7681 -170
rect 7651 -195 7681 -190
rect 8136 -170 8166 -165
rect 8136 -190 8141 -170
rect 8141 -190 8161 -170
rect 8161 -190 8166 -170
rect 8136 -195 8166 -190
rect 8381 -170 8411 -165
rect 8381 -190 8386 -170
rect 8386 -190 8406 -170
rect 8406 -190 8411 -170
rect 8381 -195 8411 -190
rect 8621 -170 8651 -165
rect 8621 -190 8626 -170
rect 8626 -190 8646 -170
rect 8646 -190 8651 -170
rect 8621 -195 8651 -190
rect 8866 -170 8896 -165
rect 8866 -190 8871 -170
rect 8871 -190 8891 -170
rect 8891 -190 8896 -170
rect 8866 -195 8896 -190
rect 9106 -170 9136 -165
rect 9106 -190 9111 -170
rect 9111 -190 9131 -170
rect 9131 -190 9136 -170
rect 9106 -195 9136 -190
rect 9351 -170 9381 -165
rect 9351 -190 9356 -170
rect 9356 -190 9376 -170
rect 9376 -190 9381 -170
rect 9351 -195 9381 -190
rect 9841 -170 9871 -165
rect 9841 -190 9846 -170
rect 9846 -190 9866 -170
rect 9866 -190 9871 -170
rect 9841 -195 9871 -190
rect 10081 -170 10111 -165
rect 10081 -190 10086 -170
rect 10086 -190 10106 -170
rect 10106 -190 10111 -170
rect 10081 -195 10111 -190
rect 10326 -170 10356 -165
rect 10326 -190 10331 -170
rect 10331 -190 10351 -170
rect 10351 -190 10356 -170
rect 10326 -195 10356 -190
rect 10566 -170 10596 -165
rect 10566 -190 10571 -170
rect 10571 -190 10591 -170
rect 10591 -190 10596 -170
rect 10566 -195 10596 -190
rect 10811 -170 10841 -165
rect 10811 -190 10816 -170
rect 10816 -190 10836 -170
rect 10836 -190 10841 -170
rect 10811 -195 10841 -190
rect 11051 -170 11081 -165
rect 11051 -190 11056 -170
rect 11056 -190 11076 -170
rect 11076 -190 11081 -170
rect 11051 -195 11081 -190
rect 11296 -170 11326 -165
rect 11296 -190 11301 -170
rect 11301 -190 11321 -170
rect 11321 -190 11326 -170
rect 11296 -195 11326 -190
rect 11536 -170 11566 -165
rect 11536 -190 11541 -170
rect 11541 -190 11561 -170
rect 11561 -190 11566 -170
rect 11536 -195 11566 -190
rect 11781 -170 11811 -165
rect 11781 -190 11786 -170
rect 11786 -190 11806 -170
rect 11806 -190 11811 -170
rect 11781 -195 11811 -190
rect 12266 -170 12296 -165
rect 12266 -190 12271 -170
rect 12271 -190 12291 -170
rect 12291 -190 12296 -170
rect 12266 -195 12296 -190
rect 12506 -170 12536 -165
rect 12506 -190 12511 -170
rect 12511 -190 12531 -170
rect 12531 -190 12536 -170
rect 12506 -195 12536 -190
rect 12751 -170 12781 -165
rect 12751 -190 12756 -170
rect 12756 -190 12776 -170
rect 12776 -190 12781 -170
rect 12751 -195 12781 -190
rect 12991 -170 13021 -165
rect 12991 -190 12996 -170
rect 12996 -190 13016 -170
rect 13016 -190 13021 -170
rect 12991 -195 13021 -190
rect 13236 -170 13266 -165
rect 13236 -190 13241 -170
rect 13241 -190 13261 -170
rect 13261 -190 13266 -170
rect 13236 -195 13266 -190
rect 13476 -170 13506 -165
rect 13476 -190 13481 -170
rect 13481 -190 13501 -170
rect 13501 -190 13506 -170
rect 13476 -195 13506 -190
rect 13721 -170 13751 -165
rect 13721 -190 13726 -170
rect 13726 -190 13746 -170
rect 13746 -190 13751 -170
rect 13721 -195 13751 -190
rect 14206 -170 14236 -165
rect 14206 -190 14211 -170
rect 14211 -190 14231 -170
rect 14231 -190 14236 -170
rect 14206 -195 14236 -190
rect 14446 -170 14476 -165
rect 14446 -190 14451 -170
rect 14451 -190 14471 -170
rect 14471 -190 14476 -170
rect 14446 -195 14476 -190
rect 14691 -170 14721 -165
rect 14691 -190 14696 -170
rect 14696 -190 14716 -170
rect 14716 -190 14721 -170
rect 14691 -195 14721 -190
rect 14931 -170 14961 -165
rect 14931 -190 14936 -170
rect 14936 -190 14956 -170
rect 14956 -190 14961 -170
rect 14931 -195 14961 -190
rect 15176 -170 15206 -165
rect 15176 -190 15181 -170
rect 15181 -190 15201 -170
rect 15201 -190 15206 -170
rect 15176 -195 15206 -190
rect 15416 -170 15446 -165
rect 15416 -190 15421 -170
rect 15421 -190 15441 -170
rect 15441 -190 15446 -170
rect 15416 -195 15446 -190
rect 15661 -170 15691 -165
rect 15661 -190 15666 -170
rect 15666 -190 15686 -170
rect 15686 -190 15691 -170
rect 15661 -195 15691 -190
rect 16146 -170 16176 -165
rect 16146 -190 16151 -170
rect 16151 -190 16171 -170
rect 16171 -190 16176 -170
rect 16146 -195 16176 -190
rect 16386 -170 16416 -165
rect 16386 -190 16391 -170
rect 16391 -190 16411 -170
rect 16411 -190 16416 -170
rect 16386 -195 16416 -190
rect 16631 -170 16661 -165
rect 16631 -190 16636 -170
rect 16636 -190 16656 -170
rect 16656 -190 16661 -170
rect 16631 -195 16661 -190
rect 16871 -170 16901 -165
rect 16871 -190 16876 -170
rect 16876 -190 16896 -170
rect 16896 -190 16901 -170
rect 16871 -195 16901 -190
rect 17116 -170 17146 -165
rect 17116 -190 17121 -170
rect 17121 -190 17141 -170
rect 17141 -190 17146 -170
rect 17116 -195 17146 -190
rect 17356 -170 17386 -165
rect 17356 -190 17361 -170
rect 17361 -190 17381 -170
rect 17381 -190 17386 -170
rect 17356 -195 17386 -190
rect 17601 -170 17631 -165
rect 17601 -190 17606 -170
rect 17606 -190 17626 -170
rect 17626 -190 17631 -170
rect 17601 -195 17631 -190
rect 17841 -170 17871 -165
rect 17841 -190 17846 -170
rect 17846 -190 17866 -170
rect 17866 -190 17871 -170
rect 17841 -195 17871 -190
rect 18086 -170 18116 -165
rect 18086 -190 18091 -170
rect 18091 -190 18111 -170
rect 18111 -190 18116 -170
rect 18086 -195 18116 -190
rect 18326 -170 18356 -165
rect 18326 -190 18331 -170
rect 18331 -190 18351 -170
rect 18351 -190 18356 -170
rect 18326 -195 18356 -190
rect 18571 -170 18601 -165
rect 18571 -190 18576 -170
rect 18576 -190 18596 -170
rect 18596 -190 18601 -170
rect 18571 -195 18601 -190
rect 18811 -170 18841 -165
rect 18811 -190 18816 -170
rect 18816 -190 18836 -170
rect 18836 -190 18841 -170
rect 18811 -195 18841 -190
rect 19056 -170 19086 -165
rect 19056 -190 19061 -170
rect 19061 -190 19081 -170
rect 19081 -190 19086 -170
rect 19056 -195 19086 -190
rect 19296 -170 19326 -165
rect 19296 -190 19301 -170
rect 19301 -190 19321 -170
rect 19321 -190 19326 -170
rect 19296 -195 19326 -190
rect 19541 -170 19571 -165
rect 19541 -190 19546 -170
rect 19546 -190 19566 -170
rect 19566 -190 19571 -170
rect 19541 -195 19571 -190
rect 19781 -170 19811 -165
rect 19781 -190 19786 -170
rect 19786 -190 19806 -170
rect 19806 -190 19811 -170
rect 19781 -195 19811 -190
rect 20026 -170 20056 -165
rect 20026 -190 20031 -170
rect 20031 -190 20051 -170
rect 20051 -190 20056 -170
rect 20026 -195 20056 -190
rect 20266 -170 20296 -165
rect 20266 -190 20271 -170
rect 20271 -190 20291 -170
rect 20291 -190 20296 -170
rect 20266 -195 20296 -190
rect 20511 -170 20541 -165
rect 20511 -190 20516 -170
rect 20516 -190 20536 -170
rect 20536 -190 20541 -170
rect 20511 -195 20541 -190
rect 20751 -170 20781 -165
rect 20751 -190 20756 -170
rect 20756 -190 20776 -170
rect 20776 -190 20781 -170
rect 20751 -195 20781 -190
rect 20996 -170 21026 -165
rect 20996 -190 21001 -170
rect 21001 -190 21021 -170
rect 21021 -190 21026 -170
rect 20996 -195 21026 -190
rect 90 -250 120 -245
rect 90 -270 95 -250
rect 95 -270 115 -250
rect 115 -270 120 -250
rect 90 -275 120 -270
rect 330 -250 360 -245
rect 330 -270 335 -250
rect 335 -270 355 -250
rect 355 -270 360 -250
rect 330 -275 360 -270
rect 570 -250 600 -245
rect 570 -270 575 -250
rect 575 -270 595 -250
rect 595 -270 600 -250
rect 570 -275 600 -270
rect 810 -250 840 -245
rect 810 -270 815 -250
rect 815 -270 835 -250
rect 835 -270 840 -250
rect 810 -275 840 -270
rect 1050 -250 1080 -245
rect 1050 -270 1055 -250
rect 1055 -270 1075 -250
rect 1075 -270 1080 -250
rect 1050 -275 1080 -270
rect 1290 -250 1320 -245
rect 1290 -270 1295 -250
rect 1295 -270 1315 -250
rect 1315 -270 1320 -250
rect 1290 -275 1320 -270
rect 1530 -250 1560 -245
rect 1530 -270 1535 -250
rect 1535 -270 1555 -250
rect 1555 -270 1560 -250
rect 1530 -275 1560 -270
rect 1770 -250 1800 -245
rect 1770 -270 1775 -250
rect 1775 -270 1795 -250
rect 1795 -270 1800 -250
rect 1770 -275 1800 -270
rect 2010 -250 2040 -245
rect 2010 -270 2015 -250
rect 2015 -270 2035 -250
rect 2035 -270 2040 -250
rect 2010 -275 2040 -270
rect 2250 -250 2280 -245
rect 2250 -270 2255 -250
rect 2255 -270 2275 -250
rect 2275 -270 2280 -250
rect 2250 -275 2280 -270
rect 2490 -250 2520 -245
rect 2490 -270 2495 -250
rect 2495 -270 2515 -250
rect 2515 -270 2520 -250
rect 2490 -275 2520 -270
rect 2730 -250 2760 -245
rect 2730 -270 2735 -250
rect 2735 -270 2755 -250
rect 2755 -270 2760 -250
rect 2730 -275 2760 -270
rect 2970 -250 3000 -245
rect 2970 -270 2975 -250
rect 2975 -270 2995 -250
rect 2995 -270 3000 -250
rect 2970 -275 3000 -270
rect 3210 -250 3240 -245
rect 3210 -270 3215 -250
rect 3215 -270 3235 -250
rect 3235 -270 3240 -250
rect 3210 -275 3240 -270
rect 3450 -250 3480 -245
rect 3450 -270 3455 -250
rect 3455 -270 3475 -250
rect 3475 -270 3480 -250
rect 3450 -275 3480 -270
rect 3690 -250 3720 -245
rect 3690 -270 3695 -250
rect 3695 -270 3715 -250
rect 3715 -270 3720 -250
rect 3690 -275 3720 -270
rect 3930 -250 3960 -245
rect 3930 -270 3935 -250
rect 3935 -270 3955 -250
rect 3955 -270 3960 -250
rect 3930 -275 3960 -270
rect 4170 -250 4200 -245
rect 4170 -270 4175 -250
rect 4175 -270 4195 -250
rect 4195 -270 4200 -250
rect 4170 -275 4200 -270
rect 4410 -250 4440 -245
rect 4410 -270 4415 -250
rect 4415 -270 4435 -250
rect 4435 -270 4440 -250
rect 4410 -275 4440 -270
rect 4650 -250 4680 -245
rect 4650 -270 4655 -250
rect 4655 -270 4675 -250
rect 4675 -270 4680 -250
rect 4650 -275 4680 -270
rect 4890 -250 4920 -245
rect 4890 -270 4895 -250
rect 4895 -270 4915 -250
rect 4915 -270 4920 -250
rect 4890 -275 4920 -270
rect 5130 -250 5160 -245
rect 5130 -270 5135 -250
rect 5135 -270 5155 -250
rect 5155 -270 5160 -250
rect 5130 -275 5160 -270
rect 5370 -250 5400 -245
rect 5370 -270 5375 -250
rect 5375 -270 5395 -250
rect 5395 -270 5400 -250
rect 5370 -275 5400 -270
rect 5610 -250 5640 -245
rect 5610 -270 5615 -250
rect 5615 -270 5635 -250
rect 5635 -270 5640 -250
rect 5610 -275 5640 -270
rect 5850 -250 5880 -245
rect 5850 -270 5855 -250
rect 5855 -270 5875 -250
rect 5875 -270 5880 -250
rect 5850 -275 5880 -270
rect 6090 -250 6120 -245
rect 6090 -270 6095 -250
rect 6095 -270 6115 -250
rect 6115 -270 6120 -250
rect 6090 -275 6120 -270
rect 6330 -250 6360 -245
rect 6330 -270 6335 -250
rect 6335 -270 6355 -250
rect 6355 -270 6360 -250
rect 6330 -275 6360 -270
rect 6455 -260 6495 -220
rect 6570 -250 6600 -245
rect 6570 -270 6575 -250
rect 6575 -270 6595 -250
rect 6595 -270 6600 -250
rect 6570 -275 6600 -270
rect 6810 -250 6840 -245
rect 6810 -270 6815 -250
rect 6815 -270 6835 -250
rect 6835 -270 6840 -250
rect 6810 -275 6840 -270
rect 7050 -250 7080 -245
rect 7050 -270 7055 -250
rect 7055 -270 7075 -250
rect 7075 -270 7080 -250
rect 7050 -275 7080 -270
rect 7290 -250 7320 -245
rect 7290 -270 7295 -250
rect 7295 -270 7315 -250
rect 7315 -270 7320 -250
rect 7290 -275 7320 -270
rect 7530 -250 7560 -245
rect 7530 -270 7535 -250
rect 7535 -270 7555 -250
rect 7555 -270 7560 -250
rect 7530 -275 7560 -270
rect 7770 -250 7800 -245
rect 7770 -270 7775 -250
rect 7775 -270 7795 -250
rect 7795 -270 7800 -250
rect 7770 -275 7800 -270
rect 7880 -260 7920 -220
rect 8010 -250 8040 -245
rect 8010 -270 8015 -250
rect 8015 -270 8035 -250
rect 8035 -270 8040 -250
rect 8010 -275 8040 -270
rect 8250 -250 8280 -245
rect 8250 -270 8255 -250
rect 8255 -270 8275 -250
rect 8275 -270 8280 -250
rect 8250 -275 8280 -270
rect 8490 -250 8520 -245
rect 8490 -270 8495 -250
rect 8495 -270 8515 -250
rect 8515 -270 8520 -250
rect 8490 -275 8520 -270
rect 8730 -250 8760 -245
rect 8730 -270 8735 -250
rect 8735 -270 8755 -250
rect 8755 -270 8760 -250
rect 8730 -275 8760 -270
rect 8970 -250 9000 -245
rect 8970 -270 8975 -250
rect 8975 -270 8995 -250
rect 8995 -270 9000 -250
rect 8970 -275 9000 -270
rect 9210 -250 9240 -245
rect 9210 -270 9215 -250
rect 9215 -270 9235 -250
rect 9235 -270 9240 -250
rect 9210 -275 9240 -270
rect 9450 -250 9480 -245
rect 9450 -270 9455 -250
rect 9455 -270 9475 -250
rect 9475 -270 9480 -250
rect 9450 -275 9480 -270
rect 9570 -250 9610 -210
rect 9690 -250 9720 -245
rect 9690 -270 9695 -250
rect 9695 -270 9715 -250
rect 9715 -270 9720 -250
rect 9690 -275 9720 -270
rect 9930 -250 9960 -245
rect 9930 -270 9935 -250
rect 9935 -270 9955 -250
rect 9955 -270 9960 -250
rect 9930 -275 9960 -270
rect 10170 -250 10200 -245
rect 10170 -270 10175 -250
rect 10175 -270 10195 -250
rect 10195 -270 10200 -250
rect 10170 -275 10200 -270
rect 10410 -250 10440 -245
rect 10410 -270 10415 -250
rect 10415 -270 10435 -250
rect 10435 -270 10440 -250
rect 10410 -275 10440 -270
rect 10650 -250 10680 -245
rect 10650 -270 10655 -250
rect 10655 -270 10675 -250
rect 10675 -270 10680 -250
rect 10650 -275 10680 -270
rect 10890 -250 10920 -245
rect 10890 -270 10895 -250
rect 10895 -270 10915 -250
rect 10915 -270 10920 -250
rect 10890 -275 10920 -270
rect 11130 -250 11160 -245
rect 11130 -270 11135 -250
rect 11135 -270 11155 -250
rect 11155 -270 11160 -250
rect 11130 -275 11160 -270
rect 11370 -250 11400 -245
rect 11370 -270 11375 -250
rect 11375 -270 11395 -250
rect 11395 -270 11400 -250
rect 11370 -275 11400 -270
rect 11610 -250 11640 -245
rect 11610 -270 11615 -250
rect 11615 -270 11635 -250
rect 11635 -270 11640 -250
rect 11610 -275 11640 -270
rect 11850 -250 11880 -245
rect 11850 -270 11855 -250
rect 11855 -270 11875 -250
rect 11875 -270 11880 -250
rect 11850 -275 11880 -270
rect 11950 -260 11990 -220
rect 12090 -250 12120 -245
rect 12090 -270 12095 -250
rect 12095 -270 12115 -250
rect 12115 -270 12120 -250
rect 12090 -275 12120 -270
rect 12330 -250 12360 -245
rect 12330 -270 12335 -250
rect 12335 -270 12355 -250
rect 12355 -270 12360 -250
rect 12330 -275 12360 -270
rect 12570 -250 12600 -245
rect 12570 -270 12575 -250
rect 12575 -270 12595 -250
rect 12595 -270 12600 -250
rect 12570 -275 12600 -270
rect 12810 -250 12840 -245
rect 12810 -270 12815 -250
rect 12815 -270 12835 -250
rect 12835 -270 12840 -250
rect 12810 -275 12840 -270
rect 13050 -250 13080 -245
rect 13050 -270 13055 -250
rect 13055 -270 13075 -250
rect 13075 -270 13080 -250
rect 13050 -275 13080 -270
rect 13290 -250 13320 -245
rect 13290 -270 13295 -250
rect 13295 -270 13315 -250
rect 13315 -270 13320 -250
rect 13290 -275 13320 -270
rect 13530 -250 13560 -245
rect 13530 -270 13535 -250
rect 13535 -270 13555 -250
rect 13555 -270 13560 -250
rect 13530 -275 13560 -270
rect 13770 -250 13800 -245
rect 13770 -270 13775 -250
rect 13775 -270 13795 -250
rect 13795 -270 13800 -250
rect 13770 -275 13800 -270
rect 13870 -260 13910 -220
rect 14010 -250 14040 -245
rect 14010 -270 14015 -250
rect 14015 -270 14035 -250
rect 14035 -270 14040 -250
rect 14010 -275 14040 -270
rect 14250 -250 14280 -245
rect 14250 -270 14255 -250
rect 14255 -270 14275 -250
rect 14275 -270 14280 -250
rect 14250 -275 14280 -270
rect 14490 -250 14520 -245
rect 14490 -270 14495 -250
rect 14495 -270 14515 -250
rect 14515 -270 14520 -250
rect 14490 -275 14520 -270
rect 14730 -250 14760 -245
rect 14730 -270 14735 -250
rect 14735 -270 14755 -250
rect 14755 -270 14760 -250
rect 14730 -275 14760 -270
rect 14970 -250 15000 -245
rect 14970 -270 14975 -250
rect 14975 -270 14995 -250
rect 14995 -270 15000 -250
rect 14970 -275 15000 -270
rect 15210 -250 15240 -245
rect 15210 -270 15215 -250
rect 15215 -270 15235 -250
rect 15235 -270 15240 -250
rect 15210 -275 15240 -270
rect 15450 -250 15480 -245
rect 15450 -270 15455 -250
rect 15455 -270 15475 -250
rect 15475 -270 15480 -250
rect 15450 -275 15480 -270
rect 15690 -250 15720 -245
rect 15690 -270 15695 -250
rect 15695 -270 15715 -250
rect 15715 -270 15720 -250
rect 15690 -275 15720 -270
rect 15815 -260 15855 -220
rect 15930 -250 15960 -245
rect 15930 -270 15935 -250
rect 15935 -270 15955 -250
rect 15955 -270 15960 -250
rect 15930 -275 15960 -270
rect 16170 -250 16200 -245
rect 16170 -270 16175 -250
rect 16175 -270 16195 -250
rect 16195 -270 16200 -250
rect 16170 -275 16200 -270
rect 16410 -250 16440 -245
rect 16410 -270 16415 -250
rect 16415 -270 16435 -250
rect 16435 -270 16440 -250
rect 16410 -275 16440 -270
rect 16650 -250 16680 -245
rect 16650 -270 16655 -250
rect 16655 -270 16675 -250
rect 16675 -270 16680 -250
rect 16650 -275 16680 -270
rect 16890 -250 16920 -245
rect 16890 -270 16895 -250
rect 16895 -270 16915 -250
rect 16915 -270 16920 -250
rect 16890 -275 16920 -270
rect 17130 -250 17160 -245
rect 17130 -270 17135 -250
rect 17135 -270 17155 -250
rect 17155 -270 17160 -250
rect 17130 -275 17160 -270
rect 17370 -250 17400 -245
rect 17370 -270 17375 -250
rect 17375 -270 17395 -250
rect 17395 -270 17400 -250
rect 17370 -275 17400 -270
rect 17610 -250 17640 -245
rect 17610 -270 17615 -250
rect 17615 -270 17635 -250
rect 17635 -270 17640 -250
rect 17610 -275 17640 -270
rect 17705 -250 17745 -210
rect 17850 -250 17880 -245
rect 17850 -270 17855 -250
rect 17855 -270 17875 -250
rect 17875 -270 17880 -250
rect 17850 -275 17880 -270
rect 18090 -250 18120 -245
rect 18090 -270 18095 -250
rect 18095 -270 18115 -250
rect 18115 -270 18120 -250
rect 18090 -275 18120 -270
rect 18330 -250 18360 -245
rect 18330 -270 18335 -250
rect 18335 -270 18355 -250
rect 18355 -270 18360 -250
rect 18330 -275 18360 -270
rect 18570 -250 18600 -245
rect 18570 -270 18575 -250
rect 18575 -270 18595 -250
rect 18595 -270 18600 -250
rect 18570 -275 18600 -270
rect 18810 -250 18840 -245
rect 18810 -270 18815 -250
rect 18815 -270 18835 -250
rect 18835 -270 18840 -250
rect 18810 -275 18840 -270
rect 19050 -250 19080 -245
rect 19050 -270 19055 -250
rect 19055 -270 19075 -250
rect 19075 -270 19080 -250
rect 19050 -275 19080 -270
rect 19290 -250 19320 -245
rect 19290 -270 19295 -250
rect 19295 -270 19315 -250
rect 19315 -270 19320 -250
rect 19290 -275 19320 -270
rect 19530 -250 19560 -245
rect 19530 -270 19535 -250
rect 19535 -270 19555 -250
rect 19555 -270 19560 -250
rect 19530 -275 19560 -270
rect 19645 -250 19685 -210
rect 19770 -250 19800 -245
rect 19770 -270 19775 -250
rect 19775 -270 19795 -250
rect 19795 -270 19800 -250
rect 19770 -275 19800 -270
rect 20010 -250 20040 -245
rect 20010 -270 20015 -250
rect 20015 -270 20035 -250
rect 20035 -270 20040 -250
rect 20010 -275 20040 -270
rect 20250 -250 20280 -245
rect 20250 -270 20255 -250
rect 20255 -270 20275 -250
rect 20275 -270 20280 -250
rect 20250 -275 20280 -270
rect 20490 -250 20520 -245
rect 20490 -270 20495 -250
rect 20495 -270 20515 -250
rect 20515 -270 20520 -250
rect 20490 -275 20520 -270
rect 20730 -250 20760 -245
rect 20730 -270 20735 -250
rect 20735 -270 20755 -250
rect 20755 -270 20760 -250
rect 20730 -275 20760 -270
rect 20970 -250 21000 -245
rect 20970 -270 20975 -250
rect 20975 -270 20995 -250
rect 20995 -270 21000 -250
rect 20970 -275 21000 -270
rect 21210 -250 21240 -245
rect 21210 -270 21215 -250
rect 21215 -270 21235 -250
rect 21235 -270 21240 -250
rect 21210 -275 21240 -270
rect 21450 -250 21480 -245
rect 21450 -270 21455 -250
rect 21455 -270 21475 -250
rect 21475 -270 21480 -250
rect 21450 -275 21480 -270
rect 21690 -250 21720 -245
rect 21690 -270 21695 -250
rect 21695 -270 21715 -250
rect 21715 -270 21720 -250
rect 21690 -275 21720 -270
rect 21930 -250 21960 -245
rect 21930 -270 21935 -250
rect 21935 -270 21955 -250
rect 21955 -270 21960 -250
rect 21930 -275 21960 -270
rect 22170 -250 22200 -245
rect 22170 -270 22175 -250
rect 22175 -270 22195 -250
rect 22195 -270 22200 -250
rect 22170 -275 22200 -270
rect 22410 -250 22440 -245
rect 22410 -270 22415 -250
rect 22415 -270 22435 -250
rect 22435 -270 22440 -250
rect 22410 -275 22440 -270
rect 22650 -250 22680 -245
rect 22650 -270 22655 -250
rect 22655 -270 22675 -250
rect 22675 -270 22680 -250
rect 22650 -275 22680 -270
rect 22890 -250 22920 -245
rect 22890 -270 22895 -250
rect 22895 -270 22915 -250
rect 22915 -270 22920 -250
rect 22890 -275 22920 -270
rect 23130 -250 23160 -245
rect 23130 -270 23135 -250
rect 23135 -270 23155 -250
rect 23155 -270 23160 -250
rect 23130 -275 23160 -270
rect 23370 -250 23400 -245
rect 23370 -270 23375 -250
rect 23375 -270 23395 -250
rect 23395 -270 23400 -250
rect 23370 -275 23400 -270
rect 23610 -250 23640 -245
rect 23610 -270 23615 -250
rect 23615 -270 23635 -250
rect 23635 -270 23640 -250
rect 23610 -275 23640 -270
rect 23850 -250 23880 -245
rect 23850 -270 23855 -250
rect 23855 -270 23875 -250
rect 23875 -270 23880 -250
rect 23850 -275 23880 -270
rect 24090 -250 24120 -245
rect 24090 -270 24095 -250
rect 24095 -270 24115 -250
rect 24115 -270 24120 -250
rect 24090 -275 24120 -270
rect 24330 -250 24360 -245
rect 24330 -270 24335 -250
rect 24335 -270 24355 -250
rect 24355 -270 24360 -250
rect 24330 -275 24360 -270
rect 24570 -250 24600 -245
rect 24570 -270 24575 -250
rect 24575 -270 24595 -250
rect 24595 -270 24600 -250
rect 24570 -275 24600 -270
rect 24810 -250 24840 -245
rect 24810 -270 24815 -250
rect 24815 -270 24835 -250
rect 24835 -270 24840 -250
rect 24810 -275 24840 -270
rect 25050 -250 25080 -245
rect 25050 -270 25055 -250
rect 25055 -270 25075 -250
rect 25075 -270 25080 -250
rect 25050 -275 25080 -270
rect 25290 -250 25320 -245
rect 25290 -270 25295 -250
rect 25295 -270 25315 -250
rect 25315 -270 25320 -250
rect 25290 -275 25320 -270
rect 25530 -250 25560 -245
rect 25530 -270 25535 -250
rect 25535 -270 25555 -250
rect 25555 -270 25560 -250
rect 25530 -275 25560 -270
rect 25770 -250 25800 -245
rect 25770 -270 25775 -250
rect 25775 -270 25795 -250
rect 25795 -270 25800 -250
rect 25770 -275 25800 -270
rect 26010 -250 26040 -245
rect 26010 -270 26015 -250
rect 26015 -270 26035 -250
rect 26035 -270 26040 -250
rect 26010 -275 26040 -270
rect 26250 -250 26280 -245
rect 26250 -270 26255 -250
rect 26255 -270 26275 -250
rect 26275 -270 26280 -250
rect 26250 -275 26280 -270
rect 26490 -250 26520 -245
rect 26490 -270 26495 -250
rect 26495 -270 26515 -250
rect 26515 -270 26520 -250
rect 26490 -275 26520 -270
rect 26730 -250 26760 -245
rect 26730 -270 26735 -250
rect 26735 -270 26755 -250
rect 26755 -270 26760 -250
rect 26730 -275 26760 -270
rect 26970 -250 27000 -245
rect 26970 -270 26975 -250
rect 26975 -270 26995 -250
rect 26995 -270 27000 -250
rect 26970 -275 27000 -270
rect 27210 -250 27240 -245
rect 27210 -270 27215 -250
rect 27215 -270 27235 -250
rect 27235 -270 27240 -250
rect 27210 -275 27240 -270
rect 27450 -250 27480 -245
rect 27450 -270 27455 -250
rect 27455 -270 27475 -250
rect 27475 -270 27480 -250
rect 27450 -275 27480 -270
rect 27690 -250 27720 -245
rect 27690 -270 27695 -250
rect 27695 -270 27715 -250
rect 27715 -270 27720 -250
rect 27690 -275 27720 -270
rect 27930 -250 27960 -245
rect 27930 -270 27935 -250
rect 27935 -270 27955 -250
rect 27955 -270 27960 -250
rect 27930 -275 27960 -270
rect 28170 -250 28200 -245
rect 28170 -270 28175 -250
rect 28175 -270 28195 -250
rect 28195 -270 28200 -250
rect 28170 -275 28200 -270
rect 28410 -250 28440 -245
rect 28410 -270 28415 -250
rect 28415 -270 28435 -250
rect 28435 -270 28440 -250
rect 28410 -275 28440 -270
rect 28650 -250 28680 -245
rect 28650 -270 28655 -250
rect 28655 -270 28675 -250
rect 28675 -270 28680 -250
rect 28650 -275 28680 -270
rect 28890 -250 28920 -245
rect 28890 -270 28895 -250
rect 28895 -270 28915 -250
rect 28915 -270 28920 -250
rect 28890 -275 28920 -270
rect 29130 -250 29160 -245
rect 29130 -270 29135 -250
rect 29135 -270 29155 -250
rect 29155 -270 29160 -250
rect 29130 -275 29160 -270
rect 29370 -250 29400 -245
rect 29370 -270 29375 -250
rect 29375 -270 29395 -250
rect 29395 -270 29400 -250
rect 29370 -275 29400 -270
rect 29610 -250 29640 -245
rect 29610 -270 29615 -250
rect 29615 -270 29635 -250
rect 29635 -270 29640 -250
rect 29610 -275 29640 -270
rect 29850 -250 29880 -245
rect 29850 -270 29855 -250
rect 29855 -270 29875 -250
rect 29875 -270 29880 -250
rect 29850 -275 29880 -270
rect 30090 -250 30120 -245
rect 30090 -270 30095 -250
rect 30095 -270 30115 -250
rect 30115 -270 30120 -250
rect 30090 -275 30120 -270
rect 30330 -250 30360 -245
rect 30330 -270 30335 -250
rect 30335 -270 30355 -250
rect 30355 -270 30360 -250
rect 30330 -275 30360 -270
rect 30570 -250 30600 -245
rect 30570 -270 30575 -250
rect 30575 -270 30595 -250
rect 30595 -270 30600 -250
rect 30570 -275 30600 -270
rect 30735 -485 30765 -480
rect 30735 -505 30740 -485
rect 30740 -505 30760 -485
rect 30760 -505 30765 -485
rect 30735 -510 30765 -505
rect 85 -825 115 -820
rect 85 -845 90 -825
rect 90 -845 110 -825
rect 110 -845 115 -825
rect 85 -850 115 -845
rect 325 -825 355 -820
rect 325 -845 330 -825
rect 330 -845 350 -825
rect 350 -845 355 -825
rect 325 -850 355 -845
rect 565 -825 595 -820
rect 565 -845 570 -825
rect 570 -845 590 -825
rect 590 -845 595 -825
rect 565 -850 595 -845
rect 800 -870 835 -835
rect 1045 -825 1075 -820
rect 1045 -845 1050 -825
rect 1050 -845 1070 -825
rect 1070 -845 1075 -825
rect 1045 -850 1075 -845
rect 1285 -825 1315 -820
rect 1285 -845 1290 -825
rect 1290 -845 1310 -825
rect 1310 -845 1315 -825
rect 1285 -850 1315 -845
rect 1525 -825 1555 -820
rect 1525 -845 1530 -825
rect 1530 -845 1550 -825
rect 1550 -845 1555 -825
rect 1525 -850 1555 -845
rect 1765 -825 1795 -820
rect 1765 -845 1770 -825
rect 1770 -845 1790 -825
rect 1790 -845 1795 -825
rect 1765 -850 1795 -845
rect 2005 -825 2035 -820
rect 2005 -845 2010 -825
rect 2010 -845 2030 -825
rect 2030 -845 2035 -825
rect 2005 -850 2035 -845
rect 2245 -825 2275 -820
rect 2245 -845 2250 -825
rect 2250 -845 2270 -825
rect 2270 -845 2275 -825
rect 2245 -850 2275 -845
rect 2485 -825 2515 -820
rect 2485 -845 2490 -825
rect 2490 -845 2510 -825
rect 2510 -845 2515 -825
rect 2485 -850 2515 -845
rect 2725 -825 2755 -820
rect 2725 -845 2730 -825
rect 2730 -845 2750 -825
rect 2750 -845 2755 -825
rect 2725 -850 2755 -845
rect 2960 -870 2995 -835
rect 3205 -825 3235 -820
rect 3205 -845 3210 -825
rect 3210 -845 3230 -825
rect 3230 -845 3235 -825
rect 3205 -850 3235 -845
rect 3445 -825 3475 -820
rect 3445 -845 3450 -825
rect 3450 -845 3470 -825
rect 3470 -845 3475 -825
rect 3445 -850 3475 -845
rect 3685 -825 3715 -820
rect 3685 -845 3690 -825
rect 3690 -845 3710 -825
rect 3710 -845 3715 -825
rect 3685 -850 3715 -845
rect 3925 -825 3955 -820
rect 3925 -845 3930 -825
rect 3930 -845 3950 -825
rect 3950 -845 3955 -825
rect 3925 -850 3955 -845
rect 4165 -825 4195 -820
rect 4165 -845 4170 -825
rect 4170 -845 4190 -825
rect 4190 -845 4195 -825
rect 4165 -850 4195 -845
rect 4405 -825 4435 -820
rect 4405 -845 4410 -825
rect 4410 -845 4430 -825
rect 4430 -845 4435 -825
rect 4405 -850 4435 -845
rect 4645 -825 4675 -820
rect 4645 -845 4650 -825
rect 4650 -845 4670 -825
rect 4670 -845 4675 -825
rect 4645 -850 4675 -845
rect 4885 -825 4915 -820
rect 4885 -845 4890 -825
rect 4890 -845 4910 -825
rect 4910 -845 4915 -825
rect 4885 -850 4915 -845
rect 5120 -870 5155 -835
rect 5365 -825 5395 -820
rect 5365 -845 5370 -825
rect 5370 -845 5390 -825
rect 5390 -845 5395 -825
rect 5365 -850 5395 -845
rect 5605 -825 5635 -820
rect 5605 -845 5610 -825
rect 5610 -845 5630 -825
rect 5630 -845 5635 -825
rect 5605 -850 5635 -845
rect 5845 -825 5875 -820
rect 5845 -845 5850 -825
rect 5850 -845 5870 -825
rect 5870 -845 5875 -825
rect 5845 -850 5875 -845
rect 6085 -825 6115 -820
rect 6085 -845 6090 -825
rect 6090 -845 6110 -825
rect 6110 -845 6115 -825
rect 6085 -850 6115 -845
rect 6325 -825 6355 -820
rect 6325 -845 6330 -825
rect 6330 -845 6350 -825
rect 6350 -845 6355 -825
rect 6325 -850 6355 -845
rect 6565 -825 6595 -820
rect 6565 -845 6570 -825
rect 6570 -845 6590 -825
rect 6590 -845 6595 -825
rect 6565 -850 6595 -845
rect 6805 -825 6835 -820
rect 6805 -845 6810 -825
rect 6810 -845 6830 -825
rect 6830 -845 6835 -825
rect 6805 -850 6835 -845
rect 7045 -825 7075 -820
rect 7045 -845 7050 -825
rect 7050 -845 7070 -825
rect 7070 -845 7075 -825
rect 7045 -850 7075 -845
rect 7280 -870 7315 -835
rect 7525 -825 7555 -820
rect 7525 -845 7530 -825
rect 7530 -845 7550 -825
rect 7550 -845 7555 -825
rect 7525 -850 7555 -845
rect 7765 -825 7795 -820
rect 7765 -845 7770 -825
rect 7770 -845 7790 -825
rect 7790 -845 7795 -825
rect 7765 -850 7795 -845
rect 8005 -825 8035 -820
rect 8005 -845 8010 -825
rect 8010 -845 8030 -825
rect 8030 -845 8035 -825
rect 8005 -850 8035 -845
rect 8245 -825 8275 -820
rect 8245 -845 8250 -825
rect 8250 -845 8270 -825
rect 8270 -845 8275 -825
rect 8245 -850 8275 -845
rect 8485 -825 8515 -820
rect 8485 -845 8490 -825
rect 8490 -845 8510 -825
rect 8510 -845 8515 -825
rect 8485 -850 8515 -845
rect 8725 -825 8755 -820
rect 8725 -845 8730 -825
rect 8730 -845 8750 -825
rect 8750 -845 8755 -825
rect 8725 -850 8755 -845
rect 8965 -825 8995 -820
rect 8965 -845 8970 -825
rect 8970 -845 8990 -825
rect 8990 -845 8995 -825
rect 8965 -850 8995 -845
rect 9205 -825 9235 -820
rect 9205 -845 9210 -825
rect 9210 -845 9230 -825
rect 9230 -845 9235 -825
rect 9205 -850 9235 -845
rect 9440 -870 9475 -835
rect 9685 -825 9715 -820
rect 9685 -845 9690 -825
rect 9690 -845 9710 -825
rect 9710 -845 9715 -825
rect 9685 -850 9715 -845
rect 9925 -825 9955 -820
rect 9925 -845 9930 -825
rect 9930 -845 9950 -825
rect 9950 -845 9955 -825
rect 9925 -850 9955 -845
rect 10165 -825 10195 -820
rect 10165 -845 10170 -825
rect 10170 -845 10190 -825
rect 10190 -845 10195 -825
rect 10165 -850 10195 -845
rect 10405 -825 10435 -820
rect 10405 -845 10410 -825
rect 10410 -845 10430 -825
rect 10430 -845 10435 -825
rect 10405 -850 10435 -845
rect 10645 -825 10675 -820
rect 10645 -845 10650 -825
rect 10650 -845 10670 -825
rect 10670 -845 10675 -825
rect 10645 -850 10675 -845
rect 10885 -825 10915 -820
rect 10885 -845 10890 -825
rect 10890 -845 10910 -825
rect 10910 -845 10915 -825
rect 10885 -850 10915 -845
rect 11125 -825 11155 -820
rect 11125 -845 11130 -825
rect 11130 -845 11150 -825
rect 11150 -845 11155 -825
rect 11125 -850 11155 -845
rect 11365 -825 11395 -820
rect 11365 -845 11370 -825
rect 11370 -845 11390 -825
rect 11390 -845 11395 -825
rect 11365 -850 11395 -845
rect 11600 -870 11635 -835
rect 11845 -825 11875 -820
rect 11845 -845 11850 -825
rect 11850 -845 11870 -825
rect 11870 -845 11875 -825
rect 11845 -850 11875 -845
rect 12085 -825 12115 -820
rect 12085 -845 12090 -825
rect 12090 -845 12110 -825
rect 12110 -845 12115 -825
rect 12085 -850 12115 -845
rect 12325 -825 12355 -820
rect 12325 -845 12330 -825
rect 12330 -845 12350 -825
rect 12350 -845 12355 -825
rect 12325 -850 12355 -845
rect 12565 -825 12595 -820
rect 12565 -845 12570 -825
rect 12570 -845 12590 -825
rect 12590 -845 12595 -825
rect 12565 -850 12595 -845
rect 12805 -825 12835 -820
rect 12805 -845 12810 -825
rect 12810 -845 12830 -825
rect 12830 -845 12835 -825
rect 12805 -850 12835 -845
rect 13045 -825 13075 -820
rect 13045 -845 13050 -825
rect 13050 -845 13070 -825
rect 13070 -845 13075 -825
rect 13045 -850 13075 -845
rect 13285 -825 13315 -820
rect 13285 -845 13290 -825
rect 13290 -845 13310 -825
rect 13310 -845 13315 -825
rect 13285 -850 13315 -845
rect 13525 -825 13555 -820
rect 13525 -845 13530 -825
rect 13530 -845 13550 -825
rect 13550 -845 13555 -825
rect 13525 -850 13555 -845
rect 13760 -870 13795 -835
rect 14005 -825 14035 -820
rect 14005 -845 14010 -825
rect 14010 -845 14030 -825
rect 14030 -845 14035 -825
rect 14005 -850 14035 -845
rect 14245 -825 14275 -820
rect 14245 -845 14250 -825
rect 14250 -845 14270 -825
rect 14270 -845 14275 -825
rect 14245 -850 14275 -845
rect 14485 -825 14515 -820
rect 14485 -845 14490 -825
rect 14490 -845 14510 -825
rect 14510 -845 14515 -825
rect 14485 -850 14515 -845
rect 14725 -825 14755 -820
rect 14725 -845 14730 -825
rect 14730 -845 14750 -825
rect 14750 -845 14755 -825
rect 14725 -850 14755 -845
rect 14965 -825 14995 -820
rect 14965 -845 14970 -825
rect 14970 -845 14990 -825
rect 14990 -845 14995 -825
rect 14965 -850 14995 -845
rect 15205 -825 15235 -820
rect 15205 -845 15210 -825
rect 15210 -845 15230 -825
rect 15230 -845 15235 -825
rect 15205 -850 15235 -845
rect 15445 -825 15475 -820
rect 15445 -845 15450 -825
rect 15450 -845 15470 -825
rect 15470 -845 15475 -825
rect 15445 -850 15475 -845
rect 15685 -825 15715 -820
rect 15685 -845 15690 -825
rect 15690 -845 15710 -825
rect 15710 -845 15715 -825
rect 15685 -850 15715 -845
rect 15920 -870 15955 -835
rect 16165 -825 16195 -820
rect 16165 -845 16170 -825
rect 16170 -845 16190 -825
rect 16190 -845 16195 -825
rect 16165 -850 16195 -845
rect 16405 -825 16435 -820
rect 16405 -845 16410 -825
rect 16410 -845 16430 -825
rect 16430 -845 16435 -825
rect 16405 -850 16435 -845
rect 16645 -825 16675 -820
rect 16645 -845 16650 -825
rect 16650 -845 16670 -825
rect 16670 -845 16675 -825
rect 16645 -850 16675 -845
rect 16885 -825 16915 -820
rect 16885 -845 16890 -825
rect 16890 -845 16910 -825
rect 16910 -845 16915 -825
rect 16885 -850 16915 -845
rect 17125 -825 17155 -820
rect 17125 -845 17130 -825
rect 17130 -845 17150 -825
rect 17150 -845 17155 -825
rect 17125 -850 17155 -845
rect 17365 -825 17395 -820
rect 17365 -845 17370 -825
rect 17370 -845 17390 -825
rect 17390 -845 17395 -825
rect 17365 -850 17395 -845
rect 17605 -825 17635 -820
rect 17605 -845 17610 -825
rect 17610 -845 17630 -825
rect 17630 -845 17635 -825
rect 17605 -850 17635 -845
rect 17845 -825 17875 -820
rect 17845 -845 17850 -825
rect 17850 -845 17870 -825
rect 17870 -845 17875 -825
rect 17845 -850 17875 -845
rect 18080 -870 18115 -835
rect 18325 -825 18355 -820
rect 18325 -845 18330 -825
rect 18330 -845 18350 -825
rect 18350 -845 18355 -825
rect 18325 -850 18355 -845
rect 18565 -825 18595 -820
rect 18565 -845 18570 -825
rect 18570 -845 18590 -825
rect 18590 -845 18595 -825
rect 18565 -850 18595 -845
rect 18805 -825 18835 -820
rect 18805 -845 18810 -825
rect 18810 -845 18830 -825
rect 18830 -845 18835 -825
rect 18805 -850 18835 -845
rect 19045 -825 19075 -820
rect 19045 -845 19050 -825
rect 19050 -845 19070 -825
rect 19070 -845 19075 -825
rect 19045 -850 19075 -845
rect 19285 -825 19315 -820
rect 19285 -845 19290 -825
rect 19290 -845 19310 -825
rect 19310 -845 19315 -825
rect 19285 -850 19315 -845
rect 19525 -825 19555 -820
rect 19525 -845 19530 -825
rect 19530 -845 19550 -825
rect 19550 -845 19555 -825
rect 19525 -850 19555 -845
rect 19765 -825 19795 -820
rect 19765 -845 19770 -825
rect 19770 -845 19790 -825
rect 19790 -845 19795 -825
rect 19765 -850 19795 -845
rect 20005 -825 20035 -820
rect 20005 -845 20010 -825
rect 20010 -845 20030 -825
rect 20030 -845 20035 -825
rect 20005 -850 20035 -845
rect 20240 -870 20275 -835
rect 20485 -825 20515 -820
rect 20485 -845 20490 -825
rect 20490 -845 20510 -825
rect 20510 -845 20515 -825
rect 20485 -850 20515 -845
rect 20725 -825 20755 -820
rect 20725 -845 20730 -825
rect 20730 -845 20750 -825
rect 20750 -845 20755 -825
rect 20725 -850 20755 -845
rect 20965 -825 20995 -820
rect 20965 -845 20970 -825
rect 20970 -845 20990 -825
rect 20990 -845 20995 -825
rect 20965 -850 20995 -845
rect 21205 -825 21235 -820
rect 21205 -845 21210 -825
rect 21210 -845 21230 -825
rect 21230 -845 21235 -825
rect 21205 -850 21235 -845
rect 21445 -825 21475 -820
rect 21445 -845 21450 -825
rect 21450 -845 21470 -825
rect 21470 -845 21475 -825
rect 21445 -850 21475 -845
rect 21685 -825 21715 -820
rect 21685 -845 21690 -825
rect 21690 -845 21710 -825
rect 21710 -845 21715 -825
rect 21685 -850 21715 -845
rect 21925 -825 21955 -820
rect 21925 -845 21930 -825
rect 21930 -845 21950 -825
rect 21950 -845 21955 -825
rect 21925 -850 21955 -845
rect 22165 -825 22195 -820
rect 22165 -845 22170 -825
rect 22170 -845 22190 -825
rect 22190 -845 22195 -825
rect 22165 -850 22195 -845
rect 22400 -870 22435 -835
rect 22645 -825 22675 -820
rect 22645 -845 22650 -825
rect 22650 -845 22670 -825
rect 22670 -845 22675 -825
rect 22645 -850 22675 -845
rect 22885 -825 22915 -820
rect 22885 -845 22890 -825
rect 22890 -845 22910 -825
rect 22910 -845 22915 -825
rect 22885 -850 22915 -845
rect 23125 -825 23155 -820
rect 23125 -845 23130 -825
rect 23130 -845 23150 -825
rect 23150 -845 23155 -825
rect 23125 -850 23155 -845
rect 23365 -825 23395 -820
rect 23365 -845 23370 -825
rect 23370 -845 23390 -825
rect 23390 -845 23395 -825
rect 23365 -850 23395 -845
rect 23605 -825 23635 -820
rect 23605 -845 23610 -825
rect 23610 -845 23630 -825
rect 23630 -845 23635 -825
rect 23605 -850 23635 -845
rect 23845 -825 23875 -820
rect 23845 -845 23850 -825
rect 23850 -845 23870 -825
rect 23870 -845 23875 -825
rect 23845 -850 23875 -845
rect 24085 -825 24115 -820
rect 24085 -845 24090 -825
rect 24090 -845 24110 -825
rect 24110 -845 24115 -825
rect 24085 -850 24115 -845
rect 24320 -870 24355 -835
rect 24565 -825 24595 -820
rect 24565 -845 24570 -825
rect 24570 -845 24590 -825
rect 24590 -845 24595 -825
rect 24565 -850 24595 -845
rect 24805 -825 24835 -820
rect 24805 -845 24810 -825
rect 24810 -845 24830 -825
rect 24830 -845 24835 -825
rect 24805 -850 24835 -845
rect 25045 -825 25075 -820
rect 25045 -845 25050 -825
rect 25050 -845 25070 -825
rect 25070 -845 25075 -825
rect 25045 -850 25075 -845
rect 25285 -825 25315 -820
rect 25285 -845 25290 -825
rect 25290 -845 25310 -825
rect 25310 -845 25315 -825
rect 25285 -850 25315 -845
rect 25525 -825 25555 -820
rect 25525 -845 25530 -825
rect 25530 -845 25550 -825
rect 25550 -845 25555 -825
rect 25525 -850 25555 -845
rect 25765 -825 25795 -820
rect 25765 -845 25770 -825
rect 25770 -845 25790 -825
rect 25790 -845 25795 -825
rect 25765 -850 25795 -845
rect 26005 -825 26035 -820
rect 26005 -845 26010 -825
rect 26010 -845 26030 -825
rect 26030 -845 26035 -825
rect 26005 -850 26035 -845
rect 26240 -870 26275 -835
rect 26485 -825 26515 -820
rect 26485 -845 26490 -825
rect 26490 -845 26510 -825
rect 26510 -845 26515 -825
rect 26485 -850 26515 -845
rect 26725 -825 26755 -820
rect 26725 -845 26730 -825
rect 26730 -845 26750 -825
rect 26750 -845 26755 -825
rect 26725 -850 26755 -845
rect 26965 -825 26995 -820
rect 26965 -845 26970 -825
rect 26970 -845 26990 -825
rect 26990 -845 26995 -825
rect 26965 -850 26995 -845
rect 27205 -825 27235 -820
rect 27205 -845 27210 -825
rect 27210 -845 27230 -825
rect 27230 -845 27235 -825
rect 27205 -850 27235 -845
rect 27445 -825 27475 -820
rect 27445 -845 27450 -825
rect 27450 -845 27470 -825
rect 27470 -845 27475 -825
rect 27445 -850 27475 -845
rect 27685 -825 27715 -820
rect 27685 -845 27690 -825
rect 27690 -845 27710 -825
rect 27710 -845 27715 -825
rect 27685 -850 27715 -845
rect 27925 -825 27955 -820
rect 27925 -845 27930 -825
rect 27930 -845 27950 -825
rect 27950 -845 27955 -825
rect 27925 -850 27955 -845
rect 28160 -870 28195 -835
rect 28405 -825 28435 -820
rect 28405 -845 28410 -825
rect 28410 -845 28430 -825
rect 28430 -845 28435 -825
rect 28405 -850 28435 -845
rect 28645 -825 28675 -820
rect 28645 -845 28650 -825
rect 28650 -845 28670 -825
rect 28670 -845 28675 -825
rect 28645 -850 28675 -845
rect 28885 -825 28915 -820
rect 28885 -845 28890 -825
rect 28890 -845 28910 -825
rect 28910 -845 28915 -825
rect 28885 -850 28915 -845
rect 29125 -825 29155 -820
rect 29125 -845 29130 -825
rect 29130 -845 29150 -825
rect 29150 -845 29155 -825
rect 29125 -850 29155 -845
rect 29365 -825 29395 -820
rect 29365 -845 29370 -825
rect 29370 -845 29390 -825
rect 29390 -845 29395 -825
rect 29365 -850 29395 -845
rect 29605 -825 29635 -820
rect 29605 -845 29610 -825
rect 29610 -845 29630 -825
rect 29630 -845 29635 -825
rect 29605 -850 29635 -845
rect 29840 -870 29875 -835
rect 30085 -825 30115 -820
rect 30085 -845 30090 -825
rect 30090 -845 30110 -825
rect 30110 -845 30115 -825
rect 30085 -850 30115 -845
rect 30325 -825 30355 -820
rect 30325 -845 30330 -825
rect 30330 -845 30350 -825
rect 30350 -845 30355 -825
rect 30325 -850 30355 -845
rect 30565 -825 30595 -820
rect 30565 -845 30570 -825
rect 30570 -845 30590 -825
rect 30590 -845 30595 -825
rect 30565 -850 30595 -845
<< metal2 >>
rect 2255 305 2310 315
rect 185 275 240 285
rect 185 240 195 275
rect 230 240 240 275
rect 185 230 240 240
rect 426 265 476 275
rect 426 235 436 265
rect 466 235 476 265
rect 426 225 476 235
rect 731 265 781 275
rect 731 235 741 265
rect 771 235 781 265
rect 731 225 781 235
rect 976 265 1026 275
rect 976 235 986 265
rect 1016 235 1026 265
rect 976 225 1026 235
rect 1216 265 1266 275
rect 1216 235 1226 265
rect 1256 235 1266 265
rect 1216 225 1266 235
rect 1461 265 1511 275
rect 1461 235 1471 265
rect 1501 235 1511 265
rect 1461 225 1511 235
rect 1766 265 1816 275
rect 1766 235 1776 265
rect 1806 235 1816 265
rect 1766 225 1816 235
rect 2011 265 2061 275
rect 2011 235 2021 265
rect 2051 235 2061 265
rect 2255 270 2265 305
rect 2300 270 2310 305
rect 4195 305 4250 315
rect 2255 260 2310 270
rect 2496 265 2546 275
rect 2011 225 2061 235
rect 2496 235 2506 265
rect 2536 235 2546 265
rect 2496 225 2546 235
rect 2736 265 2786 275
rect 2736 235 2746 265
rect 2776 235 2786 265
rect 2736 225 2786 235
rect 2981 265 3031 275
rect 2981 235 2991 265
rect 3021 235 3031 265
rect 2981 225 3031 235
rect 3221 265 3271 275
rect 3221 235 3231 265
rect 3261 235 3271 265
rect 3221 225 3271 235
rect 3466 265 3516 275
rect 3466 235 3476 265
rect 3506 235 3516 265
rect 3466 225 3516 235
rect 3706 265 3756 275
rect 3706 235 3716 265
rect 3746 235 3756 265
rect 3706 225 3756 235
rect 3951 265 4001 275
rect 3951 235 3961 265
rect 3991 235 4001 265
rect 4195 270 4205 305
rect 4240 270 4250 305
rect 6445 305 6500 315
rect 4195 260 4250 270
rect 4436 265 4486 275
rect 3951 225 4001 235
rect 4436 235 4446 265
rect 4476 235 4486 265
rect 4436 225 4486 235
rect 4676 265 4726 275
rect 4676 235 4686 265
rect 4716 235 4726 265
rect 4676 225 4726 235
rect 4921 265 4971 275
rect 4921 235 4931 265
rect 4961 235 4971 265
rect 4921 225 4971 235
rect 5161 265 5211 275
rect 5161 235 5171 265
rect 5201 235 5211 265
rect 5161 225 5211 235
rect 5406 265 5456 275
rect 5406 235 5416 265
rect 5446 235 5456 265
rect 5406 225 5456 235
rect 5711 265 5761 275
rect 5711 235 5721 265
rect 5751 235 5761 265
rect 5711 225 5761 235
rect 5956 265 6006 275
rect 5956 235 5966 265
rect 5996 235 6006 265
rect 5956 225 6006 235
rect 6196 265 6246 275
rect 6196 235 6206 265
rect 6236 235 6246 265
rect 6445 270 6455 305
rect 6490 270 6500 305
rect 9350 305 9405 315
rect 6445 260 6500 270
rect 6681 265 6731 275
rect 6196 225 6246 235
rect 6681 235 6691 265
rect 6721 235 6731 265
rect 6681 225 6731 235
rect 6926 265 6976 275
rect 6926 235 6936 265
rect 6966 235 6976 265
rect 6926 225 6976 235
rect 7166 265 7216 275
rect 7166 235 7176 265
rect 7206 235 7216 265
rect 7166 225 7216 235
rect 7406 265 7456 275
rect 7406 235 7416 265
rect 7446 235 7456 265
rect 7406 225 7456 235
rect 7646 265 7696 275
rect 7646 235 7656 265
rect 7686 235 7696 265
rect 7646 225 7696 235
rect 7891 265 7941 275
rect 7891 235 7901 265
rect 7931 235 7941 265
rect 7891 225 7941 235
rect 8131 265 8181 275
rect 8131 235 8141 265
rect 8171 235 8181 265
rect 8131 225 8181 235
rect 8376 265 8426 275
rect 8376 235 8386 265
rect 8416 235 8426 265
rect 8376 225 8426 235
rect 8616 265 8666 275
rect 8616 235 8626 265
rect 8656 235 8666 265
rect 8616 225 8666 235
rect 8861 265 8911 275
rect 8861 235 8871 265
rect 8901 235 8911 265
rect 8861 225 8911 235
rect 9101 265 9151 275
rect 9101 235 9111 265
rect 9141 235 9151 265
rect 9350 270 9360 305
rect 9395 270 9405 305
rect 11295 305 11350 315
rect 9350 260 9405 270
rect 9591 265 9641 275
rect 9101 225 9151 235
rect 9591 235 9601 265
rect 9631 235 9641 265
rect 9591 225 9641 235
rect 9836 265 9886 275
rect 9836 235 9846 265
rect 9876 235 9886 265
rect 9836 225 9886 235
rect 10076 265 10126 275
rect 10076 235 10086 265
rect 10116 235 10126 265
rect 10076 225 10126 235
rect 10321 265 10371 275
rect 10321 235 10331 265
rect 10361 235 10371 265
rect 10321 225 10371 235
rect 10561 265 10611 275
rect 10561 235 10571 265
rect 10601 235 10611 265
rect 10561 225 10611 235
rect 10806 265 10856 275
rect 10806 235 10816 265
rect 10846 235 10856 265
rect 10806 225 10856 235
rect 11046 265 11096 275
rect 11046 235 11056 265
rect 11086 235 11096 265
rect 11295 270 11305 305
rect 11340 270 11350 305
rect 12990 305 13045 315
rect 11295 260 11350 270
rect 11531 265 11581 275
rect 11046 225 11096 235
rect 11531 235 11541 265
rect 11571 235 11581 265
rect 11531 225 11581 235
rect 11776 265 11826 275
rect 11776 235 11786 265
rect 11816 235 11826 265
rect 11776 225 11826 235
rect 12016 265 12066 275
rect 12016 235 12026 265
rect 12056 235 12066 265
rect 12016 225 12066 235
rect 12261 265 12311 275
rect 12261 235 12271 265
rect 12301 235 12311 265
rect 12261 225 12311 235
rect 12501 265 12551 275
rect 12501 235 12511 265
rect 12541 235 12551 265
rect 12501 225 12551 235
rect 12746 265 12796 275
rect 12746 235 12756 265
rect 12786 235 12796 265
rect 12990 270 13000 305
rect 13035 270 13045 305
rect 15175 305 15230 315
rect 12990 260 13045 270
rect 13231 265 13281 275
rect 12746 225 12796 235
rect 13231 235 13241 265
rect 13271 235 13281 265
rect 13231 225 13281 235
rect 13471 265 13521 275
rect 13471 235 13481 265
rect 13511 235 13521 265
rect 13471 225 13521 235
rect 13716 265 13766 275
rect 13716 235 13726 265
rect 13756 235 13766 265
rect 13716 225 13766 235
rect 13956 265 14006 275
rect 13956 235 13966 265
rect 13996 235 14006 265
rect 13956 225 14006 235
rect 14201 265 14251 275
rect 14201 235 14211 265
rect 14241 235 14251 265
rect 14201 225 14251 235
rect 14441 265 14491 275
rect 14441 235 14451 265
rect 14481 235 14491 265
rect 14441 225 14491 235
rect 14686 265 14736 275
rect 14686 235 14696 265
rect 14726 235 14736 265
rect 14686 225 14736 235
rect 14926 265 14976 275
rect 14926 235 14936 265
rect 14966 235 14976 265
rect 15175 270 15185 305
rect 15220 270 15230 305
rect 17355 305 17410 315
rect 15175 260 15230 270
rect 15411 265 15461 275
rect 14926 225 14976 235
rect 15411 235 15421 265
rect 15451 235 15461 265
rect 15411 225 15461 235
rect 15656 265 15706 275
rect 15656 235 15666 265
rect 15696 235 15706 265
rect 15656 225 15706 235
rect 15896 265 15946 275
rect 15896 235 15906 265
rect 15936 235 15946 265
rect 15896 225 15946 235
rect 16141 265 16191 275
rect 16141 235 16151 265
rect 16181 235 16191 265
rect 16141 225 16191 235
rect 16381 265 16431 275
rect 16381 235 16391 265
rect 16421 235 16431 265
rect 16381 225 16431 235
rect 16626 265 16676 275
rect 16626 235 16636 265
rect 16666 235 16676 265
rect 16626 225 16676 235
rect 16866 265 16916 275
rect 16866 235 16876 265
rect 16906 235 16916 265
rect 16866 225 16916 235
rect 17111 265 17161 275
rect 17111 235 17121 265
rect 17151 235 17161 265
rect 17355 270 17365 305
rect 17400 270 17410 305
rect 19540 305 19595 315
rect 17355 260 17410 270
rect 17596 265 17646 275
rect 17111 225 17161 235
rect 17596 235 17606 265
rect 17636 235 17646 265
rect 17596 225 17646 235
rect 17836 265 17886 275
rect 17836 235 17846 265
rect 17876 235 17886 265
rect 17836 225 17886 235
rect 18081 265 18131 275
rect 18081 235 18091 265
rect 18121 235 18131 265
rect 18081 225 18131 235
rect 18321 265 18371 275
rect 18321 235 18331 265
rect 18361 235 18371 265
rect 18321 225 18371 235
rect 18566 265 18616 275
rect 18566 235 18576 265
rect 18606 235 18616 265
rect 18566 225 18616 235
rect 18806 265 18856 275
rect 18806 235 18816 265
rect 18846 235 18856 265
rect 18806 225 18856 235
rect 19051 265 19101 275
rect 19051 235 19061 265
rect 19091 235 19101 265
rect 19051 225 19101 235
rect 19291 265 19341 275
rect 19291 235 19301 265
rect 19331 235 19341 265
rect 19540 270 19550 305
rect 19585 270 19595 305
rect 20750 305 20805 315
rect 19540 260 19595 270
rect 19776 265 19826 275
rect 19291 225 19341 235
rect 19776 235 19786 265
rect 19816 235 19826 265
rect 19776 225 19826 235
rect 20021 265 20071 275
rect 20021 235 20031 265
rect 20061 235 20071 265
rect 20021 225 20071 235
rect 20261 265 20311 275
rect 20261 235 20271 265
rect 20301 235 20311 265
rect 20261 225 20311 235
rect 20506 265 20556 275
rect 20506 235 20516 265
rect 20546 235 20556 265
rect 20750 270 20760 305
rect 20795 270 20805 305
rect 20750 260 20805 270
rect 20991 265 21041 275
rect 20506 225 20556 235
rect 20991 235 21001 265
rect 21031 235 21041 265
rect 20991 225 21041 235
rect 21145 15 21195 25
rect 21145 -15 21155 15
rect 21185 -15 21195 15
rect 21145 -25 21195 -15
rect 176 -165 226 -155
rect -425 -190 -355 -180
rect -425 -240 -415 -190
rect -365 -240 -355 -190
rect 176 -195 186 -165
rect 216 -195 226 -165
rect 176 -205 226 -195
rect 421 -165 471 -155
rect 421 -195 431 -165
rect 461 -195 471 -165
rect 421 -205 471 -195
rect 726 -165 776 -155
rect 726 -195 736 -165
rect 766 -195 776 -165
rect 726 -205 776 -195
rect 971 -165 1021 -155
rect 971 -195 981 -165
rect 1011 -195 1021 -165
rect 971 -205 1021 -195
rect 1211 -165 1261 -155
rect 1211 -195 1221 -165
rect 1251 -195 1261 -165
rect 1211 -205 1261 -195
rect 1456 -165 1506 -155
rect 1456 -195 1466 -165
rect 1496 -195 1506 -165
rect 1761 -165 1811 -155
rect 1456 -205 1506 -195
rect 1625 -200 1685 -190
rect -425 -250 -355 -240
rect 80 -245 130 -235
rect 80 -275 90 -245
rect 120 -275 130 -245
rect 80 -285 130 -275
rect 320 -245 370 -235
rect 320 -275 330 -245
rect 360 -275 370 -245
rect 320 -285 370 -275
rect 560 -245 610 -235
rect 560 -275 570 -245
rect 600 -275 610 -245
rect 560 -285 610 -275
rect 800 -245 850 -235
rect 800 -275 810 -245
rect 840 -275 850 -245
rect 800 -285 850 -275
rect 1040 -245 1090 -235
rect 1040 -275 1050 -245
rect 1080 -275 1090 -245
rect 1040 -285 1090 -275
rect 1280 -245 1330 -235
rect 1280 -275 1290 -245
rect 1320 -275 1330 -245
rect 1280 -285 1330 -275
rect 1520 -245 1570 -235
rect 1520 -275 1530 -245
rect 1560 -275 1570 -245
rect 1625 -240 1635 -200
rect 1675 -240 1685 -200
rect 1761 -195 1771 -165
rect 1801 -195 1811 -165
rect 1761 -205 1811 -195
rect 2006 -165 2056 -155
rect 2006 -195 2016 -165
rect 2046 -195 2056 -165
rect 2006 -205 2056 -195
rect 2246 -165 2296 -155
rect 2246 -195 2256 -165
rect 2286 -195 2296 -165
rect 2246 -205 2296 -195
rect 2491 -165 2541 -155
rect 2491 -195 2501 -165
rect 2531 -195 2541 -165
rect 2491 -205 2541 -195
rect 2731 -165 2781 -155
rect 2731 -195 2741 -165
rect 2771 -195 2781 -165
rect 2731 -205 2781 -195
rect 2976 -165 3026 -155
rect 2976 -195 2986 -165
rect 3016 -195 3026 -165
rect 2976 -205 3026 -195
rect 3216 -165 3266 -155
rect 3216 -195 3226 -165
rect 3256 -195 3266 -165
rect 3216 -205 3266 -195
rect 3461 -165 3511 -155
rect 3461 -195 3471 -165
rect 3501 -195 3511 -165
rect 3461 -205 3511 -195
rect 3701 -165 3751 -155
rect 3701 -195 3711 -165
rect 3741 -195 3751 -165
rect 3701 -205 3751 -195
rect 3946 -165 3996 -155
rect 3946 -195 3956 -165
rect 3986 -195 3996 -165
rect 4186 -165 4236 -155
rect 3946 -205 3996 -195
rect 4050 -195 4110 -185
rect 4050 -235 4060 -195
rect 4100 -235 4110 -195
rect 4186 -195 4196 -165
rect 4226 -195 4236 -165
rect 4186 -205 4236 -195
rect 4431 -165 4481 -155
rect 4431 -195 4441 -165
rect 4471 -195 4481 -165
rect 4431 -205 4481 -195
rect 4671 -165 4721 -155
rect 4671 -195 4681 -165
rect 4711 -195 4721 -165
rect 4671 -205 4721 -195
rect 4916 -165 4966 -155
rect 4916 -195 4926 -165
rect 4956 -195 4966 -165
rect 4916 -205 4966 -195
rect 5156 -165 5206 -155
rect 5156 -195 5166 -165
rect 5196 -195 5206 -165
rect 5156 -205 5206 -195
rect 5401 -165 5451 -155
rect 5401 -195 5411 -165
rect 5441 -195 5451 -165
rect 5401 -205 5451 -195
rect 5706 -165 5756 -155
rect 5706 -195 5716 -165
rect 5746 -195 5756 -165
rect 5706 -205 5756 -195
rect 5951 -165 6001 -155
rect 5951 -195 5961 -165
rect 5991 -195 6001 -165
rect 5951 -205 6001 -195
rect 6191 -165 6241 -155
rect 6191 -195 6201 -165
rect 6231 -195 6241 -165
rect 6191 -205 6241 -195
rect 6676 -165 6726 -155
rect 6676 -195 6686 -165
rect 6716 -195 6726 -165
rect 6676 -205 6726 -195
rect 6921 -165 6971 -155
rect 6921 -195 6931 -165
rect 6961 -195 6971 -165
rect 6921 -205 6971 -195
rect 7161 -165 7211 -155
rect 7161 -195 7171 -165
rect 7201 -195 7211 -165
rect 7161 -205 7211 -195
rect 7401 -165 7451 -155
rect 7401 -195 7411 -165
rect 7441 -195 7451 -165
rect 7401 -205 7451 -195
rect 7641 -165 7691 -155
rect 7641 -195 7651 -165
rect 7681 -195 7691 -165
rect 7641 -205 7691 -195
rect 8126 -165 8176 -155
rect 8126 -195 8136 -165
rect 8166 -195 8176 -165
rect 8126 -205 8176 -195
rect 8371 -165 8421 -155
rect 8371 -195 8381 -165
rect 8411 -195 8421 -165
rect 8371 -205 8421 -195
rect 8611 -165 8661 -155
rect 8611 -195 8621 -165
rect 8651 -195 8661 -165
rect 8611 -205 8661 -195
rect 8856 -165 8906 -155
rect 8856 -195 8866 -165
rect 8896 -195 8906 -165
rect 8856 -205 8906 -195
rect 9096 -165 9146 -155
rect 9096 -195 9106 -165
rect 9136 -195 9146 -165
rect 9096 -205 9146 -195
rect 9341 -165 9391 -155
rect 9341 -195 9351 -165
rect 9381 -195 9391 -165
rect 9341 -205 9391 -195
rect 9831 -165 9881 -155
rect 9831 -195 9841 -165
rect 9871 -195 9881 -165
rect 9560 -210 9620 -200
rect 9831 -205 9881 -195
rect 10071 -165 10121 -155
rect 10071 -195 10081 -165
rect 10111 -195 10121 -165
rect 10071 -205 10121 -195
rect 10316 -165 10366 -155
rect 10316 -195 10326 -165
rect 10356 -195 10366 -165
rect 10316 -205 10366 -195
rect 10556 -165 10606 -155
rect 10556 -195 10566 -165
rect 10596 -195 10606 -165
rect 10556 -205 10606 -195
rect 10801 -165 10851 -155
rect 10801 -195 10811 -165
rect 10841 -195 10851 -165
rect 10801 -205 10851 -195
rect 11041 -165 11091 -155
rect 11041 -195 11051 -165
rect 11081 -195 11091 -165
rect 11041 -205 11091 -195
rect 11286 -165 11336 -155
rect 11286 -195 11296 -165
rect 11326 -195 11336 -165
rect 11286 -205 11336 -195
rect 11526 -165 11576 -155
rect 11526 -195 11536 -165
rect 11566 -195 11576 -165
rect 11526 -205 11576 -195
rect 11771 -165 11821 -155
rect 11771 -195 11781 -165
rect 11811 -195 11821 -165
rect 11771 -205 11821 -195
rect 12256 -165 12306 -155
rect 12256 -195 12266 -165
rect 12296 -195 12306 -165
rect 12256 -205 12306 -195
rect 12496 -165 12546 -155
rect 12496 -195 12506 -165
rect 12536 -195 12546 -165
rect 12496 -205 12546 -195
rect 12741 -165 12791 -155
rect 12741 -195 12751 -165
rect 12781 -195 12791 -165
rect 12741 -205 12791 -195
rect 12981 -165 13031 -155
rect 12981 -195 12991 -165
rect 13021 -195 13031 -165
rect 12981 -205 13031 -195
rect 13226 -165 13276 -155
rect 13226 -195 13236 -165
rect 13266 -195 13276 -165
rect 13226 -205 13276 -195
rect 13466 -165 13516 -155
rect 13466 -195 13476 -165
rect 13506 -195 13516 -165
rect 13466 -205 13516 -195
rect 13711 -165 13761 -155
rect 13711 -195 13721 -165
rect 13751 -195 13761 -165
rect 13711 -205 13761 -195
rect 14196 -165 14246 -155
rect 14196 -195 14206 -165
rect 14236 -195 14246 -165
rect 14196 -205 14246 -195
rect 14436 -165 14486 -155
rect 14436 -195 14446 -165
rect 14476 -195 14486 -165
rect 14436 -205 14486 -195
rect 14681 -165 14731 -155
rect 14681 -195 14691 -165
rect 14721 -195 14731 -165
rect 14681 -205 14731 -195
rect 14921 -165 14971 -155
rect 14921 -195 14931 -165
rect 14961 -195 14971 -165
rect 14921 -205 14971 -195
rect 15166 -165 15216 -155
rect 15166 -195 15176 -165
rect 15206 -195 15216 -165
rect 15166 -205 15216 -195
rect 15406 -165 15456 -155
rect 15406 -195 15416 -165
rect 15446 -195 15456 -165
rect 15406 -205 15456 -195
rect 15651 -165 15701 -155
rect 15651 -195 15661 -165
rect 15691 -195 15701 -165
rect 15651 -205 15701 -195
rect 16136 -165 16186 -155
rect 16136 -195 16146 -165
rect 16176 -195 16186 -165
rect 16136 -205 16186 -195
rect 16376 -165 16426 -155
rect 16376 -195 16386 -165
rect 16416 -195 16426 -165
rect 16376 -205 16426 -195
rect 16621 -165 16671 -155
rect 16621 -195 16631 -165
rect 16661 -195 16671 -165
rect 16621 -205 16671 -195
rect 16861 -165 16911 -155
rect 16861 -195 16871 -165
rect 16901 -195 16911 -165
rect 16861 -205 16911 -195
rect 17106 -165 17156 -155
rect 17106 -195 17116 -165
rect 17146 -195 17156 -165
rect 17106 -205 17156 -195
rect 17346 -165 17396 -155
rect 17346 -195 17356 -165
rect 17386 -195 17396 -165
rect 17346 -205 17396 -195
rect 17591 -165 17641 -155
rect 17591 -195 17601 -165
rect 17631 -195 17641 -165
rect 17591 -205 17641 -195
rect 17831 -165 17881 -155
rect 17831 -195 17841 -165
rect 17871 -195 17881 -165
rect 17695 -210 17755 -200
rect 17831 -205 17881 -195
rect 18076 -165 18126 -155
rect 18076 -195 18086 -165
rect 18116 -195 18126 -165
rect 18076 -205 18126 -195
rect 18316 -165 18366 -155
rect 18316 -195 18326 -165
rect 18356 -195 18366 -165
rect 18316 -205 18366 -195
rect 18561 -165 18611 -155
rect 18561 -195 18571 -165
rect 18601 -195 18611 -165
rect 18561 -205 18611 -195
rect 18801 -165 18851 -155
rect 18801 -195 18811 -165
rect 18841 -195 18851 -165
rect 18801 -205 18851 -195
rect 19046 -165 19096 -155
rect 19046 -195 19056 -165
rect 19086 -195 19096 -165
rect 19046 -205 19096 -195
rect 19286 -165 19336 -155
rect 19286 -195 19296 -165
rect 19326 -195 19336 -165
rect 19286 -205 19336 -195
rect 19531 -165 19581 -155
rect 19531 -195 19541 -165
rect 19571 -195 19581 -165
rect 19531 -205 19581 -195
rect 19771 -165 19821 -155
rect 19771 -195 19781 -165
rect 19811 -195 19821 -165
rect 6445 -220 6505 -210
rect 1625 -250 1685 -240
rect 1760 -245 1810 -235
rect 1520 -285 1570 -275
rect 1760 -275 1770 -245
rect 1800 -275 1810 -245
rect 1760 -285 1810 -275
rect 2000 -245 2050 -235
rect 2000 -275 2010 -245
rect 2040 -275 2050 -245
rect 2000 -285 2050 -275
rect 2240 -245 2290 -235
rect 2240 -275 2250 -245
rect 2280 -275 2290 -245
rect 2240 -285 2290 -275
rect 2480 -245 2530 -235
rect 2480 -275 2490 -245
rect 2520 -275 2530 -245
rect 2480 -285 2530 -275
rect 2720 -245 2770 -235
rect 2720 -275 2730 -245
rect 2760 -275 2770 -245
rect 2720 -285 2770 -275
rect 2960 -245 3010 -235
rect 2960 -275 2970 -245
rect 3000 -275 3010 -245
rect 2960 -285 3010 -275
rect 3200 -245 3250 -235
rect 3200 -275 3210 -245
rect 3240 -275 3250 -245
rect 3200 -285 3250 -275
rect 3440 -245 3490 -235
rect 3440 -275 3450 -245
rect 3480 -275 3490 -245
rect 3440 -285 3490 -275
rect 3680 -245 3730 -235
rect 3680 -275 3690 -245
rect 3720 -275 3730 -245
rect 3680 -285 3730 -275
rect 3920 -245 3970 -235
rect 4050 -245 4110 -235
rect 4160 -245 4210 -235
rect 3920 -275 3930 -245
rect 3960 -275 3970 -245
rect 3920 -285 3970 -275
rect 4160 -275 4170 -245
rect 4200 -275 4210 -245
rect 4160 -285 4210 -275
rect 4400 -245 4450 -235
rect 4400 -275 4410 -245
rect 4440 -275 4450 -245
rect 4400 -285 4450 -275
rect 4640 -245 4690 -235
rect 4640 -275 4650 -245
rect 4680 -275 4690 -245
rect 4640 -285 4690 -275
rect 4880 -245 4930 -235
rect 4880 -275 4890 -245
rect 4920 -275 4930 -245
rect 4880 -285 4930 -275
rect 5120 -245 5170 -235
rect 5120 -275 5130 -245
rect 5160 -275 5170 -245
rect 5120 -285 5170 -275
rect 5360 -245 5410 -235
rect 5360 -275 5370 -245
rect 5400 -275 5410 -245
rect 5360 -285 5410 -275
rect 5600 -245 5650 -235
rect 5600 -275 5610 -245
rect 5640 -275 5650 -245
rect 5600 -285 5650 -275
rect 5840 -245 5890 -235
rect 5840 -275 5850 -245
rect 5880 -275 5890 -245
rect 5840 -285 5890 -275
rect 6080 -245 6130 -235
rect 6080 -275 6090 -245
rect 6120 -275 6130 -245
rect 6080 -285 6130 -275
rect 6320 -245 6370 -235
rect 6320 -275 6330 -245
rect 6360 -275 6370 -245
rect 6445 -260 6455 -220
rect 6495 -260 6505 -220
rect 7870 -220 7930 -210
rect 6445 -270 6505 -260
rect 6560 -245 6610 -235
rect 6320 -285 6370 -275
rect 6560 -275 6570 -245
rect 6600 -275 6610 -245
rect 6560 -285 6610 -275
rect 6800 -245 6850 -235
rect 6800 -275 6810 -245
rect 6840 -275 6850 -245
rect 6800 -285 6850 -275
rect 7040 -245 7090 -235
rect 7040 -275 7050 -245
rect 7080 -275 7090 -245
rect 7040 -285 7090 -275
rect 7280 -245 7330 -235
rect 7280 -275 7290 -245
rect 7320 -275 7330 -245
rect 7280 -285 7330 -275
rect 7520 -245 7570 -235
rect 7520 -275 7530 -245
rect 7560 -275 7570 -245
rect 7520 -285 7570 -275
rect 7760 -245 7810 -235
rect 7760 -275 7770 -245
rect 7800 -275 7810 -245
rect 7870 -260 7880 -220
rect 7920 -260 7930 -220
rect 7870 -270 7930 -260
rect 8000 -245 8050 -235
rect 7760 -285 7810 -275
rect 8000 -275 8010 -245
rect 8040 -275 8050 -245
rect 8000 -285 8050 -275
rect 8240 -245 8290 -235
rect 8240 -275 8250 -245
rect 8280 -275 8290 -245
rect 8240 -285 8290 -275
rect 8480 -245 8530 -235
rect 8480 -275 8490 -245
rect 8520 -275 8530 -245
rect 8480 -285 8530 -275
rect 8720 -245 8770 -235
rect 8720 -275 8730 -245
rect 8760 -275 8770 -245
rect 8720 -285 8770 -275
rect 8960 -245 9010 -235
rect 8960 -275 8970 -245
rect 9000 -275 9010 -245
rect 8960 -285 9010 -275
rect 9200 -245 9250 -235
rect 9200 -275 9210 -245
rect 9240 -275 9250 -245
rect 9200 -285 9250 -275
rect 9440 -245 9490 -235
rect 9440 -275 9450 -245
rect 9480 -275 9490 -245
rect 9560 -250 9570 -210
rect 9610 -250 9620 -210
rect 11940 -220 12000 -210
rect 9560 -260 9620 -250
rect 9680 -245 9730 -235
rect 9440 -285 9490 -275
rect 9680 -275 9690 -245
rect 9720 -275 9730 -245
rect 9680 -285 9730 -275
rect 9920 -245 9970 -235
rect 9920 -275 9930 -245
rect 9960 -275 9970 -245
rect 9920 -285 9970 -275
rect 10160 -245 10210 -235
rect 10160 -275 10170 -245
rect 10200 -275 10210 -245
rect 10160 -285 10210 -275
rect 10400 -245 10450 -235
rect 10400 -275 10410 -245
rect 10440 -275 10450 -245
rect 10400 -285 10450 -275
rect 10640 -245 10690 -235
rect 10640 -275 10650 -245
rect 10680 -275 10690 -245
rect 10640 -285 10690 -275
rect 10880 -245 10930 -235
rect 10880 -275 10890 -245
rect 10920 -275 10930 -245
rect 10880 -285 10930 -275
rect 11120 -245 11170 -235
rect 11120 -275 11130 -245
rect 11160 -275 11170 -245
rect 11120 -285 11170 -275
rect 11360 -245 11410 -235
rect 11360 -275 11370 -245
rect 11400 -275 11410 -245
rect 11360 -285 11410 -275
rect 11600 -245 11650 -235
rect 11600 -275 11610 -245
rect 11640 -275 11650 -245
rect 11600 -285 11650 -275
rect 11840 -245 11890 -235
rect 11840 -275 11850 -245
rect 11880 -275 11890 -245
rect 11940 -260 11950 -220
rect 11990 -260 12000 -220
rect 13860 -220 13920 -210
rect 11940 -270 12000 -260
rect 12080 -245 12130 -235
rect 11840 -285 11890 -275
rect 12080 -275 12090 -245
rect 12120 -275 12130 -245
rect 12080 -285 12130 -275
rect 12320 -245 12370 -235
rect 12320 -275 12330 -245
rect 12360 -275 12370 -245
rect 12320 -285 12370 -275
rect 12560 -245 12610 -235
rect 12560 -275 12570 -245
rect 12600 -275 12610 -245
rect 12560 -285 12610 -275
rect 12800 -245 12850 -235
rect 12800 -275 12810 -245
rect 12840 -275 12850 -245
rect 12800 -285 12850 -275
rect 13040 -245 13090 -235
rect 13040 -275 13050 -245
rect 13080 -275 13090 -245
rect 13040 -285 13090 -275
rect 13280 -245 13330 -235
rect 13280 -275 13290 -245
rect 13320 -275 13330 -245
rect 13280 -285 13330 -275
rect 13520 -245 13570 -235
rect 13520 -275 13530 -245
rect 13560 -275 13570 -245
rect 13520 -285 13570 -275
rect 13760 -245 13810 -235
rect 13760 -275 13770 -245
rect 13800 -275 13810 -245
rect 13860 -260 13870 -220
rect 13910 -260 13920 -220
rect 15805 -220 15865 -210
rect 13860 -270 13920 -260
rect 14000 -245 14050 -235
rect 13760 -285 13810 -275
rect 14000 -275 14010 -245
rect 14040 -275 14050 -245
rect 14000 -285 14050 -275
rect 14240 -245 14290 -235
rect 14240 -275 14250 -245
rect 14280 -275 14290 -245
rect 14240 -285 14290 -275
rect 14480 -245 14530 -235
rect 14480 -275 14490 -245
rect 14520 -275 14530 -245
rect 14480 -285 14530 -275
rect 14720 -245 14770 -235
rect 14720 -275 14730 -245
rect 14760 -275 14770 -245
rect 14720 -285 14770 -275
rect 14960 -245 15010 -235
rect 14960 -275 14970 -245
rect 15000 -275 15010 -245
rect 14960 -285 15010 -275
rect 15200 -245 15250 -235
rect 15200 -275 15210 -245
rect 15240 -275 15250 -245
rect 15200 -285 15250 -275
rect 15440 -245 15490 -235
rect 15440 -275 15450 -245
rect 15480 -275 15490 -245
rect 15440 -285 15490 -275
rect 15680 -245 15730 -235
rect 15680 -275 15690 -245
rect 15720 -275 15730 -245
rect 15805 -260 15815 -220
rect 15855 -260 15865 -220
rect 15805 -270 15865 -260
rect 15920 -245 15970 -235
rect 15680 -285 15730 -275
rect 15920 -275 15930 -245
rect 15960 -275 15970 -245
rect 15920 -285 15970 -275
rect 16160 -245 16210 -235
rect 16160 -275 16170 -245
rect 16200 -275 16210 -245
rect 16160 -285 16210 -275
rect 16400 -245 16450 -235
rect 16400 -275 16410 -245
rect 16440 -275 16450 -245
rect 16400 -285 16450 -275
rect 16640 -245 16690 -235
rect 16640 -275 16650 -245
rect 16680 -275 16690 -245
rect 16640 -285 16690 -275
rect 16880 -245 16930 -235
rect 16880 -275 16890 -245
rect 16920 -275 16930 -245
rect 16880 -285 16930 -275
rect 17120 -245 17170 -235
rect 17120 -275 17130 -245
rect 17160 -275 17170 -245
rect 17120 -285 17170 -275
rect 17360 -245 17410 -235
rect 17360 -275 17370 -245
rect 17400 -275 17410 -245
rect 17360 -285 17410 -275
rect 17600 -245 17650 -235
rect 17600 -275 17610 -245
rect 17640 -275 17650 -245
rect 17695 -250 17705 -210
rect 17745 -250 17755 -210
rect 19635 -210 19695 -200
rect 19771 -205 19821 -195
rect 20016 -165 20066 -155
rect 20016 -195 20026 -165
rect 20056 -195 20066 -165
rect 20016 -205 20066 -195
rect 20256 -165 20306 -155
rect 20256 -195 20266 -165
rect 20296 -195 20306 -165
rect 20256 -205 20306 -195
rect 20501 -165 20551 -155
rect 20501 -195 20511 -165
rect 20541 -195 20551 -165
rect 20501 -205 20551 -195
rect 20741 -165 20791 -155
rect 20741 -195 20751 -165
rect 20781 -195 20791 -165
rect 20741 -205 20791 -195
rect 20986 -165 21036 -155
rect 20986 -195 20996 -165
rect 21026 -195 21036 -165
rect 21160 -185 21180 -25
rect 20986 -205 21036 -195
rect 21155 -205 30765 -185
rect 17695 -260 17755 -250
rect 17840 -245 17890 -235
rect 17600 -285 17650 -275
rect 17840 -275 17850 -245
rect 17880 -275 17890 -245
rect 17840 -285 17890 -275
rect 18080 -245 18130 -235
rect 18080 -275 18090 -245
rect 18120 -275 18130 -245
rect 18080 -285 18130 -275
rect 18320 -245 18370 -235
rect 18320 -275 18330 -245
rect 18360 -275 18370 -245
rect 18320 -285 18370 -275
rect 18560 -245 18610 -235
rect 18560 -275 18570 -245
rect 18600 -275 18610 -245
rect 18560 -285 18610 -275
rect 18800 -245 18850 -235
rect 18800 -275 18810 -245
rect 18840 -275 18850 -245
rect 18800 -285 18850 -275
rect 19040 -245 19090 -235
rect 19040 -275 19050 -245
rect 19080 -275 19090 -245
rect 19040 -285 19090 -275
rect 19280 -245 19330 -235
rect 19280 -275 19290 -245
rect 19320 -275 19330 -245
rect 19280 -285 19330 -275
rect 19520 -245 19570 -235
rect 19520 -275 19530 -245
rect 19560 -275 19570 -245
rect 19635 -250 19645 -210
rect 19685 -250 19695 -210
rect 19635 -260 19695 -250
rect 19760 -245 19810 -235
rect 19520 -285 19570 -275
rect 19760 -275 19770 -245
rect 19800 -275 19810 -245
rect 19760 -285 19810 -275
rect 20000 -245 20050 -235
rect 20000 -275 20010 -245
rect 20040 -275 20050 -245
rect 20000 -285 20050 -275
rect 20240 -245 20290 -235
rect 20240 -275 20250 -245
rect 20280 -275 20290 -245
rect 20240 -285 20290 -275
rect 20480 -245 20530 -235
rect 20480 -275 20490 -245
rect 20520 -275 20530 -245
rect 20480 -285 20530 -275
rect 20720 -245 20770 -235
rect 20720 -275 20730 -245
rect 20760 -275 20770 -245
rect 20720 -285 20770 -275
rect 20960 -245 21010 -235
rect 20960 -275 20970 -245
rect 21000 -275 21010 -245
rect 20960 -285 21010 -275
rect 21200 -245 21250 -235
rect 21200 -275 21210 -245
rect 21240 -275 21250 -245
rect 21200 -285 21250 -275
rect 21440 -245 21490 -235
rect 21440 -275 21450 -245
rect 21480 -275 21490 -245
rect 21440 -285 21490 -275
rect 21680 -245 21730 -235
rect 21680 -275 21690 -245
rect 21720 -275 21730 -245
rect 21680 -285 21730 -275
rect 21920 -245 21970 -235
rect 21920 -275 21930 -245
rect 21960 -275 21970 -245
rect 21920 -285 21970 -275
rect 22160 -245 22210 -235
rect 22160 -275 22170 -245
rect 22200 -275 22210 -245
rect 22160 -285 22210 -275
rect 22400 -245 22450 -235
rect 22400 -275 22410 -245
rect 22440 -275 22450 -245
rect 22400 -285 22450 -275
rect 22640 -245 22690 -235
rect 22640 -275 22650 -245
rect 22680 -275 22690 -245
rect 22640 -285 22690 -275
rect 22880 -245 22930 -235
rect 22880 -275 22890 -245
rect 22920 -275 22930 -245
rect 22880 -285 22930 -275
rect 23120 -245 23170 -235
rect 23120 -275 23130 -245
rect 23160 -275 23170 -245
rect 23120 -285 23170 -275
rect 23360 -245 23410 -235
rect 23360 -275 23370 -245
rect 23400 -275 23410 -245
rect 23360 -285 23410 -275
rect 23600 -245 23650 -235
rect 23600 -275 23610 -245
rect 23640 -275 23650 -245
rect 23600 -285 23650 -275
rect 23840 -245 23890 -235
rect 23840 -275 23850 -245
rect 23880 -275 23890 -245
rect 23840 -285 23890 -275
rect 24080 -245 24130 -235
rect 24080 -275 24090 -245
rect 24120 -275 24130 -245
rect 24080 -285 24130 -275
rect 24320 -245 24370 -235
rect 24320 -275 24330 -245
rect 24360 -275 24370 -245
rect 24320 -285 24370 -275
rect 24560 -245 24610 -235
rect 24560 -275 24570 -245
rect 24600 -275 24610 -245
rect 24560 -285 24610 -275
rect 24800 -245 24850 -235
rect 24800 -275 24810 -245
rect 24840 -275 24850 -245
rect 24800 -285 24850 -275
rect 25040 -245 25090 -235
rect 25040 -275 25050 -245
rect 25080 -275 25090 -245
rect 25040 -285 25090 -275
rect 25280 -245 25330 -235
rect 25280 -275 25290 -245
rect 25320 -275 25330 -245
rect 25280 -285 25330 -275
rect 25520 -245 25570 -235
rect 25520 -275 25530 -245
rect 25560 -275 25570 -245
rect 25520 -285 25570 -275
rect 25760 -245 25810 -235
rect 25760 -275 25770 -245
rect 25800 -275 25810 -245
rect 25760 -285 25810 -275
rect 26000 -245 26050 -235
rect 26000 -275 26010 -245
rect 26040 -275 26050 -245
rect 26000 -285 26050 -275
rect 26240 -245 26290 -235
rect 26240 -275 26250 -245
rect 26280 -275 26290 -245
rect 26240 -285 26290 -275
rect 26480 -245 26530 -235
rect 26480 -275 26490 -245
rect 26520 -275 26530 -245
rect 26480 -285 26530 -275
rect 26720 -245 26770 -235
rect 26720 -275 26730 -245
rect 26760 -275 26770 -245
rect 26720 -285 26770 -275
rect 26960 -245 27010 -235
rect 26960 -275 26970 -245
rect 27000 -275 27010 -245
rect 26960 -285 27010 -275
rect 27200 -245 27250 -235
rect 27200 -275 27210 -245
rect 27240 -275 27250 -245
rect 27200 -285 27250 -275
rect 27440 -245 27490 -235
rect 27440 -275 27450 -245
rect 27480 -275 27490 -245
rect 27440 -285 27490 -275
rect 27680 -245 27730 -235
rect 27680 -275 27690 -245
rect 27720 -275 27730 -245
rect 27680 -285 27730 -275
rect 27920 -245 27970 -235
rect 27920 -275 27930 -245
rect 27960 -275 27970 -245
rect 27920 -285 27970 -275
rect 28160 -245 28210 -235
rect 28160 -275 28170 -245
rect 28200 -275 28210 -245
rect 28160 -285 28210 -275
rect 28400 -245 28450 -235
rect 28400 -275 28410 -245
rect 28440 -275 28450 -245
rect 28400 -285 28450 -275
rect 28640 -245 28690 -235
rect 28640 -275 28650 -245
rect 28680 -275 28690 -245
rect 28640 -285 28690 -275
rect 28880 -245 28930 -235
rect 28880 -275 28890 -245
rect 28920 -275 28930 -245
rect 28880 -285 28930 -275
rect 29120 -245 29170 -235
rect 29120 -275 29130 -245
rect 29160 -275 29170 -245
rect 29120 -285 29170 -275
rect 29360 -245 29410 -235
rect 29360 -275 29370 -245
rect 29400 -275 29410 -245
rect 29360 -285 29410 -275
rect 29600 -245 29650 -235
rect 29600 -275 29610 -245
rect 29640 -275 29650 -245
rect 29600 -285 29650 -275
rect 29840 -245 29890 -235
rect 29840 -275 29850 -245
rect 29880 -275 29890 -245
rect 29840 -285 29890 -275
rect 30080 -245 30130 -235
rect 30080 -275 30090 -245
rect 30120 -275 30130 -245
rect 30080 -285 30130 -275
rect 30320 -245 30370 -235
rect 30320 -275 30330 -245
rect 30360 -275 30370 -245
rect 30320 -285 30370 -275
rect 30560 -245 30610 -235
rect 30560 -275 30570 -245
rect 30600 -275 30610 -245
rect 30560 -285 30610 -275
rect 30740 -470 30760 -205
rect 30725 -480 30775 -470
rect 30725 -510 30735 -480
rect 30765 -510 30775 -480
rect 30725 -520 30775 -510
rect 75 -820 125 -810
rect 75 -850 85 -820
rect 115 -850 125 -820
rect 75 -860 125 -850
rect 315 -820 365 -810
rect 315 -850 325 -820
rect 355 -850 365 -820
rect 315 -860 365 -850
rect 555 -820 605 -810
rect 555 -850 565 -820
rect 595 -850 605 -820
rect 1035 -820 1085 -810
rect 555 -860 605 -850
rect 790 -835 845 -825
rect 790 -870 800 -835
rect 835 -870 845 -835
rect 1035 -850 1045 -820
rect 1075 -850 1085 -820
rect 1035 -860 1085 -850
rect 1275 -820 1325 -810
rect 1275 -850 1285 -820
rect 1315 -850 1325 -820
rect 1275 -860 1325 -850
rect 1515 -820 1565 -810
rect 1515 -850 1525 -820
rect 1555 -850 1565 -820
rect 1515 -860 1565 -850
rect 1755 -820 1805 -810
rect 1755 -850 1765 -820
rect 1795 -850 1805 -820
rect 1755 -860 1805 -850
rect 1995 -820 2045 -810
rect 1995 -850 2005 -820
rect 2035 -850 2045 -820
rect 1995 -860 2045 -850
rect 2235 -820 2285 -810
rect 2235 -850 2245 -820
rect 2275 -850 2285 -820
rect 2235 -860 2285 -850
rect 2475 -820 2525 -810
rect 2475 -850 2485 -820
rect 2515 -850 2525 -820
rect 2475 -860 2525 -850
rect 2715 -820 2765 -810
rect 2715 -850 2725 -820
rect 2755 -850 2765 -820
rect 3195 -820 3245 -810
rect 2715 -860 2765 -850
rect 2950 -835 3005 -825
rect 790 -880 845 -870
rect 2950 -870 2960 -835
rect 2995 -870 3005 -835
rect 3195 -850 3205 -820
rect 3235 -850 3245 -820
rect 3195 -860 3245 -850
rect 3435 -820 3485 -810
rect 3435 -850 3445 -820
rect 3475 -850 3485 -820
rect 3435 -860 3485 -850
rect 3675 -820 3725 -810
rect 3675 -850 3685 -820
rect 3715 -850 3725 -820
rect 3675 -860 3725 -850
rect 3915 -820 3965 -810
rect 3915 -850 3925 -820
rect 3955 -850 3965 -820
rect 3915 -860 3965 -850
rect 4155 -820 4205 -810
rect 4155 -850 4165 -820
rect 4195 -850 4205 -820
rect 4155 -860 4205 -850
rect 4395 -820 4445 -810
rect 4395 -850 4405 -820
rect 4435 -850 4445 -820
rect 4395 -860 4445 -850
rect 4635 -820 4685 -810
rect 4635 -850 4645 -820
rect 4675 -850 4685 -820
rect 4635 -860 4685 -850
rect 4875 -820 4925 -810
rect 4875 -850 4885 -820
rect 4915 -850 4925 -820
rect 5355 -820 5405 -810
rect 4875 -860 4925 -850
rect 5110 -835 5165 -825
rect 2950 -880 3005 -870
rect 5110 -870 5120 -835
rect 5155 -870 5165 -835
rect 5355 -850 5365 -820
rect 5395 -850 5405 -820
rect 5355 -860 5405 -850
rect 5595 -820 5645 -810
rect 5595 -850 5605 -820
rect 5635 -850 5645 -820
rect 5595 -860 5645 -850
rect 5835 -820 5885 -810
rect 5835 -850 5845 -820
rect 5875 -850 5885 -820
rect 5835 -860 5885 -850
rect 6075 -820 6125 -810
rect 6075 -850 6085 -820
rect 6115 -850 6125 -820
rect 6075 -860 6125 -850
rect 6315 -820 6365 -810
rect 6315 -850 6325 -820
rect 6355 -850 6365 -820
rect 6315 -860 6365 -850
rect 6555 -820 6605 -810
rect 6555 -850 6565 -820
rect 6595 -850 6605 -820
rect 6555 -860 6605 -850
rect 6795 -820 6845 -810
rect 6795 -850 6805 -820
rect 6835 -850 6845 -820
rect 6795 -860 6845 -850
rect 7035 -820 7085 -810
rect 7035 -850 7045 -820
rect 7075 -850 7085 -820
rect 7515 -820 7565 -810
rect 7035 -860 7085 -850
rect 7270 -835 7325 -825
rect 5110 -880 5165 -870
rect 7270 -870 7280 -835
rect 7315 -870 7325 -835
rect 7515 -850 7525 -820
rect 7555 -850 7565 -820
rect 7515 -860 7565 -850
rect 7755 -820 7805 -810
rect 7755 -850 7765 -820
rect 7795 -850 7805 -820
rect 7755 -860 7805 -850
rect 7995 -820 8045 -810
rect 7995 -850 8005 -820
rect 8035 -850 8045 -820
rect 7995 -860 8045 -850
rect 8235 -820 8285 -810
rect 8235 -850 8245 -820
rect 8275 -850 8285 -820
rect 8235 -860 8285 -850
rect 8475 -820 8525 -810
rect 8475 -850 8485 -820
rect 8515 -850 8525 -820
rect 8475 -860 8525 -850
rect 8715 -820 8765 -810
rect 8715 -850 8725 -820
rect 8755 -850 8765 -820
rect 8715 -860 8765 -850
rect 8955 -820 9005 -810
rect 8955 -850 8965 -820
rect 8995 -850 9005 -820
rect 8955 -860 9005 -850
rect 9195 -820 9245 -810
rect 9195 -850 9205 -820
rect 9235 -850 9245 -820
rect 9675 -820 9725 -810
rect 9195 -860 9245 -850
rect 9430 -835 9485 -825
rect 7270 -880 7325 -870
rect 9430 -870 9440 -835
rect 9475 -870 9485 -835
rect 9675 -850 9685 -820
rect 9715 -850 9725 -820
rect 9675 -860 9725 -850
rect 9915 -820 9965 -810
rect 9915 -850 9925 -820
rect 9955 -850 9965 -820
rect 9915 -860 9965 -850
rect 10155 -820 10205 -810
rect 10155 -850 10165 -820
rect 10195 -850 10205 -820
rect 10155 -860 10205 -850
rect 10395 -820 10445 -810
rect 10395 -850 10405 -820
rect 10435 -850 10445 -820
rect 10395 -860 10445 -850
rect 10635 -820 10685 -810
rect 10635 -850 10645 -820
rect 10675 -850 10685 -820
rect 10635 -860 10685 -850
rect 10875 -820 10925 -810
rect 10875 -850 10885 -820
rect 10915 -850 10925 -820
rect 10875 -860 10925 -850
rect 11115 -820 11165 -810
rect 11115 -850 11125 -820
rect 11155 -850 11165 -820
rect 11115 -860 11165 -850
rect 11355 -820 11405 -810
rect 11355 -850 11365 -820
rect 11395 -850 11405 -820
rect 11835 -820 11885 -810
rect 11355 -860 11405 -850
rect 11590 -835 11645 -825
rect 9430 -880 9485 -870
rect 11590 -870 11600 -835
rect 11635 -870 11645 -835
rect 11835 -850 11845 -820
rect 11875 -850 11885 -820
rect 11835 -860 11885 -850
rect 12075 -820 12125 -810
rect 12075 -850 12085 -820
rect 12115 -850 12125 -820
rect 12075 -860 12125 -850
rect 12315 -820 12365 -810
rect 12315 -850 12325 -820
rect 12355 -850 12365 -820
rect 12315 -860 12365 -850
rect 12555 -820 12605 -810
rect 12555 -850 12565 -820
rect 12595 -850 12605 -820
rect 12555 -860 12605 -850
rect 12795 -820 12845 -810
rect 12795 -850 12805 -820
rect 12835 -850 12845 -820
rect 12795 -860 12845 -850
rect 13035 -820 13085 -810
rect 13035 -850 13045 -820
rect 13075 -850 13085 -820
rect 13035 -860 13085 -850
rect 13275 -820 13325 -810
rect 13275 -850 13285 -820
rect 13315 -850 13325 -820
rect 13275 -860 13325 -850
rect 13515 -820 13565 -810
rect 13515 -850 13525 -820
rect 13555 -850 13565 -820
rect 13995 -820 14045 -810
rect 13515 -860 13565 -850
rect 13750 -835 13805 -825
rect 11590 -880 11645 -870
rect 13750 -870 13760 -835
rect 13795 -870 13805 -835
rect 13995 -850 14005 -820
rect 14035 -850 14045 -820
rect 13995 -860 14045 -850
rect 14235 -820 14285 -810
rect 14235 -850 14245 -820
rect 14275 -850 14285 -820
rect 14235 -860 14285 -850
rect 14475 -820 14525 -810
rect 14475 -850 14485 -820
rect 14515 -850 14525 -820
rect 14475 -860 14525 -850
rect 14715 -820 14765 -810
rect 14715 -850 14725 -820
rect 14755 -850 14765 -820
rect 14715 -860 14765 -850
rect 14955 -820 15005 -810
rect 14955 -850 14965 -820
rect 14995 -850 15005 -820
rect 14955 -860 15005 -850
rect 15195 -820 15245 -810
rect 15195 -850 15205 -820
rect 15235 -850 15245 -820
rect 15195 -860 15245 -850
rect 15435 -820 15485 -810
rect 15435 -850 15445 -820
rect 15475 -850 15485 -820
rect 15435 -860 15485 -850
rect 15675 -820 15725 -810
rect 15675 -850 15685 -820
rect 15715 -850 15725 -820
rect 16155 -820 16205 -810
rect 15675 -860 15725 -850
rect 15910 -835 15965 -825
rect 13750 -880 13805 -870
rect 15910 -870 15920 -835
rect 15955 -870 15965 -835
rect 16155 -850 16165 -820
rect 16195 -850 16205 -820
rect 16155 -860 16205 -850
rect 16395 -820 16445 -810
rect 16395 -850 16405 -820
rect 16435 -850 16445 -820
rect 16395 -860 16445 -850
rect 16635 -820 16685 -810
rect 16635 -850 16645 -820
rect 16675 -850 16685 -820
rect 16635 -860 16685 -850
rect 16875 -820 16925 -810
rect 16875 -850 16885 -820
rect 16915 -850 16925 -820
rect 16875 -860 16925 -850
rect 17115 -820 17165 -810
rect 17115 -850 17125 -820
rect 17155 -850 17165 -820
rect 17115 -860 17165 -850
rect 17355 -820 17405 -810
rect 17355 -850 17365 -820
rect 17395 -850 17405 -820
rect 17355 -860 17405 -850
rect 17595 -820 17645 -810
rect 17595 -850 17605 -820
rect 17635 -850 17645 -820
rect 17595 -860 17645 -850
rect 17835 -820 17885 -810
rect 17835 -850 17845 -820
rect 17875 -850 17885 -820
rect 18315 -820 18365 -810
rect 17835 -860 17885 -850
rect 18070 -835 18125 -825
rect 15910 -880 15965 -870
rect 18070 -870 18080 -835
rect 18115 -870 18125 -835
rect 18315 -850 18325 -820
rect 18355 -850 18365 -820
rect 18315 -860 18365 -850
rect 18555 -820 18605 -810
rect 18555 -850 18565 -820
rect 18595 -850 18605 -820
rect 18555 -860 18605 -850
rect 18795 -820 18845 -810
rect 18795 -850 18805 -820
rect 18835 -850 18845 -820
rect 18795 -860 18845 -850
rect 19035 -820 19085 -810
rect 19035 -850 19045 -820
rect 19075 -850 19085 -820
rect 19035 -860 19085 -850
rect 19275 -820 19325 -810
rect 19275 -850 19285 -820
rect 19315 -850 19325 -820
rect 19275 -860 19325 -850
rect 19515 -820 19565 -810
rect 19515 -850 19525 -820
rect 19555 -850 19565 -820
rect 19515 -860 19565 -850
rect 19755 -820 19805 -810
rect 19755 -850 19765 -820
rect 19795 -850 19805 -820
rect 19755 -860 19805 -850
rect 19995 -820 20045 -810
rect 19995 -850 20005 -820
rect 20035 -850 20045 -820
rect 20475 -820 20525 -810
rect 19995 -860 20045 -850
rect 20230 -835 20285 -825
rect 18070 -880 18125 -870
rect 20230 -870 20240 -835
rect 20275 -870 20285 -835
rect 20475 -850 20485 -820
rect 20515 -850 20525 -820
rect 20475 -860 20525 -850
rect 20715 -820 20765 -810
rect 20715 -850 20725 -820
rect 20755 -850 20765 -820
rect 20715 -860 20765 -850
rect 20955 -820 21005 -810
rect 20955 -850 20965 -820
rect 20995 -850 21005 -820
rect 20955 -860 21005 -850
rect 21195 -820 21245 -810
rect 21195 -850 21205 -820
rect 21235 -850 21245 -820
rect 21195 -860 21245 -850
rect 21435 -820 21485 -810
rect 21435 -850 21445 -820
rect 21475 -850 21485 -820
rect 21435 -860 21485 -850
rect 21675 -820 21725 -810
rect 21675 -850 21685 -820
rect 21715 -850 21725 -820
rect 21675 -860 21725 -850
rect 21915 -820 21965 -810
rect 21915 -850 21925 -820
rect 21955 -850 21965 -820
rect 21915 -860 21965 -850
rect 22155 -820 22205 -810
rect 22155 -850 22165 -820
rect 22195 -850 22205 -820
rect 22635 -820 22685 -810
rect 22155 -860 22205 -850
rect 22390 -835 22445 -825
rect 20230 -880 20285 -870
rect 22390 -870 22400 -835
rect 22435 -870 22445 -835
rect 22635 -850 22645 -820
rect 22675 -850 22685 -820
rect 22635 -860 22685 -850
rect 22875 -820 22925 -810
rect 22875 -850 22885 -820
rect 22915 -850 22925 -820
rect 22875 -860 22925 -850
rect 23115 -820 23165 -810
rect 23115 -850 23125 -820
rect 23155 -850 23165 -820
rect 23115 -860 23165 -850
rect 23355 -820 23405 -810
rect 23355 -850 23365 -820
rect 23395 -850 23405 -820
rect 23355 -860 23405 -850
rect 23595 -820 23645 -810
rect 23595 -850 23605 -820
rect 23635 -850 23645 -820
rect 23595 -860 23645 -850
rect 23835 -820 23885 -810
rect 23835 -850 23845 -820
rect 23875 -850 23885 -820
rect 23835 -860 23885 -850
rect 24075 -820 24125 -810
rect 24075 -850 24085 -820
rect 24115 -850 24125 -820
rect 24555 -820 24605 -810
rect 24075 -860 24125 -850
rect 24310 -835 24365 -825
rect 22390 -880 22445 -870
rect 24310 -870 24320 -835
rect 24355 -870 24365 -835
rect 24555 -850 24565 -820
rect 24595 -850 24605 -820
rect 24555 -860 24605 -850
rect 24795 -820 24845 -810
rect 24795 -850 24805 -820
rect 24835 -850 24845 -820
rect 24795 -860 24845 -850
rect 25035 -820 25085 -810
rect 25035 -850 25045 -820
rect 25075 -850 25085 -820
rect 25035 -860 25085 -850
rect 25275 -820 25325 -810
rect 25275 -850 25285 -820
rect 25315 -850 25325 -820
rect 25275 -860 25325 -850
rect 25515 -820 25565 -810
rect 25515 -850 25525 -820
rect 25555 -850 25565 -820
rect 25515 -860 25565 -850
rect 25755 -820 25805 -810
rect 25755 -850 25765 -820
rect 25795 -850 25805 -820
rect 25755 -860 25805 -850
rect 25995 -820 26045 -810
rect 25995 -850 26005 -820
rect 26035 -850 26045 -820
rect 26475 -820 26525 -810
rect 25995 -860 26045 -850
rect 26230 -835 26285 -825
rect 24310 -880 24365 -870
rect 26230 -870 26240 -835
rect 26275 -870 26285 -835
rect 26475 -850 26485 -820
rect 26515 -850 26525 -820
rect 26475 -860 26525 -850
rect 26715 -820 26765 -810
rect 26715 -850 26725 -820
rect 26755 -850 26765 -820
rect 26715 -860 26765 -850
rect 26955 -820 27005 -810
rect 26955 -850 26965 -820
rect 26995 -850 27005 -820
rect 26955 -860 27005 -850
rect 27195 -820 27245 -810
rect 27195 -850 27205 -820
rect 27235 -850 27245 -820
rect 27195 -860 27245 -850
rect 27435 -820 27485 -810
rect 27435 -850 27445 -820
rect 27475 -850 27485 -820
rect 27435 -860 27485 -850
rect 27675 -820 27725 -810
rect 27675 -850 27685 -820
rect 27715 -850 27725 -820
rect 27675 -860 27725 -850
rect 27915 -820 27965 -810
rect 27915 -850 27925 -820
rect 27955 -850 27965 -820
rect 28395 -820 28445 -810
rect 27915 -860 27965 -850
rect 28150 -835 28205 -825
rect 26230 -880 26285 -870
rect 28150 -870 28160 -835
rect 28195 -870 28205 -835
rect 28395 -850 28405 -820
rect 28435 -850 28445 -820
rect 28395 -860 28445 -850
rect 28635 -820 28685 -810
rect 28635 -850 28645 -820
rect 28675 -850 28685 -820
rect 28635 -860 28685 -850
rect 28875 -820 28925 -810
rect 28875 -850 28885 -820
rect 28915 -850 28925 -820
rect 28875 -860 28925 -850
rect 29115 -820 29165 -810
rect 29115 -850 29125 -820
rect 29155 -850 29165 -820
rect 29115 -860 29165 -850
rect 29355 -820 29405 -810
rect 29355 -850 29365 -820
rect 29395 -850 29405 -820
rect 29355 -860 29405 -850
rect 29595 -820 29645 -810
rect 29595 -850 29605 -820
rect 29635 -850 29645 -820
rect 30075 -820 30125 -810
rect 29595 -860 29645 -850
rect 29830 -835 29885 -825
rect 28150 -880 28205 -870
rect 29830 -870 29840 -835
rect 29875 -870 29885 -835
rect 30075 -850 30085 -820
rect 30115 -850 30125 -820
rect 30075 -860 30125 -850
rect 30315 -820 30365 -810
rect 30315 -850 30325 -820
rect 30355 -850 30365 -820
rect 30315 -860 30365 -850
rect 30555 -820 30605 -810
rect 30555 -850 30565 -820
rect 30595 -850 30605 -820
rect 30555 -860 30605 -850
rect 29830 -880 29885 -870
<< via2 >>
rect 195 240 230 275
rect 436 235 466 265
rect 741 235 771 265
rect 986 235 1016 265
rect 1226 235 1256 265
rect 1471 235 1501 265
rect 1776 235 1806 265
rect 2021 235 2051 265
rect 2265 270 2300 305
rect 2506 235 2536 265
rect 2746 235 2776 265
rect 2991 235 3021 265
rect 3231 235 3261 265
rect 3476 235 3506 265
rect 3716 235 3746 265
rect 3961 235 3991 265
rect 4205 270 4240 305
rect 4446 235 4476 265
rect 4686 235 4716 265
rect 4931 235 4961 265
rect 5171 235 5201 265
rect 5416 235 5446 265
rect 5721 235 5751 265
rect 5966 235 5996 265
rect 6206 235 6236 265
rect 6455 270 6490 305
rect 6691 235 6721 265
rect 6936 235 6966 265
rect 7176 235 7206 265
rect 7416 235 7446 265
rect 7656 235 7686 265
rect 7901 235 7931 265
rect 8141 235 8171 265
rect 8386 235 8416 265
rect 8626 235 8656 265
rect 8871 235 8901 265
rect 9111 235 9141 265
rect 9360 270 9395 305
rect 9601 235 9631 265
rect 9846 235 9876 265
rect 10086 235 10116 265
rect 10331 235 10361 265
rect 10571 235 10601 265
rect 10816 235 10846 265
rect 11056 235 11086 265
rect 11305 270 11340 305
rect 11541 235 11571 265
rect 11786 235 11816 265
rect 12026 235 12056 265
rect 12271 235 12301 265
rect 12511 235 12541 265
rect 12756 235 12786 265
rect 13000 270 13035 305
rect 13241 235 13271 265
rect 13481 235 13511 265
rect 13726 235 13756 265
rect 13966 235 13996 265
rect 14211 235 14241 265
rect 14451 235 14481 265
rect 14696 235 14726 265
rect 14936 235 14966 265
rect 15185 270 15220 305
rect 15421 235 15451 265
rect 15666 235 15696 265
rect 15906 235 15936 265
rect 16151 235 16181 265
rect 16391 235 16421 265
rect 16636 235 16666 265
rect 16876 235 16906 265
rect 17121 235 17151 265
rect 17365 270 17400 305
rect 17606 235 17636 265
rect 17846 235 17876 265
rect 18091 235 18121 265
rect 18331 235 18361 265
rect 18576 235 18606 265
rect 18816 235 18846 265
rect 19061 235 19091 265
rect 19301 235 19331 265
rect 19550 270 19585 305
rect 19786 235 19816 265
rect 20031 235 20061 265
rect 20271 235 20301 265
rect 20516 235 20546 265
rect 20760 270 20795 305
rect 21001 235 21031 265
rect -415 -240 -365 -190
rect 186 -195 216 -165
rect 431 -195 461 -165
rect 736 -195 766 -165
rect 981 -195 1011 -165
rect 1221 -195 1251 -165
rect 1466 -195 1496 -165
rect 90 -275 120 -245
rect 330 -275 360 -245
rect 570 -275 600 -245
rect 810 -275 840 -245
rect 1050 -275 1080 -245
rect 1290 -275 1320 -245
rect 1530 -275 1560 -245
rect 1635 -240 1675 -200
rect 1771 -195 1801 -165
rect 2016 -195 2046 -165
rect 2256 -195 2286 -165
rect 2501 -195 2531 -165
rect 2741 -195 2771 -165
rect 2986 -195 3016 -165
rect 3226 -195 3256 -165
rect 3471 -195 3501 -165
rect 3711 -195 3741 -165
rect 3956 -195 3986 -165
rect 4060 -235 4100 -195
rect 4196 -195 4226 -165
rect 4441 -195 4471 -165
rect 4681 -195 4711 -165
rect 4926 -195 4956 -165
rect 5166 -195 5196 -165
rect 5411 -195 5441 -165
rect 5716 -195 5746 -165
rect 5961 -195 5991 -165
rect 6201 -195 6231 -165
rect 6686 -195 6716 -165
rect 6931 -195 6961 -165
rect 7171 -195 7201 -165
rect 7411 -195 7441 -165
rect 7651 -195 7681 -165
rect 8136 -195 8166 -165
rect 8381 -195 8411 -165
rect 8621 -195 8651 -165
rect 8866 -195 8896 -165
rect 9106 -195 9136 -165
rect 9351 -195 9381 -165
rect 9841 -195 9871 -165
rect 10081 -195 10111 -165
rect 10326 -195 10356 -165
rect 10566 -195 10596 -165
rect 10811 -195 10841 -165
rect 11051 -195 11081 -165
rect 11296 -195 11326 -165
rect 11536 -195 11566 -165
rect 11781 -195 11811 -165
rect 12266 -195 12296 -165
rect 12506 -195 12536 -165
rect 12751 -195 12781 -165
rect 12991 -195 13021 -165
rect 13236 -195 13266 -165
rect 13476 -195 13506 -165
rect 13721 -195 13751 -165
rect 14206 -195 14236 -165
rect 14446 -195 14476 -165
rect 14691 -195 14721 -165
rect 14931 -195 14961 -165
rect 15176 -195 15206 -165
rect 15416 -195 15446 -165
rect 15661 -195 15691 -165
rect 16146 -195 16176 -165
rect 16386 -195 16416 -165
rect 16631 -195 16661 -165
rect 16871 -195 16901 -165
rect 17116 -195 17146 -165
rect 17356 -195 17386 -165
rect 17601 -195 17631 -165
rect 17841 -195 17871 -165
rect 18086 -195 18116 -165
rect 18326 -195 18356 -165
rect 18571 -195 18601 -165
rect 18811 -195 18841 -165
rect 19056 -195 19086 -165
rect 19296 -195 19326 -165
rect 19541 -195 19571 -165
rect 19781 -195 19811 -165
rect 1770 -275 1800 -245
rect 2010 -275 2040 -245
rect 2250 -275 2280 -245
rect 2490 -275 2520 -245
rect 2730 -275 2760 -245
rect 2970 -275 3000 -245
rect 3210 -275 3240 -245
rect 3450 -275 3480 -245
rect 3690 -275 3720 -245
rect 3930 -275 3960 -245
rect 4170 -275 4200 -245
rect 4410 -275 4440 -245
rect 4650 -275 4680 -245
rect 4890 -275 4920 -245
rect 5130 -275 5160 -245
rect 5370 -275 5400 -245
rect 5610 -275 5640 -245
rect 5850 -275 5880 -245
rect 6090 -275 6120 -245
rect 6330 -275 6360 -245
rect 6455 -260 6495 -220
rect 6570 -275 6600 -245
rect 6810 -275 6840 -245
rect 7050 -275 7080 -245
rect 7290 -275 7320 -245
rect 7530 -275 7560 -245
rect 7770 -275 7800 -245
rect 7880 -260 7920 -220
rect 8010 -275 8040 -245
rect 8250 -275 8280 -245
rect 8490 -275 8520 -245
rect 8730 -275 8760 -245
rect 8970 -275 9000 -245
rect 9210 -275 9240 -245
rect 9450 -275 9480 -245
rect 9570 -250 9610 -210
rect 9690 -275 9720 -245
rect 9930 -275 9960 -245
rect 10170 -275 10200 -245
rect 10410 -275 10440 -245
rect 10650 -275 10680 -245
rect 10890 -275 10920 -245
rect 11130 -275 11160 -245
rect 11370 -275 11400 -245
rect 11610 -275 11640 -245
rect 11850 -275 11880 -245
rect 11950 -260 11990 -220
rect 12090 -275 12120 -245
rect 12330 -275 12360 -245
rect 12570 -275 12600 -245
rect 12810 -275 12840 -245
rect 13050 -275 13080 -245
rect 13290 -275 13320 -245
rect 13530 -275 13560 -245
rect 13770 -275 13800 -245
rect 13870 -260 13910 -220
rect 14010 -275 14040 -245
rect 14250 -275 14280 -245
rect 14490 -275 14520 -245
rect 14730 -275 14760 -245
rect 14970 -275 15000 -245
rect 15210 -275 15240 -245
rect 15450 -275 15480 -245
rect 15690 -275 15720 -245
rect 15815 -260 15855 -220
rect 15930 -275 15960 -245
rect 16170 -275 16200 -245
rect 16410 -275 16440 -245
rect 16650 -275 16680 -245
rect 16890 -275 16920 -245
rect 17130 -275 17160 -245
rect 17370 -275 17400 -245
rect 17610 -275 17640 -245
rect 17705 -250 17745 -210
rect 20026 -195 20056 -165
rect 20266 -195 20296 -165
rect 20511 -195 20541 -165
rect 20751 -195 20781 -165
rect 20996 -195 21026 -165
rect 17850 -275 17880 -245
rect 18090 -275 18120 -245
rect 18330 -275 18360 -245
rect 18570 -275 18600 -245
rect 18810 -275 18840 -245
rect 19050 -275 19080 -245
rect 19290 -275 19320 -245
rect 19530 -275 19560 -245
rect 19645 -250 19685 -210
rect 19770 -275 19800 -245
rect 20010 -275 20040 -245
rect 20250 -275 20280 -245
rect 20490 -275 20520 -245
rect 20730 -275 20760 -245
rect 20970 -275 21000 -245
rect 21210 -275 21240 -245
rect 21450 -275 21480 -245
rect 21690 -275 21720 -245
rect 21930 -275 21960 -245
rect 22170 -275 22200 -245
rect 22410 -275 22440 -245
rect 22650 -275 22680 -245
rect 22890 -275 22920 -245
rect 23130 -275 23160 -245
rect 23370 -275 23400 -245
rect 23610 -275 23640 -245
rect 23850 -275 23880 -245
rect 24090 -275 24120 -245
rect 24330 -275 24360 -245
rect 24570 -275 24600 -245
rect 24810 -275 24840 -245
rect 25050 -275 25080 -245
rect 25290 -275 25320 -245
rect 25530 -275 25560 -245
rect 25770 -275 25800 -245
rect 26010 -275 26040 -245
rect 26250 -275 26280 -245
rect 26490 -275 26520 -245
rect 26730 -275 26760 -245
rect 26970 -275 27000 -245
rect 27210 -275 27240 -245
rect 27450 -275 27480 -245
rect 27690 -275 27720 -245
rect 27930 -275 27960 -245
rect 28170 -275 28200 -245
rect 28410 -275 28440 -245
rect 28650 -275 28680 -245
rect 28890 -275 28920 -245
rect 29130 -275 29160 -245
rect 29370 -275 29400 -245
rect 29610 -275 29640 -245
rect 29850 -275 29880 -245
rect 30090 -275 30120 -245
rect 30330 -275 30360 -245
rect 30570 -275 30600 -245
rect 85 -850 115 -820
rect 325 -850 355 -820
rect 565 -850 595 -820
rect 800 -870 835 -835
rect 1045 -850 1075 -820
rect 1285 -850 1315 -820
rect 1525 -850 1555 -820
rect 1765 -850 1795 -820
rect 2005 -850 2035 -820
rect 2245 -850 2275 -820
rect 2485 -850 2515 -820
rect 2725 -850 2755 -820
rect 2960 -870 2995 -835
rect 3205 -850 3235 -820
rect 3445 -850 3475 -820
rect 3685 -850 3715 -820
rect 3925 -850 3955 -820
rect 4165 -850 4195 -820
rect 4405 -850 4435 -820
rect 4645 -850 4675 -820
rect 4885 -850 4915 -820
rect 5120 -870 5155 -835
rect 5365 -850 5395 -820
rect 5605 -850 5635 -820
rect 5845 -850 5875 -820
rect 6085 -850 6115 -820
rect 6325 -850 6355 -820
rect 6565 -850 6595 -820
rect 6805 -850 6835 -820
rect 7045 -850 7075 -820
rect 7280 -870 7315 -835
rect 7525 -850 7555 -820
rect 7765 -850 7795 -820
rect 8005 -850 8035 -820
rect 8245 -850 8275 -820
rect 8485 -850 8515 -820
rect 8725 -850 8755 -820
rect 8965 -850 8995 -820
rect 9205 -850 9235 -820
rect 9440 -870 9475 -835
rect 9685 -850 9715 -820
rect 9925 -850 9955 -820
rect 10165 -850 10195 -820
rect 10405 -850 10435 -820
rect 10645 -850 10675 -820
rect 10885 -850 10915 -820
rect 11125 -850 11155 -820
rect 11365 -850 11395 -820
rect 11600 -870 11635 -835
rect 11845 -850 11875 -820
rect 12085 -850 12115 -820
rect 12325 -850 12355 -820
rect 12565 -850 12595 -820
rect 12805 -850 12835 -820
rect 13045 -850 13075 -820
rect 13285 -850 13315 -820
rect 13525 -850 13555 -820
rect 13760 -870 13795 -835
rect 14005 -850 14035 -820
rect 14245 -850 14275 -820
rect 14485 -850 14515 -820
rect 14725 -850 14755 -820
rect 14965 -850 14995 -820
rect 15205 -850 15235 -820
rect 15445 -850 15475 -820
rect 15685 -850 15715 -820
rect 15920 -870 15955 -835
rect 16165 -850 16195 -820
rect 16405 -850 16435 -820
rect 16645 -850 16675 -820
rect 16885 -850 16915 -820
rect 17125 -850 17155 -820
rect 17365 -850 17395 -820
rect 17605 -850 17635 -820
rect 17845 -850 17875 -820
rect 18080 -870 18115 -835
rect 18325 -850 18355 -820
rect 18565 -850 18595 -820
rect 18805 -850 18835 -820
rect 19045 -850 19075 -820
rect 19285 -850 19315 -820
rect 19525 -850 19555 -820
rect 19765 -850 19795 -820
rect 20005 -850 20035 -820
rect 20240 -870 20275 -835
rect 20485 -850 20515 -820
rect 20725 -850 20755 -820
rect 20965 -850 20995 -820
rect 21205 -850 21235 -820
rect 21445 -850 21475 -820
rect 21685 -850 21715 -820
rect 21925 -850 21955 -820
rect 22165 -850 22195 -820
rect 22400 -870 22435 -835
rect 22645 -850 22675 -820
rect 22885 -850 22915 -820
rect 23125 -850 23155 -820
rect 23365 -850 23395 -820
rect 23605 -850 23635 -820
rect 23845 -850 23875 -820
rect 24085 -850 24115 -820
rect 24320 -870 24355 -835
rect 24565 -850 24595 -820
rect 24805 -850 24835 -820
rect 25045 -850 25075 -820
rect 25285 -850 25315 -820
rect 25525 -850 25555 -820
rect 25765 -850 25795 -820
rect 26005 -850 26035 -820
rect 26240 -870 26275 -835
rect 26485 -850 26515 -820
rect 26725 -850 26755 -820
rect 26965 -850 26995 -820
rect 27205 -850 27235 -820
rect 27445 -850 27475 -820
rect 27685 -850 27715 -820
rect 27925 -850 27955 -820
rect 28160 -870 28195 -835
rect 28405 -850 28435 -820
rect 28645 -850 28675 -820
rect 28885 -850 28915 -820
rect 29125 -850 29155 -820
rect 29365 -850 29395 -820
rect 29605 -850 29635 -820
rect 29840 -870 29875 -835
rect 30085 -850 30115 -820
rect 30325 -850 30355 -820
rect 30565 -850 30595 -820
<< metal3 >>
rect 2255 305 2310 315
rect 185 275 240 285
rect 185 240 195 275
rect 230 240 240 275
rect 185 230 240 240
rect 426 270 476 275
rect 426 230 431 270
rect 471 230 476 270
rect 426 225 476 230
rect 731 270 781 275
rect 731 230 736 270
rect 776 230 781 270
rect 731 225 781 230
rect 976 270 1026 275
rect 976 230 981 270
rect 1021 230 1026 270
rect 976 225 1026 230
rect 1216 270 1266 275
rect 1216 230 1221 270
rect 1261 230 1266 270
rect 1216 225 1266 230
rect 1461 270 1511 275
rect 1461 230 1466 270
rect 1506 230 1511 270
rect 1461 225 1511 230
rect 1766 270 1816 275
rect 1766 230 1771 270
rect 1811 230 1816 270
rect 1766 225 1816 230
rect 2011 270 2061 275
rect 2011 230 2016 270
rect 2056 230 2061 270
rect 2255 270 2265 305
rect 2300 270 2310 305
rect 4195 305 4250 315
rect 2255 260 2310 270
rect 2496 270 2546 275
rect 2011 225 2061 230
rect 2496 230 2501 270
rect 2541 230 2546 270
rect 2496 225 2546 230
rect 2736 270 2786 275
rect 2736 230 2741 270
rect 2781 230 2786 270
rect 2736 225 2786 230
rect 2981 270 3031 275
rect 2981 230 2986 270
rect 3026 230 3031 270
rect 2981 225 3031 230
rect 3221 270 3271 275
rect 3221 230 3226 270
rect 3266 230 3271 270
rect 3221 225 3271 230
rect 3466 270 3516 275
rect 3466 230 3471 270
rect 3511 230 3516 270
rect 3466 225 3516 230
rect 3706 270 3756 275
rect 3706 230 3711 270
rect 3751 230 3756 270
rect 3706 225 3756 230
rect 3951 270 4001 275
rect 3951 230 3956 270
rect 3996 230 4001 270
rect 4195 270 4205 305
rect 4240 270 4250 305
rect 6445 305 6500 315
rect 4195 260 4250 270
rect 4436 270 4486 275
rect 3951 225 4001 230
rect 4436 230 4441 270
rect 4481 230 4486 270
rect 4436 225 4486 230
rect 4676 270 4726 275
rect 4676 230 4681 270
rect 4721 230 4726 270
rect 4676 225 4726 230
rect 4921 270 4971 275
rect 4921 230 4926 270
rect 4966 230 4971 270
rect 4921 225 4971 230
rect 5161 270 5211 275
rect 5161 230 5166 270
rect 5206 230 5211 270
rect 5161 225 5211 230
rect 5406 270 5456 275
rect 5406 230 5411 270
rect 5451 230 5456 270
rect 5406 225 5456 230
rect 5711 270 5761 275
rect 5711 230 5716 270
rect 5756 230 5761 270
rect 5711 225 5761 230
rect 5956 270 6006 275
rect 5956 230 5961 270
rect 6001 230 6006 270
rect 5956 225 6006 230
rect 6196 270 6246 275
rect 6196 230 6201 270
rect 6241 230 6246 270
rect 6445 270 6455 305
rect 6490 270 6500 305
rect 9350 305 9405 315
rect 6445 260 6500 270
rect 6681 270 6731 275
rect 6196 225 6246 230
rect 6681 230 6686 270
rect 6726 230 6731 270
rect 6681 225 6731 230
rect 6926 270 6976 275
rect 6926 230 6931 270
rect 6971 230 6976 270
rect 6926 225 6976 230
rect 7166 270 7216 275
rect 7166 230 7171 270
rect 7211 230 7216 270
rect 7166 225 7216 230
rect 7406 270 7456 275
rect 7406 230 7411 270
rect 7451 230 7456 270
rect 7406 225 7456 230
rect 7646 270 7696 275
rect 7646 230 7651 270
rect 7691 230 7696 270
rect 7646 225 7696 230
rect 7891 270 7941 275
rect 7891 230 7896 270
rect 7936 230 7941 270
rect 7891 225 7941 230
rect 8131 270 8181 275
rect 8131 230 8136 270
rect 8176 230 8181 270
rect 8131 225 8181 230
rect 8376 270 8426 275
rect 8376 230 8381 270
rect 8421 230 8426 270
rect 8376 225 8426 230
rect 8616 270 8666 275
rect 8616 230 8621 270
rect 8661 230 8666 270
rect 8616 225 8666 230
rect 8861 270 8911 275
rect 8861 230 8866 270
rect 8906 230 8911 270
rect 8861 225 8911 230
rect 9101 270 9151 275
rect 9101 230 9106 270
rect 9146 230 9151 270
rect 9350 270 9360 305
rect 9395 270 9405 305
rect 11295 305 11350 315
rect 9350 260 9405 270
rect 9591 270 9641 275
rect 9101 225 9151 230
rect 9591 230 9596 270
rect 9636 230 9641 270
rect 9591 225 9641 230
rect 9836 270 9886 275
rect 9836 230 9841 270
rect 9881 230 9886 270
rect 9836 225 9886 230
rect 10076 270 10126 275
rect 10076 230 10081 270
rect 10121 230 10126 270
rect 10076 225 10126 230
rect 10321 270 10371 275
rect 10321 230 10326 270
rect 10366 230 10371 270
rect 10321 225 10371 230
rect 10561 270 10611 275
rect 10561 230 10566 270
rect 10606 230 10611 270
rect 10561 225 10611 230
rect 10806 270 10856 275
rect 10806 230 10811 270
rect 10851 230 10856 270
rect 10806 225 10856 230
rect 11046 270 11096 275
rect 11046 230 11051 270
rect 11091 230 11096 270
rect 11295 270 11305 305
rect 11340 270 11350 305
rect 12990 305 13045 315
rect 11295 260 11350 270
rect 11531 270 11581 275
rect 11046 225 11096 230
rect 11531 230 11536 270
rect 11576 230 11581 270
rect 11531 225 11581 230
rect 11776 270 11826 275
rect 11776 230 11781 270
rect 11821 230 11826 270
rect 11776 225 11826 230
rect 12016 270 12066 275
rect 12016 230 12021 270
rect 12061 230 12066 270
rect 12016 225 12066 230
rect 12261 270 12311 275
rect 12261 230 12266 270
rect 12306 230 12311 270
rect 12261 225 12311 230
rect 12501 270 12551 275
rect 12501 230 12506 270
rect 12546 230 12551 270
rect 12501 225 12551 230
rect 12746 270 12796 275
rect 12746 230 12751 270
rect 12791 230 12796 270
rect 12990 270 13000 305
rect 13035 270 13045 305
rect 15175 305 15230 315
rect 12990 260 13045 270
rect 13231 270 13281 275
rect 12746 225 12796 230
rect 13231 230 13236 270
rect 13276 230 13281 270
rect 13231 225 13281 230
rect 13471 270 13521 275
rect 13471 230 13476 270
rect 13516 230 13521 270
rect 13471 225 13521 230
rect 13716 270 13766 275
rect 13716 230 13721 270
rect 13761 230 13766 270
rect 13716 225 13766 230
rect 13956 270 14006 275
rect 13956 230 13961 270
rect 14001 230 14006 270
rect 13956 225 14006 230
rect 14201 270 14251 275
rect 14201 230 14206 270
rect 14246 230 14251 270
rect 14201 225 14251 230
rect 14441 270 14491 275
rect 14441 230 14446 270
rect 14486 230 14491 270
rect 14441 225 14491 230
rect 14686 270 14736 275
rect 14686 230 14691 270
rect 14731 230 14736 270
rect 14686 225 14736 230
rect 14926 270 14976 275
rect 14926 230 14931 270
rect 14971 230 14976 270
rect 15175 270 15185 305
rect 15220 270 15230 305
rect 17355 305 17410 315
rect 15175 260 15230 270
rect 15411 270 15461 275
rect 14926 225 14976 230
rect 15411 230 15416 270
rect 15456 230 15461 270
rect 15411 225 15461 230
rect 15656 270 15706 275
rect 15656 230 15661 270
rect 15701 230 15706 270
rect 15656 225 15706 230
rect 15896 270 15946 275
rect 15896 230 15901 270
rect 15941 230 15946 270
rect 15896 225 15946 230
rect 16141 270 16191 275
rect 16141 230 16146 270
rect 16186 230 16191 270
rect 16141 225 16191 230
rect 16381 270 16431 275
rect 16381 230 16386 270
rect 16426 230 16431 270
rect 16381 225 16431 230
rect 16626 270 16676 275
rect 16626 230 16631 270
rect 16671 230 16676 270
rect 16626 225 16676 230
rect 16866 270 16916 275
rect 16866 230 16871 270
rect 16911 230 16916 270
rect 16866 225 16916 230
rect 17111 270 17161 275
rect 17111 230 17116 270
rect 17156 230 17161 270
rect 17355 270 17365 305
rect 17400 270 17410 305
rect 19540 305 19595 315
rect 17355 260 17410 270
rect 17596 270 17646 275
rect 17111 225 17161 230
rect 17596 230 17601 270
rect 17641 230 17646 270
rect 17596 225 17646 230
rect 17836 270 17886 275
rect 17836 230 17841 270
rect 17881 230 17886 270
rect 17836 225 17886 230
rect 18081 270 18131 275
rect 18081 230 18086 270
rect 18126 230 18131 270
rect 18081 225 18131 230
rect 18321 270 18371 275
rect 18321 230 18326 270
rect 18366 230 18371 270
rect 18321 225 18371 230
rect 18566 270 18616 275
rect 18566 230 18571 270
rect 18611 230 18616 270
rect 18566 225 18616 230
rect 18806 270 18856 275
rect 18806 230 18811 270
rect 18851 230 18856 270
rect 18806 225 18856 230
rect 19051 270 19101 275
rect 19051 230 19056 270
rect 19096 230 19101 270
rect 19051 225 19101 230
rect 19291 270 19341 275
rect 19291 230 19296 270
rect 19336 230 19341 270
rect 19540 270 19550 305
rect 19585 270 19595 305
rect 20750 305 20805 315
rect 19540 260 19595 270
rect 19776 270 19826 275
rect 19291 225 19341 230
rect 19776 230 19781 270
rect 19821 230 19826 270
rect 19776 225 19826 230
rect 20021 270 20071 275
rect 20021 230 20026 270
rect 20066 230 20071 270
rect 20021 225 20071 230
rect 20261 270 20311 275
rect 20261 230 20266 270
rect 20306 230 20311 270
rect 20261 225 20311 230
rect 20506 270 20556 275
rect 20506 230 20511 270
rect 20551 230 20556 270
rect 20750 270 20760 305
rect 20795 270 20805 305
rect 20750 260 20805 270
rect 20991 270 21041 275
rect 20506 225 20556 230
rect 20991 230 20996 270
rect 21036 230 21041 270
rect 20991 225 21041 230
rect 176 -160 226 -155
rect -425 -190 40 -175
rect -425 -240 -415 -190
rect -365 -240 -25 -190
rect 25 -240 40 -190
rect 176 -200 181 -160
rect 221 -200 226 -160
rect 176 -205 226 -200
rect 421 -160 471 -155
rect 421 -200 426 -160
rect 466 -200 471 -160
rect 421 -205 471 -200
rect 726 -160 776 -155
rect 726 -200 731 -160
rect 771 -200 776 -160
rect 726 -205 776 -200
rect 971 -160 1021 -155
rect 971 -200 976 -160
rect 1016 -200 1021 -160
rect 971 -205 1021 -200
rect 1211 -160 1261 -155
rect 1211 -200 1216 -160
rect 1256 -200 1261 -160
rect 1211 -205 1261 -200
rect 1456 -160 1506 -155
rect 1456 -200 1461 -160
rect 1501 -200 1506 -160
rect 1761 -160 1811 -155
rect 1456 -205 1506 -200
rect 1625 -200 1685 -190
rect -425 -255 40 -240
rect 80 -240 130 -235
rect 80 -280 85 -240
rect 125 -280 130 -240
rect 80 -285 130 -280
rect 320 -240 370 -235
rect 320 -280 325 -240
rect 365 -280 370 -240
rect 320 -285 370 -280
rect 560 -240 610 -235
rect 560 -280 565 -240
rect 605 -280 610 -240
rect 560 -285 610 -280
rect 800 -240 850 -235
rect 800 -280 805 -240
rect 845 -280 850 -240
rect 800 -285 850 -280
rect 1040 -240 1090 -235
rect 1040 -280 1045 -240
rect 1085 -280 1090 -240
rect 1040 -285 1090 -280
rect 1280 -240 1330 -235
rect 1280 -280 1285 -240
rect 1325 -280 1330 -240
rect 1280 -285 1330 -280
rect 1520 -240 1570 -235
rect 1520 -280 1525 -240
rect 1565 -280 1570 -240
rect 1625 -240 1635 -200
rect 1675 -240 1685 -200
rect 1761 -200 1766 -160
rect 1806 -200 1811 -160
rect 1761 -205 1811 -200
rect 2006 -160 2056 -155
rect 2006 -200 2011 -160
rect 2051 -200 2056 -160
rect 2006 -205 2056 -200
rect 2246 -160 2296 -155
rect 2246 -200 2251 -160
rect 2291 -200 2296 -160
rect 2246 -205 2296 -200
rect 2491 -160 2541 -155
rect 2491 -200 2496 -160
rect 2536 -200 2541 -160
rect 2491 -205 2541 -200
rect 2731 -160 2781 -155
rect 2731 -200 2736 -160
rect 2776 -200 2781 -160
rect 2731 -205 2781 -200
rect 2976 -160 3026 -155
rect 2976 -200 2981 -160
rect 3021 -200 3026 -160
rect 2976 -205 3026 -200
rect 3216 -160 3266 -155
rect 3216 -200 3221 -160
rect 3261 -200 3266 -160
rect 3216 -205 3266 -200
rect 3461 -160 3511 -155
rect 3461 -200 3466 -160
rect 3506 -200 3511 -160
rect 3461 -205 3511 -200
rect 3701 -160 3751 -155
rect 3701 -200 3706 -160
rect 3746 -200 3751 -160
rect 3701 -205 3751 -200
rect 3946 -160 3996 -155
rect 3946 -200 3951 -160
rect 3991 -200 3996 -160
rect 4186 -160 4236 -155
rect 3946 -205 3996 -200
rect 4050 -195 4110 -185
rect 4050 -235 4060 -195
rect 4100 -235 4110 -195
rect 4186 -200 4191 -160
rect 4231 -200 4236 -160
rect 4186 -205 4236 -200
rect 4431 -160 4481 -155
rect 4431 -200 4436 -160
rect 4476 -200 4481 -160
rect 4431 -205 4481 -200
rect 4671 -160 4721 -155
rect 4671 -200 4676 -160
rect 4716 -200 4721 -160
rect 4671 -205 4721 -200
rect 4916 -160 4966 -155
rect 4916 -200 4921 -160
rect 4961 -200 4966 -160
rect 4916 -205 4966 -200
rect 5156 -160 5206 -155
rect 5156 -200 5161 -160
rect 5201 -200 5206 -160
rect 5156 -205 5206 -200
rect 5401 -160 5451 -155
rect 5401 -200 5406 -160
rect 5446 -200 5451 -160
rect 5401 -205 5451 -200
rect 5706 -160 5756 -155
rect 5706 -200 5711 -160
rect 5751 -200 5756 -160
rect 5706 -205 5756 -200
rect 5951 -160 6001 -155
rect 5951 -200 5956 -160
rect 5996 -200 6001 -160
rect 5951 -205 6001 -200
rect 6191 -160 6241 -155
rect 6191 -200 6196 -160
rect 6236 -200 6241 -160
rect 6191 -205 6241 -200
rect 6676 -160 6726 -155
rect 6676 -200 6681 -160
rect 6721 -200 6726 -160
rect 6676 -205 6726 -200
rect 6921 -160 6971 -155
rect 6921 -200 6926 -160
rect 6966 -200 6971 -160
rect 6921 -205 6971 -200
rect 7161 -160 7211 -155
rect 7161 -200 7166 -160
rect 7206 -200 7211 -160
rect 7161 -205 7211 -200
rect 7401 -160 7451 -155
rect 7401 -200 7406 -160
rect 7446 -200 7451 -160
rect 7401 -205 7451 -200
rect 7641 -160 7691 -155
rect 7641 -200 7646 -160
rect 7686 -200 7691 -160
rect 7641 -205 7691 -200
rect 8126 -160 8176 -155
rect 8126 -200 8131 -160
rect 8171 -200 8176 -160
rect 8126 -205 8176 -200
rect 8371 -160 8421 -155
rect 8371 -200 8376 -160
rect 8416 -200 8421 -160
rect 8371 -205 8421 -200
rect 8611 -160 8661 -155
rect 8611 -200 8616 -160
rect 8656 -200 8661 -160
rect 8611 -205 8661 -200
rect 8856 -160 8906 -155
rect 8856 -200 8861 -160
rect 8901 -200 8906 -160
rect 8856 -205 8906 -200
rect 9096 -160 9146 -155
rect 9096 -200 9101 -160
rect 9141 -200 9146 -160
rect 9096 -205 9146 -200
rect 9341 -160 9391 -155
rect 9341 -200 9346 -160
rect 9386 -200 9391 -160
rect 9831 -160 9881 -155
rect 9831 -200 9836 -160
rect 9876 -200 9881 -160
rect 9341 -205 9391 -200
rect 9560 -210 9620 -200
rect 9831 -205 9881 -200
rect 10071 -160 10121 -155
rect 10071 -200 10076 -160
rect 10116 -200 10121 -160
rect 10071 -205 10121 -200
rect 10316 -160 10366 -155
rect 10316 -200 10321 -160
rect 10361 -200 10366 -160
rect 10316 -205 10366 -200
rect 10556 -160 10606 -155
rect 10556 -200 10561 -160
rect 10601 -200 10606 -160
rect 10556 -205 10606 -200
rect 10801 -160 10851 -155
rect 10801 -200 10806 -160
rect 10846 -200 10851 -160
rect 10801 -205 10851 -200
rect 11041 -160 11091 -155
rect 11041 -200 11046 -160
rect 11086 -200 11091 -160
rect 11041 -205 11091 -200
rect 11286 -160 11336 -155
rect 11286 -200 11291 -160
rect 11331 -200 11336 -160
rect 11286 -205 11336 -200
rect 11526 -160 11576 -155
rect 11526 -200 11531 -160
rect 11571 -200 11576 -160
rect 11526 -205 11576 -200
rect 11771 -160 11821 -155
rect 11771 -200 11776 -160
rect 11816 -200 11821 -160
rect 11771 -205 11821 -200
rect 12256 -160 12306 -155
rect 12256 -200 12261 -160
rect 12301 -200 12306 -160
rect 12256 -205 12306 -200
rect 12496 -160 12546 -155
rect 12496 -200 12501 -160
rect 12541 -200 12546 -160
rect 12496 -205 12546 -200
rect 12741 -160 12791 -155
rect 12741 -200 12746 -160
rect 12786 -200 12791 -160
rect 12741 -205 12791 -200
rect 12981 -160 13031 -155
rect 12981 -200 12986 -160
rect 13026 -200 13031 -160
rect 12981 -205 13031 -200
rect 13226 -160 13276 -155
rect 13226 -200 13231 -160
rect 13271 -200 13276 -160
rect 13226 -205 13276 -200
rect 13466 -160 13516 -155
rect 13466 -200 13471 -160
rect 13511 -200 13516 -160
rect 13466 -205 13516 -200
rect 13711 -160 13761 -155
rect 13711 -200 13716 -160
rect 13756 -200 13761 -160
rect 13711 -205 13761 -200
rect 14196 -160 14246 -155
rect 14196 -200 14201 -160
rect 14241 -200 14246 -160
rect 14196 -205 14246 -200
rect 14436 -160 14486 -155
rect 14436 -200 14441 -160
rect 14481 -200 14486 -160
rect 14436 -205 14486 -200
rect 14681 -160 14731 -155
rect 14681 -200 14686 -160
rect 14726 -200 14731 -160
rect 14681 -205 14731 -200
rect 14921 -160 14971 -155
rect 14921 -200 14926 -160
rect 14966 -200 14971 -160
rect 14921 -205 14971 -200
rect 15166 -160 15216 -155
rect 15166 -200 15171 -160
rect 15211 -200 15216 -160
rect 15166 -205 15216 -200
rect 15406 -160 15456 -155
rect 15406 -200 15411 -160
rect 15451 -200 15456 -160
rect 15406 -205 15456 -200
rect 15651 -160 15701 -155
rect 15651 -200 15656 -160
rect 15696 -200 15701 -160
rect 15651 -205 15701 -200
rect 16136 -160 16186 -155
rect 16136 -200 16141 -160
rect 16181 -200 16186 -160
rect 16136 -205 16186 -200
rect 16376 -160 16426 -155
rect 16376 -200 16381 -160
rect 16421 -200 16426 -160
rect 16376 -205 16426 -200
rect 16621 -160 16671 -155
rect 16621 -200 16626 -160
rect 16666 -200 16671 -160
rect 16621 -205 16671 -200
rect 16861 -160 16911 -155
rect 16861 -200 16866 -160
rect 16906 -200 16911 -160
rect 16861 -205 16911 -200
rect 17106 -160 17156 -155
rect 17106 -200 17111 -160
rect 17151 -200 17156 -160
rect 17106 -205 17156 -200
rect 17346 -160 17396 -155
rect 17346 -200 17351 -160
rect 17391 -200 17396 -160
rect 17346 -205 17396 -200
rect 17591 -160 17641 -155
rect 17591 -200 17596 -160
rect 17636 -200 17641 -160
rect 17831 -160 17881 -155
rect 17831 -200 17836 -160
rect 17876 -200 17881 -160
rect 17591 -205 17641 -200
rect 17695 -210 17755 -200
rect 17831 -205 17881 -200
rect 18076 -160 18126 -155
rect 18076 -200 18081 -160
rect 18121 -200 18126 -160
rect 18076 -205 18126 -200
rect 18316 -160 18366 -155
rect 18316 -200 18321 -160
rect 18361 -200 18366 -160
rect 18316 -205 18366 -200
rect 18561 -160 18611 -155
rect 18561 -200 18566 -160
rect 18606 -200 18611 -160
rect 18561 -205 18611 -200
rect 18801 -160 18851 -155
rect 18801 -200 18806 -160
rect 18846 -200 18851 -160
rect 18801 -205 18851 -200
rect 19046 -160 19096 -155
rect 19046 -200 19051 -160
rect 19091 -200 19096 -160
rect 19046 -205 19096 -200
rect 19286 -160 19336 -155
rect 19286 -200 19291 -160
rect 19331 -200 19336 -160
rect 19286 -205 19336 -200
rect 19531 -160 19581 -155
rect 19531 -200 19536 -160
rect 19576 -200 19581 -160
rect 19771 -160 19821 -155
rect 19771 -200 19776 -160
rect 19816 -200 19821 -160
rect 19531 -205 19581 -200
rect 6445 -220 6505 -210
rect 1625 -250 1685 -240
rect 1760 -240 1810 -235
rect 1520 -285 1570 -280
rect 1760 -280 1765 -240
rect 1805 -280 1810 -240
rect 1760 -285 1810 -280
rect 2000 -240 2050 -235
rect 2000 -280 2005 -240
rect 2045 -280 2050 -240
rect 2000 -285 2050 -280
rect 2240 -240 2290 -235
rect 2240 -280 2245 -240
rect 2285 -280 2290 -240
rect 2240 -285 2290 -280
rect 2480 -240 2530 -235
rect 2480 -280 2485 -240
rect 2525 -280 2530 -240
rect 2480 -285 2530 -280
rect 2720 -240 2770 -235
rect 2720 -280 2725 -240
rect 2765 -280 2770 -240
rect 2720 -285 2770 -280
rect 2960 -240 3010 -235
rect 2960 -280 2965 -240
rect 3005 -280 3010 -240
rect 2960 -285 3010 -280
rect 3200 -240 3250 -235
rect 3200 -280 3205 -240
rect 3245 -280 3250 -240
rect 3200 -285 3250 -280
rect 3440 -240 3490 -235
rect 3440 -280 3445 -240
rect 3485 -280 3490 -240
rect 3440 -285 3490 -280
rect 3680 -240 3730 -235
rect 3680 -280 3685 -240
rect 3725 -280 3730 -240
rect 3680 -285 3730 -280
rect 3920 -240 3970 -235
rect 3920 -280 3925 -240
rect 3965 -280 3970 -240
rect 4050 -245 4110 -235
rect 4160 -240 4210 -235
rect 3920 -285 3970 -280
rect 4160 -280 4165 -240
rect 4205 -280 4210 -240
rect 4160 -285 4210 -280
rect 4400 -240 4450 -235
rect 4400 -280 4405 -240
rect 4445 -280 4450 -240
rect 4400 -285 4450 -280
rect 4640 -240 4690 -235
rect 4640 -280 4645 -240
rect 4685 -280 4690 -240
rect 4640 -285 4690 -280
rect 4880 -240 4930 -235
rect 4880 -280 4885 -240
rect 4925 -280 4930 -240
rect 4880 -285 4930 -280
rect 5120 -240 5170 -235
rect 5120 -280 5125 -240
rect 5165 -280 5170 -240
rect 5120 -285 5170 -280
rect 5360 -240 5410 -235
rect 5360 -280 5365 -240
rect 5405 -280 5410 -240
rect 5360 -285 5410 -280
rect 5600 -240 5650 -235
rect 5600 -280 5605 -240
rect 5645 -280 5650 -240
rect 5600 -285 5650 -280
rect 5840 -240 5890 -235
rect 5840 -280 5845 -240
rect 5885 -280 5890 -240
rect 5840 -285 5890 -280
rect 6080 -240 6130 -235
rect 6080 -280 6085 -240
rect 6125 -280 6130 -240
rect 6080 -285 6130 -280
rect 6320 -240 6370 -235
rect 6320 -280 6325 -240
rect 6365 -280 6370 -240
rect 6445 -260 6455 -220
rect 6495 -260 6505 -220
rect 7870 -220 7930 -210
rect 6445 -270 6505 -260
rect 6560 -240 6610 -235
rect 6320 -285 6370 -280
rect 6560 -280 6565 -240
rect 6605 -280 6610 -240
rect 6560 -285 6610 -280
rect 6800 -240 6850 -235
rect 6800 -280 6805 -240
rect 6845 -280 6850 -240
rect 6800 -285 6850 -280
rect 7040 -240 7090 -235
rect 7040 -280 7045 -240
rect 7085 -280 7090 -240
rect 7040 -285 7090 -280
rect 7280 -240 7330 -235
rect 7280 -280 7285 -240
rect 7325 -280 7330 -240
rect 7280 -285 7330 -280
rect 7520 -240 7570 -235
rect 7520 -280 7525 -240
rect 7565 -280 7570 -240
rect 7520 -285 7570 -280
rect 7760 -240 7810 -235
rect 7760 -280 7765 -240
rect 7805 -280 7810 -240
rect 7870 -260 7880 -220
rect 7920 -260 7930 -220
rect 7870 -270 7930 -260
rect 8000 -240 8050 -235
rect 7760 -285 7810 -280
rect 8000 -280 8005 -240
rect 8045 -280 8050 -240
rect 8000 -285 8050 -280
rect 8240 -240 8290 -235
rect 8240 -280 8245 -240
rect 8285 -280 8290 -240
rect 8240 -285 8290 -280
rect 8480 -240 8530 -235
rect 8480 -280 8485 -240
rect 8525 -280 8530 -240
rect 8480 -285 8530 -280
rect 8720 -240 8770 -235
rect 8720 -280 8725 -240
rect 8765 -280 8770 -240
rect 8720 -285 8770 -280
rect 8960 -240 9010 -235
rect 8960 -280 8965 -240
rect 9005 -280 9010 -240
rect 8960 -285 9010 -280
rect 9200 -240 9250 -235
rect 9200 -280 9205 -240
rect 9245 -280 9250 -240
rect 9200 -285 9250 -280
rect 9440 -240 9490 -235
rect 9440 -280 9445 -240
rect 9485 -280 9490 -240
rect 9560 -250 9570 -210
rect 9610 -250 9620 -210
rect 11940 -220 12000 -210
rect 9560 -260 9620 -250
rect 9680 -240 9730 -235
rect 9440 -285 9490 -280
rect 9680 -280 9685 -240
rect 9725 -280 9730 -240
rect 9680 -285 9730 -280
rect 9920 -240 9970 -235
rect 9920 -280 9925 -240
rect 9965 -280 9970 -240
rect 9920 -285 9970 -280
rect 10160 -240 10210 -235
rect 10160 -280 10165 -240
rect 10205 -280 10210 -240
rect 10160 -285 10210 -280
rect 10400 -240 10450 -235
rect 10400 -280 10405 -240
rect 10445 -280 10450 -240
rect 10400 -285 10450 -280
rect 10640 -240 10690 -235
rect 10640 -280 10645 -240
rect 10685 -280 10690 -240
rect 10640 -285 10690 -280
rect 10880 -240 10930 -235
rect 10880 -280 10885 -240
rect 10925 -280 10930 -240
rect 10880 -285 10930 -280
rect 11120 -240 11170 -235
rect 11120 -280 11125 -240
rect 11165 -280 11170 -240
rect 11120 -285 11170 -280
rect 11360 -240 11410 -235
rect 11360 -280 11365 -240
rect 11405 -280 11410 -240
rect 11360 -285 11410 -280
rect 11600 -240 11650 -235
rect 11600 -280 11605 -240
rect 11645 -280 11650 -240
rect 11600 -285 11650 -280
rect 11840 -240 11890 -235
rect 11840 -280 11845 -240
rect 11885 -280 11890 -240
rect 11940 -260 11950 -220
rect 11990 -260 12000 -220
rect 13860 -220 13920 -210
rect 11940 -270 12000 -260
rect 12080 -240 12130 -235
rect 11840 -285 11890 -280
rect 12080 -280 12085 -240
rect 12125 -280 12130 -240
rect 12080 -285 12130 -280
rect 12320 -240 12370 -235
rect 12320 -280 12325 -240
rect 12365 -280 12370 -240
rect 12320 -285 12370 -280
rect 12560 -240 12610 -235
rect 12560 -280 12565 -240
rect 12605 -280 12610 -240
rect 12560 -285 12610 -280
rect 12800 -240 12850 -235
rect 12800 -280 12805 -240
rect 12845 -280 12850 -240
rect 12800 -285 12850 -280
rect 13040 -240 13090 -235
rect 13040 -280 13045 -240
rect 13085 -280 13090 -240
rect 13040 -285 13090 -280
rect 13280 -240 13330 -235
rect 13280 -280 13285 -240
rect 13325 -280 13330 -240
rect 13280 -285 13330 -280
rect 13520 -240 13570 -235
rect 13520 -280 13525 -240
rect 13565 -280 13570 -240
rect 13520 -285 13570 -280
rect 13760 -240 13810 -235
rect 13760 -280 13765 -240
rect 13805 -280 13810 -240
rect 13860 -260 13870 -220
rect 13910 -260 13920 -220
rect 15805 -220 15865 -210
rect 13860 -270 13920 -260
rect 14000 -240 14050 -235
rect 13760 -285 13810 -280
rect 14000 -280 14005 -240
rect 14045 -280 14050 -240
rect 14000 -285 14050 -280
rect 14240 -240 14290 -235
rect 14240 -280 14245 -240
rect 14285 -280 14290 -240
rect 14240 -285 14290 -280
rect 14480 -240 14530 -235
rect 14480 -280 14485 -240
rect 14525 -280 14530 -240
rect 14480 -285 14530 -280
rect 14720 -240 14770 -235
rect 14720 -280 14725 -240
rect 14765 -280 14770 -240
rect 14720 -285 14770 -280
rect 14960 -240 15010 -235
rect 14960 -280 14965 -240
rect 15005 -280 15010 -240
rect 14960 -285 15010 -280
rect 15200 -240 15250 -235
rect 15200 -280 15205 -240
rect 15245 -280 15250 -240
rect 15200 -285 15250 -280
rect 15440 -240 15490 -235
rect 15440 -280 15445 -240
rect 15485 -280 15490 -240
rect 15440 -285 15490 -280
rect 15680 -240 15730 -235
rect 15680 -280 15685 -240
rect 15725 -280 15730 -240
rect 15805 -260 15815 -220
rect 15855 -260 15865 -220
rect 15805 -270 15865 -260
rect 15920 -240 15970 -235
rect 15680 -285 15730 -280
rect 15920 -280 15925 -240
rect 15965 -280 15970 -240
rect 15920 -285 15970 -280
rect 16160 -240 16210 -235
rect 16160 -280 16165 -240
rect 16205 -280 16210 -240
rect 16160 -285 16210 -280
rect 16400 -240 16450 -235
rect 16400 -280 16405 -240
rect 16445 -280 16450 -240
rect 16400 -285 16450 -280
rect 16640 -240 16690 -235
rect 16640 -280 16645 -240
rect 16685 -280 16690 -240
rect 16640 -285 16690 -280
rect 16880 -240 16930 -235
rect 16880 -280 16885 -240
rect 16925 -280 16930 -240
rect 16880 -285 16930 -280
rect 17120 -240 17170 -235
rect 17120 -280 17125 -240
rect 17165 -280 17170 -240
rect 17120 -285 17170 -280
rect 17360 -240 17410 -235
rect 17360 -280 17365 -240
rect 17405 -280 17410 -240
rect 17360 -285 17410 -280
rect 17600 -240 17650 -235
rect 17600 -280 17605 -240
rect 17645 -280 17650 -240
rect 17695 -250 17705 -210
rect 17745 -250 17755 -210
rect 19635 -210 19695 -200
rect 19771 -205 19821 -200
rect 20016 -160 20066 -155
rect 20016 -200 20021 -160
rect 20061 -200 20066 -160
rect 20016 -205 20066 -200
rect 20256 -160 20306 -155
rect 20256 -200 20261 -160
rect 20301 -200 20306 -160
rect 20256 -205 20306 -200
rect 20501 -160 20551 -155
rect 20501 -200 20506 -160
rect 20546 -200 20551 -160
rect 20501 -205 20551 -200
rect 20741 -160 20791 -155
rect 20741 -200 20746 -160
rect 20786 -200 20791 -160
rect 20741 -205 20791 -200
rect 20986 -160 21036 -155
rect 20986 -200 20991 -160
rect 21031 -200 21036 -160
rect 20986 -205 21036 -200
rect 17695 -260 17755 -250
rect 17840 -240 17890 -235
rect 17600 -285 17650 -280
rect 17840 -280 17845 -240
rect 17885 -280 17890 -240
rect 17840 -285 17890 -280
rect 18080 -240 18130 -235
rect 18080 -280 18085 -240
rect 18125 -280 18130 -240
rect 18080 -285 18130 -280
rect 18320 -240 18370 -235
rect 18320 -280 18325 -240
rect 18365 -280 18370 -240
rect 18320 -285 18370 -280
rect 18560 -240 18610 -235
rect 18560 -280 18565 -240
rect 18605 -280 18610 -240
rect 18560 -285 18610 -280
rect 18800 -240 18850 -235
rect 18800 -280 18805 -240
rect 18845 -280 18850 -240
rect 18800 -285 18850 -280
rect 19040 -240 19090 -235
rect 19040 -280 19045 -240
rect 19085 -280 19090 -240
rect 19040 -285 19090 -280
rect 19280 -240 19330 -235
rect 19280 -280 19285 -240
rect 19325 -280 19330 -240
rect 19280 -285 19330 -280
rect 19520 -240 19570 -235
rect 19520 -280 19525 -240
rect 19565 -280 19570 -240
rect 19635 -250 19645 -210
rect 19685 -250 19695 -210
rect 19635 -260 19695 -250
rect 19760 -240 19810 -235
rect 19520 -285 19570 -280
rect 19760 -280 19765 -240
rect 19805 -280 19810 -240
rect 19760 -285 19810 -280
rect 20000 -240 20050 -235
rect 20000 -280 20005 -240
rect 20045 -280 20050 -240
rect 20000 -285 20050 -280
rect 20240 -240 20290 -235
rect 20240 -280 20245 -240
rect 20285 -280 20290 -240
rect 20240 -285 20290 -280
rect 20480 -240 20530 -235
rect 20480 -280 20485 -240
rect 20525 -280 20530 -240
rect 20480 -285 20530 -280
rect 20720 -240 20770 -235
rect 20720 -280 20725 -240
rect 20765 -280 20770 -240
rect 20720 -285 20770 -280
rect 20960 -240 21010 -235
rect 20960 -280 20965 -240
rect 21005 -280 21010 -240
rect 20960 -285 21010 -280
rect 21200 -240 21250 -235
rect 21200 -280 21205 -240
rect 21245 -280 21250 -240
rect 21200 -285 21250 -280
rect 21440 -240 21490 -235
rect 21440 -280 21445 -240
rect 21485 -280 21490 -240
rect 21440 -285 21490 -280
rect 21680 -240 21730 -235
rect 21680 -280 21685 -240
rect 21725 -280 21730 -240
rect 21680 -285 21730 -280
rect 21920 -240 21970 -235
rect 21920 -280 21925 -240
rect 21965 -280 21970 -240
rect 21920 -285 21970 -280
rect 22160 -240 22210 -235
rect 22160 -280 22165 -240
rect 22205 -280 22210 -240
rect 22160 -285 22210 -280
rect 22400 -240 22450 -235
rect 22400 -280 22405 -240
rect 22445 -280 22450 -240
rect 22400 -285 22450 -280
rect 22640 -240 22690 -235
rect 22640 -280 22645 -240
rect 22685 -280 22690 -240
rect 22640 -285 22690 -280
rect 22880 -240 22930 -235
rect 22880 -280 22885 -240
rect 22925 -280 22930 -240
rect 22880 -285 22930 -280
rect 23120 -240 23170 -235
rect 23120 -280 23125 -240
rect 23165 -280 23170 -240
rect 23120 -285 23170 -280
rect 23360 -240 23410 -235
rect 23360 -280 23365 -240
rect 23405 -280 23410 -240
rect 23360 -285 23410 -280
rect 23600 -240 23650 -235
rect 23600 -280 23605 -240
rect 23645 -280 23650 -240
rect 23600 -285 23650 -280
rect 23840 -240 23890 -235
rect 23840 -280 23845 -240
rect 23885 -280 23890 -240
rect 23840 -285 23890 -280
rect 24080 -240 24130 -235
rect 24080 -280 24085 -240
rect 24125 -280 24130 -240
rect 24080 -285 24130 -280
rect 24320 -240 24370 -235
rect 24320 -280 24325 -240
rect 24365 -280 24370 -240
rect 24320 -285 24370 -280
rect 24560 -240 24610 -235
rect 24560 -280 24565 -240
rect 24605 -280 24610 -240
rect 24560 -285 24610 -280
rect 24800 -240 24850 -235
rect 24800 -280 24805 -240
rect 24845 -280 24850 -240
rect 24800 -285 24850 -280
rect 25040 -240 25090 -235
rect 25040 -280 25045 -240
rect 25085 -280 25090 -240
rect 25040 -285 25090 -280
rect 25280 -240 25330 -235
rect 25280 -280 25285 -240
rect 25325 -280 25330 -240
rect 25280 -285 25330 -280
rect 25520 -240 25570 -235
rect 25520 -280 25525 -240
rect 25565 -280 25570 -240
rect 25520 -285 25570 -280
rect 25760 -240 25810 -235
rect 25760 -280 25765 -240
rect 25805 -280 25810 -240
rect 25760 -285 25810 -280
rect 26000 -240 26050 -235
rect 26000 -280 26005 -240
rect 26045 -280 26050 -240
rect 26000 -285 26050 -280
rect 26240 -240 26290 -235
rect 26240 -280 26245 -240
rect 26285 -280 26290 -240
rect 26240 -285 26290 -280
rect 26480 -240 26530 -235
rect 26480 -280 26485 -240
rect 26525 -280 26530 -240
rect 26480 -285 26530 -280
rect 26720 -240 26770 -235
rect 26720 -280 26725 -240
rect 26765 -280 26770 -240
rect 26720 -285 26770 -280
rect 26960 -240 27010 -235
rect 26960 -280 26965 -240
rect 27005 -280 27010 -240
rect 26960 -285 27010 -280
rect 27200 -240 27250 -235
rect 27200 -280 27205 -240
rect 27245 -280 27250 -240
rect 27200 -285 27250 -280
rect 27440 -240 27490 -235
rect 27440 -280 27445 -240
rect 27485 -280 27490 -240
rect 27440 -285 27490 -280
rect 27680 -240 27730 -235
rect 27680 -280 27685 -240
rect 27725 -280 27730 -240
rect 27680 -285 27730 -280
rect 27920 -240 27970 -235
rect 27920 -280 27925 -240
rect 27965 -280 27970 -240
rect 27920 -285 27970 -280
rect 28160 -240 28210 -235
rect 28160 -280 28165 -240
rect 28205 -280 28210 -240
rect 28160 -285 28210 -280
rect 28400 -240 28450 -235
rect 28400 -280 28405 -240
rect 28445 -280 28450 -240
rect 28400 -285 28450 -280
rect 28640 -240 28690 -235
rect 28640 -280 28645 -240
rect 28685 -280 28690 -240
rect 28640 -285 28690 -280
rect 28880 -240 28930 -235
rect 28880 -280 28885 -240
rect 28925 -280 28930 -240
rect 28880 -285 28930 -280
rect 29120 -240 29170 -235
rect 29120 -280 29125 -240
rect 29165 -280 29170 -240
rect 29120 -285 29170 -280
rect 29360 -240 29410 -235
rect 29360 -280 29365 -240
rect 29405 -280 29410 -240
rect 29360 -285 29410 -280
rect 29600 -240 29650 -235
rect 29600 -280 29605 -240
rect 29645 -280 29650 -240
rect 29600 -285 29650 -280
rect 29840 -240 29890 -235
rect 29840 -280 29845 -240
rect 29885 -280 29890 -240
rect 29840 -285 29890 -280
rect 30080 -240 30130 -235
rect 30080 -280 30085 -240
rect 30125 -280 30130 -240
rect 30080 -285 30130 -280
rect 30320 -240 30370 -235
rect 30320 -280 30325 -240
rect 30365 -280 30370 -240
rect 30320 -285 30370 -280
rect 30560 -240 30610 -235
rect 30560 -280 30565 -240
rect 30605 -280 30610 -240
rect 30560 -285 30610 -280
rect 75 -815 125 -810
rect 75 -855 80 -815
rect 120 -855 125 -815
rect 75 -860 125 -855
rect 315 -815 365 -810
rect 315 -855 320 -815
rect 360 -855 365 -815
rect 315 -860 365 -855
rect 555 -815 605 -810
rect 555 -855 560 -815
rect 600 -855 605 -815
rect 1035 -815 1085 -810
rect 555 -860 605 -855
rect 790 -835 845 -825
rect 790 -870 800 -835
rect 835 -870 845 -835
rect 1035 -855 1040 -815
rect 1080 -855 1085 -815
rect 1035 -860 1085 -855
rect 1275 -815 1325 -810
rect 1275 -855 1280 -815
rect 1320 -855 1325 -815
rect 1275 -860 1325 -855
rect 1515 -815 1565 -810
rect 1515 -855 1520 -815
rect 1560 -855 1565 -815
rect 1515 -860 1565 -855
rect 1755 -815 1805 -810
rect 1755 -855 1760 -815
rect 1800 -855 1805 -815
rect 1755 -860 1805 -855
rect 1995 -815 2045 -810
rect 1995 -855 2000 -815
rect 2040 -855 2045 -815
rect 1995 -860 2045 -855
rect 2235 -815 2285 -810
rect 2235 -855 2240 -815
rect 2280 -855 2285 -815
rect 2235 -860 2285 -855
rect 2475 -815 2525 -810
rect 2475 -855 2480 -815
rect 2520 -855 2525 -815
rect 2475 -860 2525 -855
rect 2715 -815 2765 -810
rect 2715 -855 2720 -815
rect 2760 -855 2765 -815
rect 3195 -815 3245 -810
rect 2715 -860 2765 -855
rect 2950 -835 3005 -825
rect 790 -880 845 -870
rect 2950 -870 2960 -835
rect 2995 -870 3005 -835
rect 3195 -855 3200 -815
rect 3240 -855 3245 -815
rect 3195 -860 3245 -855
rect 3435 -815 3485 -810
rect 3435 -855 3440 -815
rect 3480 -855 3485 -815
rect 3435 -860 3485 -855
rect 3675 -815 3725 -810
rect 3675 -855 3680 -815
rect 3720 -855 3725 -815
rect 3675 -860 3725 -855
rect 3915 -815 3965 -810
rect 3915 -855 3920 -815
rect 3960 -855 3965 -815
rect 3915 -860 3965 -855
rect 4155 -815 4205 -810
rect 4155 -855 4160 -815
rect 4200 -855 4205 -815
rect 4155 -860 4205 -855
rect 4395 -815 4445 -810
rect 4395 -855 4400 -815
rect 4440 -855 4445 -815
rect 4395 -860 4445 -855
rect 4635 -815 4685 -810
rect 4635 -855 4640 -815
rect 4680 -855 4685 -815
rect 4635 -860 4685 -855
rect 4875 -815 4925 -810
rect 4875 -855 4880 -815
rect 4920 -855 4925 -815
rect 5355 -815 5405 -810
rect 4875 -860 4925 -855
rect 5110 -835 5165 -825
rect 2950 -880 3005 -870
rect 5110 -870 5120 -835
rect 5155 -870 5165 -835
rect 5355 -855 5360 -815
rect 5400 -855 5405 -815
rect 5355 -860 5405 -855
rect 5595 -815 5645 -810
rect 5595 -855 5600 -815
rect 5640 -855 5645 -815
rect 5595 -860 5645 -855
rect 5835 -815 5885 -810
rect 5835 -855 5840 -815
rect 5880 -855 5885 -815
rect 5835 -860 5885 -855
rect 6075 -815 6125 -810
rect 6075 -855 6080 -815
rect 6120 -855 6125 -815
rect 6075 -860 6125 -855
rect 6315 -815 6365 -810
rect 6315 -855 6320 -815
rect 6360 -855 6365 -815
rect 6315 -860 6365 -855
rect 6555 -815 6605 -810
rect 6555 -855 6560 -815
rect 6600 -855 6605 -815
rect 6555 -860 6605 -855
rect 6795 -815 6845 -810
rect 6795 -855 6800 -815
rect 6840 -855 6845 -815
rect 6795 -860 6845 -855
rect 7035 -815 7085 -810
rect 7035 -855 7040 -815
rect 7080 -855 7085 -815
rect 7515 -815 7565 -810
rect 7035 -860 7085 -855
rect 7270 -835 7325 -825
rect 5110 -880 5165 -870
rect 7270 -870 7280 -835
rect 7315 -870 7325 -835
rect 7515 -855 7520 -815
rect 7560 -855 7565 -815
rect 7515 -860 7565 -855
rect 7755 -815 7805 -810
rect 7755 -855 7760 -815
rect 7800 -855 7805 -815
rect 7755 -860 7805 -855
rect 7995 -815 8045 -810
rect 7995 -855 8000 -815
rect 8040 -855 8045 -815
rect 7995 -860 8045 -855
rect 8235 -815 8285 -810
rect 8235 -855 8240 -815
rect 8280 -855 8285 -815
rect 8235 -860 8285 -855
rect 8475 -815 8525 -810
rect 8475 -855 8480 -815
rect 8520 -855 8525 -815
rect 8475 -860 8525 -855
rect 8715 -815 8765 -810
rect 8715 -855 8720 -815
rect 8760 -855 8765 -815
rect 8715 -860 8765 -855
rect 8955 -815 9005 -810
rect 8955 -855 8960 -815
rect 9000 -855 9005 -815
rect 8955 -860 9005 -855
rect 9195 -815 9245 -810
rect 9195 -855 9200 -815
rect 9240 -855 9245 -815
rect 9675 -815 9725 -810
rect 9195 -860 9245 -855
rect 9430 -835 9485 -825
rect 7270 -880 7325 -870
rect 9430 -870 9440 -835
rect 9475 -870 9485 -835
rect 9675 -855 9680 -815
rect 9720 -855 9725 -815
rect 9675 -860 9725 -855
rect 9915 -815 9965 -810
rect 9915 -855 9920 -815
rect 9960 -855 9965 -815
rect 9915 -860 9965 -855
rect 10155 -815 10205 -810
rect 10155 -855 10160 -815
rect 10200 -855 10205 -815
rect 10155 -860 10205 -855
rect 10395 -815 10445 -810
rect 10395 -855 10400 -815
rect 10440 -855 10445 -815
rect 10395 -860 10445 -855
rect 10635 -815 10685 -810
rect 10635 -855 10640 -815
rect 10680 -855 10685 -815
rect 10635 -860 10685 -855
rect 10875 -815 10925 -810
rect 10875 -855 10880 -815
rect 10920 -855 10925 -815
rect 10875 -860 10925 -855
rect 11115 -815 11165 -810
rect 11115 -855 11120 -815
rect 11160 -855 11165 -815
rect 11115 -860 11165 -855
rect 11355 -815 11405 -810
rect 11355 -855 11360 -815
rect 11400 -855 11405 -815
rect 11835 -815 11885 -810
rect 11355 -860 11405 -855
rect 11590 -835 11645 -825
rect 9430 -880 9485 -870
rect 11590 -870 11600 -835
rect 11635 -870 11645 -835
rect 11835 -855 11840 -815
rect 11880 -855 11885 -815
rect 11835 -860 11885 -855
rect 12075 -815 12125 -810
rect 12075 -855 12080 -815
rect 12120 -855 12125 -815
rect 12075 -860 12125 -855
rect 12315 -815 12365 -810
rect 12315 -855 12320 -815
rect 12360 -855 12365 -815
rect 12315 -860 12365 -855
rect 12555 -815 12605 -810
rect 12555 -855 12560 -815
rect 12600 -855 12605 -815
rect 12555 -860 12605 -855
rect 12795 -815 12845 -810
rect 12795 -855 12800 -815
rect 12840 -855 12845 -815
rect 12795 -860 12845 -855
rect 13035 -815 13085 -810
rect 13035 -855 13040 -815
rect 13080 -855 13085 -815
rect 13035 -860 13085 -855
rect 13275 -815 13325 -810
rect 13275 -855 13280 -815
rect 13320 -855 13325 -815
rect 13275 -860 13325 -855
rect 13515 -815 13565 -810
rect 13515 -855 13520 -815
rect 13560 -855 13565 -815
rect 13995 -815 14045 -810
rect 13515 -860 13565 -855
rect 13750 -835 13805 -825
rect 11590 -880 11645 -870
rect 13750 -870 13760 -835
rect 13795 -870 13805 -835
rect 13995 -855 14000 -815
rect 14040 -855 14045 -815
rect 13995 -860 14045 -855
rect 14235 -815 14285 -810
rect 14235 -855 14240 -815
rect 14280 -855 14285 -815
rect 14235 -860 14285 -855
rect 14475 -815 14525 -810
rect 14475 -855 14480 -815
rect 14520 -855 14525 -815
rect 14475 -860 14525 -855
rect 14715 -815 14765 -810
rect 14715 -855 14720 -815
rect 14760 -855 14765 -815
rect 14715 -860 14765 -855
rect 14955 -815 15005 -810
rect 14955 -855 14960 -815
rect 15000 -855 15005 -815
rect 14955 -860 15005 -855
rect 15195 -815 15245 -810
rect 15195 -855 15200 -815
rect 15240 -855 15245 -815
rect 15195 -860 15245 -855
rect 15435 -815 15485 -810
rect 15435 -855 15440 -815
rect 15480 -855 15485 -815
rect 15435 -860 15485 -855
rect 15675 -815 15725 -810
rect 15675 -855 15680 -815
rect 15720 -855 15725 -815
rect 16155 -815 16205 -810
rect 15675 -860 15725 -855
rect 15910 -835 15965 -825
rect 13750 -880 13805 -870
rect 15910 -870 15920 -835
rect 15955 -870 15965 -835
rect 16155 -855 16160 -815
rect 16200 -855 16205 -815
rect 16155 -860 16205 -855
rect 16395 -815 16445 -810
rect 16395 -855 16400 -815
rect 16440 -855 16445 -815
rect 16395 -860 16445 -855
rect 16635 -815 16685 -810
rect 16635 -855 16640 -815
rect 16680 -855 16685 -815
rect 16635 -860 16685 -855
rect 16875 -815 16925 -810
rect 16875 -855 16880 -815
rect 16920 -855 16925 -815
rect 16875 -860 16925 -855
rect 17115 -815 17165 -810
rect 17115 -855 17120 -815
rect 17160 -855 17165 -815
rect 17115 -860 17165 -855
rect 17355 -815 17405 -810
rect 17355 -855 17360 -815
rect 17400 -855 17405 -815
rect 17355 -860 17405 -855
rect 17595 -815 17645 -810
rect 17595 -855 17600 -815
rect 17640 -855 17645 -815
rect 17595 -860 17645 -855
rect 17835 -815 17885 -810
rect 17835 -855 17840 -815
rect 17880 -855 17885 -815
rect 18315 -815 18365 -810
rect 17835 -860 17885 -855
rect 18070 -835 18125 -825
rect 15910 -880 15965 -870
rect 18070 -870 18080 -835
rect 18115 -870 18125 -835
rect 18315 -855 18320 -815
rect 18360 -855 18365 -815
rect 18315 -860 18365 -855
rect 18555 -815 18605 -810
rect 18555 -855 18560 -815
rect 18600 -855 18605 -815
rect 18555 -860 18605 -855
rect 18795 -815 18845 -810
rect 18795 -855 18800 -815
rect 18840 -855 18845 -815
rect 18795 -860 18845 -855
rect 19035 -815 19085 -810
rect 19035 -855 19040 -815
rect 19080 -855 19085 -815
rect 19035 -860 19085 -855
rect 19275 -815 19325 -810
rect 19275 -855 19280 -815
rect 19320 -855 19325 -815
rect 19275 -860 19325 -855
rect 19515 -815 19565 -810
rect 19515 -855 19520 -815
rect 19560 -855 19565 -815
rect 19515 -860 19565 -855
rect 19755 -815 19805 -810
rect 19755 -855 19760 -815
rect 19800 -855 19805 -815
rect 19755 -860 19805 -855
rect 19995 -815 20045 -810
rect 19995 -855 20000 -815
rect 20040 -855 20045 -815
rect 20475 -815 20525 -810
rect 19995 -860 20045 -855
rect 20230 -835 20285 -825
rect 18070 -880 18125 -870
rect 20230 -870 20240 -835
rect 20275 -870 20285 -835
rect 20475 -855 20480 -815
rect 20520 -855 20525 -815
rect 20475 -860 20525 -855
rect 20715 -815 20765 -810
rect 20715 -855 20720 -815
rect 20760 -855 20765 -815
rect 20715 -860 20765 -855
rect 20955 -815 21005 -810
rect 20955 -855 20960 -815
rect 21000 -855 21005 -815
rect 20955 -860 21005 -855
rect 21195 -815 21245 -810
rect 21195 -855 21200 -815
rect 21240 -855 21245 -815
rect 21195 -860 21245 -855
rect 21435 -815 21485 -810
rect 21435 -855 21440 -815
rect 21480 -855 21485 -815
rect 21435 -860 21485 -855
rect 21675 -815 21725 -810
rect 21675 -855 21680 -815
rect 21720 -855 21725 -815
rect 21675 -860 21725 -855
rect 21915 -815 21965 -810
rect 21915 -855 21920 -815
rect 21960 -855 21965 -815
rect 21915 -860 21965 -855
rect 22155 -815 22205 -810
rect 22155 -855 22160 -815
rect 22200 -855 22205 -815
rect 22635 -815 22685 -810
rect 22155 -860 22205 -855
rect 22390 -835 22445 -825
rect 20230 -880 20285 -870
rect 22390 -870 22400 -835
rect 22435 -870 22445 -835
rect 22635 -855 22640 -815
rect 22680 -855 22685 -815
rect 22635 -860 22685 -855
rect 22875 -815 22925 -810
rect 22875 -855 22880 -815
rect 22920 -855 22925 -815
rect 22875 -860 22925 -855
rect 23115 -815 23165 -810
rect 23115 -855 23120 -815
rect 23160 -855 23165 -815
rect 23115 -860 23165 -855
rect 23355 -815 23405 -810
rect 23355 -855 23360 -815
rect 23400 -855 23405 -815
rect 23355 -860 23405 -855
rect 23595 -815 23645 -810
rect 23595 -855 23600 -815
rect 23640 -855 23645 -815
rect 23595 -860 23645 -855
rect 23835 -815 23885 -810
rect 23835 -855 23840 -815
rect 23880 -855 23885 -815
rect 23835 -860 23885 -855
rect 24075 -815 24125 -810
rect 24075 -855 24080 -815
rect 24120 -855 24125 -815
rect 24555 -815 24605 -810
rect 24075 -860 24125 -855
rect 24310 -835 24365 -825
rect 22390 -880 22445 -870
rect 24310 -870 24320 -835
rect 24355 -870 24365 -835
rect 24555 -855 24560 -815
rect 24600 -855 24605 -815
rect 24555 -860 24605 -855
rect 24795 -815 24845 -810
rect 24795 -855 24800 -815
rect 24840 -855 24845 -815
rect 24795 -860 24845 -855
rect 25035 -815 25085 -810
rect 25035 -855 25040 -815
rect 25080 -855 25085 -815
rect 25035 -860 25085 -855
rect 25275 -815 25325 -810
rect 25275 -855 25280 -815
rect 25320 -855 25325 -815
rect 25275 -860 25325 -855
rect 25515 -815 25565 -810
rect 25515 -855 25520 -815
rect 25560 -855 25565 -815
rect 25515 -860 25565 -855
rect 25755 -815 25805 -810
rect 25755 -855 25760 -815
rect 25800 -855 25805 -815
rect 25755 -860 25805 -855
rect 25995 -815 26045 -810
rect 25995 -855 26000 -815
rect 26040 -855 26045 -815
rect 26475 -815 26525 -810
rect 25995 -860 26045 -855
rect 26230 -835 26285 -825
rect 24310 -880 24365 -870
rect 26230 -870 26240 -835
rect 26275 -870 26285 -835
rect 26475 -855 26480 -815
rect 26520 -855 26525 -815
rect 26475 -860 26525 -855
rect 26715 -815 26765 -810
rect 26715 -855 26720 -815
rect 26760 -855 26765 -815
rect 26715 -860 26765 -855
rect 26955 -815 27005 -810
rect 26955 -855 26960 -815
rect 27000 -855 27005 -815
rect 26955 -860 27005 -855
rect 27195 -815 27245 -810
rect 27195 -855 27200 -815
rect 27240 -855 27245 -815
rect 27195 -860 27245 -855
rect 27435 -815 27485 -810
rect 27435 -855 27440 -815
rect 27480 -855 27485 -815
rect 27435 -860 27485 -855
rect 27675 -815 27725 -810
rect 27675 -855 27680 -815
rect 27720 -855 27725 -815
rect 27675 -860 27725 -855
rect 27915 -815 27965 -810
rect 27915 -855 27920 -815
rect 27960 -855 27965 -815
rect 28395 -815 28445 -810
rect 27915 -860 27965 -855
rect 28150 -835 28205 -825
rect 26230 -880 26285 -870
rect 28150 -870 28160 -835
rect 28195 -870 28205 -835
rect 28395 -855 28400 -815
rect 28440 -855 28445 -815
rect 28395 -860 28445 -855
rect 28635 -815 28685 -810
rect 28635 -855 28640 -815
rect 28680 -855 28685 -815
rect 28635 -860 28685 -855
rect 28875 -815 28925 -810
rect 28875 -855 28880 -815
rect 28920 -855 28925 -815
rect 28875 -860 28925 -855
rect 29115 -815 29165 -810
rect 29115 -855 29120 -815
rect 29160 -855 29165 -815
rect 29115 -860 29165 -855
rect 29355 -815 29405 -810
rect 29355 -855 29360 -815
rect 29400 -855 29405 -815
rect 29355 -860 29405 -855
rect 29595 -815 29645 -810
rect 29595 -855 29600 -815
rect 29640 -855 29645 -815
rect 30075 -815 30125 -810
rect 29595 -860 29645 -855
rect 29830 -835 29885 -825
rect 28150 -880 28205 -870
rect 29830 -870 29840 -835
rect 29875 -870 29885 -835
rect 30075 -855 30080 -815
rect 30120 -855 30125 -815
rect 30075 -860 30125 -855
rect 30315 -815 30365 -810
rect 30315 -855 30320 -815
rect 30360 -855 30365 -815
rect 30315 -860 30365 -855
rect 30555 -815 30605 -810
rect 30555 -855 30560 -815
rect 30600 -855 30605 -815
rect 30555 -860 30605 -855
rect 29830 -880 29885 -870
<< via3 >>
rect 195 240 230 275
rect 431 265 471 270
rect 431 235 436 265
rect 436 235 466 265
rect 466 235 471 265
rect 431 230 471 235
rect 736 265 776 270
rect 736 235 741 265
rect 741 235 771 265
rect 771 235 776 265
rect 736 230 776 235
rect 981 265 1021 270
rect 981 235 986 265
rect 986 235 1016 265
rect 1016 235 1021 265
rect 981 230 1021 235
rect 1221 265 1261 270
rect 1221 235 1226 265
rect 1226 235 1256 265
rect 1256 235 1261 265
rect 1221 230 1261 235
rect 1466 265 1506 270
rect 1466 235 1471 265
rect 1471 235 1501 265
rect 1501 235 1506 265
rect 1466 230 1506 235
rect 1771 265 1811 270
rect 1771 235 1776 265
rect 1776 235 1806 265
rect 1806 235 1811 265
rect 1771 230 1811 235
rect 2016 265 2056 270
rect 2016 235 2021 265
rect 2021 235 2051 265
rect 2051 235 2056 265
rect 2016 230 2056 235
rect 2265 270 2300 305
rect 2501 265 2541 270
rect 2501 235 2506 265
rect 2506 235 2536 265
rect 2536 235 2541 265
rect 2501 230 2541 235
rect 2741 265 2781 270
rect 2741 235 2746 265
rect 2746 235 2776 265
rect 2776 235 2781 265
rect 2741 230 2781 235
rect 2986 265 3026 270
rect 2986 235 2991 265
rect 2991 235 3021 265
rect 3021 235 3026 265
rect 2986 230 3026 235
rect 3226 265 3266 270
rect 3226 235 3231 265
rect 3231 235 3261 265
rect 3261 235 3266 265
rect 3226 230 3266 235
rect 3471 265 3511 270
rect 3471 235 3476 265
rect 3476 235 3506 265
rect 3506 235 3511 265
rect 3471 230 3511 235
rect 3711 265 3751 270
rect 3711 235 3716 265
rect 3716 235 3746 265
rect 3746 235 3751 265
rect 3711 230 3751 235
rect 3956 265 3996 270
rect 3956 235 3961 265
rect 3961 235 3991 265
rect 3991 235 3996 265
rect 3956 230 3996 235
rect 4205 270 4240 305
rect 4441 265 4481 270
rect 4441 235 4446 265
rect 4446 235 4476 265
rect 4476 235 4481 265
rect 4441 230 4481 235
rect 4681 265 4721 270
rect 4681 235 4686 265
rect 4686 235 4716 265
rect 4716 235 4721 265
rect 4681 230 4721 235
rect 4926 265 4966 270
rect 4926 235 4931 265
rect 4931 235 4961 265
rect 4961 235 4966 265
rect 4926 230 4966 235
rect 5166 265 5206 270
rect 5166 235 5171 265
rect 5171 235 5201 265
rect 5201 235 5206 265
rect 5166 230 5206 235
rect 5411 265 5451 270
rect 5411 235 5416 265
rect 5416 235 5446 265
rect 5446 235 5451 265
rect 5411 230 5451 235
rect 5716 265 5756 270
rect 5716 235 5721 265
rect 5721 235 5751 265
rect 5751 235 5756 265
rect 5716 230 5756 235
rect 5961 265 6001 270
rect 5961 235 5966 265
rect 5966 235 5996 265
rect 5996 235 6001 265
rect 5961 230 6001 235
rect 6201 265 6241 270
rect 6201 235 6206 265
rect 6206 235 6236 265
rect 6236 235 6241 265
rect 6201 230 6241 235
rect 6455 270 6490 305
rect 6686 265 6726 270
rect 6686 235 6691 265
rect 6691 235 6721 265
rect 6721 235 6726 265
rect 6686 230 6726 235
rect 6931 265 6971 270
rect 6931 235 6936 265
rect 6936 235 6966 265
rect 6966 235 6971 265
rect 6931 230 6971 235
rect 7171 265 7211 270
rect 7171 235 7176 265
rect 7176 235 7206 265
rect 7206 235 7211 265
rect 7171 230 7211 235
rect 7411 265 7451 270
rect 7411 235 7416 265
rect 7416 235 7446 265
rect 7446 235 7451 265
rect 7411 230 7451 235
rect 7651 265 7691 270
rect 7651 235 7656 265
rect 7656 235 7686 265
rect 7686 235 7691 265
rect 7651 230 7691 235
rect 7896 265 7936 270
rect 7896 235 7901 265
rect 7901 235 7931 265
rect 7931 235 7936 265
rect 7896 230 7936 235
rect 8136 265 8176 270
rect 8136 235 8141 265
rect 8141 235 8171 265
rect 8171 235 8176 265
rect 8136 230 8176 235
rect 8381 265 8421 270
rect 8381 235 8386 265
rect 8386 235 8416 265
rect 8416 235 8421 265
rect 8381 230 8421 235
rect 8621 265 8661 270
rect 8621 235 8626 265
rect 8626 235 8656 265
rect 8656 235 8661 265
rect 8621 230 8661 235
rect 8866 265 8906 270
rect 8866 235 8871 265
rect 8871 235 8901 265
rect 8901 235 8906 265
rect 8866 230 8906 235
rect 9106 265 9146 270
rect 9106 235 9111 265
rect 9111 235 9141 265
rect 9141 235 9146 265
rect 9106 230 9146 235
rect 9360 270 9395 305
rect 9596 265 9636 270
rect 9596 235 9601 265
rect 9601 235 9631 265
rect 9631 235 9636 265
rect 9596 230 9636 235
rect 9841 265 9881 270
rect 9841 235 9846 265
rect 9846 235 9876 265
rect 9876 235 9881 265
rect 9841 230 9881 235
rect 10081 265 10121 270
rect 10081 235 10086 265
rect 10086 235 10116 265
rect 10116 235 10121 265
rect 10081 230 10121 235
rect 10326 265 10366 270
rect 10326 235 10331 265
rect 10331 235 10361 265
rect 10361 235 10366 265
rect 10326 230 10366 235
rect 10566 265 10606 270
rect 10566 235 10571 265
rect 10571 235 10601 265
rect 10601 235 10606 265
rect 10566 230 10606 235
rect 10811 265 10851 270
rect 10811 235 10816 265
rect 10816 235 10846 265
rect 10846 235 10851 265
rect 10811 230 10851 235
rect 11051 265 11091 270
rect 11051 235 11056 265
rect 11056 235 11086 265
rect 11086 235 11091 265
rect 11051 230 11091 235
rect 11305 270 11340 305
rect 11536 265 11576 270
rect 11536 235 11541 265
rect 11541 235 11571 265
rect 11571 235 11576 265
rect 11536 230 11576 235
rect 11781 265 11821 270
rect 11781 235 11786 265
rect 11786 235 11816 265
rect 11816 235 11821 265
rect 11781 230 11821 235
rect 12021 265 12061 270
rect 12021 235 12026 265
rect 12026 235 12056 265
rect 12056 235 12061 265
rect 12021 230 12061 235
rect 12266 265 12306 270
rect 12266 235 12271 265
rect 12271 235 12301 265
rect 12301 235 12306 265
rect 12266 230 12306 235
rect 12506 265 12546 270
rect 12506 235 12511 265
rect 12511 235 12541 265
rect 12541 235 12546 265
rect 12506 230 12546 235
rect 12751 265 12791 270
rect 12751 235 12756 265
rect 12756 235 12786 265
rect 12786 235 12791 265
rect 12751 230 12791 235
rect 13000 270 13035 305
rect 13236 265 13276 270
rect 13236 235 13241 265
rect 13241 235 13271 265
rect 13271 235 13276 265
rect 13236 230 13276 235
rect 13476 265 13516 270
rect 13476 235 13481 265
rect 13481 235 13511 265
rect 13511 235 13516 265
rect 13476 230 13516 235
rect 13721 265 13761 270
rect 13721 235 13726 265
rect 13726 235 13756 265
rect 13756 235 13761 265
rect 13721 230 13761 235
rect 13961 265 14001 270
rect 13961 235 13966 265
rect 13966 235 13996 265
rect 13996 235 14001 265
rect 13961 230 14001 235
rect 14206 265 14246 270
rect 14206 235 14211 265
rect 14211 235 14241 265
rect 14241 235 14246 265
rect 14206 230 14246 235
rect 14446 265 14486 270
rect 14446 235 14451 265
rect 14451 235 14481 265
rect 14481 235 14486 265
rect 14446 230 14486 235
rect 14691 265 14731 270
rect 14691 235 14696 265
rect 14696 235 14726 265
rect 14726 235 14731 265
rect 14691 230 14731 235
rect 14931 265 14971 270
rect 14931 235 14936 265
rect 14936 235 14966 265
rect 14966 235 14971 265
rect 14931 230 14971 235
rect 15185 270 15220 305
rect 15416 265 15456 270
rect 15416 235 15421 265
rect 15421 235 15451 265
rect 15451 235 15456 265
rect 15416 230 15456 235
rect 15661 265 15701 270
rect 15661 235 15666 265
rect 15666 235 15696 265
rect 15696 235 15701 265
rect 15661 230 15701 235
rect 15901 265 15941 270
rect 15901 235 15906 265
rect 15906 235 15936 265
rect 15936 235 15941 265
rect 15901 230 15941 235
rect 16146 265 16186 270
rect 16146 235 16151 265
rect 16151 235 16181 265
rect 16181 235 16186 265
rect 16146 230 16186 235
rect 16386 265 16426 270
rect 16386 235 16391 265
rect 16391 235 16421 265
rect 16421 235 16426 265
rect 16386 230 16426 235
rect 16631 265 16671 270
rect 16631 235 16636 265
rect 16636 235 16666 265
rect 16666 235 16671 265
rect 16631 230 16671 235
rect 16871 265 16911 270
rect 16871 235 16876 265
rect 16876 235 16906 265
rect 16906 235 16911 265
rect 16871 230 16911 235
rect 17116 265 17156 270
rect 17116 235 17121 265
rect 17121 235 17151 265
rect 17151 235 17156 265
rect 17116 230 17156 235
rect 17365 270 17400 305
rect 17601 265 17641 270
rect 17601 235 17606 265
rect 17606 235 17636 265
rect 17636 235 17641 265
rect 17601 230 17641 235
rect 17841 265 17881 270
rect 17841 235 17846 265
rect 17846 235 17876 265
rect 17876 235 17881 265
rect 17841 230 17881 235
rect 18086 265 18126 270
rect 18086 235 18091 265
rect 18091 235 18121 265
rect 18121 235 18126 265
rect 18086 230 18126 235
rect 18326 265 18366 270
rect 18326 235 18331 265
rect 18331 235 18361 265
rect 18361 235 18366 265
rect 18326 230 18366 235
rect 18571 265 18611 270
rect 18571 235 18576 265
rect 18576 235 18606 265
rect 18606 235 18611 265
rect 18571 230 18611 235
rect 18811 265 18851 270
rect 18811 235 18816 265
rect 18816 235 18846 265
rect 18846 235 18851 265
rect 18811 230 18851 235
rect 19056 265 19096 270
rect 19056 235 19061 265
rect 19061 235 19091 265
rect 19091 235 19096 265
rect 19056 230 19096 235
rect 19296 265 19336 270
rect 19296 235 19301 265
rect 19301 235 19331 265
rect 19331 235 19336 265
rect 19296 230 19336 235
rect 19550 270 19585 305
rect 19781 265 19821 270
rect 19781 235 19786 265
rect 19786 235 19816 265
rect 19816 235 19821 265
rect 19781 230 19821 235
rect 20026 265 20066 270
rect 20026 235 20031 265
rect 20031 235 20061 265
rect 20061 235 20066 265
rect 20026 230 20066 235
rect 20266 265 20306 270
rect 20266 235 20271 265
rect 20271 235 20301 265
rect 20301 235 20306 265
rect 20266 230 20306 235
rect 20511 265 20551 270
rect 20511 235 20516 265
rect 20516 235 20546 265
rect 20546 235 20551 265
rect 20511 230 20551 235
rect 20760 270 20795 305
rect 20996 265 21036 270
rect 20996 235 21001 265
rect 21001 235 21031 265
rect 21031 235 21036 265
rect 20996 230 21036 235
rect -25 -240 25 -190
rect 181 -165 221 -160
rect 181 -195 186 -165
rect 186 -195 216 -165
rect 216 -195 221 -165
rect 181 -200 221 -195
rect 426 -165 466 -160
rect 426 -195 431 -165
rect 431 -195 461 -165
rect 461 -195 466 -165
rect 426 -200 466 -195
rect 731 -165 771 -160
rect 731 -195 736 -165
rect 736 -195 766 -165
rect 766 -195 771 -165
rect 731 -200 771 -195
rect 976 -165 1016 -160
rect 976 -195 981 -165
rect 981 -195 1011 -165
rect 1011 -195 1016 -165
rect 976 -200 1016 -195
rect 1216 -165 1256 -160
rect 1216 -195 1221 -165
rect 1221 -195 1251 -165
rect 1251 -195 1256 -165
rect 1216 -200 1256 -195
rect 1461 -165 1501 -160
rect 1461 -195 1466 -165
rect 1466 -195 1496 -165
rect 1496 -195 1501 -165
rect 1461 -200 1501 -195
rect 85 -245 125 -240
rect 85 -275 90 -245
rect 90 -275 120 -245
rect 120 -275 125 -245
rect 85 -280 125 -275
rect 325 -245 365 -240
rect 325 -275 330 -245
rect 330 -275 360 -245
rect 360 -275 365 -245
rect 325 -280 365 -275
rect 565 -245 605 -240
rect 565 -275 570 -245
rect 570 -275 600 -245
rect 600 -275 605 -245
rect 565 -280 605 -275
rect 805 -245 845 -240
rect 805 -275 810 -245
rect 810 -275 840 -245
rect 840 -275 845 -245
rect 805 -280 845 -275
rect 1045 -245 1085 -240
rect 1045 -275 1050 -245
rect 1050 -275 1080 -245
rect 1080 -275 1085 -245
rect 1045 -280 1085 -275
rect 1285 -245 1325 -240
rect 1285 -275 1290 -245
rect 1290 -275 1320 -245
rect 1320 -275 1325 -245
rect 1285 -280 1325 -275
rect 1525 -245 1565 -240
rect 1525 -275 1530 -245
rect 1530 -275 1560 -245
rect 1560 -275 1565 -245
rect 1525 -280 1565 -275
rect 1635 -240 1675 -200
rect 1766 -165 1806 -160
rect 1766 -195 1771 -165
rect 1771 -195 1801 -165
rect 1801 -195 1806 -165
rect 1766 -200 1806 -195
rect 2011 -165 2051 -160
rect 2011 -195 2016 -165
rect 2016 -195 2046 -165
rect 2046 -195 2051 -165
rect 2011 -200 2051 -195
rect 2251 -165 2291 -160
rect 2251 -195 2256 -165
rect 2256 -195 2286 -165
rect 2286 -195 2291 -165
rect 2251 -200 2291 -195
rect 2496 -165 2536 -160
rect 2496 -195 2501 -165
rect 2501 -195 2531 -165
rect 2531 -195 2536 -165
rect 2496 -200 2536 -195
rect 2736 -165 2776 -160
rect 2736 -195 2741 -165
rect 2741 -195 2771 -165
rect 2771 -195 2776 -165
rect 2736 -200 2776 -195
rect 2981 -165 3021 -160
rect 2981 -195 2986 -165
rect 2986 -195 3016 -165
rect 3016 -195 3021 -165
rect 2981 -200 3021 -195
rect 3221 -165 3261 -160
rect 3221 -195 3226 -165
rect 3226 -195 3256 -165
rect 3256 -195 3261 -165
rect 3221 -200 3261 -195
rect 3466 -165 3506 -160
rect 3466 -195 3471 -165
rect 3471 -195 3501 -165
rect 3501 -195 3506 -165
rect 3466 -200 3506 -195
rect 3706 -165 3746 -160
rect 3706 -195 3711 -165
rect 3711 -195 3741 -165
rect 3741 -195 3746 -165
rect 3706 -200 3746 -195
rect 3951 -165 3991 -160
rect 3951 -195 3956 -165
rect 3956 -195 3986 -165
rect 3986 -195 3991 -165
rect 3951 -200 3991 -195
rect 4060 -235 4100 -195
rect 4191 -165 4231 -160
rect 4191 -195 4196 -165
rect 4196 -195 4226 -165
rect 4226 -195 4231 -165
rect 4191 -200 4231 -195
rect 4436 -165 4476 -160
rect 4436 -195 4441 -165
rect 4441 -195 4471 -165
rect 4471 -195 4476 -165
rect 4436 -200 4476 -195
rect 4676 -165 4716 -160
rect 4676 -195 4681 -165
rect 4681 -195 4711 -165
rect 4711 -195 4716 -165
rect 4676 -200 4716 -195
rect 4921 -165 4961 -160
rect 4921 -195 4926 -165
rect 4926 -195 4956 -165
rect 4956 -195 4961 -165
rect 4921 -200 4961 -195
rect 5161 -165 5201 -160
rect 5161 -195 5166 -165
rect 5166 -195 5196 -165
rect 5196 -195 5201 -165
rect 5161 -200 5201 -195
rect 5406 -165 5446 -160
rect 5406 -195 5411 -165
rect 5411 -195 5441 -165
rect 5441 -195 5446 -165
rect 5406 -200 5446 -195
rect 5711 -165 5751 -160
rect 5711 -195 5716 -165
rect 5716 -195 5746 -165
rect 5746 -195 5751 -165
rect 5711 -200 5751 -195
rect 5956 -165 5996 -160
rect 5956 -195 5961 -165
rect 5961 -195 5991 -165
rect 5991 -195 5996 -165
rect 5956 -200 5996 -195
rect 6196 -165 6236 -160
rect 6196 -195 6201 -165
rect 6201 -195 6231 -165
rect 6231 -195 6236 -165
rect 6196 -200 6236 -195
rect 6681 -165 6721 -160
rect 6681 -195 6686 -165
rect 6686 -195 6716 -165
rect 6716 -195 6721 -165
rect 6681 -200 6721 -195
rect 6926 -165 6966 -160
rect 6926 -195 6931 -165
rect 6931 -195 6961 -165
rect 6961 -195 6966 -165
rect 6926 -200 6966 -195
rect 7166 -165 7206 -160
rect 7166 -195 7171 -165
rect 7171 -195 7201 -165
rect 7201 -195 7206 -165
rect 7166 -200 7206 -195
rect 7406 -165 7446 -160
rect 7406 -195 7411 -165
rect 7411 -195 7441 -165
rect 7441 -195 7446 -165
rect 7406 -200 7446 -195
rect 7646 -165 7686 -160
rect 7646 -195 7651 -165
rect 7651 -195 7681 -165
rect 7681 -195 7686 -165
rect 7646 -200 7686 -195
rect 8131 -165 8171 -160
rect 8131 -195 8136 -165
rect 8136 -195 8166 -165
rect 8166 -195 8171 -165
rect 8131 -200 8171 -195
rect 8376 -165 8416 -160
rect 8376 -195 8381 -165
rect 8381 -195 8411 -165
rect 8411 -195 8416 -165
rect 8376 -200 8416 -195
rect 8616 -165 8656 -160
rect 8616 -195 8621 -165
rect 8621 -195 8651 -165
rect 8651 -195 8656 -165
rect 8616 -200 8656 -195
rect 8861 -165 8901 -160
rect 8861 -195 8866 -165
rect 8866 -195 8896 -165
rect 8896 -195 8901 -165
rect 8861 -200 8901 -195
rect 9101 -165 9141 -160
rect 9101 -195 9106 -165
rect 9106 -195 9136 -165
rect 9136 -195 9141 -165
rect 9101 -200 9141 -195
rect 9346 -165 9386 -160
rect 9346 -195 9351 -165
rect 9351 -195 9381 -165
rect 9381 -195 9386 -165
rect 9346 -200 9386 -195
rect 9836 -165 9876 -160
rect 9836 -195 9841 -165
rect 9841 -195 9871 -165
rect 9871 -195 9876 -165
rect 9836 -200 9876 -195
rect 10076 -165 10116 -160
rect 10076 -195 10081 -165
rect 10081 -195 10111 -165
rect 10111 -195 10116 -165
rect 10076 -200 10116 -195
rect 10321 -165 10361 -160
rect 10321 -195 10326 -165
rect 10326 -195 10356 -165
rect 10356 -195 10361 -165
rect 10321 -200 10361 -195
rect 10561 -165 10601 -160
rect 10561 -195 10566 -165
rect 10566 -195 10596 -165
rect 10596 -195 10601 -165
rect 10561 -200 10601 -195
rect 10806 -165 10846 -160
rect 10806 -195 10811 -165
rect 10811 -195 10841 -165
rect 10841 -195 10846 -165
rect 10806 -200 10846 -195
rect 11046 -165 11086 -160
rect 11046 -195 11051 -165
rect 11051 -195 11081 -165
rect 11081 -195 11086 -165
rect 11046 -200 11086 -195
rect 11291 -165 11331 -160
rect 11291 -195 11296 -165
rect 11296 -195 11326 -165
rect 11326 -195 11331 -165
rect 11291 -200 11331 -195
rect 11531 -165 11571 -160
rect 11531 -195 11536 -165
rect 11536 -195 11566 -165
rect 11566 -195 11571 -165
rect 11531 -200 11571 -195
rect 11776 -165 11816 -160
rect 11776 -195 11781 -165
rect 11781 -195 11811 -165
rect 11811 -195 11816 -165
rect 11776 -200 11816 -195
rect 12261 -165 12301 -160
rect 12261 -195 12266 -165
rect 12266 -195 12296 -165
rect 12296 -195 12301 -165
rect 12261 -200 12301 -195
rect 12501 -165 12541 -160
rect 12501 -195 12506 -165
rect 12506 -195 12536 -165
rect 12536 -195 12541 -165
rect 12501 -200 12541 -195
rect 12746 -165 12786 -160
rect 12746 -195 12751 -165
rect 12751 -195 12781 -165
rect 12781 -195 12786 -165
rect 12746 -200 12786 -195
rect 12986 -165 13026 -160
rect 12986 -195 12991 -165
rect 12991 -195 13021 -165
rect 13021 -195 13026 -165
rect 12986 -200 13026 -195
rect 13231 -165 13271 -160
rect 13231 -195 13236 -165
rect 13236 -195 13266 -165
rect 13266 -195 13271 -165
rect 13231 -200 13271 -195
rect 13471 -165 13511 -160
rect 13471 -195 13476 -165
rect 13476 -195 13506 -165
rect 13506 -195 13511 -165
rect 13471 -200 13511 -195
rect 13716 -165 13756 -160
rect 13716 -195 13721 -165
rect 13721 -195 13751 -165
rect 13751 -195 13756 -165
rect 13716 -200 13756 -195
rect 14201 -165 14241 -160
rect 14201 -195 14206 -165
rect 14206 -195 14236 -165
rect 14236 -195 14241 -165
rect 14201 -200 14241 -195
rect 14441 -165 14481 -160
rect 14441 -195 14446 -165
rect 14446 -195 14476 -165
rect 14476 -195 14481 -165
rect 14441 -200 14481 -195
rect 14686 -165 14726 -160
rect 14686 -195 14691 -165
rect 14691 -195 14721 -165
rect 14721 -195 14726 -165
rect 14686 -200 14726 -195
rect 14926 -165 14966 -160
rect 14926 -195 14931 -165
rect 14931 -195 14961 -165
rect 14961 -195 14966 -165
rect 14926 -200 14966 -195
rect 15171 -165 15211 -160
rect 15171 -195 15176 -165
rect 15176 -195 15206 -165
rect 15206 -195 15211 -165
rect 15171 -200 15211 -195
rect 15411 -165 15451 -160
rect 15411 -195 15416 -165
rect 15416 -195 15446 -165
rect 15446 -195 15451 -165
rect 15411 -200 15451 -195
rect 15656 -165 15696 -160
rect 15656 -195 15661 -165
rect 15661 -195 15691 -165
rect 15691 -195 15696 -165
rect 15656 -200 15696 -195
rect 16141 -165 16181 -160
rect 16141 -195 16146 -165
rect 16146 -195 16176 -165
rect 16176 -195 16181 -165
rect 16141 -200 16181 -195
rect 16381 -165 16421 -160
rect 16381 -195 16386 -165
rect 16386 -195 16416 -165
rect 16416 -195 16421 -165
rect 16381 -200 16421 -195
rect 16626 -165 16666 -160
rect 16626 -195 16631 -165
rect 16631 -195 16661 -165
rect 16661 -195 16666 -165
rect 16626 -200 16666 -195
rect 16866 -165 16906 -160
rect 16866 -195 16871 -165
rect 16871 -195 16901 -165
rect 16901 -195 16906 -165
rect 16866 -200 16906 -195
rect 17111 -165 17151 -160
rect 17111 -195 17116 -165
rect 17116 -195 17146 -165
rect 17146 -195 17151 -165
rect 17111 -200 17151 -195
rect 17351 -165 17391 -160
rect 17351 -195 17356 -165
rect 17356 -195 17386 -165
rect 17386 -195 17391 -165
rect 17351 -200 17391 -195
rect 17596 -165 17636 -160
rect 17596 -195 17601 -165
rect 17601 -195 17631 -165
rect 17631 -195 17636 -165
rect 17596 -200 17636 -195
rect 17836 -165 17876 -160
rect 17836 -195 17841 -165
rect 17841 -195 17871 -165
rect 17871 -195 17876 -165
rect 17836 -200 17876 -195
rect 18081 -165 18121 -160
rect 18081 -195 18086 -165
rect 18086 -195 18116 -165
rect 18116 -195 18121 -165
rect 18081 -200 18121 -195
rect 18321 -165 18361 -160
rect 18321 -195 18326 -165
rect 18326 -195 18356 -165
rect 18356 -195 18361 -165
rect 18321 -200 18361 -195
rect 18566 -165 18606 -160
rect 18566 -195 18571 -165
rect 18571 -195 18601 -165
rect 18601 -195 18606 -165
rect 18566 -200 18606 -195
rect 18806 -165 18846 -160
rect 18806 -195 18811 -165
rect 18811 -195 18841 -165
rect 18841 -195 18846 -165
rect 18806 -200 18846 -195
rect 19051 -165 19091 -160
rect 19051 -195 19056 -165
rect 19056 -195 19086 -165
rect 19086 -195 19091 -165
rect 19051 -200 19091 -195
rect 19291 -165 19331 -160
rect 19291 -195 19296 -165
rect 19296 -195 19326 -165
rect 19326 -195 19331 -165
rect 19291 -200 19331 -195
rect 19536 -165 19576 -160
rect 19536 -195 19541 -165
rect 19541 -195 19571 -165
rect 19571 -195 19576 -165
rect 19536 -200 19576 -195
rect 19776 -165 19816 -160
rect 19776 -195 19781 -165
rect 19781 -195 19811 -165
rect 19811 -195 19816 -165
rect 19776 -200 19816 -195
rect 1765 -245 1805 -240
rect 1765 -275 1770 -245
rect 1770 -275 1800 -245
rect 1800 -275 1805 -245
rect 1765 -280 1805 -275
rect 2005 -245 2045 -240
rect 2005 -275 2010 -245
rect 2010 -275 2040 -245
rect 2040 -275 2045 -245
rect 2005 -280 2045 -275
rect 2245 -245 2285 -240
rect 2245 -275 2250 -245
rect 2250 -275 2280 -245
rect 2280 -275 2285 -245
rect 2245 -280 2285 -275
rect 2485 -245 2525 -240
rect 2485 -275 2490 -245
rect 2490 -275 2520 -245
rect 2520 -275 2525 -245
rect 2485 -280 2525 -275
rect 2725 -245 2765 -240
rect 2725 -275 2730 -245
rect 2730 -275 2760 -245
rect 2760 -275 2765 -245
rect 2725 -280 2765 -275
rect 2965 -245 3005 -240
rect 2965 -275 2970 -245
rect 2970 -275 3000 -245
rect 3000 -275 3005 -245
rect 2965 -280 3005 -275
rect 3205 -245 3245 -240
rect 3205 -275 3210 -245
rect 3210 -275 3240 -245
rect 3240 -275 3245 -245
rect 3205 -280 3245 -275
rect 3445 -245 3485 -240
rect 3445 -275 3450 -245
rect 3450 -275 3480 -245
rect 3480 -275 3485 -245
rect 3445 -280 3485 -275
rect 3685 -245 3725 -240
rect 3685 -275 3690 -245
rect 3690 -275 3720 -245
rect 3720 -275 3725 -245
rect 3685 -280 3725 -275
rect 3925 -245 3965 -240
rect 3925 -275 3930 -245
rect 3930 -275 3960 -245
rect 3960 -275 3965 -245
rect 3925 -280 3965 -275
rect 4165 -245 4205 -240
rect 4165 -275 4170 -245
rect 4170 -275 4200 -245
rect 4200 -275 4205 -245
rect 4165 -280 4205 -275
rect 4405 -245 4445 -240
rect 4405 -275 4410 -245
rect 4410 -275 4440 -245
rect 4440 -275 4445 -245
rect 4405 -280 4445 -275
rect 4645 -245 4685 -240
rect 4645 -275 4650 -245
rect 4650 -275 4680 -245
rect 4680 -275 4685 -245
rect 4645 -280 4685 -275
rect 4885 -245 4925 -240
rect 4885 -275 4890 -245
rect 4890 -275 4920 -245
rect 4920 -275 4925 -245
rect 4885 -280 4925 -275
rect 5125 -245 5165 -240
rect 5125 -275 5130 -245
rect 5130 -275 5160 -245
rect 5160 -275 5165 -245
rect 5125 -280 5165 -275
rect 5365 -245 5405 -240
rect 5365 -275 5370 -245
rect 5370 -275 5400 -245
rect 5400 -275 5405 -245
rect 5365 -280 5405 -275
rect 5605 -245 5645 -240
rect 5605 -275 5610 -245
rect 5610 -275 5640 -245
rect 5640 -275 5645 -245
rect 5605 -280 5645 -275
rect 5845 -245 5885 -240
rect 5845 -275 5850 -245
rect 5850 -275 5880 -245
rect 5880 -275 5885 -245
rect 5845 -280 5885 -275
rect 6085 -245 6125 -240
rect 6085 -275 6090 -245
rect 6090 -275 6120 -245
rect 6120 -275 6125 -245
rect 6085 -280 6125 -275
rect 6325 -245 6365 -240
rect 6325 -275 6330 -245
rect 6330 -275 6360 -245
rect 6360 -275 6365 -245
rect 6325 -280 6365 -275
rect 6455 -260 6495 -220
rect 6565 -245 6605 -240
rect 6565 -275 6570 -245
rect 6570 -275 6600 -245
rect 6600 -275 6605 -245
rect 6565 -280 6605 -275
rect 6805 -245 6845 -240
rect 6805 -275 6810 -245
rect 6810 -275 6840 -245
rect 6840 -275 6845 -245
rect 6805 -280 6845 -275
rect 7045 -245 7085 -240
rect 7045 -275 7050 -245
rect 7050 -275 7080 -245
rect 7080 -275 7085 -245
rect 7045 -280 7085 -275
rect 7285 -245 7325 -240
rect 7285 -275 7290 -245
rect 7290 -275 7320 -245
rect 7320 -275 7325 -245
rect 7285 -280 7325 -275
rect 7525 -245 7565 -240
rect 7525 -275 7530 -245
rect 7530 -275 7560 -245
rect 7560 -275 7565 -245
rect 7525 -280 7565 -275
rect 7765 -245 7805 -240
rect 7765 -275 7770 -245
rect 7770 -275 7800 -245
rect 7800 -275 7805 -245
rect 7765 -280 7805 -275
rect 7880 -260 7920 -220
rect 8005 -245 8045 -240
rect 8005 -275 8010 -245
rect 8010 -275 8040 -245
rect 8040 -275 8045 -245
rect 8005 -280 8045 -275
rect 8245 -245 8285 -240
rect 8245 -275 8250 -245
rect 8250 -275 8280 -245
rect 8280 -275 8285 -245
rect 8245 -280 8285 -275
rect 8485 -245 8525 -240
rect 8485 -275 8490 -245
rect 8490 -275 8520 -245
rect 8520 -275 8525 -245
rect 8485 -280 8525 -275
rect 8725 -245 8765 -240
rect 8725 -275 8730 -245
rect 8730 -275 8760 -245
rect 8760 -275 8765 -245
rect 8725 -280 8765 -275
rect 8965 -245 9005 -240
rect 8965 -275 8970 -245
rect 8970 -275 9000 -245
rect 9000 -275 9005 -245
rect 8965 -280 9005 -275
rect 9205 -245 9245 -240
rect 9205 -275 9210 -245
rect 9210 -275 9240 -245
rect 9240 -275 9245 -245
rect 9205 -280 9245 -275
rect 9445 -245 9485 -240
rect 9445 -275 9450 -245
rect 9450 -275 9480 -245
rect 9480 -275 9485 -245
rect 9445 -280 9485 -275
rect 9570 -250 9610 -210
rect 9685 -245 9725 -240
rect 9685 -275 9690 -245
rect 9690 -275 9720 -245
rect 9720 -275 9725 -245
rect 9685 -280 9725 -275
rect 9925 -245 9965 -240
rect 9925 -275 9930 -245
rect 9930 -275 9960 -245
rect 9960 -275 9965 -245
rect 9925 -280 9965 -275
rect 10165 -245 10205 -240
rect 10165 -275 10170 -245
rect 10170 -275 10200 -245
rect 10200 -275 10205 -245
rect 10165 -280 10205 -275
rect 10405 -245 10445 -240
rect 10405 -275 10410 -245
rect 10410 -275 10440 -245
rect 10440 -275 10445 -245
rect 10405 -280 10445 -275
rect 10645 -245 10685 -240
rect 10645 -275 10650 -245
rect 10650 -275 10680 -245
rect 10680 -275 10685 -245
rect 10645 -280 10685 -275
rect 10885 -245 10925 -240
rect 10885 -275 10890 -245
rect 10890 -275 10920 -245
rect 10920 -275 10925 -245
rect 10885 -280 10925 -275
rect 11125 -245 11165 -240
rect 11125 -275 11130 -245
rect 11130 -275 11160 -245
rect 11160 -275 11165 -245
rect 11125 -280 11165 -275
rect 11365 -245 11405 -240
rect 11365 -275 11370 -245
rect 11370 -275 11400 -245
rect 11400 -275 11405 -245
rect 11365 -280 11405 -275
rect 11605 -245 11645 -240
rect 11605 -275 11610 -245
rect 11610 -275 11640 -245
rect 11640 -275 11645 -245
rect 11605 -280 11645 -275
rect 11845 -245 11885 -240
rect 11845 -275 11850 -245
rect 11850 -275 11880 -245
rect 11880 -275 11885 -245
rect 11845 -280 11885 -275
rect 11950 -260 11990 -220
rect 12085 -245 12125 -240
rect 12085 -275 12090 -245
rect 12090 -275 12120 -245
rect 12120 -275 12125 -245
rect 12085 -280 12125 -275
rect 12325 -245 12365 -240
rect 12325 -275 12330 -245
rect 12330 -275 12360 -245
rect 12360 -275 12365 -245
rect 12325 -280 12365 -275
rect 12565 -245 12605 -240
rect 12565 -275 12570 -245
rect 12570 -275 12600 -245
rect 12600 -275 12605 -245
rect 12565 -280 12605 -275
rect 12805 -245 12845 -240
rect 12805 -275 12810 -245
rect 12810 -275 12840 -245
rect 12840 -275 12845 -245
rect 12805 -280 12845 -275
rect 13045 -245 13085 -240
rect 13045 -275 13050 -245
rect 13050 -275 13080 -245
rect 13080 -275 13085 -245
rect 13045 -280 13085 -275
rect 13285 -245 13325 -240
rect 13285 -275 13290 -245
rect 13290 -275 13320 -245
rect 13320 -275 13325 -245
rect 13285 -280 13325 -275
rect 13525 -245 13565 -240
rect 13525 -275 13530 -245
rect 13530 -275 13560 -245
rect 13560 -275 13565 -245
rect 13525 -280 13565 -275
rect 13765 -245 13805 -240
rect 13765 -275 13770 -245
rect 13770 -275 13800 -245
rect 13800 -275 13805 -245
rect 13765 -280 13805 -275
rect 13870 -260 13910 -220
rect 14005 -245 14045 -240
rect 14005 -275 14010 -245
rect 14010 -275 14040 -245
rect 14040 -275 14045 -245
rect 14005 -280 14045 -275
rect 14245 -245 14285 -240
rect 14245 -275 14250 -245
rect 14250 -275 14280 -245
rect 14280 -275 14285 -245
rect 14245 -280 14285 -275
rect 14485 -245 14525 -240
rect 14485 -275 14490 -245
rect 14490 -275 14520 -245
rect 14520 -275 14525 -245
rect 14485 -280 14525 -275
rect 14725 -245 14765 -240
rect 14725 -275 14730 -245
rect 14730 -275 14760 -245
rect 14760 -275 14765 -245
rect 14725 -280 14765 -275
rect 14965 -245 15005 -240
rect 14965 -275 14970 -245
rect 14970 -275 15000 -245
rect 15000 -275 15005 -245
rect 14965 -280 15005 -275
rect 15205 -245 15245 -240
rect 15205 -275 15210 -245
rect 15210 -275 15240 -245
rect 15240 -275 15245 -245
rect 15205 -280 15245 -275
rect 15445 -245 15485 -240
rect 15445 -275 15450 -245
rect 15450 -275 15480 -245
rect 15480 -275 15485 -245
rect 15445 -280 15485 -275
rect 15685 -245 15725 -240
rect 15685 -275 15690 -245
rect 15690 -275 15720 -245
rect 15720 -275 15725 -245
rect 15685 -280 15725 -275
rect 15815 -260 15855 -220
rect 15925 -245 15965 -240
rect 15925 -275 15930 -245
rect 15930 -275 15960 -245
rect 15960 -275 15965 -245
rect 15925 -280 15965 -275
rect 16165 -245 16205 -240
rect 16165 -275 16170 -245
rect 16170 -275 16200 -245
rect 16200 -275 16205 -245
rect 16165 -280 16205 -275
rect 16405 -245 16445 -240
rect 16405 -275 16410 -245
rect 16410 -275 16440 -245
rect 16440 -275 16445 -245
rect 16405 -280 16445 -275
rect 16645 -245 16685 -240
rect 16645 -275 16650 -245
rect 16650 -275 16680 -245
rect 16680 -275 16685 -245
rect 16645 -280 16685 -275
rect 16885 -245 16925 -240
rect 16885 -275 16890 -245
rect 16890 -275 16920 -245
rect 16920 -275 16925 -245
rect 16885 -280 16925 -275
rect 17125 -245 17165 -240
rect 17125 -275 17130 -245
rect 17130 -275 17160 -245
rect 17160 -275 17165 -245
rect 17125 -280 17165 -275
rect 17365 -245 17405 -240
rect 17365 -275 17370 -245
rect 17370 -275 17400 -245
rect 17400 -275 17405 -245
rect 17365 -280 17405 -275
rect 17605 -245 17645 -240
rect 17605 -275 17610 -245
rect 17610 -275 17640 -245
rect 17640 -275 17645 -245
rect 17605 -280 17645 -275
rect 17705 -250 17745 -210
rect 20021 -165 20061 -160
rect 20021 -195 20026 -165
rect 20026 -195 20056 -165
rect 20056 -195 20061 -165
rect 20021 -200 20061 -195
rect 20261 -165 20301 -160
rect 20261 -195 20266 -165
rect 20266 -195 20296 -165
rect 20296 -195 20301 -165
rect 20261 -200 20301 -195
rect 20506 -165 20546 -160
rect 20506 -195 20511 -165
rect 20511 -195 20541 -165
rect 20541 -195 20546 -165
rect 20506 -200 20546 -195
rect 20746 -165 20786 -160
rect 20746 -195 20751 -165
rect 20751 -195 20781 -165
rect 20781 -195 20786 -165
rect 20746 -200 20786 -195
rect 20991 -165 21031 -160
rect 20991 -195 20996 -165
rect 20996 -195 21026 -165
rect 21026 -195 21031 -165
rect 20991 -200 21031 -195
rect 17845 -245 17885 -240
rect 17845 -275 17850 -245
rect 17850 -275 17880 -245
rect 17880 -275 17885 -245
rect 17845 -280 17885 -275
rect 18085 -245 18125 -240
rect 18085 -275 18090 -245
rect 18090 -275 18120 -245
rect 18120 -275 18125 -245
rect 18085 -280 18125 -275
rect 18325 -245 18365 -240
rect 18325 -275 18330 -245
rect 18330 -275 18360 -245
rect 18360 -275 18365 -245
rect 18325 -280 18365 -275
rect 18565 -245 18605 -240
rect 18565 -275 18570 -245
rect 18570 -275 18600 -245
rect 18600 -275 18605 -245
rect 18565 -280 18605 -275
rect 18805 -245 18845 -240
rect 18805 -275 18810 -245
rect 18810 -275 18840 -245
rect 18840 -275 18845 -245
rect 18805 -280 18845 -275
rect 19045 -245 19085 -240
rect 19045 -275 19050 -245
rect 19050 -275 19080 -245
rect 19080 -275 19085 -245
rect 19045 -280 19085 -275
rect 19285 -245 19325 -240
rect 19285 -275 19290 -245
rect 19290 -275 19320 -245
rect 19320 -275 19325 -245
rect 19285 -280 19325 -275
rect 19525 -245 19565 -240
rect 19525 -275 19530 -245
rect 19530 -275 19560 -245
rect 19560 -275 19565 -245
rect 19525 -280 19565 -275
rect 19645 -250 19685 -210
rect 19765 -245 19805 -240
rect 19765 -275 19770 -245
rect 19770 -275 19800 -245
rect 19800 -275 19805 -245
rect 19765 -280 19805 -275
rect 20005 -245 20045 -240
rect 20005 -275 20010 -245
rect 20010 -275 20040 -245
rect 20040 -275 20045 -245
rect 20005 -280 20045 -275
rect 20245 -245 20285 -240
rect 20245 -275 20250 -245
rect 20250 -275 20280 -245
rect 20280 -275 20285 -245
rect 20245 -280 20285 -275
rect 20485 -245 20525 -240
rect 20485 -275 20490 -245
rect 20490 -275 20520 -245
rect 20520 -275 20525 -245
rect 20485 -280 20525 -275
rect 20725 -245 20765 -240
rect 20725 -275 20730 -245
rect 20730 -275 20760 -245
rect 20760 -275 20765 -245
rect 20725 -280 20765 -275
rect 20965 -245 21005 -240
rect 20965 -275 20970 -245
rect 20970 -275 21000 -245
rect 21000 -275 21005 -245
rect 20965 -280 21005 -275
rect 21205 -245 21245 -240
rect 21205 -275 21210 -245
rect 21210 -275 21240 -245
rect 21240 -275 21245 -245
rect 21205 -280 21245 -275
rect 21445 -245 21485 -240
rect 21445 -275 21450 -245
rect 21450 -275 21480 -245
rect 21480 -275 21485 -245
rect 21445 -280 21485 -275
rect 21685 -245 21725 -240
rect 21685 -275 21690 -245
rect 21690 -275 21720 -245
rect 21720 -275 21725 -245
rect 21685 -280 21725 -275
rect 21925 -245 21965 -240
rect 21925 -275 21930 -245
rect 21930 -275 21960 -245
rect 21960 -275 21965 -245
rect 21925 -280 21965 -275
rect 22165 -245 22205 -240
rect 22165 -275 22170 -245
rect 22170 -275 22200 -245
rect 22200 -275 22205 -245
rect 22165 -280 22205 -275
rect 22405 -245 22445 -240
rect 22405 -275 22410 -245
rect 22410 -275 22440 -245
rect 22440 -275 22445 -245
rect 22405 -280 22445 -275
rect 22645 -245 22685 -240
rect 22645 -275 22650 -245
rect 22650 -275 22680 -245
rect 22680 -275 22685 -245
rect 22645 -280 22685 -275
rect 22885 -245 22925 -240
rect 22885 -275 22890 -245
rect 22890 -275 22920 -245
rect 22920 -275 22925 -245
rect 22885 -280 22925 -275
rect 23125 -245 23165 -240
rect 23125 -275 23130 -245
rect 23130 -275 23160 -245
rect 23160 -275 23165 -245
rect 23125 -280 23165 -275
rect 23365 -245 23405 -240
rect 23365 -275 23370 -245
rect 23370 -275 23400 -245
rect 23400 -275 23405 -245
rect 23365 -280 23405 -275
rect 23605 -245 23645 -240
rect 23605 -275 23610 -245
rect 23610 -275 23640 -245
rect 23640 -275 23645 -245
rect 23605 -280 23645 -275
rect 23845 -245 23885 -240
rect 23845 -275 23850 -245
rect 23850 -275 23880 -245
rect 23880 -275 23885 -245
rect 23845 -280 23885 -275
rect 24085 -245 24125 -240
rect 24085 -275 24090 -245
rect 24090 -275 24120 -245
rect 24120 -275 24125 -245
rect 24085 -280 24125 -275
rect 24325 -245 24365 -240
rect 24325 -275 24330 -245
rect 24330 -275 24360 -245
rect 24360 -275 24365 -245
rect 24325 -280 24365 -275
rect 24565 -245 24605 -240
rect 24565 -275 24570 -245
rect 24570 -275 24600 -245
rect 24600 -275 24605 -245
rect 24565 -280 24605 -275
rect 24805 -245 24845 -240
rect 24805 -275 24810 -245
rect 24810 -275 24840 -245
rect 24840 -275 24845 -245
rect 24805 -280 24845 -275
rect 25045 -245 25085 -240
rect 25045 -275 25050 -245
rect 25050 -275 25080 -245
rect 25080 -275 25085 -245
rect 25045 -280 25085 -275
rect 25285 -245 25325 -240
rect 25285 -275 25290 -245
rect 25290 -275 25320 -245
rect 25320 -275 25325 -245
rect 25285 -280 25325 -275
rect 25525 -245 25565 -240
rect 25525 -275 25530 -245
rect 25530 -275 25560 -245
rect 25560 -275 25565 -245
rect 25525 -280 25565 -275
rect 25765 -245 25805 -240
rect 25765 -275 25770 -245
rect 25770 -275 25800 -245
rect 25800 -275 25805 -245
rect 25765 -280 25805 -275
rect 26005 -245 26045 -240
rect 26005 -275 26010 -245
rect 26010 -275 26040 -245
rect 26040 -275 26045 -245
rect 26005 -280 26045 -275
rect 26245 -245 26285 -240
rect 26245 -275 26250 -245
rect 26250 -275 26280 -245
rect 26280 -275 26285 -245
rect 26245 -280 26285 -275
rect 26485 -245 26525 -240
rect 26485 -275 26490 -245
rect 26490 -275 26520 -245
rect 26520 -275 26525 -245
rect 26485 -280 26525 -275
rect 26725 -245 26765 -240
rect 26725 -275 26730 -245
rect 26730 -275 26760 -245
rect 26760 -275 26765 -245
rect 26725 -280 26765 -275
rect 26965 -245 27005 -240
rect 26965 -275 26970 -245
rect 26970 -275 27000 -245
rect 27000 -275 27005 -245
rect 26965 -280 27005 -275
rect 27205 -245 27245 -240
rect 27205 -275 27210 -245
rect 27210 -275 27240 -245
rect 27240 -275 27245 -245
rect 27205 -280 27245 -275
rect 27445 -245 27485 -240
rect 27445 -275 27450 -245
rect 27450 -275 27480 -245
rect 27480 -275 27485 -245
rect 27445 -280 27485 -275
rect 27685 -245 27725 -240
rect 27685 -275 27690 -245
rect 27690 -275 27720 -245
rect 27720 -275 27725 -245
rect 27685 -280 27725 -275
rect 27925 -245 27965 -240
rect 27925 -275 27930 -245
rect 27930 -275 27960 -245
rect 27960 -275 27965 -245
rect 27925 -280 27965 -275
rect 28165 -245 28205 -240
rect 28165 -275 28170 -245
rect 28170 -275 28200 -245
rect 28200 -275 28205 -245
rect 28165 -280 28205 -275
rect 28405 -245 28445 -240
rect 28405 -275 28410 -245
rect 28410 -275 28440 -245
rect 28440 -275 28445 -245
rect 28405 -280 28445 -275
rect 28645 -245 28685 -240
rect 28645 -275 28650 -245
rect 28650 -275 28680 -245
rect 28680 -275 28685 -245
rect 28645 -280 28685 -275
rect 28885 -245 28925 -240
rect 28885 -275 28890 -245
rect 28890 -275 28920 -245
rect 28920 -275 28925 -245
rect 28885 -280 28925 -275
rect 29125 -245 29165 -240
rect 29125 -275 29130 -245
rect 29130 -275 29160 -245
rect 29160 -275 29165 -245
rect 29125 -280 29165 -275
rect 29365 -245 29405 -240
rect 29365 -275 29370 -245
rect 29370 -275 29400 -245
rect 29400 -275 29405 -245
rect 29365 -280 29405 -275
rect 29605 -245 29645 -240
rect 29605 -275 29610 -245
rect 29610 -275 29640 -245
rect 29640 -275 29645 -245
rect 29605 -280 29645 -275
rect 29845 -245 29885 -240
rect 29845 -275 29850 -245
rect 29850 -275 29880 -245
rect 29880 -275 29885 -245
rect 29845 -280 29885 -275
rect 30085 -245 30125 -240
rect 30085 -275 30090 -245
rect 30090 -275 30120 -245
rect 30120 -275 30125 -245
rect 30085 -280 30125 -275
rect 30325 -245 30365 -240
rect 30325 -275 30330 -245
rect 30330 -275 30360 -245
rect 30360 -275 30365 -245
rect 30325 -280 30365 -275
rect 30565 -245 30605 -240
rect 30565 -275 30570 -245
rect 30570 -275 30600 -245
rect 30600 -275 30605 -245
rect 30565 -280 30605 -275
rect 80 -820 120 -815
rect 80 -850 85 -820
rect 85 -850 115 -820
rect 115 -850 120 -820
rect 80 -855 120 -850
rect 320 -820 360 -815
rect 320 -850 325 -820
rect 325 -850 355 -820
rect 355 -850 360 -820
rect 320 -855 360 -850
rect 560 -820 600 -815
rect 560 -850 565 -820
rect 565 -850 595 -820
rect 595 -850 600 -820
rect 560 -855 600 -850
rect 800 -870 835 -835
rect 1040 -820 1080 -815
rect 1040 -850 1045 -820
rect 1045 -850 1075 -820
rect 1075 -850 1080 -820
rect 1040 -855 1080 -850
rect 1280 -820 1320 -815
rect 1280 -850 1285 -820
rect 1285 -850 1315 -820
rect 1315 -850 1320 -820
rect 1280 -855 1320 -850
rect 1520 -820 1560 -815
rect 1520 -850 1525 -820
rect 1525 -850 1555 -820
rect 1555 -850 1560 -820
rect 1520 -855 1560 -850
rect 1760 -820 1800 -815
rect 1760 -850 1765 -820
rect 1765 -850 1795 -820
rect 1795 -850 1800 -820
rect 1760 -855 1800 -850
rect 2000 -820 2040 -815
rect 2000 -850 2005 -820
rect 2005 -850 2035 -820
rect 2035 -850 2040 -820
rect 2000 -855 2040 -850
rect 2240 -820 2280 -815
rect 2240 -850 2245 -820
rect 2245 -850 2275 -820
rect 2275 -850 2280 -820
rect 2240 -855 2280 -850
rect 2480 -820 2520 -815
rect 2480 -850 2485 -820
rect 2485 -850 2515 -820
rect 2515 -850 2520 -820
rect 2480 -855 2520 -850
rect 2720 -820 2760 -815
rect 2720 -850 2725 -820
rect 2725 -850 2755 -820
rect 2755 -850 2760 -820
rect 2720 -855 2760 -850
rect 2960 -870 2995 -835
rect 3200 -820 3240 -815
rect 3200 -850 3205 -820
rect 3205 -850 3235 -820
rect 3235 -850 3240 -820
rect 3200 -855 3240 -850
rect 3440 -820 3480 -815
rect 3440 -850 3445 -820
rect 3445 -850 3475 -820
rect 3475 -850 3480 -820
rect 3440 -855 3480 -850
rect 3680 -820 3720 -815
rect 3680 -850 3685 -820
rect 3685 -850 3715 -820
rect 3715 -850 3720 -820
rect 3680 -855 3720 -850
rect 3920 -820 3960 -815
rect 3920 -850 3925 -820
rect 3925 -850 3955 -820
rect 3955 -850 3960 -820
rect 3920 -855 3960 -850
rect 4160 -820 4200 -815
rect 4160 -850 4165 -820
rect 4165 -850 4195 -820
rect 4195 -850 4200 -820
rect 4160 -855 4200 -850
rect 4400 -820 4440 -815
rect 4400 -850 4405 -820
rect 4405 -850 4435 -820
rect 4435 -850 4440 -820
rect 4400 -855 4440 -850
rect 4640 -820 4680 -815
rect 4640 -850 4645 -820
rect 4645 -850 4675 -820
rect 4675 -850 4680 -820
rect 4640 -855 4680 -850
rect 4880 -820 4920 -815
rect 4880 -850 4885 -820
rect 4885 -850 4915 -820
rect 4915 -850 4920 -820
rect 4880 -855 4920 -850
rect 5120 -870 5155 -835
rect 5360 -820 5400 -815
rect 5360 -850 5365 -820
rect 5365 -850 5395 -820
rect 5395 -850 5400 -820
rect 5360 -855 5400 -850
rect 5600 -820 5640 -815
rect 5600 -850 5605 -820
rect 5605 -850 5635 -820
rect 5635 -850 5640 -820
rect 5600 -855 5640 -850
rect 5840 -820 5880 -815
rect 5840 -850 5845 -820
rect 5845 -850 5875 -820
rect 5875 -850 5880 -820
rect 5840 -855 5880 -850
rect 6080 -820 6120 -815
rect 6080 -850 6085 -820
rect 6085 -850 6115 -820
rect 6115 -850 6120 -820
rect 6080 -855 6120 -850
rect 6320 -820 6360 -815
rect 6320 -850 6325 -820
rect 6325 -850 6355 -820
rect 6355 -850 6360 -820
rect 6320 -855 6360 -850
rect 6560 -820 6600 -815
rect 6560 -850 6565 -820
rect 6565 -850 6595 -820
rect 6595 -850 6600 -820
rect 6560 -855 6600 -850
rect 6800 -820 6840 -815
rect 6800 -850 6805 -820
rect 6805 -850 6835 -820
rect 6835 -850 6840 -820
rect 6800 -855 6840 -850
rect 7040 -820 7080 -815
rect 7040 -850 7045 -820
rect 7045 -850 7075 -820
rect 7075 -850 7080 -820
rect 7040 -855 7080 -850
rect 7280 -870 7315 -835
rect 7520 -820 7560 -815
rect 7520 -850 7525 -820
rect 7525 -850 7555 -820
rect 7555 -850 7560 -820
rect 7520 -855 7560 -850
rect 7760 -820 7800 -815
rect 7760 -850 7765 -820
rect 7765 -850 7795 -820
rect 7795 -850 7800 -820
rect 7760 -855 7800 -850
rect 8000 -820 8040 -815
rect 8000 -850 8005 -820
rect 8005 -850 8035 -820
rect 8035 -850 8040 -820
rect 8000 -855 8040 -850
rect 8240 -820 8280 -815
rect 8240 -850 8245 -820
rect 8245 -850 8275 -820
rect 8275 -850 8280 -820
rect 8240 -855 8280 -850
rect 8480 -820 8520 -815
rect 8480 -850 8485 -820
rect 8485 -850 8515 -820
rect 8515 -850 8520 -820
rect 8480 -855 8520 -850
rect 8720 -820 8760 -815
rect 8720 -850 8725 -820
rect 8725 -850 8755 -820
rect 8755 -850 8760 -820
rect 8720 -855 8760 -850
rect 8960 -820 9000 -815
rect 8960 -850 8965 -820
rect 8965 -850 8995 -820
rect 8995 -850 9000 -820
rect 8960 -855 9000 -850
rect 9200 -820 9240 -815
rect 9200 -850 9205 -820
rect 9205 -850 9235 -820
rect 9235 -850 9240 -820
rect 9200 -855 9240 -850
rect 9440 -870 9475 -835
rect 9680 -820 9720 -815
rect 9680 -850 9685 -820
rect 9685 -850 9715 -820
rect 9715 -850 9720 -820
rect 9680 -855 9720 -850
rect 9920 -820 9960 -815
rect 9920 -850 9925 -820
rect 9925 -850 9955 -820
rect 9955 -850 9960 -820
rect 9920 -855 9960 -850
rect 10160 -820 10200 -815
rect 10160 -850 10165 -820
rect 10165 -850 10195 -820
rect 10195 -850 10200 -820
rect 10160 -855 10200 -850
rect 10400 -820 10440 -815
rect 10400 -850 10405 -820
rect 10405 -850 10435 -820
rect 10435 -850 10440 -820
rect 10400 -855 10440 -850
rect 10640 -820 10680 -815
rect 10640 -850 10645 -820
rect 10645 -850 10675 -820
rect 10675 -850 10680 -820
rect 10640 -855 10680 -850
rect 10880 -820 10920 -815
rect 10880 -850 10885 -820
rect 10885 -850 10915 -820
rect 10915 -850 10920 -820
rect 10880 -855 10920 -850
rect 11120 -820 11160 -815
rect 11120 -850 11125 -820
rect 11125 -850 11155 -820
rect 11155 -850 11160 -820
rect 11120 -855 11160 -850
rect 11360 -820 11400 -815
rect 11360 -850 11365 -820
rect 11365 -850 11395 -820
rect 11395 -850 11400 -820
rect 11360 -855 11400 -850
rect 11600 -870 11635 -835
rect 11840 -820 11880 -815
rect 11840 -850 11845 -820
rect 11845 -850 11875 -820
rect 11875 -850 11880 -820
rect 11840 -855 11880 -850
rect 12080 -820 12120 -815
rect 12080 -850 12085 -820
rect 12085 -850 12115 -820
rect 12115 -850 12120 -820
rect 12080 -855 12120 -850
rect 12320 -820 12360 -815
rect 12320 -850 12325 -820
rect 12325 -850 12355 -820
rect 12355 -850 12360 -820
rect 12320 -855 12360 -850
rect 12560 -820 12600 -815
rect 12560 -850 12565 -820
rect 12565 -850 12595 -820
rect 12595 -850 12600 -820
rect 12560 -855 12600 -850
rect 12800 -820 12840 -815
rect 12800 -850 12805 -820
rect 12805 -850 12835 -820
rect 12835 -850 12840 -820
rect 12800 -855 12840 -850
rect 13040 -820 13080 -815
rect 13040 -850 13045 -820
rect 13045 -850 13075 -820
rect 13075 -850 13080 -820
rect 13040 -855 13080 -850
rect 13280 -820 13320 -815
rect 13280 -850 13285 -820
rect 13285 -850 13315 -820
rect 13315 -850 13320 -820
rect 13280 -855 13320 -850
rect 13520 -820 13560 -815
rect 13520 -850 13525 -820
rect 13525 -850 13555 -820
rect 13555 -850 13560 -820
rect 13520 -855 13560 -850
rect 13760 -870 13795 -835
rect 14000 -820 14040 -815
rect 14000 -850 14005 -820
rect 14005 -850 14035 -820
rect 14035 -850 14040 -820
rect 14000 -855 14040 -850
rect 14240 -820 14280 -815
rect 14240 -850 14245 -820
rect 14245 -850 14275 -820
rect 14275 -850 14280 -820
rect 14240 -855 14280 -850
rect 14480 -820 14520 -815
rect 14480 -850 14485 -820
rect 14485 -850 14515 -820
rect 14515 -850 14520 -820
rect 14480 -855 14520 -850
rect 14720 -820 14760 -815
rect 14720 -850 14725 -820
rect 14725 -850 14755 -820
rect 14755 -850 14760 -820
rect 14720 -855 14760 -850
rect 14960 -820 15000 -815
rect 14960 -850 14965 -820
rect 14965 -850 14995 -820
rect 14995 -850 15000 -820
rect 14960 -855 15000 -850
rect 15200 -820 15240 -815
rect 15200 -850 15205 -820
rect 15205 -850 15235 -820
rect 15235 -850 15240 -820
rect 15200 -855 15240 -850
rect 15440 -820 15480 -815
rect 15440 -850 15445 -820
rect 15445 -850 15475 -820
rect 15475 -850 15480 -820
rect 15440 -855 15480 -850
rect 15680 -820 15720 -815
rect 15680 -850 15685 -820
rect 15685 -850 15715 -820
rect 15715 -850 15720 -820
rect 15680 -855 15720 -850
rect 15920 -870 15955 -835
rect 16160 -820 16200 -815
rect 16160 -850 16165 -820
rect 16165 -850 16195 -820
rect 16195 -850 16200 -820
rect 16160 -855 16200 -850
rect 16400 -820 16440 -815
rect 16400 -850 16405 -820
rect 16405 -850 16435 -820
rect 16435 -850 16440 -820
rect 16400 -855 16440 -850
rect 16640 -820 16680 -815
rect 16640 -850 16645 -820
rect 16645 -850 16675 -820
rect 16675 -850 16680 -820
rect 16640 -855 16680 -850
rect 16880 -820 16920 -815
rect 16880 -850 16885 -820
rect 16885 -850 16915 -820
rect 16915 -850 16920 -820
rect 16880 -855 16920 -850
rect 17120 -820 17160 -815
rect 17120 -850 17125 -820
rect 17125 -850 17155 -820
rect 17155 -850 17160 -820
rect 17120 -855 17160 -850
rect 17360 -820 17400 -815
rect 17360 -850 17365 -820
rect 17365 -850 17395 -820
rect 17395 -850 17400 -820
rect 17360 -855 17400 -850
rect 17600 -820 17640 -815
rect 17600 -850 17605 -820
rect 17605 -850 17635 -820
rect 17635 -850 17640 -820
rect 17600 -855 17640 -850
rect 17840 -820 17880 -815
rect 17840 -850 17845 -820
rect 17845 -850 17875 -820
rect 17875 -850 17880 -820
rect 17840 -855 17880 -850
rect 18080 -870 18115 -835
rect 18320 -820 18360 -815
rect 18320 -850 18325 -820
rect 18325 -850 18355 -820
rect 18355 -850 18360 -820
rect 18320 -855 18360 -850
rect 18560 -820 18600 -815
rect 18560 -850 18565 -820
rect 18565 -850 18595 -820
rect 18595 -850 18600 -820
rect 18560 -855 18600 -850
rect 18800 -820 18840 -815
rect 18800 -850 18805 -820
rect 18805 -850 18835 -820
rect 18835 -850 18840 -820
rect 18800 -855 18840 -850
rect 19040 -820 19080 -815
rect 19040 -850 19045 -820
rect 19045 -850 19075 -820
rect 19075 -850 19080 -820
rect 19040 -855 19080 -850
rect 19280 -820 19320 -815
rect 19280 -850 19285 -820
rect 19285 -850 19315 -820
rect 19315 -850 19320 -820
rect 19280 -855 19320 -850
rect 19520 -820 19560 -815
rect 19520 -850 19525 -820
rect 19525 -850 19555 -820
rect 19555 -850 19560 -820
rect 19520 -855 19560 -850
rect 19760 -820 19800 -815
rect 19760 -850 19765 -820
rect 19765 -850 19795 -820
rect 19795 -850 19800 -820
rect 19760 -855 19800 -850
rect 20000 -820 20040 -815
rect 20000 -850 20005 -820
rect 20005 -850 20035 -820
rect 20035 -850 20040 -820
rect 20000 -855 20040 -850
rect 20240 -870 20275 -835
rect 20480 -820 20520 -815
rect 20480 -850 20485 -820
rect 20485 -850 20515 -820
rect 20515 -850 20520 -820
rect 20480 -855 20520 -850
rect 20720 -820 20760 -815
rect 20720 -850 20725 -820
rect 20725 -850 20755 -820
rect 20755 -850 20760 -820
rect 20720 -855 20760 -850
rect 20960 -820 21000 -815
rect 20960 -850 20965 -820
rect 20965 -850 20995 -820
rect 20995 -850 21000 -820
rect 20960 -855 21000 -850
rect 21200 -820 21240 -815
rect 21200 -850 21205 -820
rect 21205 -850 21235 -820
rect 21235 -850 21240 -820
rect 21200 -855 21240 -850
rect 21440 -820 21480 -815
rect 21440 -850 21445 -820
rect 21445 -850 21475 -820
rect 21475 -850 21480 -820
rect 21440 -855 21480 -850
rect 21680 -820 21720 -815
rect 21680 -850 21685 -820
rect 21685 -850 21715 -820
rect 21715 -850 21720 -820
rect 21680 -855 21720 -850
rect 21920 -820 21960 -815
rect 21920 -850 21925 -820
rect 21925 -850 21955 -820
rect 21955 -850 21960 -820
rect 21920 -855 21960 -850
rect 22160 -820 22200 -815
rect 22160 -850 22165 -820
rect 22165 -850 22195 -820
rect 22195 -850 22200 -820
rect 22160 -855 22200 -850
rect 22400 -870 22435 -835
rect 22640 -820 22680 -815
rect 22640 -850 22645 -820
rect 22645 -850 22675 -820
rect 22675 -850 22680 -820
rect 22640 -855 22680 -850
rect 22880 -820 22920 -815
rect 22880 -850 22885 -820
rect 22885 -850 22915 -820
rect 22915 -850 22920 -820
rect 22880 -855 22920 -850
rect 23120 -820 23160 -815
rect 23120 -850 23125 -820
rect 23125 -850 23155 -820
rect 23155 -850 23160 -820
rect 23120 -855 23160 -850
rect 23360 -820 23400 -815
rect 23360 -850 23365 -820
rect 23365 -850 23395 -820
rect 23395 -850 23400 -820
rect 23360 -855 23400 -850
rect 23600 -820 23640 -815
rect 23600 -850 23605 -820
rect 23605 -850 23635 -820
rect 23635 -850 23640 -820
rect 23600 -855 23640 -850
rect 23840 -820 23880 -815
rect 23840 -850 23845 -820
rect 23845 -850 23875 -820
rect 23875 -850 23880 -820
rect 23840 -855 23880 -850
rect 24080 -820 24120 -815
rect 24080 -850 24085 -820
rect 24085 -850 24115 -820
rect 24115 -850 24120 -820
rect 24080 -855 24120 -850
rect 24320 -870 24355 -835
rect 24560 -820 24600 -815
rect 24560 -850 24565 -820
rect 24565 -850 24595 -820
rect 24595 -850 24600 -820
rect 24560 -855 24600 -850
rect 24800 -820 24840 -815
rect 24800 -850 24805 -820
rect 24805 -850 24835 -820
rect 24835 -850 24840 -820
rect 24800 -855 24840 -850
rect 25040 -820 25080 -815
rect 25040 -850 25045 -820
rect 25045 -850 25075 -820
rect 25075 -850 25080 -820
rect 25040 -855 25080 -850
rect 25280 -820 25320 -815
rect 25280 -850 25285 -820
rect 25285 -850 25315 -820
rect 25315 -850 25320 -820
rect 25280 -855 25320 -850
rect 25520 -820 25560 -815
rect 25520 -850 25525 -820
rect 25525 -850 25555 -820
rect 25555 -850 25560 -820
rect 25520 -855 25560 -850
rect 25760 -820 25800 -815
rect 25760 -850 25765 -820
rect 25765 -850 25795 -820
rect 25795 -850 25800 -820
rect 25760 -855 25800 -850
rect 26000 -820 26040 -815
rect 26000 -850 26005 -820
rect 26005 -850 26035 -820
rect 26035 -850 26040 -820
rect 26000 -855 26040 -850
rect 26240 -870 26275 -835
rect 26480 -820 26520 -815
rect 26480 -850 26485 -820
rect 26485 -850 26515 -820
rect 26515 -850 26520 -820
rect 26480 -855 26520 -850
rect 26720 -820 26760 -815
rect 26720 -850 26725 -820
rect 26725 -850 26755 -820
rect 26755 -850 26760 -820
rect 26720 -855 26760 -850
rect 26960 -820 27000 -815
rect 26960 -850 26965 -820
rect 26965 -850 26995 -820
rect 26995 -850 27000 -820
rect 26960 -855 27000 -850
rect 27200 -820 27240 -815
rect 27200 -850 27205 -820
rect 27205 -850 27235 -820
rect 27235 -850 27240 -820
rect 27200 -855 27240 -850
rect 27440 -820 27480 -815
rect 27440 -850 27445 -820
rect 27445 -850 27475 -820
rect 27475 -850 27480 -820
rect 27440 -855 27480 -850
rect 27680 -820 27720 -815
rect 27680 -850 27685 -820
rect 27685 -850 27715 -820
rect 27715 -850 27720 -820
rect 27680 -855 27720 -850
rect 27920 -820 27960 -815
rect 27920 -850 27925 -820
rect 27925 -850 27955 -820
rect 27955 -850 27960 -820
rect 27920 -855 27960 -850
rect 28160 -870 28195 -835
rect 28400 -820 28440 -815
rect 28400 -850 28405 -820
rect 28405 -850 28435 -820
rect 28435 -850 28440 -820
rect 28400 -855 28440 -850
rect 28640 -820 28680 -815
rect 28640 -850 28645 -820
rect 28645 -850 28675 -820
rect 28675 -850 28680 -820
rect 28640 -855 28680 -850
rect 28880 -820 28920 -815
rect 28880 -850 28885 -820
rect 28885 -850 28915 -820
rect 28915 -850 28920 -820
rect 28880 -855 28920 -850
rect 29120 -820 29160 -815
rect 29120 -850 29125 -820
rect 29125 -850 29155 -820
rect 29155 -850 29160 -820
rect 29120 -855 29160 -850
rect 29360 -820 29400 -815
rect 29360 -850 29365 -820
rect 29365 -850 29395 -820
rect 29395 -850 29400 -820
rect 29360 -855 29400 -850
rect 29600 -820 29640 -815
rect 29600 -850 29605 -820
rect 29605 -850 29635 -820
rect 29635 -850 29640 -820
rect 29600 -855 29640 -850
rect 29840 -870 29875 -835
rect 30080 -820 30120 -815
rect 30080 -850 30085 -820
rect 30085 -850 30115 -820
rect 30115 -850 30120 -820
rect 30080 -855 30120 -850
rect 30320 -820 30360 -815
rect 30320 -850 30325 -820
rect 30325 -850 30355 -820
rect 30355 -850 30360 -820
rect 30320 -855 30360 -850
rect 30560 -820 30600 -815
rect 30560 -850 30565 -820
rect 30565 -850 30595 -820
rect 30595 -850 30600 -820
rect 30560 -855 30600 -850
<< metal4 >>
rect 2255 305 2310 315
rect 2255 300 2265 305
rect 185 275 240 285
rect 185 270 195 275
rect -145 240 195 270
rect 230 270 240 275
rect 426 270 476 275
rect 731 270 781 275
rect 976 270 1026 275
rect 1216 270 1266 275
rect 1461 270 1511 275
rect 1766 270 1816 275
rect 2011 270 2061 275
rect 2250 270 2265 300
rect 2300 300 2310 305
rect 4195 305 4250 315
rect 4195 300 4205 305
rect 2300 270 2315 300
rect 2496 270 2546 275
rect 2736 270 2786 275
rect 2981 270 3031 275
rect 3221 270 3271 275
rect 3466 270 3516 275
rect 3706 270 3756 275
rect 3951 270 4001 275
rect 4190 270 4205 300
rect 4240 300 4250 305
rect 6445 305 6500 315
rect 6445 300 6455 305
rect 4240 270 4255 300
rect 4436 270 4486 275
rect 4676 270 4726 275
rect 4921 270 4971 275
rect 5161 270 5211 275
rect 5406 270 5456 275
rect 5711 270 5761 275
rect 5956 270 6006 275
rect 6196 270 6246 275
rect 6440 270 6455 300
rect 6490 300 6500 305
rect 9350 305 9405 315
rect 9350 300 9360 305
rect 6490 270 6505 300
rect 6681 270 6731 275
rect 6926 270 6976 275
rect 7166 270 7216 275
rect 7406 270 7456 275
rect 7646 270 7696 275
rect 7891 270 7941 275
rect 8131 270 8181 275
rect 8376 270 8426 275
rect 8616 270 8666 275
rect 8861 270 8911 275
rect 9101 270 9151 275
rect 9345 270 9360 300
rect 9395 300 9405 305
rect 11295 305 11350 315
rect 11295 300 11305 305
rect 9395 270 9410 300
rect 9591 270 9641 275
rect 9836 270 9886 275
rect 10076 270 10126 275
rect 10321 270 10371 275
rect 10561 270 10611 275
rect 10806 270 10856 275
rect 11046 270 11096 275
rect 11290 270 11305 300
rect 11340 300 11350 305
rect 12990 305 13045 315
rect 12990 300 13000 305
rect 11340 270 11355 300
rect 11531 270 11581 275
rect 11776 270 11826 275
rect 12016 270 12066 275
rect 12261 270 12311 275
rect 12501 270 12551 275
rect 12746 270 12796 275
rect 12985 270 13000 300
rect 13035 300 13045 305
rect 15175 305 15230 315
rect 15175 300 15185 305
rect 13035 270 13050 300
rect 13231 270 13281 275
rect 13471 270 13521 275
rect 13716 270 13766 275
rect 13956 270 14006 275
rect 14201 270 14251 275
rect 14441 270 14491 275
rect 14686 270 14736 275
rect 14926 270 14976 275
rect 15170 270 15185 300
rect 15220 300 15230 305
rect 17355 305 17410 315
rect 17355 300 17365 305
rect 15220 270 15235 300
rect 15411 270 15461 275
rect 15656 270 15706 275
rect 15896 270 15946 275
rect 16141 270 16191 275
rect 16381 270 16431 275
rect 16626 270 16676 275
rect 16866 270 16916 275
rect 17111 270 17161 275
rect 17350 270 17365 300
rect 17400 300 17410 305
rect 19540 305 19595 315
rect 19540 300 19550 305
rect 17400 270 17415 300
rect 17596 270 17646 275
rect 17836 270 17886 275
rect 18081 270 18131 275
rect 18321 270 18371 275
rect 18566 270 18616 275
rect 18806 270 18856 275
rect 19051 270 19101 275
rect 19291 270 19341 275
rect 19535 270 19550 300
rect 19585 300 19595 305
rect 20750 305 20805 315
rect 20750 300 20760 305
rect 19585 270 19600 300
rect 19776 270 19826 275
rect 20021 270 20071 275
rect 20261 270 20311 275
rect 20506 270 20556 275
rect 20745 270 20760 300
rect 20795 300 20805 305
rect 20795 270 20810 300
rect 20991 270 21041 275
rect 230 240 431 270
rect -145 -825 -110 240
rect 185 230 240 240
rect 426 230 431 240
rect 471 240 736 270
rect 471 230 476 240
rect 426 225 476 230
rect 731 230 736 240
rect 776 240 981 270
rect 776 230 781 240
rect 731 225 781 230
rect 976 230 981 240
rect 1021 240 1221 270
rect 1021 230 1026 240
rect 976 225 1026 230
rect 1216 230 1221 240
rect 1261 240 1466 270
rect 1261 230 1266 240
rect 1216 225 1266 230
rect 1461 230 1466 240
rect 1506 240 1771 270
rect 1506 230 1511 240
rect 1461 225 1511 230
rect 1766 230 1771 240
rect 1811 240 2016 270
rect 1811 230 1816 240
rect 1766 225 1816 230
rect 2011 230 2016 240
rect 2056 240 2501 270
rect 2056 230 2061 240
rect 2011 225 2061 230
rect 2496 230 2501 240
rect 2541 240 2741 270
rect 2541 230 2546 240
rect 2496 225 2546 230
rect 2736 230 2741 240
rect 2781 240 2986 270
rect 2781 230 2786 240
rect 2736 225 2786 230
rect 2981 230 2986 240
rect 3026 240 3226 270
rect 3026 230 3031 240
rect 2981 225 3031 230
rect 3221 230 3226 240
rect 3266 240 3471 270
rect 3266 230 3271 240
rect 3221 225 3271 230
rect 3466 230 3471 240
rect 3511 240 3711 270
rect 3511 230 3516 240
rect 3466 225 3516 230
rect 3706 230 3711 240
rect 3751 240 3956 270
rect 3751 230 3756 240
rect 3706 225 3756 230
rect 3951 230 3956 240
rect 3996 240 4441 270
rect 3996 230 4001 240
rect 3951 225 4001 230
rect 4436 230 4441 240
rect 4481 240 4681 270
rect 4481 230 4486 240
rect 4436 225 4486 230
rect 4676 230 4681 240
rect 4721 240 4926 270
rect 4721 230 4726 240
rect 4676 225 4726 230
rect 4921 230 4926 240
rect 4966 240 5166 270
rect 4966 230 4971 240
rect 4921 225 4971 230
rect 5161 230 5166 240
rect 5206 240 5411 270
rect 5206 230 5211 240
rect 5161 225 5211 230
rect 5406 230 5411 240
rect 5451 240 5716 270
rect 5451 230 5456 240
rect 5406 225 5456 230
rect 5711 230 5716 240
rect 5756 240 5961 270
rect 5756 230 5761 240
rect 5711 225 5761 230
rect 5956 230 5961 240
rect 6001 240 6201 270
rect 6001 230 6006 240
rect 5956 225 6006 230
rect 6196 230 6201 240
rect 6241 240 6686 270
rect 6241 230 6246 240
rect 6196 225 6246 230
rect 6681 230 6686 240
rect 6726 240 6931 270
rect 6726 230 6731 240
rect 6681 225 6731 230
rect 6926 230 6931 240
rect 6971 240 7171 270
rect 6971 230 6976 240
rect 6926 225 6976 230
rect 7166 230 7171 240
rect 7211 240 7411 270
rect 7211 230 7216 240
rect 7166 225 7216 230
rect 7406 230 7411 240
rect 7451 240 7651 270
rect 7451 230 7456 240
rect 7406 225 7456 230
rect 7646 230 7651 240
rect 7691 240 7896 270
rect 7691 230 7696 240
rect 7646 225 7696 230
rect 7891 230 7896 240
rect 7936 240 8136 270
rect 7936 230 7941 240
rect 7891 225 7941 230
rect 8131 230 8136 240
rect 8176 240 8381 270
rect 8176 230 8181 240
rect 8131 225 8181 230
rect 8376 230 8381 240
rect 8421 240 8621 270
rect 8421 230 8426 240
rect 8376 225 8426 230
rect 8616 230 8621 240
rect 8661 240 8866 270
rect 8661 230 8666 240
rect 8616 225 8666 230
rect 8861 230 8866 240
rect 8906 240 9106 270
rect 8906 230 8911 240
rect 8861 225 8911 230
rect 9101 230 9106 240
rect 9146 240 9596 270
rect 9146 230 9151 240
rect 9101 225 9151 230
rect 9591 230 9596 240
rect 9636 240 9841 270
rect 9636 230 9641 240
rect 9591 225 9641 230
rect 9836 230 9841 240
rect 9881 240 10081 270
rect 9881 230 9886 240
rect 9836 225 9886 230
rect 10076 230 10081 240
rect 10121 240 10326 270
rect 10121 230 10126 240
rect 10076 225 10126 230
rect 10321 230 10326 240
rect 10366 240 10566 270
rect 10366 230 10371 240
rect 10321 225 10371 230
rect 10561 230 10566 240
rect 10606 240 10811 270
rect 10606 230 10611 240
rect 10561 225 10611 230
rect 10806 230 10811 240
rect 10851 240 11051 270
rect 10851 230 10856 240
rect 10806 225 10856 230
rect 11046 230 11051 240
rect 11091 240 11536 270
rect 11091 230 11096 240
rect 11046 225 11096 230
rect 11531 230 11536 240
rect 11576 240 11781 270
rect 11576 230 11581 240
rect 11531 225 11581 230
rect 11776 230 11781 240
rect 11821 240 12021 270
rect 11821 230 11826 240
rect 11776 225 11826 230
rect 12016 230 12021 240
rect 12061 240 12266 270
rect 12061 230 12066 240
rect 12016 225 12066 230
rect 12261 230 12266 240
rect 12306 240 12506 270
rect 12306 230 12311 240
rect 12261 225 12311 230
rect 12501 230 12506 240
rect 12546 240 12751 270
rect 12546 230 12551 240
rect 12501 225 12551 230
rect 12746 230 12751 240
rect 12791 240 13236 270
rect 12791 230 12796 240
rect 12746 225 12796 230
rect 13231 230 13236 240
rect 13276 240 13476 270
rect 13276 230 13281 240
rect 13231 225 13281 230
rect 13471 230 13476 240
rect 13516 240 13721 270
rect 13516 230 13521 240
rect 13471 225 13521 230
rect 13716 230 13721 240
rect 13761 240 13961 270
rect 13761 230 13766 240
rect 13716 225 13766 230
rect 13956 230 13961 240
rect 14001 240 14206 270
rect 14001 230 14006 240
rect 13956 225 14006 230
rect 14201 230 14206 240
rect 14246 240 14446 270
rect 14246 230 14251 240
rect 14201 225 14251 230
rect 14441 230 14446 240
rect 14486 240 14691 270
rect 14486 230 14491 240
rect 14441 225 14491 230
rect 14686 230 14691 240
rect 14731 240 14931 270
rect 14731 230 14736 240
rect 14686 225 14736 230
rect 14926 230 14931 240
rect 14971 240 15416 270
rect 14971 230 14976 240
rect 14926 225 14976 230
rect 15411 230 15416 240
rect 15456 240 15661 270
rect 15456 230 15461 240
rect 15411 225 15461 230
rect 15656 230 15661 240
rect 15701 240 15901 270
rect 15701 230 15706 240
rect 15656 225 15706 230
rect 15896 230 15901 240
rect 15941 240 16146 270
rect 15941 230 15946 240
rect 15896 225 15946 230
rect 16141 230 16146 240
rect 16186 240 16386 270
rect 16186 230 16191 240
rect 16141 225 16191 230
rect 16381 230 16386 240
rect 16426 240 16631 270
rect 16426 230 16431 240
rect 16381 225 16431 230
rect 16626 230 16631 240
rect 16671 240 16871 270
rect 16671 230 16676 240
rect 16626 225 16676 230
rect 16866 230 16871 240
rect 16911 240 17116 270
rect 16911 230 16916 240
rect 16866 225 16916 230
rect 17111 230 17116 240
rect 17156 240 17601 270
rect 17156 230 17161 240
rect 17111 225 17161 230
rect 17596 230 17601 240
rect 17641 240 17841 270
rect 17641 230 17646 240
rect 17596 225 17646 230
rect 17836 230 17841 240
rect 17881 240 18086 270
rect 17881 230 17886 240
rect 17836 225 17886 230
rect 18081 230 18086 240
rect 18126 240 18326 270
rect 18126 230 18131 240
rect 18081 225 18131 230
rect 18321 230 18326 240
rect 18366 240 18571 270
rect 18366 230 18371 240
rect 18321 225 18371 230
rect 18566 230 18571 240
rect 18611 240 18811 270
rect 18611 230 18616 240
rect 18566 225 18616 230
rect 18806 230 18811 240
rect 18851 240 19056 270
rect 18851 230 18856 240
rect 18806 225 18856 230
rect 19051 230 19056 240
rect 19096 240 19296 270
rect 19096 230 19101 240
rect 19051 225 19101 230
rect 19291 230 19296 240
rect 19336 240 19781 270
rect 19336 230 19341 240
rect 19291 225 19341 230
rect 19776 230 19781 240
rect 19821 240 20026 270
rect 19821 230 19826 240
rect 19776 225 19826 230
rect 20021 230 20026 240
rect 20066 240 20266 270
rect 20066 230 20071 240
rect 20021 225 20071 230
rect 20261 230 20266 240
rect 20306 240 20511 270
rect 20306 230 20311 240
rect 20261 225 20311 230
rect 20506 230 20511 240
rect 20551 240 20996 270
rect 20551 230 20556 240
rect 20506 225 20556 230
rect 20991 230 20996 240
rect 21036 240 21156 270
rect 21036 230 21041 240
rect 20991 225 21041 230
rect 176 -160 226 -155
rect 176 -165 181 -160
rect -40 -190 181 -165
rect -40 -240 -25 -190
rect 25 -200 181 -190
rect 221 -165 226 -160
rect 421 -160 471 -155
rect 421 -165 426 -160
rect 221 -200 426 -165
rect 466 -165 471 -160
rect 726 -160 776 -155
rect 726 -165 731 -160
rect 466 -200 731 -165
rect 771 -165 776 -160
rect 971 -160 1021 -155
rect 971 -165 976 -160
rect 771 -200 976 -165
rect 1016 -165 1021 -160
rect 1211 -160 1261 -155
rect 1211 -165 1216 -160
rect 1016 -200 1216 -165
rect 1256 -165 1261 -160
rect 1456 -160 1506 -155
rect 1456 -165 1461 -160
rect 1256 -200 1461 -165
rect 1501 -165 1506 -160
rect 1761 -160 1811 -155
rect 1761 -165 1766 -160
rect 1501 -200 1766 -165
rect 1806 -165 1811 -160
rect 2006 -160 2056 -155
rect 2006 -165 2011 -160
rect 1806 -200 2011 -165
rect 2051 -165 2056 -160
rect 2246 -160 2296 -155
rect 2246 -165 2251 -160
rect 2051 -200 2251 -165
rect 2291 -165 2296 -160
rect 2491 -160 2541 -155
rect 2491 -165 2496 -160
rect 2291 -200 2496 -165
rect 2536 -165 2541 -160
rect 2731 -160 2781 -155
rect 2731 -165 2736 -160
rect 2536 -200 2736 -165
rect 2776 -165 2781 -160
rect 2976 -160 3026 -155
rect 2976 -165 2981 -160
rect 2776 -200 2981 -165
rect 3021 -165 3026 -160
rect 3216 -160 3266 -155
rect 3216 -165 3221 -160
rect 3021 -200 3221 -165
rect 3261 -165 3266 -160
rect 3461 -160 3511 -155
rect 3461 -165 3466 -160
rect 3261 -200 3466 -165
rect 3506 -165 3511 -160
rect 3701 -160 3751 -155
rect 3701 -165 3706 -160
rect 3506 -200 3706 -165
rect 3746 -165 3751 -160
rect 3946 -160 3996 -155
rect 3946 -165 3951 -160
rect 3746 -200 3951 -165
rect 3991 -165 3996 -160
rect 4186 -160 4236 -155
rect 4186 -165 4191 -160
rect 3991 -195 4191 -165
rect 3991 -200 4060 -195
rect 25 -240 1635 -200
rect 1675 -235 4060 -200
rect 4100 -200 4191 -195
rect 4231 -165 4236 -160
rect 4431 -160 4481 -155
rect 4431 -165 4436 -160
rect 4231 -200 4436 -165
rect 4476 -165 4481 -160
rect 4671 -160 4721 -155
rect 4671 -165 4676 -160
rect 4476 -200 4676 -165
rect 4716 -165 4721 -160
rect 4916 -160 4966 -155
rect 4916 -165 4921 -160
rect 4716 -200 4921 -165
rect 4961 -165 4966 -160
rect 5156 -160 5206 -155
rect 5156 -165 5161 -160
rect 4961 -200 5161 -165
rect 5201 -165 5206 -160
rect 5401 -160 5451 -155
rect 5401 -165 5406 -160
rect 5201 -200 5406 -165
rect 5446 -165 5451 -160
rect 5706 -160 5756 -155
rect 5706 -165 5711 -160
rect 5446 -200 5711 -165
rect 5751 -165 5756 -160
rect 5951 -160 6001 -155
rect 5951 -165 5956 -160
rect 5751 -200 5956 -165
rect 5996 -165 6001 -160
rect 6191 -160 6241 -155
rect 6191 -165 6196 -160
rect 5996 -200 6196 -165
rect 6236 -165 6241 -160
rect 6676 -160 6726 -155
rect 6676 -165 6681 -160
rect 6236 -170 6335 -165
rect 6430 -170 6681 -165
rect 6236 -200 6681 -170
rect 6721 -165 6726 -160
rect 6921 -160 6971 -155
rect 6921 -165 6926 -160
rect 6721 -200 6926 -165
rect 6966 -165 6971 -160
rect 7161 -160 7211 -155
rect 7161 -165 7166 -160
rect 6966 -200 7166 -165
rect 7206 -165 7211 -160
rect 7401 -160 7451 -155
rect 7401 -165 7406 -160
rect 7206 -200 7406 -165
rect 7446 -165 7451 -160
rect 7641 -160 7691 -155
rect 7641 -165 7646 -160
rect 7446 -200 7646 -165
rect 7686 -165 7691 -160
rect 8126 -160 8176 -155
rect 8126 -165 8131 -160
rect 7686 -170 7775 -165
rect 7920 -170 8131 -165
rect 7686 -200 8131 -170
rect 8171 -165 8176 -160
rect 8371 -160 8421 -155
rect 8371 -165 8376 -160
rect 8171 -200 8376 -165
rect 8416 -165 8421 -160
rect 8611 -160 8661 -155
rect 8611 -165 8616 -160
rect 8416 -200 8616 -165
rect 8656 -165 8661 -160
rect 8856 -160 8906 -155
rect 8856 -165 8861 -160
rect 8656 -200 8861 -165
rect 8901 -165 8906 -160
rect 9096 -160 9146 -155
rect 9096 -165 9101 -160
rect 8901 -200 9101 -165
rect 9141 -165 9146 -160
rect 9341 -160 9391 -155
rect 9341 -165 9346 -160
rect 9141 -200 9346 -165
rect 9386 -165 9391 -160
rect 9831 -160 9881 -155
rect 9831 -165 9836 -160
rect 9386 -200 9836 -165
rect 9876 -165 9881 -160
rect 10071 -160 10121 -155
rect 10071 -165 10076 -160
rect 9876 -200 10076 -165
rect 10116 -165 10121 -160
rect 10316 -160 10366 -155
rect 10316 -165 10321 -160
rect 10116 -200 10321 -165
rect 10361 -165 10366 -160
rect 10556 -160 10606 -155
rect 10556 -165 10561 -160
rect 10361 -200 10561 -165
rect 10601 -165 10606 -160
rect 10801 -160 10851 -155
rect 10801 -165 10806 -160
rect 10601 -200 10806 -165
rect 10846 -165 10851 -160
rect 11041 -160 11091 -155
rect 11041 -165 11046 -160
rect 10846 -200 11046 -165
rect 11086 -165 11091 -160
rect 11286 -160 11336 -155
rect 11286 -165 11291 -160
rect 11086 -200 11291 -165
rect 11331 -165 11336 -160
rect 11526 -160 11576 -155
rect 11526 -165 11531 -160
rect 11331 -200 11531 -165
rect 11571 -165 11576 -160
rect 11771 -160 11821 -155
rect 11771 -165 11776 -160
rect 11571 -200 11776 -165
rect 11816 -165 11821 -160
rect 12256 -160 12306 -155
rect 12256 -165 12261 -160
rect 11816 -200 12261 -165
rect 12301 -165 12306 -160
rect 12496 -160 12546 -155
rect 12496 -165 12501 -160
rect 12301 -200 12501 -165
rect 12541 -165 12546 -160
rect 12741 -160 12791 -155
rect 12741 -165 12746 -160
rect 12541 -200 12746 -165
rect 12786 -165 12791 -160
rect 12981 -160 13031 -155
rect 12981 -165 12986 -160
rect 12786 -200 12986 -165
rect 13026 -165 13031 -160
rect 13226 -160 13276 -155
rect 13226 -165 13231 -160
rect 13026 -200 13231 -165
rect 13271 -165 13276 -160
rect 13466 -160 13516 -155
rect 13466 -165 13471 -160
rect 13271 -200 13471 -165
rect 13511 -165 13516 -160
rect 13711 -160 13761 -155
rect 13711 -165 13716 -160
rect 13511 -200 13716 -165
rect 13756 -165 13761 -160
rect 14196 -160 14246 -155
rect 14196 -165 14201 -160
rect 13756 -200 14201 -165
rect 14241 -165 14246 -160
rect 14436 -160 14486 -155
rect 14436 -165 14441 -160
rect 14241 -200 14441 -165
rect 14481 -165 14486 -160
rect 14681 -160 14731 -155
rect 14681 -165 14686 -160
rect 14481 -200 14686 -165
rect 14726 -165 14731 -160
rect 14921 -160 14971 -155
rect 14921 -165 14926 -160
rect 14726 -200 14926 -165
rect 14966 -165 14971 -160
rect 15166 -160 15216 -155
rect 15166 -165 15171 -160
rect 14966 -200 15171 -165
rect 15211 -165 15216 -160
rect 15406 -160 15456 -155
rect 15406 -165 15411 -160
rect 15211 -200 15411 -165
rect 15451 -165 15456 -160
rect 15651 -160 15701 -155
rect 15651 -165 15656 -160
rect 15451 -200 15656 -165
rect 15696 -165 15701 -160
rect 16136 -160 16186 -155
rect 16136 -165 16141 -160
rect 15696 -200 16141 -165
rect 16181 -165 16186 -160
rect 16376 -160 16426 -155
rect 16376 -165 16381 -160
rect 16181 -200 16381 -165
rect 16421 -165 16426 -160
rect 16621 -160 16671 -155
rect 16621 -165 16626 -160
rect 16421 -200 16626 -165
rect 16666 -165 16671 -160
rect 16861 -160 16911 -155
rect 16861 -165 16866 -160
rect 16666 -200 16866 -165
rect 16906 -165 16911 -160
rect 17106 -160 17156 -155
rect 17106 -165 17111 -160
rect 16906 -200 17111 -165
rect 17151 -165 17156 -160
rect 17346 -160 17396 -155
rect 17346 -165 17351 -160
rect 17151 -200 17351 -165
rect 17391 -165 17396 -160
rect 17591 -160 17641 -155
rect 17591 -165 17596 -160
rect 17391 -200 17596 -165
rect 17636 -165 17641 -160
rect 17831 -160 17881 -155
rect 17831 -165 17836 -160
rect 17636 -200 17836 -165
rect 17876 -165 17881 -160
rect 18076 -160 18126 -155
rect 18076 -165 18081 -160
rect 17876 -200 18081 -165
rect 18121 -165 18126 -160
rect 18316 -160 18366 -155
rect 18316 -165 18321 -160
rect 18121 -200 18321 -165
rect 18361 -165 18366 -160
rect 18561 -160 18611 -155
rect 18561 -165 18566 -160
rect 18361 -200 18566 -165
rect 18606 -165 18611 -160
rect 18801 -160 18851 -155
rect 18801 -165 18806 -160
rect 18606 -200 18806 -165
rect 18846 -165 18851 -160
rect 19046 -160 19096 -155
rect 19046 -165 19051 -160
rect 18846 -200 19051 -165
rect 19091 -165 19096 -160
rect 19286 -160 19336 -155
rect 19286 -165 19291 -160
rect 19091 -200 19291 -165
rect 19331 -165 19336 -160
rect 19531 -160 19581 -155
rect 19531 -165 19536 -160
rect 19331 -200 19536 -165
rect 19576 -165 19581 -160
rect 19771 -160 19821 -155
rect 19771 -165 19776 -160
rect 19576 -200 19776 -165
rect 19816 -165 19821 -160
rect 20016 -160 20066 -155
rect 20016 -165 20021 -160
rect 19816 -200 20021 -165
rect 20061 -165 20066 -160
rect 20256 -160 20306 -155
rect 20256 -165 20261 -160
rect 20061 -200 20261 -165
rect 20301 -165 20306 -160
rect 20501 -160 20551 -155
rect 20501 -165 20506 -160
rect 20301 -200 20506 -165
rect 20546 -165 20551 -160
rect 20741 -160 20791 -155
rect 20741 -165 20746 -160
rect 20546 -200 20746 -165
rect 20786 -165 20791 -160
rect 20986 -160 21036 -155
rect 20986 -165 20991 -160
rect 20786 -200 20991 -165
rect 21031 -165 21036 -160
rect 21031 -195 21156 -165
rect 21031 -200 21155 -195
rect 4100 -210 21155 -200
rect 4100 -220 9570 -210
rect 4100 -235 6455 -220
rect 1675 -240 6455 -235
rect -40 -280 85 -240
rect 125 -280 325 -240
rect 365 -280 565 -240
rect 605 -280 805 -240
rect 845 -280 1045 -240
rect 1085 -280 1285 -240
rect 1325 -280 1525 -240
rect 1565 -280 1765 -240
rect 1805 -280 2005 -240
rect 2045 -280 2245 -240
rect 2285 -280 2485 -240
rect 2525 -280 2725 -240
rect 2765 -280 2965 -240
rect 3005 -280 3205 -240
rect 3245 -280 3445 -240
rect 3485 -280 3685 -240
rect 3725 -280 3925 -240
rect 3965 -280 4165 -240
rect 4205 -280 4405 -240
rect 4445 -280 4645 -240
rect 4685 -280 4885 -240
rect 4925 -280 5125 -240
rect 5165 -280 5365 -240
rect 5405 -280 5605 -240
rect 5645 -280 5845 -240
rect 5885 -280 6085 -240
rect 6125 -280 6325 -240
rect 6365 -260 6455 -240
rect 6495 -240 7880 -220
rect 6495 -260 6565 -240
rect 6365 -280 6565 -260
rect 6605 -280 6805 -240
rect 6845 -280 7045 -240
rect 7085 -280 7285 -240
rect 7325 -280 7525 -240
rect 7565 -280 7765 -240
rect 7805 -260 7880 -240
rect 7920 -240 9570 -220
rect 7920 -260 8005 -240
rect 7805 -280 8005 -260
rect 8045 -280 8245 -240
rect 8285 -280 8485 -240
rect 8525 -280 8725 -240
rect 8765 -280 8965 -240
rect 9005 -280 9205 -240
rect 9245 -280 9445 -240
rect 9485 -250 9570 -240
rect 9610 -220 17705 -210
rect 9610 -240 11950 -220
rect 9610 -250 9685 -240
rect 9485 -280 9685 -250
rect 9725 -280 9925 -240
rect 9965 -280 10165 -240
rect 10205 -280 10405 -240
rect 10445 -280 10645 -240
rect 10685 -280 10885 -240
rect 10925 -280 11125 -240
rect 11165 -280 11365 -240
rect 11405 -280 11605 -240
rect 11645 -280 11845 -240
rect 11885 -260 11950 -240
rect 11990 -240 13870 -220
rect 11990 -260 12085 -240
rect 11885 -280 12085 -260
rect 12125 -280 12325 -240
rect 12365 -280 12565 -240
rect 12605 -280 12805 -240
rect 12845 -280 13045 -240
rect 13085 -280 13285 -240
rect 13325 -280 13525 -240
rect 13565 -280 13765 -240
rect 13805 -260 13870 -240
rect 13910 -240 15815 -220
rect 13910 -260 14005 -240
rect 13805 -280 14005 -260
rect 14045 -280 14245 -240
rect 14285 -280 14485 -240
rect 14525 -280 14725 -240
rect 14765 -280 14965 -240
rect 15005 -280 15205 -240
rect 15245 -280 15445 -240
rect 15485 -280 15685 -240
rect 15725 -260 15815 -240
rect 15855 -240 17705 -220
rect 15855 -260 15925 -240
rect 15725 -280 15925 -260
rect 15965 -280 16165 -240
rect 16205 -280 16405 -240
rect 16445 -280 16645 -240
rect 16685 -280 16885 -240
rect 16925 -280 17125 -240
rect 17165 -280 17365 -240
rect 17405 -280 17605 -240
rect 17645 -250 17705 -240
rect 17745 -240 19645 -210
rect 17745 -250 17845 -240
rect 17645 -280 17845 -250
rect 17885 -280 18085 -240
rect 18125 -280 18325 -240
rect 18365 -280 18565 -240
rect 18605 -280 18805 -240
rect 18845 -280 19045 -240
rect 19085 -280 19285 -240
rect 19325 -280 19525 -240
rect 19565 -250 19645 -240
rect 19685 -240 21155 -210
rect 21200 -240 21250 -235
rect 21440 -240 21490 -235
rect 21680 -240 21730 -235
rect 21920 -240 21970 -235
rect 22160 -240 22210 -235
rect 22400 -240 22450 -235
rect 22640 -240 22690 -235
rect 22880 -240 22930 -235
rect 23120 -240 23170 -235
rect 23360 -240 23410 -235
rect 23600 -240 23650 -235
rect 23840 -240 23890 -235
rect 24080 -240 24130 -235
rect 24320 -240 24370 -235
rect 24560 -240 24610 -235
rect 24800 -240 24850 -235
rect 25040 -240 25090 -235
rect 25280 -240 25330 -235
rect 25520 -240 25570 -235
rect 25760 -240 25810 -235
rect 26000 -240 26050 -235
rect 26240 -240 26290 -235
rect 26480 -240 26530 -235
rect 26720 -240 26770 -235
rect 26960 -240 27010 -235
rect 27200 -240 27250 -235
rect 27440 -240 27490 -235
rect 27680 -240 27730 -235
rect 27920 -240 27970 -235
rect 28160 -240 28210 -235
rect 28400 -240 28450 -235
rect 28640 -240 28690 -235
rect 28880 -240 28930 -235
rect 29120 -240 29170 -235
rect 29360 -240 29410 -235
rect 29600 -240 29650 -235
rect 29840 -240 29890 -235
rect 30080 -240 30130 -235
rect 30320 -240 30370 -235
rect 30560 -240 30610 -235
rect 19685 -250 19765 -240
rect 19565 -280 19765 -250
rect 19805 -280 20005 -240
rect 20045 -280 20245 -240
rect 20285 -280 20485 -240
rect 20525 -280 20725 -240
rect 20765 -280 20965 -240
rect 21005 -280 21205 -240
rect 21245 -280 21445 -240
rect 21485 -280 21685 -240
rect 21725 -280 21925 -240
rect 21965 -280 22165 -240
rect 22205 -280 22405 -240
rect 22445 -280 22645 -240
rect 22685 -280 22885 -240
rect 22925 -280 23125 -240
rect 23165 -280 23365 -240
rect 23405 -280 23605 -240
rect 23645 -280 23845 -240
rect 23885 -280 24085 -240
rect 24125 -280 24325 -240
rect 24365 -280 24565 -240
rect 24605 -280 24805 -240
rect 24845 -280 25045 -240
rect 25085 -280 25285 -240
rect 25325 -280 25525 -240
rect 25565 -280 25765 -240
rect 25805 -280 26005 -240
rect 26045 -280 26245 -240
rect 26285 -280 26485 -240
rect 26525 -280 26725 -240
rect 26765 -280 26965 -240
rect 27005 -280 27205 -240
rect 27245 -280 27445 -240
rect 27485 -280 27685 -240
rect 27725 -280 27925 -240
rect 27965 -280 28165 -240
rect 28205 -280 28405 -240
rect 28445 -280 28645 -240
rect 28685 -280 28885 -240
rect 28925 -280 29125 -240
rect 29165 -280 29365 -240
rect 29405 -280 29605 -240
rect 29645 -280 29845 -240
rect 29885 -280 30085 -240
rect 30125 -280 30325 -240
rect 30365 -280 30565 -240
rect 30605 -280 30720 -240
rect 80 -285 130 -280
rect 320 -285 370 -280
rect 560 -285 610 -280
rect 800 -285 850 -280
rect 1040 -285 1090 -280
rect 1280 -285 1330 -280
rect 1520 -285 1570 -280
rect 1760 -285 1810 -280
rect 2000 -285 2050 -280
rect 2240 -285 2290 -280
rect 2480 -285 2530 -280
rect 2720 -285 2770 -280
rect 2960 -285 3010 -280
rect 3200 -285 3250 -280
rect 3440 -285 3490 -280
rect 3680 -285 3730 -280
rect 3920 -285 3970 -280
rect 4160 -285 4210 -280
rect 4400 -285 4450 -280
rect 4640 -285 4690 -280
rect 4880 -285 4930 -280
rect 5120 -285 5170 -280
rect 5360 -285 5410 -280
rect 5600 -285 5650 -280
rect 5840 -285 5890 -280
rect 6080 -285 6130 -280
rect 6320 -285 6370 -280
rect 6560 -285 6610 -280
rect 6800 -285 6850 -280
rect 7040 -285 7090 -280
rect 7280 -285 7330 -280
rect 7520 -285 7570 -280
rect 7760 -285 7810 -280
rect 8000 -285 8050 -280
rect 8240 -285 8290 -280
rect 8480 -285 8530 -280
rect 8720 -285 8770 -280
rect 8960 -285 9010 -280
rect 9200 -285 9250 -280
rect 9440 -285 9490 -280
rect 9680 -285 9730 -280
rect 9920 -285 9970 -280
rect 10160 -285 10210 -280
rect 10400 -285 10450 -280
rect 10640 -285 10690 -280
rect 10880 -285 10930 -280
rect 11120 -285 11170 -280
rect 11360 -285 11410 -280
rect 11600 -285 11650 -280
rect 11840 -285 11890 -280
rect 12080 -285 12130 -280
rect 12320 -285 12370 -280
rect 12560 -285 12610 -280
rect 12800 -285 12850 -280
rect 13040 -285 13090 -280
rect 13280 -285 13330 -280
rect 13520 -285 13570 -280
rect 13760 -285 13810 -280
rect 14000 -285 14050 -280
rect 14240 -285 14290 -280
rect 14480 -285 14530 -280
rect 14720 -285 14770 -280
rect 14960 -285 15010 -280
rect 15200 -285 15250 -280
rect 15440 -285 15490 -280
rect 15680 -285 15730 -280
rect 15920 -285 15970 -280
rect 16160 -285 16210 -280
rect 16400 -285 16450 -280
rect 16640 -285 16690 -280
rect 16880 -285 16930 -280
rect 17120 -285 17170 -280
rect 17360 -285 17410 -280
rect 17600 -285 17650 -280
rect 17840 -285 17890 -280
rect 18080 -285 18130 -280
rect 18320 -285 18370 -280
rect 18560 -285 18610 -280
rect 18800 -285 18850 -280
rect 19040 -285 19090 -280
rect 19280 -285 19330 -280
rect 19520 -285 19570 -280
rect 19760 -285 19810 -280
rect 20000 -285 20050 -280
rect 20240 -285 20290 -280
rect 20480 -285 20530 -280
rect 20720 -285 20770 -280
rect 20960 -285 21010 -280
rect 21200 -285 21250 -280
rect 21440 -285 21490 -280
rect 21680 -285 21730 -280
rect 21920 -285 21970 -280
rect 22160 -285 22210 -280
rect 22400 -285 22450 -280
rect 22640 -285 22690 -280
rect 22880 -285 22930 -280
rect 23120 -285 23170 -280
rect 23360 -285 23410 -280
rect 23600 -285 23650 -280
rect 23840 -285 23890 -280
rect 24080 -285 24130 -280
rect 24320 -285 24370 -280
rect 24560 -285 24610 -280
rect 24800 -285 24850 -280
rect 25040 -285 25090 -280
rect 25280 -285 25330 -280
rect 25520 -285 25570 -280
rect 25760 -285 25810 -280
rect 26000 -285 26050 -280
rect 26240 -285 26290 -280
rect 26480 -285 26530 -280
rect 26720 -285 26770 -280
rect 26960 -285 27010 -280
rect 27200 -285 27250 -280
rect 27440 -285 27490 -280
rect 27680 -285 27730 -280
rect 27920 -285 27970 -280
rect 28160 -285 28210 -280
rect 28400 -285 28450 -280
rect 28640 -285 28690 -280
rect 28880 -285 28930 -280
rect 29120 -285 29170 -280
rect 29360 -285 29410 -280
rect 29600 -285 29650 -280
rect 29840 -285 29890 -280
rect 30080 -285 30130 -280
rect 30320 -285 30370 -280
rect 30560 -285 30610 -280
rect 75 -815 125 -810
rect 75 -825 80 -815
rect -145 -855 80 -825
rect 120 -825 125 -815
rect 315 -815 365 -810
rect 315 -825 320 -815
rect 120 -855 320 -825
rect 360 -825 365 -815
rect 555 -815 605 -810
rect 555 -825 560 -815
rect 360 -855 560 -825
rect 600 -825 605 -815
rect 1035 -815 1085 -810
rect 785 -825 850 -820
rect 1035 -825 1040 -815
rect 600 -835 1040 -825
rect 600 -855 800 -835
rect 75 -860 125 -855
rect 315 -860 365 -855
rect 555 -860 605 -855
rect 785 -870 800 -855
rect 835 -855 1040 -835
rect 1080 -825 1085 -815
rect 1275 -815 1325 -810
rect 1275 -825 1280 -815
rect 1080 -855 1280 -825
rect 1320 -825 1325 -815
rect 1515 -815 1565 -810
rect 1515 -825 1520 -815
rect 1320 -855 1520 -825
rect 1560 -825 1565 -815
rect 1755 -815 1805 -810
rect 1755 -825 1760 -815
rect 1560 -855 1760 -825
rect 1800 -825 1805 -815
rect 1995 -815 2045 -810
rect 1995 -825 2000 -815
rect 1800 -855 2000 -825
rect 2040 -825 2045 -815
rect 2235 -815 2285 -810
rect 2235 -825 2240 -815
rect 2040 -855 2240 -825
rect 2280 -825 2285 -815
rect 2475 -815 2525 -810
rect 2475 -825 2480 -815
rect 2280 -855 2480 -825
rect 2520 -825 2525 -815
rect 2715 -815 2765 -810
rect 2715 -825 2720 -815
rect 2520 -855 2720 -825
rect 2760 -825 2765 -815
rect 3195 -815 3245 -810
rect 2945 -825 3010 -820
rect 3195 -825 3200 -815
rect 2760 -835 3200 -825
rect 2760 -855 2960 -835
rect 835 -870 850 -855
rect 1035 -860 1085 -855
rect 1275 -860 1325 -855
rect 1515 -860 1565 -855
rect 1755 -860 1805 -855
rect 1995 -860 2045 -855
rect 2235 -860 2285 -855
rect 2475 -860 2525 -855
rect 2715 -860 2765 -855
rect 785 -885 850 -870
rect 2945 -870 2960 -855
rect 2995 -855 3200 -835
rect 3240 -825 3245 -815
rect 3435 -815 3485 -810
rect 3435 -825 3440 -815
rect 3240 -855 3440 -825
rect 3480 -825 3485 -815
rect 3675 -815 3725 -810
rect 3675 -825 3680 -815
rect 3480 -855 3680 -825
rect 3720 -825 3725 -815
rect 3915 -815 3965 -810
rect 3915 -825 3920 -815
rect 3720 -855 3920 -825
rect 3960 -825 3965 -815
rect 4155 -815 4205 -810
rect 4155 -825 4160 -815
rect 3960 -855 4160 -825
rect 4200 -825 4205 -815
rect 4395 -815 4445 -810
rect 4395 -825 4400 -815
rect 4200 -855 4400 -825
rect 4440 -825 4445 -815
rect 4635 -815 4685 -810
rect 4635 -825 4640 -815
rect 4440 -855 4640 -825
rect 4680 -825 4685 -815
rect 4875 -815 4925 -810
rect 4875 -825 4880 -815
rect 4680 -855 4880 -825
rect 4920 -825 4925 -815
rect 5355 -815 5405 -810
rect 5105 -825 5170 -820
rect 5355 -825 5360 -815
rect 4920 -835 5360 -825
rect 4920 -855 5120 -835
rect 2995 -870 3010 -855
rect 3195 -860 3245 -855
rect 3435 -860 3485 -855
rect 3675 -860 3725 -855
rect 3915 -860 3965 -855
rect 4155 -860 4205 -855
rect 4395 -860 4445 -855
rect 4635 -860 4685 -855
rect 4875 -860 4925 -855
rect 2945 -885 3010 -870
rect 5105 -870 5120 -855
rect 5155 -855 5360 -835
rect 5400 -825 5405 -815
rect 5595 -815 5645 -810
rect 5595 -825 5600 -815
rect 5400 -855 5600 -825
rect 5640 -825 5645 -815
rect 5835 -815 5885 -810
rect 5835 -825 5840 -815
rect 5640 -855 5840 -825
rect 5880 -825 5885 -815
rect 6075 -815 6125 -810
rect 6075 -825 6080 -815
rect 5880 -855 6080 -825
rect 6120 -825 6125 -815
rect 6315 -815 6365 -810
rect 6315 -825 6320 -815
rect 6120 -855 6320 -825
rect 6360 -825 6365 -815
rect 6555 -815 6605 -810
rect 6555 -825 6560 -815
rect 6360 -855 6560 -825
rect 6600 -825 6605 -815
rect 6795 -815 6845 -810
rect 6795 -825 6800 -815
rect 6600 -855 6800 -825
rect 6840 -825 6845 -815
rect 7035 -815 7085 -810
rect 7035 -825 7040 -815
rect 6840 -855 7040 -825
rect 7080 -825 7085 -815
rect 7515 -815 7565 -810
rect 7265 -825 7330 -820
rect 7515 -825 7520 -815
rect 7080 -835 7520 -825
rect 7080 -855 7280 -835
rect 5155 -870 5170 -855
rect 5355 -860 5405 -855
rect 5595 -860 5645 -855
rect 5835 -860 5885 -855
rect 6075 -860 6125 -855
rect 6315 -860 6365 -855
rect 6555 -860 6605 -855
rect 6795 -860 6845 -855
rect 7035 -860 7085 -855
rect 5105 -885 5170 -870
rect 7265 -870 7280 -855
rect 7315 -855 7520 -835
rect 7560 -825 7565 -815
rect 7755 -815 7805 -810
rect 7755 -825 7760 -815
rect 7560 -855 7760 -825
rect 7800 -825 7805 -815
rect 7995 -815 8045 -810
rect 7995 -825 8000 -815
rect 7800 -855 8000 -825
rect 8040 -825 8045 -815
rect 8235 -815 8285 -810
rect 8235 -825 8240 -815
rect 8040 -855 8240 -825
rect 8280 -825 8285 -815
rect 8475 -815 8525 -810
rect 8475 -825 8480 -815
rect 8280 -855 8480 -825
rect 8520 -825 8525 -815
rect 8715 -815 8765 -810
rect 8715 -825 8720 -815
rect 8520 -855 8720 -825
rect 8760 -825 8765 -815
rect 8955 -815 9005 -810
rect 8955 -825 8960 -815
rect 8760 -855 8960 -825
rect 9000 -825 9005 -815
rect 9195 -815 9245 -810
rect 9195 -825 9200 -815
rect 9000 -855 9200 -825
rect 9240 -825 9245 -815
rect 9675 -815 9725 -810
rect 9425 -825 9490 -820
rect 9675 -825 9680 -815
rect 9240 -835 9680 -825
rect 9240 -855 9440 -835
rect 7315 -870 7330 -855
rect 7515 -860 7565 -855
rect 7755 -860 7805 -855
rect 7995 -860 8045 -855
rect 8235 -860 8285 -855
rect 8475 -860 8525 -855
rect 8715 -860 8765 -855
rect 8955 -860 9005 -855
rect 9195 -860 9245 -855
rect 7265 -885 7330 -870
rect 9425 -870 9440 -855
rect 9475 -855 9680 -835
rect 9720 -825 9725 -815
rect 9915 -815 9965 -810
rect 9915 -825 9920 -815
rect 9720 -855 9920 -825
rect 9960 -825 9965 -815
rect 10155 -815 10205 -810
rect 10155 -825 10160 -815
rect 9960 -855 10160 -825
rect 10200 -825 10205 -815
rect 10395 -815 10445 -810
rect 10395 -825 10400 -815
rect 10200 -855 10400 -825
rect 10440 -825 10445 -815
rect 10635 -815 10685 -810
rect 10635 -825 10640 -815
rect 10440 -855 10640 -825
rect 10680 -825 10685 -815
rect 10875 -815 10925 -810
rect 10875 -825 10880 -815
rect 10680 -855 10880 -825
rect 10920 -825 10925 -815
rect 11115 -815 11165 -810
rect 11115 -825 11120 -815
rect 10920 -855 11120 -825
rect 11160 -825 11165 -815
rect 11355 -815 11405 -810
rect 11355 -825 11360 -815
rect 11160 -855 11360 -825
rect 11400 -825 11405 -815
rect 11835 -815 11885 -810
rect 11585 -825 11650 -820
rect 11835 -825 11840 -815
rect 11400 -835 11840 -825
rect 11400 -855 11600 -835
rect 9475 -870 9490 -855
rect 9675 -860 9725 -855
rect 9915 -860 9965 -855
rect 10155 -860 10205 -855
rect 10395 -860 10445 -855
rect 10635 -860 10685 -855
rect 10875 -860 10925 -855
rect 11115 -860 11165 -855
rect 11355 -860 11405 -855
rect 9425 -885 9490 -870
rect 11585 -870 11600 -855
rect 11635 -855 11840 -835
rect 11880 -825 11885 -815
rect 12075 -815 12125 -810
rect 12075 -825 12080 -815
rect 11880 -855 12080 -825
rect 12120 -825 12125 -815
rect 12315 -815 12365 -810
rect 12315 -825 12320 -815
rect 12120 -855 12320 -825
rect 12360 -825 12365 -815
rect 12555 -815 12605 -810
rect 12555 -825 12560 -815
rect 12360 -855 12560 -825
rect 12600 -825 12605 -815
rect 12795 -815 12845 -810
rect 12795 -825 12800 -815
rect 12600 -855 12800 -825
rect 12840 -825 12845 -815
rect 13035 -815 13085 -810
rect 13035 -825 13040 -815
rect 12840 -855 13040 -825
rect 13080 -825 13085 -815
rect 13275 -815 13325 -810
rect 13275 -825 13280 -815
rect 13080 -855 13280 -825
rect 13320 -825 13325 -815
rect 13515 -815 13565 -810
rect 13515 -825 13520 -815
rect 13320 -855 13520 -825
rect 13560 -825 13565 -815
rect 13995 -815 14045 -810
rect 13745 -825 13810 -820
rect 13995 -825 14000 -815
rect 13560 -835 14000 -825
rect 13560 -855 13760 -835
rect 11635 -870 11650 -855
rect 11835 -860 11885 -855
rect 12075 -860 12125 -855
rect 12315 -860 12365 -855
rect 12555 -860 12605 -855
rect 12795 -860 12845 -855
rect 13035 -860 13085 -855
rect 13275 -860 13325 -855
rect 13515 -860 13565 -855
rect 11585 -885 11650 -870
rect 13745 -870 13760 -855
rect 13795 -855 14000 -835
rect 14040 -825 14045 -815
rect 14235 -815 14285 -810
rect 14235 -825 14240 -815
rect 14040 -855 14240 -825
rect 14280 -825 14285 -815
rect 14475 -815 14525 -810
rect 14475 -825 14480 -815
rect 14280 -855 14480 -825
rect 14520 -825 14525 -815
rect 14715 -815 14765 -810
rect 14715 -825 14720 -815
rect 14520 -855 14720 -825
rect 14760 -825 14765 -815
rect 14955 -815 15005 -810
rect 14955 -825 14960 -815
rect 14760 -855 14960 -825
rect 15000 -825 15005 -815
rect 15195 -815 15245 -810
rect 15195 -825 15200 -815
rect 15000 -855 15200 -825
rect 15240 -825 15245 -815
rect 15435 -815 15485 -810
rect 15435 -825 15440 -815
rect 15240 -855 15440 -825
rect 15480 -825 15485 -815
rect 15675 -815 15725 -810
rect 15675 -825 15680 -815
rect 15480 -855 15680 -825
rect 15720 -825 15725 -815
rect 16155 -815 16205 -810
rect 15905 -825 15970 -820
rect 16155 -825 16160 -815
rect 15720 -835 16160 -825
rect 15720 -855 15920 -835
rect 13795 -870 13810 -855
rect 13995 -860 14045 -855
rect 14235 -860 14285 -855
rect 14475 -860 14525 -855
rect 14715 -860 14765 -855
rect 14955 -860 15005 -855
rect 15195 -860 15245 -855
rect 15435 -860 15485 -855
rect 15675 -860 15725 -855
rect 13745 -885 13810 -870
rect 15905 -870 15920 -855
rect 15955 -855 16160 -835
rect 16200 -825 16205 -815
rect 16395 -815 16445 -810
rect 16395 -825 16400 -815
rect 16200 -855 16400 -825
rect 16440 -825 16445 -815
rect 16635 -815 16685 -810
rect 16635 -825 16640 -815
rect 16440 -855 16640 -825
rect 16680 -825 16685 -815
rect 16875 -815 16925 -810
rect 16875 -825 16880 -815
rect 16680 -855 16880 -825
rect 16920 -825 16925 -815
rect 17115 -815 17165 -810
rect 17115 -825 17120 -815
rect 16920 -855 17120 -825
rect 17160 -825 17165 -815
rect 17355 -815 17405 -810
rect 17355 -825 17360 -815
rect 17160 -855 17360 -825
rect 17400 -825 17405 -815
rect 17595 -815 17645 -810
rect 17595 -825 17600 -815
rect 17400 -855 17600 -825
rect 17640 -825 17645 -815
rect 17835 -815 17885 -810
rect 17835 -825 17840 -815
rect 17640 -855 17840 -825
rect 17880 -825 17885 -815
rect 18315 -815 18365 -810
rect 18065 -825 18130 -820
rect 18315 -825 18320 -815
rect 17880 -835 18320 -825
rect 17880 -855 18080 -835
rect 15955 -870 15970 -855
rect 16155 -860 16205 -855
rect 16395 -860 16445 -855
rect 16635 -860 16685 -855
rect 16875 -860 16925 -855
rect 17115 -860 17165 -855
rect 17355 -860 17405 -855
rect 17595 -860 17645 -855
rect 17835 -860 17885 -855
rect 15905 -885 15970 -870
rect 18065 -870 18080 -855
rect 18115 -855 18320 -835
rect 18360 -825 18365 -815
rect 18555 -815 18605 -810
rect 18555 -825 18560 -815
rect 18360 -855 18560 -825
rect 18600 -825 18605 -815
rect 18795 -815 18845 -810
rect 18795 -825 18800 -815
rect 18600 -855 18800 -825
rect 18840 -825 18845 -815
rect 19035 -815 19085 -810
rect 19035 -825 19040 -815
rect 18840 -855 19040 -825
rect 19080 -825 19085 -815
rect 19275 -815 19325 -810
rect 19275 -825 19280 -815
rect 19080 -855 19280 -825
rect 19320 -825 19325 -815
rect 19515 -815 19565 -810
rect 19515 -825 19520 -815
rect 19320 -855 19520 -825
rect 19560 -825 19565 -815
rect 19755 -815 19805 -810
rect 19755 -825 19760 -815
rect 19560 -855 19760 -825
rect 19800 -825 19805 -815
rect 19995 -815 20045 -810
rect 19995 -825 20000 -815
rect 19800 -855 20000 -825
rect 20040 -825 20045 -815
rect 20475 -815 20525 -810
rect 20225 -825 20290 -820
rect 20475 -825 20480 -815
rect 20040 -835 20480 -825
rect 20040 -855 20240 -835
rect 18115 -870 18130 -855
rect 18315 -860 18365 -855
rect 18555 -860 18605 -855
rect 18795 -860 18845 -855
rect 19035 -860 19085 -855
rect 19275 -860 19325 -855
rect 19515 -860 19565 -855
rect 19755 -860 19805 -855
rect 19995 -860 20045 -855
rect 18065 -885 18130 -870
rect 20225 -870 20240 -855
rect 20275 -855 20480 -835
rect 20520 -825 20525 -815
rect 20715 -815 20765 -810
rect 20715 -825 20720 -815
rect 20520 -855 20720 -825
rect 20760 -825 20765 -815
rect 20955 -815 21005 -810
rect 20955 -825 20960 -815
rect 20760 -855 20960 -825
rect 21000 -825 21005 -815
rect 21195 -815 21245 -810
rect 21195 -825 21200 -815
rect 21000 -855 21200 -825
rect 21240 -825 21245 -815
rect 21435 -815 21485 -810
rect 21435 -825 21440 -815
rect 21240 -855 21440 -825
rect 21480 -825 21485 -815
rect 21675 -815 21725 -810
rect 21675 -825 21680 -815
rect 21480 -855 21680 -825
rect 21720 -825 21725 -815
rect 21915 -815 21965 -810
rect 21915 -825 21920 -815
rect 21720 -855 21920 -825
rect 21960 -825 21965 -815
rect 22155 -815 22205 -810
rect 22155 -825 22160 -815
rect 21960 -855 22160 -825
rect 22200 -825 22205 -815
rect 22635 -815 22685 -810
rect 22385 -825 22450 -820
rect 22635 -825 22640 -815
rect 22200 -835 22640 -825
rect 22200 -855 22400 -835
rect 20275 -870 20290 -855
rect 20475 -860 20525 -855
rect 20715 -860 20765 -855
rect 20955 -860 21005 -855
rect 21195 -860 21245 -855
rect 21435 -860 21485 -855
rect 21675 -860 21725 -855
rect 21915 -860 21965 -855
rect 22155 -860 22205 -855
rect 20225 -885 20290 -870
rect 22385 -870 22400 -855
rect 22435 -855 22640 -835
rect 22680 -825 22685 -815
rect 22875 -815 22925 -810
rect 22875 -825 22880 -815
rect 22680 -855 22880 -825
rect 22920 -825 22925 -815
rect 23115 -815 23165 -810
rect 23115 -825 23120 -815
rect 22920 -855 23120 -825
rect 23160 -825 23165 -815
rect 23355 -815 23405 -810
rect 23355 -825 23360 -815
rect 23160 -855 23360 -825
rect 23400 -825 23405 -815
rect 23595 -815 23645 -810
rect 23595 -825 23600 -815
rect 23400 -855 23600 -825
rect 23640 -825 23645 -815
rect 23835 -815 23885 -810
rect 23835 -825 23840 -815
rect 23640 -855 23840 -825
rect 23880 -825 23885 -815
rect 24075 -815 24125 -810
rect 24075 -825 24080 -815
rect 23880 -855 24080 -825
rect 24120 -825 24125 -815
rect 24555 -815 24605 -810
rect 24305 -825 24370 -820
rect 24555 -825 24560 -815
rect 24120 -835 24560 -825
rect 24120 -855 24320 -835
rect 22435 -870 22450 -855
rect 22635 -860 22685 -855
rect 22875 -860 22925 -855
rect 23115 -860 23165 -855
rect 23355 -860 23405 -855
rect 23595 -860 23645 -855
rect 23835 -860 23885 -855
rect 24075 -860 24125 -855
rect 22385 -885 22450 -870
rect 24305 -870 24320 -855
rect 24355 -855 24560 -835
rect 24600 -825 24605 -815
rect 24795 -815 24845 -810
rect 24795 -825 24800 -815
rect 24600 -855 24800 -825
rect 24840 -825 24845 -815
rect 25035 -815 25085 -810
rect 25035 -825 25040 -815
rect 24840 -855 25040 -825
rect 25080 -825 25085 -815
rect 25275 -815 25325 -810
rect 25275 -825 25280 -815
rect 25080 -855 25280 -825
rect 25320 -825 25325 -815
rect 25515 -815 25565 -810
rect 25515 -825 25520 -815
rect 25320 -855 25520 -825
rect 25560 -825 25565 -815
rect 25755 -815 25805 -810
rect 25755 -825 25760 -815
rect 25560 -855 25760 -825
rect 25800 -825 25805 -815
rect 25995 -815 26045 -810
rect 25995 -825 26000 -815
rect 25800 -855 26000 -825
rect 26040 -825 26045 -815
rect 26475 -815 26525 -810
rect 26225 -825 26290 -820
rect 26475 -825 26480 -815
rect 26040 -835 26480 -825
rect 26040 -855 26240 -835
rect 24355 -870 24370 -855
rect 24555 -860 24605 -855
rect 24795 -860 24845 -855
rect 25035 -860 25085 -855
rect 25275 -860 25325 -855
rect 25515 -860 25565 -855
rect 25755 -860 25805 -855
rect 25995 -860 26045 -855
rect 24305 -885 24370 -870
rect 26225 -870 26240 -855
rect 26275 -855 26480 -835
rect 26520 -825 26525 -815
rect 26715 -815 26765 -810
rect 26715 -825 26720 -815
rect 26520 -855 26720 -825
rect 26760 -825 26765 -815
rect 26955 -815 27005 -810
rect 26955 -825 26960 -815
rect 26760 -855 26960 -825
rect 27000 -825 27005 -815
rect 27195 -815 27245 -810
rect 27195 -825 27200 -815
rect 27000 -855 27200 -825
rect 27240 -825 27245 -815
rect 27435 -815 27485 -810
rect 27435 -825 27440 -815
rect 27240 -855 27440 -825
rect 27480 -825 27485 -815
rect 27675 -815 27725 -810
rect 27675 -825 27680 -815
rect 27480 -855 27680 -825
rect 27720 -825 27725 -815
rect 27915 -815 27965 -810
rect 27915 -825 27920 -815
rect 27720 -855 27920 -825
rect 27960 -825 27965 -815
rect 28395 -815 28445 -810
rect 28145 -825 28210 -820
rect 28395 -825 28400 -815
rect 27960 -835 28400 -825
rect 27960 -855 28160 -835
rect 26275 -870 26290 -855
rect 26475 -860 26525 -855
rect 26715 -860 26765 -855
rect 26955 -860 27005 -855
rect 27195 -860 27245 -855
rect 27435 -860 27485 -855
rect 27675 -860 27725 -855
rect 27915 -860 27965 -855
rect 26225 -885 26290 -870
rect 28145 -870 28160 -855
rect 28195 -855 28400 -835
rect 28440 -825 28445 -815
rect 28635 -815 28685 -810
rect 28635 -825 28640 -815
rect 28440 -855 28640 -825
rect 28680 -825 28685 -815
rect 28875 -815 28925 -810
rect 28875 -825 28880 -815
rect 28680 -855 28880 -825
rect 28920 -825 28925 -815
rect 29115 -815 29165 -810
rect 29115 -825 29120 -815
rect 28920 -855 29120 -825
rect 29160 -825 29165 -815
rect 29355 -815 29405 -810
rect 29355 -825 29360 -815
rect 29160 -855 29360 -825
rect 29400 -825 29405 -815
rect 29595 -815 29645 -810
rect 29595 -825 29600 -815
rect 29400 -855 29600 -825
rect 29640 -825 29645 -815
rect 30075 -815 30125 -810
rect 29825 -825 29890 -820
rect 30075 -825 30080 -815
rect 29640 -835 30080 -825
rect 29640 -855 29840 -835
rect 28195 -870 28210 -855
rect 28395 -860 28445 -855
rect 28635 -860 28685 -855
rect 28875 -860 28925 -855
rect 29115 -860 29165 -855
rect 29355 -860 29405 -855
rect 29595 -860 29645 -855
rect 28145 -885 28210 -870
rect 29825 -870 29840 -855
rect 29875 -855 30080 -835
rect 30120 -825 30125 -815
rect 30315 -815 30365 -810
rect 30315 -825 30320 -815
rect 30120 -855 30320 -825
rect 30360 -825 30365 -815
rect 30555 -815 30605 -810
rect 30555 -825 30560 -815
rect 30360 -855 30560 -825
rect 30600 -825 30605 -815
rect 30600 -855 30725 -825
rect 29875 -870 29890 -855
rect 30075 -860 30125 -855
rect 30315 -860 30365 -855
rect 30555 -860 30605 -855
rect 29825 -885 29890 -870
<< labels >>
rlabel space -45 -280 80 -165 1 GND
rlabel nwell 185 240 510 270 1 VDD
rlabel metal4 -45 240 90 270 1 VDD
rlabel locali -55 -5 45 15 1 IN
rlabel locali -105 -515 -55 -495 1 OUT
rlabel locali 145 -5 230 15 1 IN
rlabel space 255 -5 355 15 1 OUT1
rlabel locali 560 -5 660 15 1 OUT2
rlabel locali 1590 -5 1690 15 1 OUT3
rlabel locali 5535 -5 5635 15 1 OUT4
rlabel locali 21120 -10 21180 10 1 OUT5
rlabel locali 30685 -505 30760 -485 1 OUT5
rlabel metal4 21155 -280 30720 -240 1 GND
rlabel metal4 -145 -825 -110 270 1 VDD
rlabel metal4 -110 240 21155 270 1 VDD
rlabel metal4 -145 -855 30725 -825 1 VDD
rlabel space -40 -280 21155 -165 1 GND
<< end >>
