magic
tech sky130A
timestamp 1643048518
<< nwell >>
rect 2885 1480 3070 1620
rect 3370 1480 4310 1620
rect -70 760 290 1460
rect 1395 1260 1995 1480
rect 1390 990 1995 1260
rect 2415 990 4310 1480
rect 1390 960 4310 990
rect 1549 941 1642 960
rect 1800 460 1990 960
rect 2730 460 2780 960
rect 3370 955 4310 960
rect 3520 460 3570 955
rect 3650 934 3711 955
<< psubdiff >>
rect -205 2115 -75 2130
rect -205 2015 -190 2115
rect -90 2015 -75 2115
rect -205 2000 -75 2015
rect 370 2115 500 2130
rect 370 2015 385 2115
rect 485 2015 500 2115
rect 370 2000 500 2015
rect 945 2115 1075 2130
rect 945 2015 960 2115
rect 1060 2015 1075 2115
rect 945 2000 1075 2015
rect 1520 2115 1650 2130
rect 1520 2015 1535 2115
rect 1635 2015 1650 2115
rect 1520 2000 1650 2015
rect 2095 2115 2225 2130
rect 2095 2015 2110 2115
rect 2210 2015 2225 2115
rect 2095 2000 2225 2015
rect 2670 2115 2800 2130
rect 2670 2015 2685 2115
rect 2785 2015 2800 2115
rect 2670 2000 2800 2015
rect 3245 2115 3375 2130
rect 3245 2015 3260 2115
rect 3360 2015 3375 2115
rect 3245 2000 3375 2015
rect 3820 2115 3950 2130
rect 3820 2015 3835 2115
rect 3935 2015 3950 2115
rect 3820 2000 3950 2015
rect 4395 2115 4525 2130
rect 4395 2015 4410 2115
rect 4510 2015 4525 2115
rect 4395 2000 4525 2015
rect -470 1830 -340 1845
rect -470 1730 -455 1830
rect -355 1730 -340 1830
rect -470 1715 -340 1730
rect 4540 1830 4670 1845
rect 4540 1730 4555 1830
rect 4655 1730 4670 1830
rect 4540 1715 4670 1730
rect -470 1255 -340 1270
rect -470 1155 -455 1255
rect -355 1155 -340 1255
rect -470 1140 -340 1155
rect 4540 1255 4670 1270
rect 4540 1155 4555 1255
rect 4655 1155 4670 1255
rect 4540 1140 4670 1155
rect -470 680 -340 695
rect -470 580 -455 680
rect -355 580 -340 680
rect -470 565 -340 580
rect 4540 680 4670 695
rect 4540 580 4555 680
rect 4655 580 4670 680
rect 4540 565 4670 580
rect -470 105 -340 120
rect -470 5 -455 105
rect -355 5 -340 105
rect -470 -10 -340 5
rect 4540 105 4670 120
rect 4540 5 4555 105
rect 4655 5 4670 105
rect 4540 -10 4670 5
rect -195 -100 -65 -85
rect -195 -200 -180 -100
rect -80 -200 -65 -100
rect -195 -215 -65 -200
rect 380 -100 510 -85
rect 380 -200 395 -100
rect 495 -200 510 -100
rect 380 -215 510 -200
rect 955 -100 1085 -85
rect 955 -200 970 -100
rect 1070 -200 1085 -100
rect 955 -215 1085 -200
rect 1530 -100 1660 -85
rect 1530 -200 1545 -100
rect 1645 -200 1660 -100
rect 1530 -215 1660 -200
rect 2105 -100 2235 -85
rect 2105 -200 2120 -100
rect 2220 -200 2235 -100
rect 2105 -215 2235 -200
rect 2680 -100 2810 -85
rect 2680 -200 2695 -100
rect 2795 -200 2810 -100
rect 2680 -215 2810 -200
rect 3255 -100 3385 -85
rect 3255 -200 3270 -100
rect 3370 -200 3385 -100
rect 3255 -215 3385 -200
rect 3830 -100 3960 -85
rect 3830 -200 3845 -100
rect 3945 -200 3960 -100
rect 3830 -215 3960 -200
rect 4405 -100 4535 -85
rect 4405 -200 4420 -100
rect 4520 -200 4535 -100
rect 4405 -215 4535 -200
<< nsubdiff >>
rect 3705 1334 3880 1370
rect 60 1229 235 1265
rect 60 1125 90 1229
rect 193 1125 235 1229
rect 3705 1230 3735 1334
rect 3838 1230 3880 1334
rect 3705 1195 3880 1230
rect 60 1090 235 1125
rect 1520 1159 1695 1195
rect 1520 1055 1550 1159
rect 1653 1055 1695 1159
rect 1520 1020 1695 1055
<< psubdiffcont >>
rect -190 2015 -90 2115
rect 385 2015 485 2115
rect 960 2015 1060 2115
rect 1535 2015 1635 2115
rect 2110 2015 2210 2115
rect 2685 2015 2785 2115
rect 3260 2015 3360 2115
rect 3835 2015 3935 2115
rect 4410 2015 4510 2115
rect -455 1730 -355 1830
rect 4555 1730 4655 1830
rect -455 1155 -355 1255
rect 4555 1155 4655 1255
rect -455 580 -355 680
rect 4555 580 4655 680
rect -455 5 -355 105
rect 4555 5 4655 105
rect -180 -200 -80 -100
rect 395 -200 495 -100
rect 970 -200 1070 -100
rect 1545 -200 1645 -100
rect 2120 -200 2220 -100
rect 2695 -200 2795 -100
rect 3270 -200 3370 -100
rect 3845 -200 3945 -100
rect 4420 -200 4520 -100
<< nsubdiffcont >>
rect 90 1125 193 1229
rect 3735 1230 3838 1334
rect 1550 1055 1653 1159
<< locali >>
rect -490 2115 4690 2150
rect -490 2015 -190 2115
rect -90 2015 385 2115
rect 485 2015 960 2115
rect 1060 2015 1535 2115
rect 1635 2015 2110 2115
rect 2210 2015 2685 2115
rect 2785 2015 3260 2115
rect 3360 2015 3835 2115
rect 3935 2015 4410 2115
rect 4510 2015 4690 2115
rect -490 1980 4690 2015
rect -490 1830 -320 1980
rect -490 1730 -455 1830
rect -355 1730 -320 1830
rect 4520 1830 4690 1980
rect -490 1255 -320 1730
rect 1975 1355 1995 1585
rect 2565 1570 2585 1695
rect 3400 1645 3420 1780
rect 3370 1625 3420 1645
rect 4520 1730 4555 1830
rect 4655 1730 4690 1830
rect 2415 1550 2585 1570
rect 1435 1335 1995 1355
rect -490 1155 -455 1255
rect -355 1155 -320 1255
rect 3724 1334 3854 1346
rect -490 680 -320 1155
rect 79 1229 209 1241
rect 79 1125 90 1229
rect 193 1228 209 1229
rect 79 1123 91 1125
rect 194 1123 209 1228
rect 3724 1230 3735 1334
rect 3838 1333 3854 1334
rect 3724 1228 3736 1230
rect 3839 1228 3854 1333
rect 3724 1217 3854 1228
rect 4520 1255 4690 1730
rect 79 1112 209 1123
rect 1539 1159 1669 1171
rect 1539 1055 1550 1159
rect 1653 1158 1669 1159
rect 1539 1053 1551 1055
rect 1654 1053 1669 1158
rect 1539 1042 1669 1053
rect 4520 1155 4555 1255
rect 4655 1155 4690 1255
rect 1655 945 2060 965
rect 1655 905 1675 945
rect 2035 850 2060 945
rect -490 580 -455 680
rect -355 580 -320 680
rect -490 105 -320 580
rect 4520 680 4690 1155
rect 4520 580 4555 680
rect 4655 580 4690 680
rect 4330 410 4395 435
rect -490 5 -455 105
rect -355 5 -320 105
rect -490 -65 -320 5
rect 4520 105 4690 580
rect 4520 5 4555 105
rect 4655 5 4690 105
rect 4520 -65 4690 5
rect -490 -100 4690 -65
rect -490 -200 -180 -100
rect -80 -200 395 -100
rect 495 -200 970 -100
rect 1070 -200 1545 -100
rect 1645 -200 2120 -100
rect 2220 -200 2695 -100
rect 2795 -200 3270 -100
rect 3370 -200 3845 -100
rect 3945 -200 4420 -100
rect 4520 -200 4690 -100
rect -490 -235 4690 -200
<< viali >>
rect 3400 1780 3420 1800
rect 3065 1675 3085 1695
rect 2870 1625 2890 1645
rect 91 1125 193 1228
rect 193 1125 194 1228
rect 91 1123 194 1125
rect 3736 1230 3838 1333
rect 3838 1230 3839 1333
rect 3736 1228 3839 1230
rect 1551 1055 1653 1158
rect 1653 1055 1654 1158
rect 1551 1053 1654 1055
rect 2730 410 2750 430
rect 3520 410 3540 430
rect 1990 340 2010 360
rect 2780 340 2800 360
rect 3570 340 3590 360
rect 970 -200 1070 -100
<< metal1 >>
rect 3390 1805 3430 1810
rect 3390 1775 3395 1805
rect 3425 1775 3430 1805
rect 3390 1770 3430 1775
rect 2970 1710 3010 1715
rect 2970 1695 2975 1710
rect 2885 1680 2975 1695
rect 3005 1680 3010 1710
rect 2970 1675 3010 1680
rect 3055 1695 3095 1705
rect 3055 1675 3065 1695
rect 3085 1675 3095 1695
rect 3370 1680 4330 1695
rect 3055 1665 3095 1675
rect 2860 1650 2900 1655
rect 2860 1620 2865 1650
rect 2895 1620 2900 1650
rect 2860 1615 2900 1620
rect 3070 1525 3085 1665
rect 2415 1510 3085 1525
rect 2970 1355 3010 1360
rect 2970 1345 2975 1355
rect 2965 1330 2975 1345
rect 2970 1325 2975 1330
rect 3005 1335 3010 1355
rect 3005 1325 3490 1335
rect 2970 1320 3490 1325
rect 79 1228 209 1241
rect 79 1123 91 1228
rect 194 1123 209 1228
rect 79 1112 209 1123
rect 1539 1158 1669 1171
rect 1539 1053 1551 1158
rect 1654 1053 1669 1158
rect 1539 1042 1669 1053
rect 2730 595 2770 600
rect 2730 585 2735 595
rect 2685 570 2735 585
rect 1980 360 2020 370
rect 1980 340 1990 360
rect 2010 340 2020 360
rect 2685 340 2700 570
rect 2730 565 2735 570
rect 2765 565 2770 595
rect 2730 560 2770 565
rect 2720 435 2760 440
rect 2720 405 2725 435
rect 2755 405 2760 435
rect 2720 400 2760 405
rect 2765 360 2810 370
rect 2730 340 2750 355
rect 1980 330 2020 340
rect 1990 290 2005 330
rect 1955 275 2005 290
rect 1955 30 1970 275
rect 2735 30 2750 340
rect 2765 340 2780 360
rect 2800 340 2810 360
rect 3475 340 3490 1320
rect 3724 1333 3854 1346
rect 3724 1228 3736 1333
rect 3839 1228 3854 1333
rect 3724 1217 3854 1228
rect 3510 435 3550 440
rect 3510 405 3515 435
rect 3545 405 3550 435
rect 3510 400 3550 405
rect 3560 360 3600 370
rect 2765 330 2810 340
rect 2765 125 2780 330
rect 2765 110 2855 125
rect 1955 15 2750 30
rect 2840 30 2855 110
rect 3530 30 3545 355
rect 3560 340 3570 360
rect 3590 340 3600 360
rect 3560 330 3600 340
rect 3575 140 3590 330
rect 3575 125 3650 140
rect 2840 15 3545 30
rect 3635 30 3650 125
rect 4315 30 4330 1680
rect 3635 15 4330 30
rect 961 -100 1080 -90
rect 961 -200 970 -100
rect 1070 -200 1080 -100
rect 961 -209 1080 -200
<< via1 >>
rect 3395 1800 3425 1805
rect 3395 1780 3400 1800
rect 3400 1780 3420 1800
rect 3420 1780 3425 1800
rect 3395 1775 3425 1780
rect 2975 1680 3005 1710
rect 2865 1645 2895 1650
rect 2865 1625 2870 1645
rect 2870 1625 2890 1645
rect 2890 1625 2895 1645
rect 2865 1620 2895 1625
rect 2975 1325 3005 1355
rect 91 1123 194 1228
rect 1551 1053 1654 1158
rect 2735 565 2765 595
rect 2725 430 2755 435
rect 2725 410 2730 430
rect 2730 410 2750 430
rect 2750 410 2755 430
rect 2725 405 2755 410
rect 3736 1228 3839 1333
rect 3515 430 3545 435
rect 3515 410 3520 430
rect 3520 410 3540 430
rect 3540 410 3545 430
rect 3515 405 3545 410
rect 970 -200 1070 -100
<< metal2 >>
rect 3385 1805 3435 1820
rect -185 1790 3395 1805
rect 3385 1775 3395 1790
rect 3425 1775 3435 1805
rect 3385 1765 3435 1775
rect 2965 1710 3015 1720
rect 2965 1680 2975 1710
rect 3005 1680 3015 1710
rect 2965 1670 3015 1680
rect 2855 1650 2905 1660
rect 2855 1620 2865 1650
rect 2895 1645 2905 1650
rect 2895 1620 2915 1645
rect 2855 1610 2915 1620
rect 79 1228 209 1241
rect 79 1123 91 1228
rect 194 1123 209 1228
rect 79 1112 209 1123
rect 1539 1158 1669 1171
rect 1539 1053 1551 1158
rect 1654 1053 1669 1158
rect 1539 1042 1669 1053
rect 2900 995 2915 1610
rect 2985 1365 3000 1670
rect 2965 1355 3015 1365
rect 2965 1325 2975 1355
rect 3005 1325 3015 1355
rect 2965 1315 3015 1325
rect 3724 1333 3854 1346
rect 3724 1228 3736 1333
rect 3839 1228 3854 1333
rect 3724 1217 3854 1228
rect 2745 980 2915 995
rect 2745 605 2760 980
rect 2725 595 2775 605
rect 2725 565 2735 595
rect 2765 565 2775 595
rect 2725 555 2775 565
rect -185 430 -155 450
rect 1955 430 1990 450
rect 2735 445 2780 450
rect 3520 445 3570 450
rect 2715 435 2780 445
rect 1955 340 1970 430
rect 2715 405 2725 435
rect 2755 430 2780 435
rect 3505 435 3570 445
rect 2755 405 2765 430
rect 2715 395 2765 405
rect 3505 405 3515 435
rect 3545 430 3570 435
rect 3545 405 3555 430
rect 3505 395 3555 405
rect 961 -100 1080 -90
rect 961 -200 970 -100
rect 1070 -200 1080 -100
rect 961 -209 1080 -200
<< via2 >>
rect 91 1123 194 1228
rect 1551 1053 1654 1158
rect 3736 1228 3839 1333
rect 970 -200 1070 -100
<< metal3 >>
rect 3724 1333 3854 1346
rect 79 1228 209 1241
rect 79 1123 91 1228
rect 194 1123 209 1228
rect 3724 1228 3736 1333
rect 3839 1228 3854 1333
rect 3724 1217 3854 1228
rect 79 1112 209 1123
rect 1539 1158 1669 1171
rect 1539 1053 1551 1158
rect 1654 1053 1669 1158
rect 1539 1042 1669 1053
rect 961 -100 1080 -90
rect 961 -200 970 -100
rect 1070 -200 1080 -100
rect 961 -209 1080 -200
<< via3 >>
rect 91 1123 194 1228
rect 3736 1228 3839 1333
rect 1551 1053 1654 1158
rect 970 -200 1070 -100
<< metal4 >>
rect 1885 1850 2040 1885
rect 2345 1865 2590 1895
rect 2885 1865 3070 1895
rect 1885 1530 1915 1850
rect 3645 1333 3940 1420
rect 129 1241 279 1278
rect 79 1228 279 1241
rect 79 1161 91 1228
rect 78 1123 91 1161
rect 194 1123 279 1228
rect 3645 1228 3736 1333
rect 3839 1228 3940 1333
rect 1589 1171 1705 1208
rect 78 1096 279 1123
rect 1539 1158 1705 1171
rect 78 1095 171 1096
rect 216 964 273 1096
rect 1539 1091 1551 1158
rect 1538 1053 1551 1091
rect 1654 1053 1705 1158
rect 2350 1080 2785 1110
rect 2885 1080 3070 1110
rect 3645 1065 3940 1228
rect 1538 1050 1705 1053
rect 1538 1025 1710 1050
rect 1549 975 1710 1025
rect 1549 941 1642 975
rect 1995 960 2415 995
rect 2725 930 2815 960
rect 3515 930 3605 960
rect 3650 934 3711 1065
rect 969 -90 1073 29
rect 1915 15 2005 45
rect 2715 15 2810 45
rect 3510 15 3600 45
rect 961 -100 1080 -90
rect 961 -200 970 -100
rect 1070 -200 1080 -100
rect 961 -209 1080 -200
use tspc  tspc_2
timestamp 1640956963
transform 1 0 3640 0 1 495
box -70 -490 690 465
use tspc  tspc_1
timestamp 1640956963
transform 1 0 2850 0 1 495
box -70 -490 690 465
use tspc  tspc_0
timestamp 1640956963
transform 1 0 2060 0 1 495
box -70 -490 690 465
use prescaler  prescaler_0
timestamp 1643048518
transform 1 0 25 0 1 200
box -210 -195 1930 1715
use and  and_0
timestamp 1640957225
transform -1 0 2330 0 -1 1465
box -85 -435 335 475
use nor  nor_0
timestamp 1640957264
transform -1 0 2830 0 -1 1605
box -55 -300 245 610
use nor  nor_1
timestamp 1640957264
transform -1 0 3315 0 -1 1605
box -55 -300 245 610
<< labels >>
rlabel metal4 1915 15 2005 45 1 gnd
rlabel metal4 2715 15 2810 45 1 gnd
rlabel space 3510 15 3605 45 1 gnd
rlabel space 3515 930 3610 960 1 vdd
rlabel metal4 2725 930 2815 960 1 vdd
rlabel metal4 1995 965 2415 995 1 vdd
rlabel metal4 2350 1080 2585 1110 1 vdd
rlabel metal4 2885 1080 3070 1110 1 vdd
rlabel metal4 1885 1560 1915 1885 1 gnd
rlabel metal4 1915 1850 2035 1885 1 gnd
rlabel locali 4330 410 4395 435 1 Out
rlabel metal2 -185 430 -155 450 1 clk
rlabel metal2 -185 1790 225 1805 1 mc2
<< end >>
