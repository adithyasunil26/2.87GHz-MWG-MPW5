magic
tech sky130A
timestamp 1647861083
<< locali >>
rect 74 11286 277 11316
rect 74 11148 100 11286
rect 247 11148 277 11286
rect 74 11113 277 11148
<< viali >>
rect 100 11148 247 11286
<< metal1 >>
rect 74 11286 277 11316
rect 74 11148 100 11286
rect 247 11148 277 11286
rect 74 11113 277 11148
rect 4144 10873 4266 10923
rect 4144 10778 4149 10873
rect 4257 10778 4266 10873
rect 4144 10406 4266 10778
rect 4141 10358 4266 10406
rect 4141 9841 4263 10358
<< via1 >>
rect 100 11148 247 11286
rect 4149 10778 4257 10873
<< metal2 >>
rect 225 14044 716 14120
rect 230 13223 395 14044
rect 225 12982 395 13223
rect 493 13171 696 13227
rect 493 13039 527 13171
rect 664 13039 696 13171
rect 225 12491 400 12982
rect 493 12653 696 13039
rect 230 12268 400 12491
rect 506 12268 685 12290
rect 230 12254 685 12268
rect 230 12138 529 12254
rect 645 12138 685 12254
rect 230 12125 685 12138
rect 506 12094 685 12125
rect 828 11598 930 12714
rect 826 11482 4275 11598
rect 74 11286 277 11316
rect 74 11148 100 11286
rect 247 11148 277 11286
rect 74 11113 277 11148
rect 4136 10873 4275 11482
rect 4136 10778 4149 10873
rect 4257 10778 4275 10873
rect 4136 10744 4275 10778
<< via2 >>
rect 527 13039 664 13171
rect 529 12138 645 12254
rect 100 11148 247 11286
<< metal3 >>
rect 511 13171 683 13187
rect 511 13039 527 13171
rect 664 13039 683 13171
rect 511 13017 683 13039
rect 506 12254 685 12290
rect 506 12138 529 12254
rect 645 12138 685 12254
rect 506 12094 685 12138
rect 74 11286 277 11316
rect 74 11148 100 11286
rect 247 11148 277 11286
rect 74 11113 277 11148
<< via3 >>
rect 527 13039 664 13171
rect 529 12138 645 12254
rect 100 11148 247 11286
<< metal4 >>
rect 70 13964 750 13966
rect 70 13835 1017 13964
rect 70 13833 750 13835
rect 72 12567 286 13833
rect 495 13171 695 13660
rect 495 13039 527 13171
rect 664 13039 695 13171
rect 495 12970 695 13039
rect 72 12552 1015 12567
rect 73 12438 1015 12552
rect 74 11286 282 12438
rect 506 12254 685 12290
rect 506 12138 529 12254
rect 645 12138 685 12254
rect 506 12094 685 12138
rect 74 11148 100 11286
rect 247 11148 282 11286
rect 74 11113 282 11148
<< metal5 >>
rect 849 13034 1059 13173
use tapered_buf  tapered_buf_1
timestamp 1647818295
transform 1 0 1130 0 1 14049
box -470 -910 43675 401
use tapered_buf  tapered_buf_0
timestamp 1647818295
transform 1 0 1128 0 1 12652
box -470 -910 43675 401
use filter  filter_0
timestamp 1640983258
transform 1 0 1799 0 1 11005
box -1800 -11005 6240 390
<< labels >>
rlabel space 1528 12972 1528 12972 1 vdd!
rlabel metal4 184 11701 184 11701 1 gnd!
rlabel space 1530 14369 1530 14369 1 vdd!
rlabel metal2 347 14081 347 14081 1 v
<< end >>
