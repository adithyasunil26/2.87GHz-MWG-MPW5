magic
tech sky130A
timestamp 1647791355
<< locali >>
rect -665 7851 -464 7889
rect -665 7720 -635 7851
rect -504 7720 -464 7851
rect -665 7690 -464 7720
rect -177 6992 19 6995
rect -177 6973 560 6992
rect -177 6827 -153 6973
rect -5 6827 560 6973
rect -177 6820 560 6827
rect -177 6809 19 6820
rect -573 613 -389 616
rect -573 595 161 613
rect -573 444 -555 595
rect -408 444 161 595
rect -573 430 -389 444
rect 1446 -30 1498 1375
rect 1931 0 1983 1359
rect 2426 93 2478 1401
rect 1440 -111 1500 -30
rect 1386 -119 1500 -111
rect -2173 -245 1500 -119
rect -2173 -249 1495 -245
rect -2173 -9118 -2064 -249
rect 1386 -250 1495 -249
rect 1927 -335 1983 0
rect 2421 -58 2478 93
rect -1869 -336 1987 -335
rect -1926 -431 1987 -336
rect -1926 -1977 -1839 -431
rect -1702 -512 -1576 -502
rect 2421 -512 2474 -58
rect 2901 -62 2953 1365
rect 3396 -34 3448 1370
rect 3999 190 4051 1437
rect -1702 -596 2479 -512
rect -1934 -8213 -1830 -1977
rect -1702 -6898 -1576 -596
rect -1450 -665 -1239 -661
rect 2895 -665 2953 -62
rect -1450 -675 2963 -665
rect -1452 -770 2963 -675
rect -1452 -772 1200 -770
rect -1452 -781 -1239 -772
rect -1452 -5319 -1336 -781
rect -1206 -880 -1122 -877
rect -1206 -885 2992 -880
rect 3395 -885 3455 -34
rect -1206 -963 3455 -885
rect -1206 -968 3453 -963
rect -1206 -1455 -1122 -968
rect 3998 -1039 4055 190
rect -1213 -1495 -1122 -1455
rect -1012 -1044 -937 -1040
rect -144 -1044 4060 -1039
rect -1012 -1137 4060 -1044
rect -1012 -1147 -113 -1137
rect -1213 -3202 -1124 -1495
rect -1012 -2032 -937 -1147
rect -1012 -2058 -732 -2032
rect -1012 -2162 -872 -2058
rect -750 -2162 -732 -2058
rect -1012 -2180 -732 -2162
rect -1213 -3648 -1125 -3202
rect -1213 -3663 -718 -3648
rect -1213 -3778 -880 -3663
rect -766 -3778 -718 -3663
rect -1213 -3796 -718 -3778
rect -898 -3802 -749 -3796
rect -1458 -5343 -862 -5319
rect -1458 -5462 -1206 -5343
rect -1081 -5462 -862 -5343
rect -1458 -5483 -862 -5462
rect -1702 -6935 -757 -6898
rect -1702 -7065 -1136 -6935
rect -994 -7065 -757 -6935
rect -1702 -7093 -757 -7065
rect -1934 -8708 -1824 -8213
rect -1934 -8735 -877 -8708
rect -1934 -8842 -1301 -8735
rect -1183 -8842 -877 -8735
rect -1934 -8870 -877 -8842
rect -2178 -9225 -2064 -9118
rect -2178 -10307 -2068 -9225
rect -1455 -10307 -1236 -10296
rect -2183 -10323 -1083 -10307
rect -2183 -10493 -1433 -10323
rect -1263 -10493 -1083 -10323
rect -2183 -10509 -1083 -10493
rect -1455 -10515 -1236 -10509
<< viali >>
rect -635 7720 -504 7851
rect -153 6827 -5 6973
rect 33 3154 137 3250
rect -555 444 -408 595
rect -872 -2162 -750 -2058
rect -880 -3778 -766 -3663
rect -1206 -5462 -1081 -5343
rect -1136 -7065 -994 -6935
rect -1301 -8842 -1183 -8735
rect -1433 -10493 -1263 -10323
<< metal1 >>
rect -665 7851 -464 7889
rect -665 7720 -635 7851
rect -504 7720 -464 7851
rect -665 7690 -464 7720
rect -628 6149 -528 7690
rect -177 6973 19 6995
rect -177 6827 -153 6973
rect -5 6827 19 6973
rect -177 6809 19 6827
rect -628 6114 -504 6149
rect 183 6114 956 6116
rect -628 6022 956 6114
rect -628 6016 239 6022
rect -628 6015 128 6016
rect 14 3250 156 3280
rect 14 3154 33 3250
rect 137 3154 156 3250
rect 14 3122 156 3154
rect -573 595 -389 616
rect -573 444 -555 595
rect -408 444 -389 595
rect -573 430 -389 444
rect -890 -2058 -719 -2030
rect -890 -2162 -872 -2058
rect -750 -2162 -719 -2058
rect -890 -2186 -719 -2162
rect -898 -3663 -749 -3648
rect -898 -3778 -880 -3663
rect -766 -3778 -749 -3663
rect -898 -3802 -749 -3778
rect -1234 -5343 -1050 -5322
rect -1234 -5462 -1206 -5343
rect -1081 -5462 -1050 -5343
rect -1234 -5480 -1050 -5462
rect -1157 -6935 -973 -6910
rect -1157 -7065 -1136 -6935
rect -994 -7065 -973 -6935
rect -1157 -7086 -973 -7065
rect -1320 -8735 -1161 -8712
rect -1320 -8842 -1301 -8735
rect -1183 -8842 -1161 -8735
rect -1320 -8866 -1161 -8842
rect -1455 -10323 -1236 -10296
rect -1455 -10493 -1433 -10323
rect -1263 -10493 -1236 -10323
rect -1455 -10515 -1236 -10493
<< via1 >>
rect -635 7720 -504 7851
rect -153 6827 -5 6973
rect 33 3154 137 3250
rect -555 444 -408 595
rect -872 -2162 -750 -2058
rect -880 -3778 -766 -3663
rect -1206 -5462 -1081 -5343
rect -1136 -7065 -994 -6935
rect -1301 -8842 -1183 -8735
rect -1433 -10493 -1263 -10323
<< metal2 >>
rect -1357 9938 -1213 9939
rect -1357 9872 -351 9938
rect -1357 7369 -1213 9872
rect -665 7851 -464 7889
rect -665 7720 -635 7851
rect -504 7720 -464 7851
rect -665 7690 -464 7720
rect -854 7369 4474 7372
rect -1357 7228 4474 7369
rect -1357 7223 1825 7228
rect -1357 7220 -765 7223
rect -177 6973 19 6995
rect -177 6827 -153 6973
rect -5 6827 19 6973
rect -177 6809 19 6827
rect 4349 6343 4469 7228
rect 14 3250 156 3280
rect 14 3154 33 3250
rect 137 3154 156 3250
rect 14 3122 156 3154
rect -573 595 -389 616
rect -573 444 -555 595
rect -408 444 -389 595
rect -573 430 -389 444
rect -890 -2058 -719 -2030
rect -890 -2162 -872 -2058
rect -750 -2162 -719 -2058
rect -890 -2186 -719 -2162
rect -898 -3663 -749 -3648
rect -898 -3778 -880 -3663
rect -766 -3778 -749 -3663
rect -898 -3802 -749 -3778
rect -1234 -5343 -1050 -5322
rect -1234 -5462 -1206 -5343
rect -1081 -5462 -1050 -5343
rect -1234 -5480 -1050 -5462
rect -1157 -6935 -973 -6910
rect -1157 -7065 -1136 -6935
rect -994 -7065 -973 -6935
rect -1157 -7086 -973 -7065
rect -1320 -8735 -1161 -8712
rect -1320 -8842 -1301 -8735
rect -1183 -8842 -1161 -8735
rect -1320 -8866 -1161 -8842
rect -1455 -10323 -1236 -10296
rect -1455 -10493 -1433 -10323
rect -1263 -10493 -1236 -10323
rect -1455 -10515 -1236 -10493
<< via2 >>
rect -635 7720 -504 7851
rect -153 6827 -5 6973
rect 33 3154 137 3250
rect -555 444 -408 595
rect -872 -2162 -750 -2058
rect -880 -3778 -766 -3663
rect -1206 -5462 -1081 -5343
rect -1136 -7065 -994 -6935
rect -1301 -8842 -1183 -8735
rect -1433 -10493 -1263 -10323
<< metal3 >>
rect -665 7851 -464 7889
rect -665 7720 -635 7851
rect -504 7720 -464 7851
rect -665 7690 -464 7720
rect -177 6973 19 6995
rect -177 6827 -153 6973
rect -5 6827 19 6973
rect -177 6809 19 6827
rect 14 3250 156 3280
rect 14 3154 33 3250
rect 137 3154 156 3250
rect 14 3122 156 3154
rect -573 595 -389 616
rect -573 444 -555 595
rect -408 444 -389 595
rect -573 430 -389 444
rect -890 -2058 -719 -2030
rect -890 -2162 -872 -2058
rect -750 -2162 -719 -2058
rect -890 -2186 -719 -2162
rect -898 -3663 -749 -3648
rect -898 -3778 -880 -3663
rect -766 -3778 -749 -3663
rect -898 -3802 -749 -3778
rect -1234 -5343 -1050 -5322
rect -1234 -5462 -1206 -5343
rect -1081 -5462 -1050 -5343
rect -1234 -5480 -1050 -5462
rect -1157 -6935 -973 -6910
rect -1157 -7065 -1136 -6935
rect -994 -7065 -973 -6935
rect -1157 -7086 -973 -7065
rect -1320 -8735 -1161 -8712
rect -1320 -8842 -1301 -8735
rect -1183 -8842 -1161 -8735
rect -1320 -8866 -1161 -8842
rect -1455 -10323 -1236 -10296
rect -1455 -10493 -1433 -10323
rect -1263 -10493 -1236 -10323
rect -1455 -10515 -1236 -10493
<< via3 >>
rect -635 7720 -504 7851
rect -153 6827 -5 6973
rect 33 3154 137 3250
rect -555 444 -408 595
rect -872 -2162 -750 -2058
rect -880 -3778 -766 -3663
rect -1206 -5462 -1081 -5343
rect -1136 -7065 -994 -6935
rect -1301 -8842 -1183 -8735
rect -1433 -10493 -1263 -10323
<< metal4 >>
rect -2962 9651 -69 9791
rect -2962 8149 -2652 9651
rect -702 8149 -417 8152
rect -2962 8009 -64 8149
rect -2962 3370 -2652 8009
rect -702 8003 -417 8009
rect -665 7859 -464 7889
rect -665 7851 -324 7859
rect -665 7720 -635 7851
rect -504 7728 -324 7851
rect -504 7720 -464 7728
rect -665 7690 -464 7720
rect -177 6973 19 6995
rect -177 6827 -153 6973
rect -5 6827 19 6973
rect -177 6809 19 6827
rect -2962 3250 167 3370
rect -2962 3154 33 3250
rect 137 3154 167 3250
rect -2962 3037 167 3154
rect -2962 -1749 -2652 3037
rect -573 595 -389 616
rect -573 444 -555 595
rect -408 444 -389 595
rect -573 430 -389 444
rect -2962 -1880 -364 -1749
rect -2962 -3367 -2652 -1880
rect -937 -2058 -654 -2014
rect -937 -2162 -872 -2058
rect -750 -2162 -654 -2058
rect -937 -2188 -654 -2162
rect -1305 -3367 -1213 -3361
rect -2962 -3498 -1213 -3367
rect -2962 -5020 -2652 -3498
rect -1305 -3502 -1213 -3498
rect -1125 -3367 -1002 -3361
rect -1125 -3498 -340 -3367
rect -1125 -3502 -1002 -3498
rect -950 -3663 -643 -3645
rect -950 -3778 -880 -3663
rect -766 -3778 -643 -3663
rect -950 -3799 -643 -3778
rect -898 -3802 -749 -3799
rect -2962 -5151 -450 -5020
rect -2962 -6646 -2652 -5151
rect -1338 -5343 -713 -5319
rect -1338 -5462 -1206 -5343
rect -1081 -5462 -713 -5343
rect -1338 -5483 -713 -5462
rect -2962 -6777 -412 -6646
rect -2962 -8426 -2652 -6777
rect -1383 -6935 -672 -6888
rect -1383 -7065 -1136 -6935
rect -994 -7065 -672 -6935
rect -1383 -7103 -672 -7065
rect -2962 -8557 -485 -8426
rect -2962 -10044 -2652 -8557
rect -1663 -8735 -844 -8692
rect -1663 -8842 -1301 -8735
rect -1183 -8842 -844 -8735
rect -1663 -8880 -844 -8842
rect -2962 -10174 -471 -10044
rect -2527 -10175 -471 -10174
rect -1576 -10323 -771 -10296
rect -1576 -10493 -1433 -10323
rect -1263 -10493 -771 -10323
rect -1576 -10504 -771 -10493
rect -1455 -10515 -1236 -10504
<< via4 >>
rect -153 6827 -5 6973
rect -555 444 -408 595
<< metal5 >>
rect -222 8629 23 8999
rect -186 6973 30 7474
rect -186 6827 -153 6973
rect -5 6827 30 6973
rect -186 6788 30 6827
rect -605 595 -369 655
rect -605 444 -555 595
rect -408 444 -369 595
rect -605 376 -369 444
rect -605 61 -367 376
rect -605 -29 -369 61
rect -606 -1262 -369 -29
rect -606 -1515 -555 -1262
rect -606 -2520 -363 -2506
rect -606 -2877 -318 -2520
rect -606 -3116 -496 -2877
rect -611 -4103 -519 -4023
rect -642 -4552 -338 -4103
rect -655 -5993 -360 -5805
rect -685 -6161 -360 -5993
rect -685 -6395 -575 -6161
rect -703 -7680 -381 -7419
rect -737 -7941 -381 -7680
rect -737 -8082 -627 -7941
rect -716 -9196 -596 -9189
rect -716 -9424 -449 -9196
rect -711 -9559 -449 -9424
rect -711 -9700 -601 -9559
use tapered_buf  tapered_buf_2
timestamp 1647784636
transform 1 0 -296 0 1 -1652
box -470 -910 43675 400
use tapered_buf  tapered_buf_3
timestamp 1647784636
transform 1 0 -256 0 1 -3271
box -470 -910 43675 400
use tapered_buf  tapered_buf_4
timestamp 1647784636
transform 1 0 -375 0 1 -4929
box -470 -910 43675 400
use tapered_buf  tapered_buf_5
timestamp 1647784636
transform 1 0 -335 0 1 -6548
box -470 -910 43675 400
use tapered_buf  tapered_buf_6
timestamp 1647784636
transform 1 0 -414 0 1 -8329
box -470 -910 43675 400
use tapered_buf  tapered_buf_7
timestamp 1647784636
transform 1 0 -374 0 1 -9948
box -470 -910 43675 400
use ro_complete  ro_complete_0
timestamp 1647788658
transform 1 0 348 0 1 5690
box -348 -5690 4661 1440
use tapered_buf  tapered_buf_1
timestamp 1647784636
transform 1 0 60 0 1 9871
box -470 -910 43675 400
use tapered_buf  tapered_buf_0
timestamp 1647784636
transform 1 0 100 0 1 8252
box -470 -910 43675 400
<< labels >>
rlabel space -112 10260 -112 10260 1 vdd!
rlabel space -324 8284 -324 8284 1 vcont
rlabel space -338 9409 -338 9409 1 out
rlabel metal4 -2844 3190 -2844 3190 1 gnd!
rlabel space -819 -9903 -819 -9903 1 a0
rlabel space -854 -8280 -854 -8280 1 a1
rlabel space -779 -6505 -779 -6505 1 a2
rlabel space -798 -4893 -798 -4893 1 a3
rlabel space -701 -3231 -701 -3231 1 a4
rlabel space -728 -1606 -728 -1606 1 a5
<< end >>
