magic
tech sky130A
timestamp 1640776259
<< nwell >>
rect -80 -35 335 265
<< nmos >>
rect 10 -235 25 -145
rect 135 -235 150 -145
rect 260 -235 275 -145
<< pmos >>
rect 10 -15 25 165
rect 135 -15 150 165
rect 260 -15 275 165
<< ndiff >>
rect -30 -155 10 -145
rect -30 -180 -25 -155
rect 0 -180 10 -155
rect -30 -200 10 -180
rect -30 -225 -25 -200
rect 0 -225 10 -200
rect -30 -235 10 -225
rect 25 -155 65 -145
rect 25 -180 35 -155
rect 60 -180 65 -155
rect 25 -200 65 -180
rect 25 -225 35 -200
rect 60 -225 65 -200
rect 25 -235 65 -225
rect 95 -155 135 -145
rect 95 -180 100 -155
rect 125 -180 135 -155
rect 95 -200 135 -180
rect 95 -225 100 -200
rect 125 -225 135 -200
rect 95 -235 135 -225
rect 150 -155 190 -145
rect 150 -180 160 -155
rect 185 -180 190 -155
rect 150 -200 190 -180
rect 150 -225 160 -200
rect 185 -225 190 -200
rect 150 -235 190 -225
rect 220 -155 260 -145
rect 220 -180 225 -155
rect 250 -180 260 -155
rect 220 -200 260 -180
rect 220 -225 225 -200
rect 250 -225 260 -200
rect 220 -235 260 -225
rect 275 -155 315 -145
rect 275 -180 285 -155
rect 310 -180 315 -155
rect 275 -200 315 -180
rect 275 -225 285 -200
rect 310 -225 315 -200
rect 275 -235 315 -225
<< pdiff >>
rect -30 155 10 165
rect -30 130 -25 155
rect 0 130 10 155
rect -30 110 10 130
rect -30 85 -25 110
rect 0 85 10 110
rect -30 65 10 85
rect -30 40 -25 65
rect 0 40 10 65
rect -30 20 10 40
rect -30 -5 -25 20
rect 0 -5 10 20
rect -30 -15 10 -5
rect 25 155 65 165
rect 25 130 35 155
rect 60 130 65 155
rect 25 110 65 130
rect 25 85 35 110
rect 60 85 65 110
rect 25 65 65 85
rect 25 40 35 65
rect 60 40 65 65
rect 25 20 65 40
rect 25 -5 35 20
rect 60 -5 65 20
rect 25 -15 65 -5
rect 95 155 135 165
rect 95 130 100 155
rect 125 130 135 155
rect 95 110 135 130
rect 95 85 100 110
rect 125 85 135 110
rect 95 65 135 85
rect 95 40 100 65
rect 125 40 135 65
rect 95 20 135 40
rect 95 -5 100 20
rect 125 -5 135 20
rect 95 -15 135 -5
rect 150 155 190 165
rect 150 130 160 155
rect 185 130 190 155
rect 150 110 190 130
rect 150 85 160 110
rect 185 85 190 110
rect 150 65 190 85
rect 150 40 160 65
rect 185 40 190 65
rect 150 20 190 40
rect 150 -5 160 20
rect 185 -5 190 20
rect 150 -15 190 -5
rect 220 155 260 165
rect 220 130 225 155
rect 250 130 260 155
rect 220 110 260 130
rect 220 85 225 110
rect 250 85 260 110
rect 220 65 260 85
rect 220 40 225 65
rect 250 40 260 65
rect 220 20 260 40
rect 220 -5 225 20
rect 250 -5 260 20
rect 220 -15 260 -5
rect 275 155 315 165
rect 275 130 285 155
rect 310 130 315 155
rect 275 110 315 130
rect 275 85 285 110
rect 310 85 315 110
rect 275 65 315 85
rect 275 40 285 65
rect 310 40 315 65
rect 275 20 315 40
rect 275 -5 285 20
rect 310 -5 315 20
rect 275 -15 315 -5
<< ndiffc >>
rect -25 -180 0 -155
rect -25 -225 0 -200
rect 35 -180 60 -155
rect 35 -225 60 -200
rect 100 -180 125 -155
rect 100 -225 125 -200
rect 160 -180 185 -155
rect 160 -225 185 -200
rect 225 -180 250 -155
rect 225 -225 250 -200
rect 285 -180 310 -155
rect 285 -225 310 -200
<< pdiffc >>
rect -25 130 0 155
rect -25 85 0 110
rect -25 40 0 65
rect -25 -5 0 20
rect 35 130 60 155
rect 35 85 60 110
rect 35 40 60 65
rect 35 -5 60 20
rect 100 130 125 155
rect 100 85 125 110
rect 100 40 125 65
rect 100 -5 125 20
rect 160 130 185 155
rect 160 85 185 110
rect 160 40 185 65
rect 160 -5 185 20
rect 225 130 250 155
rect 225 85 250 110
rect 225 40 250 65
rect 225 -5 250 20
rect 285 130 310 155
rect 285 85 310 110
rect 285 40 310 65
rect 285 -5 310 20
<< poly >>
rect 10 165 25 180
rect 135 165 150 180
rect 260 165 275 180
rect 10 -85 25 -15
rect 135 -85 150 -15
rect 260 -85 275 -15
rect -30 -95 25 -85
rect -30 -115 -20 -95
rect 0 -115 25 -95
rect -30 -125 25 -115
rect 95 -95 150 -85
rect 95 -115 105 -95
rect 125 -115 150 -95
rect 95 -125 150 -115
rect 220 -95 275 -85
rect 220 -115 230 -95
rect 250 -115 275 -95
rect 220 -125 275 -115
rect 10 -145 25 -125
rect 135 -145 150 -125
rect 260 -145 275 -125
rect 10 -255 25 -235
rect 135 -255 150 -235
rect 260 -255 275 -235
<< polycont >>
rect -20 -115 0 -95
rect 105 -115 125 -95
rect 230 -115 250 -95
<< locali >>
rect -25 165 -5 200
rect 100 165 120 200
rect 220 165 240 200
rect -30 155 5 165
rect -30 130 -25 155
rect 0 130 5 155
rect -30 110 5 130
rect -30 85 -25 110
rect 0 85 5 110
rect -30 65 5 85
rect -30 40 -25 65
rect 0 40 5 65
rect -30 20 5 40
rect -30 -5 -25 20
rect 0 -5 5 20
rect -30 -15 5 -5
rect 30 155 65 165
rect 30 130 35 155
rect 60 130 65 155
rect 30 110 65 130
rect 30 85 35 110
rect 60 85 65 110
rect 30 65 65 85
rect 30 40 35 65
rect 60 40 65 65
rect 30 20 65 40
rect 30 -5 35 20
rect 60 -5 65 20
rect 30 -15 65 -5
rect 95 155 130 165
rect 95 130 100 155
rect 125 130 130 155
rect 95 110 130 130
rect 95 85 100 110
rect 125 85 130 110
rect 95 65 130 85
rect 95 40 100 65
rect 125 40 130 65
rect 95 20 130 40
rect 95 -5 100 20
rect 125 -5 130 20
rect 95 -15 130 -5
rect 155 155 190 165
rect 155 130 160 155
rect 185 130 190 155
rect 155 110 190 130
rect 155 85 160 110
rect 185 85 190 110
rect 155 65 190 85
rect 155 40 160 65
rect 185 40 190 65
rect 155 20 190 40
rect 155 -5 160 20
rect 185 -5 190 20
rect 155 -15 190 -5
rect 220 155 255 165
rect 220 130 225 155
rect 250 130 255 155
rect 220 110 255 130
rect 220 85 225 110
rect 250 85 255 110
rect 220 65 255 85
rect 220 40 225 65
rect 250 40 255 65
rect 220 20 255 40
rect 220 -5 225 20
rect 250 -5 255 20
rect 220 -15 255 -5
rect 280 155 315 165
rect 280 130 285 155
rect 310 130 315 155
rect 280 110 315 130
rect 280 85 285 110
rect 310 85 315 110
rect 280 65 315 85
rect 280 40 285 65
rect 310 40 315 65
rect 280 20 315 40
rect 280 -5 285 20
rect 310 -5 315 20
rect 280 -15 315 -5
rect 35 -35 60 -15
rect 160 -35 185 -15
rect 35 -55 185 -35
rect -30 -95 10 -85
rect -50 -115 -20 -95
rect 0 -115 10 -95
rect -30 -125 10 -115
rect 95 -95 135 -85
rect 95 -115 105 -95
rect 125 -115 135 -95
rect 95 -125 135 -115
rect 160 -95 185 -55
rect 220 -95 260 -85
rect 160 -115 230 -95
rect 250 -115 260 -95
rect 160 -145 185 -115
rect 220 -125 260 -115
rect 285 -95 310 -15
rect 285 -115 335 -95
rect 285 -145 310 -115
rect -30 -155 5 -145
rect -30 -180 -25 -155
rect 0 -180 5 -155
rect -30 -200 5 -180
rect -30 -225 -25 -200
rect 0 -225 5 -200
rect -30 -235 5 -225
rect 30 -155 65 -145
rect 30 -180 35 -155
rect 60 -180 65 -155
rect 95 -155 130 -145
rect 95 -180 100 -155
rect 125 -180 130 -155
rect 30 -200 130 -180
rect 30 -225 35 -200
rect 60 -225 65 -200
rect 30 -235 65 -225
rect 95 -225 100 -200
rect 125 -225 130 -200
rect 95 -235 130 -225
rect 155 -155 190 -145
rect 155 -180 160 -155
rect 185 -180 190 -155
rect 155 -200 190 -180
rect 155 -225 160 -200
rect 185 -225 190 -200
rect 155 -235 190 -225
rect 220 -155 255 -145
rect 220 -180 225 -155
rect 250 -180 255 -155
rect 220 -200 255 -180
rect 220 -225 225 -200
rect 250 -225 255 -200
rect 220 -235 255 -225
rect 280 -155 315 -145
rect 280 -180 285 -155
rect 310 -180 315 -155
rect 280 -200 315 -180
rect 280 -225 285 -200
rect 310 -225 315 -200
rect 280 -235 315 -225
rect -25 -285 0 -235
rect -5 -295 0 -285
rect 225 -285 250 -235
rect 245 -295 250 -285
<< viali >>
rect -25 200 -5 220
rect 100 200 120 220
rect 220 200 240 220
rect 105 -115 125 -95
rect -25 -305 -5 -285
rect 225 -305 245 -285
<< metal1 >>
rect -35 225 5 230
rect -35 195 -30 225
rect 0 195 5 225
rect -35 190 5 195
rect 90 225 130 230
rect 90 195 95 225
rect 125 195 130 225
rect 90 190 130 195
rect 210 225 250 230
rect 210 195 215 225
rect 245 195 250 225
rect 210 190 250 195
rect -50 -60 120 -45
rect 105 -85 120 -60
rect 95 -95 135 -85
rect 95 -115 105 -95
rect 125 -115 135 -95
rect 95 -125 135 -115
rect -35 -280 5 -275
rect -35 -310 -30 -280
rect 0 -310 5 -280
rect -35 -315 5 -310
rect 215 -280 255 -275
rect 215 -310 220 -280
rect 250 -310 255 -280
rect 215 -315 255 -310
<< via1 >>
rect -30 220 0 225
rect -30 200 -25 220
rect -25 200 -5 220
rect -5 200 0 220
rect -30 195 0 200
rect 95 220 125 225
rect 95 200 100 220
rect 100 200 120 220
rect 120 200 125 220
rect 95 195 125 200
rect 215 220 245 225
rect 215 200 220 220
rect 220 200 240 220
rect 240 200 245 220
rect 215 195 245 200
rect -30 -285 0 -280
rect -30 -305 -25 -285
rect -25 -305 -5 -285
rect -5 -305 0 -285
rect -30 -310 0 -305
rect 220 -285 250 -280
rect 220 -305 225 -285
rect 225 -305 245 -285
rect 245 -305 250 -285
rect 220 -310 250 -305
<< metal2 >>
rect -40 225 10 235
rect -40 195 -30 225
rect 0 195 10 225
rect -40 185 10 195
rect 85 225 135 235
rect 85 195 95 225
rect 125 195 135 225
rect 85 185 135 195
rect 205 225 255 235
rect 205 195 215 225
rect 245 195 255 225
rect 205 185 255 195
rect -40 -280 10 -270
rect -40 -310 -30 -280
rect 0 -310 10 -280
rect -40 -320 10 -310
rect 210 -280 260 -270
rect 210 -310 220 -280
rect 250 -310 260 -280
rect 210 -320 260 -310
<< via2 >>
rect -30 195 0 225
rect 95 195 125 225
rect 215 195 245 225
rect -30 -310 0 -280
rect 220 -310 250 -280
<< metal3 >>
rect -40 230 10 235
rect -40 190 -35 230
rect 5 190 10 230
rect -40 185 10 190
rect 85 230 135 235
rect 85 190 90 230
rect 130 190 135 230
rect 85 185 135 190
rect 205 230 255 235
rect 205 190 210 230
rect 250 190 255 230
rect 205 185 255 190
rect -40 -275 10 -270
rect -40 -315 -35 -275
rect 5 -315 10 -275
rect -40 -320 10 -315
rect 210 -275 260 -270
rect 210 -315 215 -275
rect 255 -315 260 -275
rect 210 -320 260 -315
<< via3 >>
rect -35 225 5 230
rect -35 195 -30 225
rect -30 195 0 225
rect 0 195 5 225
rect -35 190 5 195
rect 90 225 130 230
rect 90 195 95 225
rect 95 195 125 225
rect 125 195 130 225
rect 90 190 130 195
rect 210 225 250 230
rect 210 195 215 225
rect 215 195 245 225
rect 245 195 250 225
rect 210 190 250 195
rect -35 -280 5 -275
rect -35 -310 -30 -280
rect -30 -310 0 -280
rect 0 -310 5 -280
rect -35 -315 5 -310
rect 215 -280 255 -275
rect 215 -310 220 -280
rect 220 -310 250 -280
rect 250 -310 255 -280
rect 215 -315 255 -310
<< metal4 >>
rect -120 235 -80 275
rect -45 235 15 240
rect 80 235 140 240
rect 200 235 260 240
rect -120 230 335 235
rect -120 205 -35 230
rect -45 190 -35 205
rect 5 205 90 230
rect 5 190 15 205
rect -45 180 15 190
rect 80 190 90 205
rect 130 205 210 230
rect 130 190 140 205
rect 80 180 140 190
rect 200 190 210 205
rect 250 205 335 230
rect 250 190 260 205
rect 200 180 260 190
rect -45 -275 15 -265
rect 205 -275 265 -265
rect -115 -310 -35 -275
rect -115 -375 -80 -310
rect -45 -315 -35 -310
rect 5 -310 215 -275
rect 5 -315 15 -310
rect -45 -325 15 -315
rect 205 -315 215 -310
rect 255 -310 335 -275
rect 255 -315 265 -310
rect 205 -325 265 -315
<< labels >>
rlabel nwell -50 205 335 235 1 VDD
rlabel metal4 -50 -310 335 -275 1 GND
rlabel locali 65 -200 95 -180 1 Z1
rlabel locali 160 -115 260 -95 1 Out1
rlabel locali 285 -115 335 -95 1 Out
rlabel locali -50 -115 0 -95 1 A
rlabel metal1 -50 -60 10 -45 1 B
<< end >>
