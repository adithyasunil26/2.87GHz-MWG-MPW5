magic
tech sky130A
timestamp 1640544842
<< nwell >>
rect 75 0 310 455
<< nmos >>
rect 185 -210 200 -60
<< pmos >>
rect 185 40 200 420
<< ndiff >>
rect 130 -75 185 -60
rect 130 -105 140 -75
rect 170 -105 185 -75
rect 130 -125 185 -105
rect 130 -155 140 -125
rect 170 -155 185 -125
rect 130 -175 185 -155
rect 130 -205 140 -175
rect 170 -205 185 -175
rect 130 -210 185 -205
rect 200 -75 255 -60
rect 200 -105 215 -75
rect 245 -105 255 -75
rect 200 -125 255 -105
rect 200 -155 215 -125
rect 245 -155 255 -125
rect 200 -175 255 -155
rect 200 -205 215 -175
rect 245 -205 255 -175
rect 200 -210 255 -205
<< pdiff >>
rect 130 415 185 420
rect 130 395 140 415
rect 170 395 185 415
rect 130 375 185 395
rect 130 345 140 375
rect 170 345 185 375
rect 130 325 185 345
rect 130 295 140 325
rect 170 295 185 325
rect 130 275 185 295
rect 130 245 140 275
rect 170 245 185 275
rect 130 225 185 245
rect 130 195 140 225
rect 170 195 185 225
rect 130 175 185 195
rect 130 145 140 175
rect 170 145 185 175
rect 130 125 185 145
rect 130 95 140 125
rect 170 95 185 125
rect 130 75 185 95
rect 130 45 140 75
rect 170 45 185 75
rect 130 40 185 45
rect 200 415 255 420
rect 200 395 215 415
rect 245 395 255 415
rect 200 375 255 395
rect 200 345 215 375
rect 245 345 255 375
rect 200 325 255 345
rect 200 295 215 325
rect 245 295 255 325
rect 200 275 255 295
rect 200 245 215 275
rect 245 245 255 275
rect 200 225 255 245
rect 200 195 215 225
rect 245 195 255 225
rect 200 175 255 195
rect 200 145 215 175
rect 245 145 255 175
rect 200 125 255 145
rect 200 95 215 125
rect 245 95 255 125
rect 200 75 255 95
rect 200 45 215 75
rect 245 45 255 75
rect 200 40 255 45
<< ndiffc >>
rect 140 -105 170 -75
rect 140 -155 170 -125
rect 140 -205 170 -175
rect 215 -105 245 -75
rect 215 -155 245 -125
rect 215 -205 245 -175
<< pdiffc >>
rect 140 395 170 415
rect 140 345 170 375
rect 140 295 170 325
rect 140 245 170 275
rect 140 195 170 225
rect 140 145 170 175
rect 140 95 170 125
rect 140 45 170 75
rect 215 395 245 415
rect 215 345 245 375
rect 215 295 245 325
rect 215 245 245 275
rect 215 195 245 225
rect 215 145 245 175
rect 215 95 245 125
rect 215 45 245 75
<< poly >>
rect 185 420 200 445
rect 185 0 200 40
rect 150 -10 200 0
rect 150 -30 160 -10
rect 180 -30 200 -10
rect 150 -40 200 -30
rect 185 -60 200 -40
rect 185 -245 200 -210
<< polycont >>
rect 160 -30 180 -10
<< locali >>
rect 140 420 170 490
rect 130 415 180 420
rect 130 395 140 415
rect 170 395 180 415
rect 130 375 180 395
rect 130 345 140 375
rect 170 345 180 375
rect 130 325 180 345
rect 130 295 140 325
rect 170 295 180 325
rect 130 275 180 295
rect 130 245 140 275
rect 170 245 180 275
rect 130 225 180 245
rect 130 195 140 225
rect 170 195 180 225
rect 130 175 180 195
rect 130 145 140 175
rect 170 145 180 175
rect 130 125 180 145
rect 130 95 140 125
rect 170 95 180 125
rect 130 75 180 95
rect 130 45 140 75
rect 170 45 180 75
rect 130 40 180 45
rect 205 415 255 420
rect 205 395 215 415
rect 245 395 255 415
rect 205 375 255 395
rect 205 345 215 375
rect 245 345 255 375
rect 205 325 255 345
rect 205 295 215 325
rect 245 295 255 325
rect 205 275 255 295
rect 205 245 215 275
rect 245 245 255 275
rect 205 225 255 245
rect 205 195 215 225
rect 245 195 255 225
rect 205 175 255 195
rect 205 145 215 175
rect 245 145 255 175
rect 205 125 255 145
rect 205 95 215 125
rect 245 95 255 125
rect 205 75 255 95
rect 205 45 215 75
rect 245 45 255 75
rect 205 40 255 45
rect 150 -10 190 0
rect 75 -30 160 -10
rect 180 -30 190 -10
rect 150 -40 190 -30
rect 225 -10 255 40
rect 225 -30 310 -10
rect 225 -60 255 -30
rect 130 -75 180 -60
rect 130 -105 140 -75
rect 170 -105 180 -75
rect 130 -125 180 -105
rect 130 -155 140 -125
rect 170 -155 180 -125
rect 130 -175 180 -155
rect 130 -205 140 -175
rect 170 -205 180 -175
rect 130 -210 180 -205
rect 205 -75 255 -60
rect 205 -105 215 -75
rect 245 -105 255 -75
rect 205 -125 255 -105
rect 205 -155 215 -125
rect 245 -155 255 -125
rect 205 -175 255 -155
rect 205 -205 215 -175
rect 245 -205 255 -175
rect 205 -210 255 -205
rect 140 -265 170 -210
<< rlocali >>
rect 140 490 170 520
rect 140 -295 170 -265
<< metal1 >>
rect 75 490 315 520
rect 75 -295 310 -265
<< labels >>
rlabel metal1 75 -295 310 -265 1 GND
rlabel locali 75 -30 180 -10 1 IN
rlabel locali 225 -30 310 -10 1 OUT
rlabel metal1 75 490 315 520 1 VDD
<< end >>
