magic
tech sky130A
timestamp 1640956963
<< nwell >>
rect -70 -35 670 465
<< nmos >>
rect -20 -340 -5 -295
rect 105 -340 120 -160
rect 230 -340 245 -160
rect 355 -340 370 -240
rect 480 -340 495 -240
rect 605 -340 620 -140
<< pmos >>
rect 10 -10 25 270
rect 150 -10 165 270
rect 290 -10 305 280
rect 430 -10 445 140
rect 565 -10 580 390
<< ndiff >>
rect 65 -170 105 -160
rect 65 -195 70 -170
rect 95 -195 105 -170
rect 65 -215 105 -195
rect 65 -240 70 -215
rect 95 -240 105 -215
rect 65 -260 105 -240
rect 65 -285 70 -260
rect 95 -285 105 -260
rect -60 -305 -20 -295
rect -60 -330 -55 -305
rect -30 -330 -20 -305
rect -60 -340 -20 -330
rect -5 -305 35 -295
rect -5 -330 5 -305
rect 30 -330 35 -305
rect -5 -340 35 -330
rect 65 -305 105 -285
rect 65 -330 70 -305
rect 95 -330 105 -305
rect 65 -340 105 -330
rect 120 -170 160 -160
rect 120 -195 130 -170
rect 155 -195 160 -170
rect 120 -215 160 -195
rect 120 -240 130 -215
rect 155 -240 160 -215
rect 120 -260 160 -240
rect 120 -285 130 -260
rect 155 -285 160 -260
rect 120 -305 160 -285
rect 120 -330 130 -305
rect 155 -330 160 -305
rect 120 -340 160 -330
rect 190 -170 230 -160
rect 190 -195 195 -170
rect 220 -195 230 -170
rect 190 -215 230 -195
rect 190 -240 195 -215
rect 220 -240 230 -215
rect 190 -260 230 -240
rect 190 -285 195 -260
rect 220 -285 230 -260
rect 190 -305 230 -285
rect 190 -330 195 -305
rect 220 -330 230 -305
rect 190 -340 230 -330
rect 245 -170 285 -160
rect 245 -195 255 -170
rect 280 -195 285 -170
rect 245 -215 285 -195
rect 245 -240 255 -215
rect 280 -240 285 -215
rect 565 -170 605 -140
rect 565 -195 570 -170
rect 595 -195 605 -170
rect 565 -215 605 -195
rect 565 -240 570 -215
rect 595 -240 605 -215
rect 245 -260 285 -240
rect 245 -285 255 -260
rect 280 -285 285 -260
rect 245 -305 285 -285
rect 245 -330 255 -305
rect 280 -330 285 -305
rect 245 -340 285 -330
rect 315 -260 355 -240
rect 315 -285 320 -260
rect 345 -285 355 -260
rect 315 -305 355 -285
rect 315 -330 320 -305
rect 345 -330 355 -305
rect 315 -340 355 -330
rect 370 -260 410 -240
rect 370 -285 380 -260
rect 405 -285 410 -260
rect 370 -305 410 -285
rect 370 -330 380 -305
rect 405 -330 410 -305
rect 370 -340 410 -330
rect 440 -260 480 -240
rect 440 -285 445 -260
rect 470 -285 480 -260
rect 440 -305 480 -285
rect 440 -330 445 -305
rect 470 -330 480 -305
rect 440 -340 480 -330
rect 495 -260 535 -240
rect 495 -285 505 -260
rect 530 -285 535 -260
rect 495 -305 535 -285
rect 495 -330 505 -305
rect 530 -330 535 -305
rect 495 -340 535 -330
rect 565 -260 605 -240
rect 565 -285 570 -260
rect 595 -285 605 -260
rect 565 -305 605 -285
rect 565 -330 570 -305
rect 595 -330 605 -305
rect 565 -340 605 -330
rect 620 -170 660 -140
rect 620 -195 630 -170
rect 655 -195 660 -170
rect 620 -215 660 -195
rect 620 -240 630 -215
rect 655 -240 660 -215
rect 620 -260 660 -240
rect 620 -285 630 -260
rect 655 -285 660 -260
rect 620 -305 660 -285
rect 620 -330 630 -305
rect 655 -330 660 -305
rect 620 -340 660 -330
<< pdiff >>
rect 525 380 565 390
rect 525 360 530 380
rect 555 360 565 380
rect 525 340 565 360
rect 525 315 530 340
rect 555 315 565 340
rect 525 295 565 315
rect -30 250 10 270
rect -30 225 -25 250
rect 0 225 10 250
rect -30 205 10 225
rect -30 180 -25 205
rect 0 180 10 205
rect -30 160 10 180
rect -30 135 -25 160
rect 0 135 10 160
rect -30 115 10 135
rect -30 90 -25 115
rect 0 90 10 115
rect -30 70 10 90
rect -30 45 -25 70
rect 0 45 10 70
rect -30 25 10 45
rect -30 0 -25 25
rect 0 0 10 25
rect -30 -10 10 0
rect 25 250 65 270
rect 25 225 35 250
rect 60 225 65 250
rect 25 205 65 225
rect 25 180 35 205
rect 60 180 65 205
rect 25 160 65 180
rect 25 135 35 160
rect 60 135 65 160
rect 25 115 65 135
rect 25 90 35 115
rect 60 90 65 115
rect 25 70 65 90
rect 25 45 35 70
rect 60 45 65 70
rect 25 25 65 45
rect 25 0 35 25
rect 60 0 65 25
rect 25 -10 65 0
rect 110 250 150 270
rect 110 225 115 250
rect 140 225 150 250
rect 110 205 150 225
rect 110 180 115 205
rect 140 180 150 205
rect 110 160 150 180
rect 110 135 115 160
rect 140 135 150 160
rect 110 115 150 135
rect 110 90 115 115
rect 140 90 150 115
rect 110 70 150 90
rect 110 45 115 70
rect 140 45 150 70
rect 110 25 150 45
rect 110 0 115 25
rect 140 0 150 25
rect 110 -10 150 0
rect 165 250 205 270
rect 165 225 175 250
rect 200 225 205 250
rect 165 205 205 225
rect 165 180 175 205
rect 200 180 205 205
rect 165 160 205 180
rect 165 135 175 160
rect 200 135 205 160
rect 165 115 205 135
rect 165 90 175 115
rect 200 90 205 115
rect 165 70 205 90
rect 165 45 175 70
rect 200 45 205 70
rect 165 25 205 45
rect 165 0 175 25
rect 200 0 205 25
rect 165 -10 205 0
rect 250 250 290 280
rect 250 225 255 250
rect 280 225 290 250
rect 250 205 290 225
rect 250 180 255 205
rect 280 180 290 205
rect 250 160 290 180
rect 250 135 255 160
rect 280 135 290 160
rect 250 115 290 135
rect 250 90 255 115
rect 280 90 290 115
rect 250 70 290 90
rect 250 45 255 70
rect 280 45 290 70
rect 250 25 290 45
rect 250 0 255 25
rect 280 0 290 25
rect 250 -10 290 0
rect 305 250 345 280
rect 305 225 315 250
rect 340 225 345 250
rect 305 205 345 225
rect 305 180 315 205
rect 340 180 345 205
rect 305 160 345 180
rect 525 270 530 295
rect 555 270 565 295
rect 525 250 565 270
rect 525 225 530 250
rect 555 225 565 250
rect 525 205 565 225
rect 525 180 530 205
rect 555 180 565 205
rect 525 160 565 180
rect 305 135 315 160
rect 340 135 345 160
rect 305 115 345 135
rect 305 90 315 115
rect 340 90 345 115
rect 305 70 345 90
rect 305 45 315 70
rect 340 45 345 70
rect 305 25 345 45
rect 305 0 315 25
rect 340 0 345 25
rect 305 -10 345 0
rect 390 115 430 140
rect 390 90 395 115
rect 420 90 430 115
rect 390 70 430 90
rect 390 45 395 70
rect 420 45 430 70
rect 390 25 430 45
rect 390 0 395 25
rect 420 0 430 25
rect 390 -10 430 0
rect 445 115 485 140
rect 445 90 455 115
rect 480 90 485 115
rect 445 70 485 90
rect 445 45 455 70
rect 480 45 485 70
rect 445 25 485 45
rect 445 0 455 25
rect 480 0 485 25
rect 445 -10 485 0
rect 525 135 530 160
rect 555 135 565 160
rect 525 115 565 135
rect 525 90 530 115
rect 555 90 565 115
rect 525 70 565 90
rect 525 45 530 70
rect 555 45 565 70
rect 525 25 565 45
rect 525 0 530 25
rect 555 0 565 25
rect 525 -10 565 0
rect 580 380 620 390
rect 580 360 590 380
rect 615 360 620 380
rect 580 340 620 360
rect 580 315 590 340
rect 615 315 620 340
rect 580 295 620 315
rect 580 270 590 295
rect 615 270 620 295
rect 580 250 620 270
rect 580 225 590 250
rect 615 225 620 250
rect 580 205 620 225
rect 580 180 590 205
rect 615 180 620 205
rect 580 160 620 180
rect 580 135 590 160
rect 615 135 620 160
rect 580 115 620 135
rect 580 90 590 115
rect 615 90 620 115
rect 580 70 620 90
rect 580 45 590 70
rect 615 45 620 70
rect 580 25 620 45
rect 580 0 590 25
rect 615 0 620 25
rect 580 -10 620 0
<< ndiffc >>
rect 70 -195 95 -170
rect 70 -240 95 -215
rect 70 -285 95 -260
rect -55 -330 -30 -305
rect 5 -330 30 -305
rect 70 -330 95 -305
rect 130 -195 155 -170
rect 130 -240 155 -215
rect 130 -285 155 -260
rect 130 -330 155 -305
rect 195 -195 220 -170
rect 195 -240 220 -215
rect 195 -285 220 -260
rect 195 -330 220 -305
rect 255 -195 280 -170
rect 255 -240 280 -215
rect 570 -195 595 -170
rect 570 -240 595 -215
rect 255 -285 280 -260
rect 255 -330 280 -305
rect 320 -285 345 -260
rect 320 -330 345 -305
rect 380 -285 405 -260
rect 380 -330 405 -305
rect 445 -285 470 -260
rect 445 -330 470 -305
rect 505 -285 530 -260
rect 505 -330 530 -305
rect 570 -285 595 -260
rect 570 -330 595 -305
rect 630 -195 655 -170
rect 630 -240 655 -215
rect 630 -285 655 -260
rect 630 -330 655 -305
<< pdiffc >>
rect 530 360 555 380
rect 530 315 555 340
rect -25 225 0 250
rect -25 180 0 205
rect -25 135 0 160
rect -25 90 0 115
rect -25 45 0 70
rect -25 0 0 25
rect 35 225 60 250
rect 35 180 60 205
rect 35 135 60 160
rect 35 90 60 115
rect 35 45 60 70
rect 35 0 60 25
rect 115 225 140 250
rect 115 180 140 205
rect 115 135 140 160
rect 115 90 140 115
rect 115 45 140 70
rect 115 0 140 25
rect 175 225 200 250
rect 175 180 200 205
rect 175 135 200 160
rect 175 90 200 115
rect 175 45 200 70
rect 175 0 200 25
rect 255 225 280 250
rect 255 180 280 205
rect 255 135 280 160
rect 255 90 280 115
rect 255 45 280 70
rect 255 0 280 25
rect 315 225 340 250
rect 315 180 340 205
rect 530 270 555 295
rect 530 225 555 250
rect 530 180 555 205
rect 315 135 340 160
rect 315 90 340 115
rect 315 45 340 70
rect 315 0 340 25
rect 395 90 420 115
rect 395 45 420 70
rect 395 0 420 25
rect 455 90 480 115
rect 455 45 480 70
rect 455 0 480 25
rect 530 135 555 160
rect 530 90 555 115
rect 530 45 555 70
rect 530 0 555 25
rect 590 360 615 380
rect 590 315 615 340
rect 590 270 615 295
rect 590 225 615 250
rect 590 180 615 205
rect 590 135 615 160
rect 590 90 615 115
rect 590 45 615 70
rect 590 0 615 25
<< poly >>
rect 565 390 580 410
rect 10 270 25 290
rect 150 270 165 290
rect 290 280 305 295
rect 430 140 445 160
rect 10 -35 25 -10
rect 150 -35 165 -10
rect 290 -20 305 -10
rect 240 -35 305 -20
rect 430 -35 445 -10
rect 565 -35 580 -10
rect 10 -45 50 -35
rect 10 -65 20 -45
rect 40 -65 50 -45
rect 10 -75 50 -65
rect 150 -45 190 -35
rect 150 -65 160 -45
rect 180 -65 190 -45
rect 150 -75 190 -65
rect 240 -90 255 -35
rect 430 -45 470 -35
rect 430 -65 440 -45
rect 460 -65 470 -45
rect 430 -75 470 -65
rect 540 -45 580 -35
rect 540 -65 550 -45
rect 570 -65 580 -45
rect 540 -75 580 -65
rect 230 -100 270 -90
rect 230 -120 240 -100
rect 260 -120 270 -100
rect 555 -105 570 -75
rect 555 -120 620 -105
rect 230 -130 270 -120
rect 105 -160 120 -140
rect 230 -160 245 -130
rect 355 -145 395 -135
rect 605 -140 620 -120
rect -20 -235 20 -225
rect -20 -255 -10 -235
rect 10 -255 20 -235
rect -20 -265 20 -255
rect -20 -295 -5 -265
rect 355 -165 365 -145
rect 385 -165 395 -145
rect 355 -175 395 -165
rect 355 -240 370 -175
rect 480 -185 520 -175
rect 480 -205 490 -185
rect 510 -205 520 -185
rect 480 -215 520 -205
rect 480 -240 495 -215
rect -20 -360 -5 -340
rect 105 -360 120 -340
rect 230 -360 245 -340
rect 355 -360 370 -340
rect 480 -360 495 -340
rect 605 -360 620 -340
rect 105 -370 145 -360
rect 105 -390 115 -370
rect 135 -390 145 -370
rect 105 -400 145 -390
<< polycont >>
rect 20 -65 40 -45
rect 160 -65 180 -45
rect 440 -65 460 -45
rect 550 -65 570 -45
rect 240 -120 260 -100
rect -10 -255 10 -235
rect 365 -165 385 -145
rect 490 -205 510 -185
rect 115 -390 135 -370
<< locali >>
rect 525 390 550 400
rect 525 380 560 390
rect -25 270 0 360
rect 175 300 180 320
rect 175 270 200 300
rect 255 280 280 360
rect -30 250 5 270
rect -30 225 -25 250
rect 0 225 5 250
rect -30 205 5 225
rect -30 180 -25 205
rect 0 180 5 205
rect -30 160 5 180
rect -30 135 -25 160
rect 0 135 5 160
rect -30 115 5 135
rect -30 90 -25 115
rect 0 90 5 115
rect -30 70 5 90
rect -30 45 -25 70
rect 0 45 5 70
rect -30 25 5 45
rect -30 0 -25 25
rect 0 0 5 25
rect -30 -10 5 0
rect 30 250 65 270
rect 30 225 35 250
rect 60 225 65 250
rect 30 205 65 225
rect 30 180 35 205
rect 60 180 65 205
rect 30 160 65 180
rect 30 135 35 160
rect 60 135 65 160
rect 30 115 65 135
rect 110 250 145 270
rect 110 225 115 250
rect 140 225 145 250
rect 110 205 145 225
rect 110 180 115 205
rect 140 180 145 205
rect 110 160 145 180
rect 110 135 115 160
rect 140 135 145 160
rect 110 115 145 135
rect 30 90 35 115
rect 60 90 115 115
rect 140 90 145 115
rect 30 70 65 90
rect 30 45 35 70
rect 60 45 65 70
rect 30 25 65 45
rect 30 0 35 25
rect 60 0 65 25
rect 30 -10 65 0
rect 110 70 145 90
rect 110 45 115 70
rect 140 45 145 70
rect 110 25 145 45
rect 110 0 115 25
rect 140 0 145 25
rect 110 -10 145 0
rect 170 250 205 270
rect 170 225 175 250
rect 200 225 205 250
rect 170 205 205 225
rect 170 180 175 205
rect 200 180 205 205
rect 170 160 205 180
rect 170 135 175 160
rect 200 135 205 160
rect 170 115 205 135
rect 170 90 175 115
rect 200 90 205 115
rect 170 70 205 90
rect 170 45 175 70
rect 200 45 205 70
rect 170 25 205 45
rect 170 0 175 25
rect 200 0 205 25
rect 170 -10 205 0
rect 250 250 285 280
rect 250 225 255 250
rect 280 225 285 250
rect 250 205 285 225
rect 250 180 255 205
rect 280 180 285 205
rect 250 160 285 180
rect 250 135 255 160
rect 280 135 285 160
rect 250 115 285 135
rect 250 90 255 115
rect 280 90 285 115
rect 250 70 285 90
rect 250 45 255 70
rect 280 45 285 70
rect 250 25 285 45
rect 250 0 255 25
rect 280 0 285 25
rect 250 -10 285 0
rect 310 250 345 280
rect 310 225 315 250
rect 340 225 345 250
rect 310 205 345 225
rect 310 180 315 205
rect 340 180 345 205
rect 310 160 345 180
rect 310 135 315 160
rect 340 135 345 160
rect 395 140 420 365
rect 525 360 530 380
rect 555 360 560 380
rect 525 340 560 360
rect 525 315 530 340
rect 555 315 560 340
rect 525 295 560 315
rect 525 270 530 295
rect 555 270 560 295
rect 525 250 560 270
rect 525 225 530 250
rect 555 225 560 250
rect 525 205 560 225
rect 455 140 480 185
rect 525 180 530 205
rect 555 180 560 205
rect 525 160 560 180
rect 310 115 345 135
rect 310 90 315 115
rect 340 90 345 115
rect 310 70 345 90
rect 310 45 315 70
rect 340 45 345 70
rect 310 25 345 45
rect 310 0 315 25
rect 340 0 345 25
rect 310 -10 345 0
rect 390 115 425 140
rect 390 90 395 115
rect 420 90 425 115
rect 390 70 425 90
rect 390 45 395 70
rect 420 45 425 70
rect 390 25 425 45
rect 390 0 395 25
rect 420 0 425 25
rect 390 -10 425 0
rect 450 115 485 140
rect 450 90 455 115
rect 480 90 485 115
rect 450 70 485 90
rect 450 45 455 70
rect 480 45 485 70
rect 450 25 485 45
rect 450 0 455 25
rect 480 0 485 25
rect 450 -10 485 0
rect 525 135 530 160
rect 555 135 560 160
rect 525 115 560 135
rect 525 90 530 115
rect 555 90 560 115
rect 525 70 560 90
rect 525 45 530 70
rect 555 45 560 70
rect 525 25 560 45
rect 525 0 530 25
rect 555 0 560 25
rect 525 -10 560 0
rect 585 380 620 390
rect 585 360 590 380
rect 615 360 620 380
rect 585 340 620 360
rect 585 315 590 340
rect 615 315 620 340
rect 585 295 620 315
rect 585 270 590 295
rect 615 270 620 295
rect 585 250 620 270
rect 585 225 590 250
rect 615 225 620 250
rect 585 205 620 225
rect 585 180 590 205
rect 615 180 620 205
rect 585 160 620 180
rect 585 135 590 160
rect 615 135 620 160
rect 585 115 620 135
rect 585 90 590 115
rect 615 90 620 115
rect 585 70 620 90
rect 585 45 590 70
rect 615 45 620 70
rect 585 25 620 45
rect 585 0 590 25
rect 615 0 655 25
rect 585 -10 655 0
rect 10 -45 50 -35
rect -10 -65 20 -45
rect 40 -65 50 -45
rect -10 -75 50 -65
rect 150 -45 190 -35
rect 315 -45 340 -10
rect 430 -45 470 -35
rect 540 -45 580 -35
rect 150 -65 160 -45
rect 180 -65 260 -45
rect 335 -65 440 -45
rect 460 -65 510 -45
rect 150 -75 190 -65
rect -10 -135 10 -75
rect 240 -90 260 -65
rect 430 -75 470 -65
rect 230 -100 270 -90
rect -70 -155 10 -135
rect -10 -225 10 -155
rect 70 -160 95 -125
rect 130 -160 155 -125
rect 230 -120 240 -100
rect 260 -120 385 -100
rect 230 -130 270 -120
rect 355 -135 385 -120
rect 355 -145 395 -135
rect 65 -170 100 -160
rect 65 -195 70 -170
rect 95 -195 100 -170
rect 65 -215 100 -195
rect -20 -235 20 -225
rect -20 -255 -10 -235
rect 10 -255 20 -235
rect -20 -265 20 -255
rect 65 -240 70 -215
rect 95 -240 100 -215
rect 65 -260 100 -240
rect 65 -285 70 -260
rect 95 -285 100 -260
rect -60 -305 -25 -295
rect -60 -330 -55 -305
rect -30 -330 -25 -305
rect -60 -340 -25 -330
rect 0 -305 35 -295
rect 0 -330 5 -305
rect 30 -330 35 -305
rect 0 -340 35 -330
rect 65 -305 100 -285
rect 65 -330 70 -305
rect 95 -330 100 -305
rect 65 -340 100 -330
rect 125 -170 160 -160
rect 125 -195 130 -170
rect 155 -195 160 -170
rect 125 -215 160 -195
rect 125 -240 130 -215
rect 155 -240 160 -215
rect 125 -260 160 -240
rect 125 -285 130 -260
rect 155 -285 160 -260
rect 125 -305 160 -285
rect 125 -330 130 -305
rect 155 -330 160 -305
rect 125 -340 160 -330
rect 190 -170 225 -160
rect 190 -195 195 -170
rect 220 -195 225 -170
rect 190 -215 225 -195
rect 190 -240 195 -215
rect 220 -240 225 -215
rect 190 -260 225 -240
rect 190 -285 195 -260
rect 220 -285 225 -260
rect 190 -305 225 -285
rect 190 -330 195 -305
rect 220 -330 225 -305
rect 190 -340 225 -330
rect 250 -170 305 -160
rect 250 -195 255 -170
rect 280 -180 305 -170
rect 355 -165 365 -145
rect 385 -165 395 -145
rect 355 -175 395 -165
rect 490 -175 510 -65
rect 540 -65 550 -45
rect 570 -65 580 -45
rect 540 -75 580 -65
rect 550 -80 580 -75
rect 630 -60 655 -10
rect 630 -85 690 -60
rect 630 -140 655 -85
rect 565 -170 600 -140
rect 280 -195 285 -180
rect 250 -215 285 -195
rect 480 -185 520 -175
rect 480 -205 490 -185
rect 510 -205 520 -185
rect 480 -215 520 -205
rect 565 -195 570 -170
rect 595 -195 600 -170
rect 565 -215 600 -195
rect 250 -240 255 -215
rect 280 -240 285 -215
rect 565 -240 570 -215
rect 595 -240 600 -215
rect 250 -260 285 -240
rect 250 -285 255 -260
rect 280 -285 285 -260
rect 250 -305 285 -285
rect 250 -330 255 -305
rect 280 -330 285 -305
rect 250 -340 285 -330
rect 315 -260 350 -240
rect 315 -285 320 -260
rect 345 -285 350 -260
rect 315 -305 350 -285
rect 315 -330 320 -305
rect 345 -330 350 -305
rect 315 -340 350 -330
rect 375 -260 410 -240
rect 375 -285 380 -260
rect 405 -285 410 -260
rect 375 -305 410 -285
rect 375 -330 380 -305
rect 405 -330 410 -305
rect 375 -340 410 -330
rect 440 -260 475 -240
rect 440 -285 445 -260
rect 470 -285 475 -260
rect 440 -305 475 -285
rect 440 -330 445 -305
rect 470 -330 475 -305
rect 440 -340 475 -330
rect 500 -260 535 -240
rect 500 -285 505 -260
rect 530 -285 535 -260
rect 500 -305 535 -285
rect 500 -330 505 -305
rect 530 -330 535 -305
rect 500 -340 535 -330
rect 565 -260 600 -240
rect 565 -285 570 -260
rect 595 -285 600 -260
rect 565 -305 600 -285
rect 565 -330 570 -305
rect 595 -330 600 -305
rect 565 -340 600 -330
rect 625 -170 660 -140
rect 625 -195 630 -170
rect 655 -195 660 -170
rect 625 -215 660 -195
rect 625 -240 630 -215
rect 655 -240 660 -215
rect 625 -260 660 -240
rect 625 -285 630 -260
rect 655 -285 660 -260
rect 625 -305 660 -285
rect 625 -330 630 -305
rect 655 -330 660 -305
rect 625 -340 660 -330
rect -55 -420 -30 -340
rect 5 -370 30 -340
rect 105 -370 145 -360
rect 5 -390 35 -370
rect 55 -390 115 -370
rect 135 -390 145 -370
rect 105 -400 145 -390
rect -35 -440 -30 -420
rect 195 -420 220 -340
rect 320 -375 345 -340
rect 215 -440 220 -420
rect 445 -400 470 -340
rect 505 -375 530 -340
rect 570 -400 595 -340
rect 445 -415 475 -400
rect 445 -435 450 -415
rect 470 -435 475 -415
rect 570 -415 600 -400
rect 570 -435 575 -415
rect 595 -435 600 -415
rect 445 -440 470 -435
rect 570 -440 595 -435
<< viali >>
rect 525 400 545 420
rect -25 360 -5 380
rect 255 360 275 380
rect 395 365 415 385
rect 180 300 200 320
rect 455 185 475 205
rect 160 -65 180 -45
rect 315 -65 335 -45
rect 75 -125 95 -105
rect 135 -125 155 -105
rect 305 -180 325 -160
rect 550 -100 570 -80
rect 385 -240 405 -220
rect 35 -390 55 -370
rect -55 -440 -35 -420
rect 320 -395 340 -375
rect 195 -440 215 -420
rect 510 -395 530 -375
rect 450 -435 470 -415
rect 575 -435 595 -415
<< metal1 >>
rect 515 400 520 430
rect 550 400 555 430
rect 515 395 555 400
rect -35 360 -30 390
rect 0 360 5 390
rect -35 355 5 360
rect 245 360 250 390
rect 280 360 285 390
rect 385 365 390 395
rect 420 365 425 395
rect 385 360 425 365
rect 245 355 285 360
rect 170 320 210 330
rect 35 305 180 320
rect 35 -355 50 305
rect 170 300 180 305
rect 200 300 210 320
rect 170 290 210 300
rect 445 205 510 215
rect 445 185 455 205
rect 475 185 510 205
rect 445 180 510 185
rect 150 -40 190 -35
rect 150 -70 155 -40
rect 185 -70 190 -40
rect 150 -75 190 -70
rect 305 -45 345 -40
rect 305 -65 315 -45
rect 335 -65 345 -45
rect 305 -85 345 -65
rect 305 -95 335 -85
rect 495 -90 510 180
rect 540 -80 575 -70
rect 540 -90 550 -80
rect 65 -105 105 -100
rect 65 -125 75 -105
rect 95 -125 105 -105
rect 65 -135 105 -125
rect 125 -105 335 -95
rect 125 -125 135 -105
rect 155 -110 335 -105
rect 425 -100 550 -90
rect 570 -100 575 -80
rect 425 -105 575 -100
rect 155 -125 165 -110
rect 125 -130 165 -125
rect 75 -205 90 -135
rect 425 -140 440 -105
rect 540 -110 575 -105
rect 425 -155 690 -140
rect 295 -160 335 -155
rect 295 -180 305 -160
rect 325 -180 335 -160
rect 295 -205 335 -180
rect 75 -220 335 -205
rect 425 -210 440 -155
rect 375 -220 440 -210
rect 375 -240 385 -220
rect 405 -225 440 -220
rect 405 -240 420 -225
rect 375 -250 420 -240
rect 25 -370 65 -355
rect 25 -390 35 -370
rect 55 -390 65 -370
rect 25 -395 65 -390
rect 315 -375 350 -365
rect 500 -375 540 -365
rect 315 -395 320 -375
rect 340 -390 510 -375
rect 340 -395 350 -390
rect 315 -405 350 -395
rect 500 -395 510 -390
rect 530 -395 540 -375
rect 500 -405 540 -395
rect 440 -410 480 -405
rect -65 -415 -25 -410
rect -65 -445 -60 -415
rect -30 -445 -25 -415
rect -65 -450 -25 -445
rect 185 -415 225 -410
rect 185 -445 190 -415
rect 220 -445 225 -415
rect 440 -440 445 -410
rect 475 -440 480 -410
rect 440 -445 480 -440
rect 565 -410 605 -405
rect 565 -440 570 -410
rect 600 -440 605 -410
rect 565 -445 605 -440
rect 185 -450 225 -445
<< via1 >>
rect 520 420 550 430
rect 520 400 525 420
rect 525 400 545 420
rect 545 400 550 420
rect -30 380 0 390
rect -30 360 -25 380
rect -25 360 -5 380
rect -5 360 0 380
rect 250 380 280 390
rect 250 360 255 380
rect 255 360 275 380
rect 275 360 280 380
rect 390 385 420 395
rect 390 365 395 385
rect 395 365 415 385
rect 415 365 420 385
rect 155 -45 185 -40
rect 155 -65 160 -45
rect 160 -65 180 -45
rect 180 -65 185 -45
rect 155 -70 185 -65
rect -60 -420 -30 -415
rect -60 -440 -55 -420
rect -55 -440 -35 -420
rect -35 -440 -30 -420
rect -60 -445 -30 -440
rect 190 -420 220 -415
rect 190 -440 195 -420
rect 195 -440 215 -420
rect 215 -440 220 -420
rect 190 -445 220 -440
rect 445 -415 475 -410
rect 445 -435 450 -415
rect 450 -435 470 -415
rect 470 -435 475 -415
rect 445 -440 475 -435
rect 570 -415 600 -410
rect 570 -435 575 -415
rect 575 -435 595 -415
rect 595 -435 600 -415
rect 570 -440 600 -435
<< metal2 >>
rect 510 400 515 435
rect 555 400 560 435
rect -40 360 -35 395
rect 5 360 10 395
rect -40 355 10 360
rect 240 360 245 395
rect 285 360 290 395
rect 380 365 385 400
rect 425 365 430 400
rect 510 395 560 400
rect 380 360 430 365
rect 240 355 290 360
rect 145 -40 195 -30
rect 145 -45 155 -40
rect -70 -65 155 -45
rect 145 -70 155 -65
rect 185 -70 195 -40
rect 145 -80 195 -70
rect 440 -410 480 -405
rect -65 -415 -25 -410
rect -65 -445 -60 -415
rect -30 -445 -25 -415
rect -65 -450 -25 -445
rect 185 -415 225 -410
rect 185 -445 190 -415
rect 220 -445 225 -415
rect 440 -440 445 -410
rect 475 -440 480 -410
rect 440 -445 480 -440
rect 565 -410 605 -405
rect 565 -440 570 -410
rect 600 -440 605 -410
rect 565 -445 605 -440
rect 185 -450 225 -445
<< via2 >>
rect 515 430 555 435
rect 515 400 520 430
rect 520 400 550 430
rect 550 400 555 430
rect -35 390 5 395
rect -35 360 -30 390
rect -30 360 0 390
rect 0 360 5 390
rect 245 390 285 395
rect 245 360 250 390
rect 250 360 280 390
rect 280 360 285 390
rect 385 395 425 400
rect 385 365 390 395
rect 390 365 420 395
rect 420 365 425 395
rect -60 -445 -30 -415
rect 190 -445 220 -415
rect 445 -440 475 -410
rect 570 -440 600 -410
<< metal3 >>
rect 505 435 565 440
rect 375 400 435 405
rect -45 395 15 400
rect -45 355 -40 395
rect 10 355 15 395
rect 235 395 295 400
rect 235 355 240 395
rect 290 355 295 395
rect 375 360 380 400
rect 430 360 435 400
rect 505 395 510 435
rect 560 395 565 435
rect 435 -405 485 -400
rect -70 -410 -20 -405
rect -70 -450 -65 -410
rect -25 -450 -20 -410
rect -70 -455 -20 -450
rect 180 -410 230 -405
rect 180 -450 185 -410
rect 225 -450 230 -410
rect 435 -445 440 -405
rect 480 -445 485 -405
rect 435 -450 485 -445
rect 560 -405 610 -400
rect 560 -445 565 -405
rect 605 -445 610 -405
rect 560 -450 610 -445
rect 180 -455 230 -450
<< via3 >>
rect -40 360 -35 395
rect -35 360 5 395
rect 5 360 10 395
rect -40 355 10 360
rect 240 360 245 395
rect 245 360 285 395
rect 285 360 290 395
rect 240 355 290 360
rect 380 365 385 400
rect 385 365 425 400
rect 425 365 430 400
rect 380 360 430 365
rect 510 400 515 435
rect 515 400 555 435
rect 555 400 560 435
rect 510 395 560 400
rect -65 -415 -25 -410
rect -65 -445 -60 -415
rect -60 -445 -30 -415
rect -30 -445 -25 -415
rect -65 -450 -25 -445
rect 185 -415 225 -410
rect 185 -445 190 -415
rect 190 -445 220 -415
rect 220 -445 225 -415
rect 185 -450 225 -445
rect 440 -410 480 -405
rect 440 -440 445 -410
rect 445 -440 475 -410
rect 475 -440 480 -410
rect 440 -445 480 -440
rect 565 -410 605 -405
rect 565 -440 570 -410
rect 570 -440 600 -410
rect 600 -440 605 -410
rect 565 -445 605 -440
<< metal4 >>
rect -70 435 670 465
rect -25 400 5 435
rect 250 400 280 435
rect 390 405 420 435
rect 375 400 435 405
rect -45 395 15 400
rect -45 355 -40 395
rect 10 355 15 395
rect -45 350 15 355
rect 235 395 295 400
rect 235 355 240 395
rect 290 355 295 395
rect 375 360 380 400
rect 430 360 435 400
rect 505 395 510 435
rect 560 395 565 435
rect 505 390 565 395
rect 375 355 435 360
rect 235 350 295 355
rect 435 -405 485 -400
rect -70 -410 -20 -405
rect -70 -450 -65 -410
rect -25 -450 -20 -410
rect 180 -410 230 -405
rect 180 -450 185 -410
rect 225 -450 230 -410
rect 435 -445 440 -405
rect 480 -445 485 -405
rect 435 -450 485 -445
rect 560 -405 610 -400
rect 560 -445 565 -405
rect 605 -445 610 -405
rect 560 -450 610 -445
rect -70 -455 660 -450
rect -60 -490 660 -455
<< labels >>
rlabel locali -10 -255 10 -45 1 D
rlabel locali -10 -65 40 -45 1 D
rlabel locali 65 90 110 115 1 Z1
rlabel metal1 130 -110 335 -95 1 Z3
rlabel locali 490 -205 510 -45 1 Z3
rlabel metal1 75 -220 330 -205 1 Z4
rlabel space 320 -405 530 -390 1 Z5
rlabel locali 630 -85 690 -60 1 Q
rlabel space 425 -105 580 -90 1 Qbar
rlabel locali 315 -65 510 -45 1 Z3
rlabel locali 5 -390 135 -370 1 Z2
rlabel space 70 -160 95 -95 1 Z4
rlabel space 285 -180 335 -160 1 Z4
rlabel metal4 -55 -470 660 -455 1 GND
rlabel locali 269 336 269 336 1 vdd!
rlabel locali 202 -379 202 -379 1 gnd!
<< end >>
