magic
tech sky130A
timestamp 1640737585
<< nwell >>
rect -80 125 450 1955
<< nmos >>
rect 0 -10 15 40
rect 175 -160 190 40
rect 355 -160 370 40
<< pmos >>
rect 0 145 15 245
rect 175 145 190 545
rect 355 145 370 1745
<< ndiff >>
rect -55 30 0 40
rect -55 5 -40 30
rect -15 5 0 30
rect -55 -10 0 5
rect 15 30 70 40
rect 15 5 30 30
rect 55 5 70 30
rect 15 -10 70 5
rect 120 30 175 40
rect 120 5 135 30
rect 160 5 175 30
rect 120 -20 175 5
rect 120 -45 135 -20
rect 160 -45 175 -20
rect 120 -70 175 -45
rect 120 -95 135 -70
rect 160 -95 175 -70
rect 120 -120 175 -95
rect 120 -145 135 -120
rect 160 -145 175 -120
rect 120 -160 175 -145
rect 190 30 245 40
rect 190 5 205 30
rect 230 5 245 30
rect 190 -20 245 5
rect 190 -45 205 -20
rect 230 -45 245 -20
rect 190 -70 245 -45
rect 190 -95 205 -70
rect 230 -95 245 -70
rect 190 -120 245 -95
rect 190 -145 205 -120
rect 230 -145 245 -120
rect 190 -160 245 -145
rect 300 30 355 40
rect 300 5 315 30
rect 340 5 355 30
rect 300 -20 355 5
rect 300 -45 315 -20
rect 340 -45 355 -20
rect 300 -70 355 -45
rect 300 -95 315 -70
rect 340 -95 355 -70
rect 300 -120 355 -95
rect 300 -145 315 -120
rect 340 -145 355 -120
rect 300 -160 355 -145
rect 370 30 425 40
rect 370 5 385 30
rect 410 5 425 30
rect 370 -20 425 5
rect 370 -45 385 -20
rect 410 -45 425 -20
rect 370 -70 425 -45
rect 370 -95 385 -70
rect 410 -95 425 -70
rect 370 -120 425 -95
rect 370 -145 385 -120
rect 410 -145 425 -120
rect 370 -160 425 -145
<< pdiff >>
rect 300 1730 355 1745
rect 300 1705 315 1730
rect 340 1705 355 1730
rect 300 1685 355 1705
rect 300 1660 315 1685
rect 340 1660 355 1685
rect 300 1630 355 1660
rect 300 1605 315 1630
rect 340 1605 355 1630
rect 300 1585 355 1605
rect 300 1560 315 1585
rect 340 1560 355 1585
rect 300 1530 355 1560
rect 300 1505 315 1530
rect 340 1505 355 1530
rect 300 1485 355 1505
rect 300 1460 315 1485
rect 340 1460 355 1485
rect 300 1430 355 1460
rect 300 1405 315 1430
rect 340 1405 355 1430
rect 300 1385 355 1405
rect 300 1360 315 1385
rect 340 1360 355 1385
rect 300 1330 355 1360
rect 300 1305 315 1330
rect 340 1305 355 1330
rect 300 1285 355 1305
rect 300 1260 315 1285
rect 340 1260 355 1285
rect 300 1230 355 1260
rect 300 1205 315 1230
rect 340 1205 355 1230
rect 300 1185 355 1205
rect 300 1160 315 1185
rect 340 1160 355 1185
rect 300 1130 355 1160
rect 300 1105 315 1130
rect 340 1105 355 1130
rect 300 1085 355 1105
rect 300 1060 315 1085
rect 340 1060 355 1085
rect 300 1030 355 1060
rect 300 1005 315 1030
rect 340 1005 355 1030
rect 300 985 355 1005
rect 300 960 315 985
rect 340 960 355 985
rect 300 930 355 960
rect 300 905 315 930
rect 340 905 355 930
rect 300 885 355 905
rect 300 860 315 885
rect 340 860 355 885
rect 300 830 355 860
rect 300 805 315 830
rect 340 805 355 830
rect 300 785 355 805
rect 300 760 315 785
rect 340 760 355 785
rect 300 730 355 760
rect 300 705 315 730
rect 340 705 355 730
rect 300 685 355 705
rect 300 660 315 685
rect 340 660 355 685
rect 300 630 355 660
rect 300 605 315 630
rect 340 605 355 630
rect 300 585 355 605
rect 300 560 315 585
rect 340 560 355 585
rect 120 530 175 545
rect 120 505 135 530
rect 160 505 175 530
rect 120 485 175 505
rect 120 460 135 485
rect 160 460 175 485
rect 120 430 175 460
rect 120 405 135 430
rect 160 405 175 430
rect 120 385 175 405
rect 120 360 135 385
rect 160 360 175 385
rect 120 330 175 360
rect 120 305 135 330
rect 160 305 175 330
rect 120 285 175 305
rect 120 260 135 285
rect 160 260 175 285
rect -55 230 0 245
rect -55 205 -40 230
rect -15 205 0 230
rect -55 185 0 205
rect -55 160 -40 185
rect -15 160 0 185
rect -55 145 0 160
rect 15 230 70 245
rect 15 205 30 230
rect 55 205 70 230
rect 15 185 70 205
rect 15 160 30 185
rect 55 160 70 185
rect 15 145 70 160
rect 120 230 175 260
rect 120 205 135 230
rect 160 205 175 230
rect 120 185 175 205
rect 120 160 135 185
rect 160 160 175 185
rect 120 145 175 160
rect 190 530 245 545
rect 190 505 205 530
rect 230 505 245 530
rect 190 485 245 505
rect 190 460 205 485
rect 230 460 245 485
rect 190 430 245 460
rect 190 405 205 430
rect 230 405 245 430
rect 190 385 245 405
rect 190 360 205 385
rect 230 360 245 385
rect 190 330 245 360
rect 190 305 205 330
rect 230 305 245 330
rect 190 285 245 305
rect 190 260 205 285
rect 230 260 245 285
rect 190 230 245 260
rect 190 205 205 230
rect 230 205 245 230
rect 190 185 245 205
rect 190 160 205 185
rect 230 160 245 185
rect 190 145 245 160
rect 300 530 355 560
rect 300 505 315 530
rect 340 505 355 530
rect 300 485 355 505
rect 300 460 315 485
rect 340 460 355 485
rect 300 430 355 460
rect 300 405 315 430
rect 340 405 355 430
rect 300 385 355 405
rect 300 360 315 385
rect 340 360 355 385
rect 300 330 355 360
rect 300 305 315 330
rect 340 305 355 330
rect 300 285 355 305
rect 300 260 315 285
rect 340 260 355 285
rect 300 230 355 260
rect 300 205 315 230
rect 340 205 355 230
rect 300 185 355 205
rect 300 160 315 185
rect 340 160 355 185
rect 300 145 355 160
rect 370 1730 425 1745
rect 370 1705 385 1730
rect 410 1705 425 1730
rect 370 1685 425 1705
rect 370 1660 385 1685
rect 410 1660 425 1685
rect 370 1630 425 1660
rect 370 1605 385 1630
rect 410 1605 425 1630
rect 370 1585 425 1605
rect 370 1560 385 1585
rect 410 1560 425 1585
rect 370 1530 425 1560
rect 370 1505 385 1530
rect 410 1505 425 1530
rect 370 1485 425 1505
rect 370 1460 385 1485
rect 410 1460 425 1485
rect 370 1430 425 1460
rect 370 1405 385 1430
rect 410 1405 425 1430
rect 370 1385 425 1405
rect 370 1360 385 1385
rect 410 1360 425 1385
rect 370 1330 425 1360
rect 370 1305 385 1330
rect 410 1305 425 1330
rect 370 1285 425 1305
rect 370 1260 385 1285
rect 410 1260 425 1285
rect 370 1230 425 1260
rect 370 1205 385 1230
rect 410 1205 425 1230
rect 370 1185 425 1205
rect 370 1160 385 1185
rect 410 1160 425 1185
rect 370 1130 425 1160
rect 370 1105 385 1130
rect 410 1105 425 1130
rect 370 1085 425 1105
rect 370 1060 385 1085
rect 410 1060 425 1085
rect 370 1030 425 1060
rect 370 1005 385 1030
rect 410 1005 425 1030
rect 370 985 425 1005
rect 370 960 385 985
rect 410 960 425 985
rect 370 930 425 960
rect 370 905 385 930
rect 410 905 425 930
rect 370 885 425 905
rect 370 860 385 885
rect 410 860 425 885
rect 370 830 425 860
rect 370 805 385 830
rect 410 805 425 830
rect 370 785 425 805
rect 370 760 385 785
rect 410 760 425 785
rect 370 730 425 760
rect 370 705 385 730
rect 410 705 425 730
rect 370 685 425 705
rect 370 660 385 685
rect 410 660 425 685
rect 370 630 425 660
rect 370 605 385 630
rect 410 605 425 630
rect 370 585 425 605
rect 370 560 385 585
rect 410 560 425 585
rect 370 530 425 560
rect 370 505 385 530
rect 410 505 425 530
rect 370 485 425 505
rect 370 460 385 485
rect 410 460 425 485
rect 370 430 425 460
rect 370 405 385 430
rect 410 405 425 430
rect 370 385 425 405
rect 370 360 385 385
rect 410 360 425 385
rect 370 330 425 360
rect 370 305 385 330
rect 410 305 425 330
rect 370 285 425 305
rect 370 260 385 285
rect 410 260 425 285
rect 370 230 425 260
rect 370 205 385 230
rect 410 205 425 230
rect 370 185 425 205
rect 370 160 385 185
rect 410 160 425 185
rect 370 145 425 160
<< ndiffc >>
rect -40 5 -15 30
rect 30 5 55 30
rect 135 5 160 30
rect 135 -45 160 -20
rect 135 -95 160 -70
rect 135 -145 160 -120
rect 205 5 230 30
rect 205 -45 230 -20
rect 205 -95 230 -70
rect 205 -145 230 -120
rect 315 5 340 30
rect 315 -45 340 -20
rect 315 -95 340 -70
rect 315 -145 340 -120
rect 385 5 410 30
rect 385 -45 410 -20
rect 385 -95 410 -70
rect 385 -145 410 -120
<< pdiffc >>
rect 315 1705 340 1730
rect 315 1660 340 1685
rect 315 1605 340 1630
rect 315 1560 340 1585
rect 315 1505 340 1530
rect 315 1460 340 1485
rect 315 1405 340 1430
rect 315 1360 340 1385
rect 315 1305 340 1330
rect 315 1260 340 1285
rect 315 1205 340 1230
rect 315 1160 340 1185
rect 315 1105 340 1130
rect 315 1060 340 1085
rect 315 1005 340 1030
rect 315 960 340 985
rect 315 905 340 930
rect 315 860 340 885
rect 315 805 340 830
rect 315 760 340 785
rect 315 705 340 730
rect 315 660 340 685
rect 315 605 340 630
rect 315 560 340 585
rect 135 505 160 530
rect 135 460 160 485
rect 135 405 160 430
rect 135 360 160 385
rect 135 305 160 330
rect 135 260 160 285
rect -40 205 -15 230
rect -40 160 -15 185
rect 30 205 55 230
rect 30 160 55 185
rect 135 205 160 230
rect 135 160 160 185
rect 205 505 230 530
rect 205 460 230 485
rect 205 405 230 430
rect 205 360 230 385
rect 205 305 230 330
rect 205 260 230 285
rect 205 205 230 230
rect 205 160 230 185
rect 315 505 340 530
rect 315 460 340 485
rect 315 405 340 430
rect 315 360 340 385
rect 315 305 340 330
rect 315 260 340 285
rect 315 205 340 230
rect 315 160 340 185
rect 385 1705 410 1730
rect 385 1660 410 1685
rect 385 1605 410 1630
rect 385 1560 410 1585
rect 385 1505 410 1530
rect 385 1460 410 1485
rect 385 1405 410 1430
rect 385 1360 410 1385
rect 385 1305 410 1330
rect 385 1260 410 1285
rect 385 1205 410 1230
rect 385 1160 410 1185
rect 385 1105 410 1130
rect 385 1060 410 1085
rect 385 1005 410 1030
rect 385 960 410 985
rect 385 905 410 930
rect 385 860 410 885
rect 385 805 410 830
rect 385 760 410 785
rect 385 705 410 730
rect 385 660 410 685
rect 385 605 410 630
rect 385 560 410 585
rect 385 505 410 530
rect 385 460 410 485
rect 385 405 410 430
rect 385 360 410 385
rect 385 305 410 330
rect 385 260 410 285
rect 385 205 410 230
rect 385 160 410 185
<< poly >>
rect 355 1745 370 1760
rect 175 545 190 560
rect 0 245 15 260
rect 0 110 15 145
rect 175 110 190 145
rect 355 110 370 145
rect -50 100 15 110
rect -50 70 -40 100
rect -10 70 15 100
rect -50 60 15 70
rect 125 100 190 110
rect 125 70 135 100
rect 165 70 190 100
rect 125 60 190 70
rect 305 100 370 110
rect 305 70 315 100
rect 345 70 370 100
rect 305 60 370 70
rect 0 40 15 60
rect 175 40 190 60
rect 355 40 370 60
rect 0 -30 15 -10
rect 175 -180 190 -160
rect 355 -180 370 -160
<< polycont >>
rect -40 70 -10 100
rect 135 70 165 100
rect 315 70 345 100
<< locali >>
rect -60 1935 10 1945
rect -60 1885 -50 1935
rect 0 1885 10 1935
rect -60 1875 10 1885
rect 115 1935 185 1945
rect 115 1885 125 1935
rect 175 1885 185 1935
rect 115 1875 185 1885
rect 295 1935 365 1945
rect 295 1885 305 1935
rect 355 1885 365 1935
rect 295 1875 365 1885
rect -50 230 -5 1875
rect 125 530 170 1875
rect 305 1730 350 1875
rect 305 1705 315 1730
rect 340 1705 350 1730
rect 305 1685 350 1705
rect 305 1660 315 1685
rect 340 1660 350 1685
rect 305 1630 350 1660
rect 305 1605 315 1630
rect 340 1605 350 1630
rect 305 1585 350 1605
rect 305 1560 315 1585
rect 340 1560 350 1585
rect 305 1530 350 1560
rect 305 1505 315 1530
rect 340 1505 350 1530
rect 305 1485 350 1505
rect 305 1460 315 1485
rect 340 1460 350 1485
rect 305 1430 350 1460
rect 305 1405 315 1430
rect 340 1405 350 1430
rect 305 1385 350 1405
rect 305 1360 315 1385
rect 340 1360 350 1385
rect 305 1330 350 1360
rect 305 1305 315 1330
rect 340 1305 350 1330
rect 305 1285 350 1305
rect 305 1260 315 1285
rect 340 1260 350 1285
rect 305 1230 350 1260
rect 305 1205 315 1230
rect 340 1205 350 1230
rect 305 1185 350 1205
rect 305 1160 315 1185
rect 340 1160 350 1185
rect 305 1130 350 1160
rect 305 1105 315 1130
rect 340 1105 350 1130
rect 305 1085 350 1105
rect 305 1060 315 1085
rect 340 1060 350 1085
rect 305 1030 350 1060
rect 305 1005 315 1030
rect 340 1005 350 1030
rect 305 985 350 1005
rect 305 960 315 985
rect 340 960 350 985
rect 305 930 350 960
rect 305 905 315 930
rect 340 905 350 930
rect 305 885 350 905
rect 305 860 315 885
rect 340 860 350 885
rect 305 830 350 860
rect 305 805 315 830
rect 340 805 350 830
rect 305 785 350 805
rect 305 760 315 785
rect 340 760 350 785
rect 305 730 350 760
rect 305 705 315 730
rect 340 705 350 730
rect 305 685 350 705
rect 305 660 315 685
rect 340 660 350 685
rect 305 630 350 660
rect 305 605 315 630
rect 340 605 350 630
rect 305 585 350 605
rect 305 560 315 585
rect 340 560 350 585
rect 125 505 135 530
rect 160 505 170 530
rect 125 485 170 505
rect 125 460 135 485
rect 160 460 170 485
rect 125 430 170 460
rect 125 405 135 430
rect 160 405 170 430
rect 125 385 170 405
rect 125 360 135 385
rect 160 360 170 385
rect 125 330 170 360
rect 125 305 135 330
rect 160 305 170 330
rect 125 285 170 305
rect 125 260 135 285
rect 160 260 170 285
rect -50 205 -40 230
rect -15 205 -5 230
rect -50 185 -5 205
rect -50 160 -40 185
rect -15 160 -5 185
rect -50 150 -5 160
rect 20 230 65 240
rect 20 205 30 230
rect 55 205 65 230
rect 20 185 65 205
rect 20 160 30 185
rect 55 160 65 185
rect -50 100 0 110
rect -50 70 -40 100
rect -10 70 0 100
rect -50 60 0 70
rect -50 30 -5 40
rect -50 5 -40 30
rect -15 5 -5 30
rect -50 -1170 -5 5
rect 20 30 65 160
rect 125 230 170 260
rect 125 205 135 230
rect 160 205 170 230
rect 125 185 170 205
rect 125 160 135 185
rect 160 160 170 185
rect 125 150 170 160
rect 195 530 240 540
rect 195 505 205 530
rect 230 505 240 530
rect 195 485 240 505
rect 195 460 205 485
rect 230 460 240 485
rect 195 430 240 460
rect 195 405 205 430
rect 230 405 240 430
rect 195 385 240 405
rect 195 360 205 385
rect 230 360 240 385
rect 195 330 240 360
rect 195 305 205 330
rect 230 305 240 330
rect 195 285 240 305
rect 195 260 205 285
rect 230 260 240 285
rect 195 230 240 260
rect 195 205 205 230
rect 230 205 240 230
rect 195 185 240 205
rect 195 160 205 185
rect 230 160 240 185
rect 125 100 175 110
rect 125 70 135 100
rect 165 70 175 100
rect 125 60 175 70
rect 20 5 30 30
rect 55 5 65 30
rect 20 -5 65 5
rect 125 30 170 40
rect 125 5 135 30
rect 160 5 170 30
rect 125 -20 170 5
rect 125 -45 135 -20
rect 160 -45 170 -20
rect 125 -70 170 -45
rect 125 -95 135 -70
rect 160 -95 170 -70
rect 125 -120 170 -95
rect 125 -145 135 -120
rect 160 -145 170 -120
rect 125 -1170 170 -145
rect 195 30 240 160
rect 305 530 350 560
rect 305 505 315 530
rect 340 505 350 530
rect 305 485 350 505
rect 305 460 315 485
rect 340 460 350 485
rect 305 430 350 460
rect 305 405 315 430
rect 340 405 350 430
rect 305 385 350 405
rect 305 360 315 385
rect 340 360 350 385
rect 305 330 350 360
rect 305 305 315 330
rect 340 305 350 330
rect 305 285 350 305
rect 305 260 315 285
rect 340 260 350 285
rect 305 230 350 260
rect 305 205 315 230
rect 340 205 350 230
rect 305 185 350 205
rect 305 160 315 185
rect 340 160 350 185
rect 305 150 350 160
rect 375 1730 420 1740
rect 375 1705 385 1730
rect 410 1705 420 1730
rect 375 1685 420 1705
rect 375 1660 385 1685
rect 410 1660 420 1685
rect 375 1630 420 1660
rect 375 1605 385 1630
rect 410 1605 420 1630
rect 375 1585 420 1605
rect 375 1560 385 1585
rect 410 1560 420 1585
rect 375 1530 420 1560
rect 375 1505 385 1530
rect 410 1505 420 1530
rect 375 1485 420 1505
rect 375 1460 385 1485
rect 410 1460 420 1485
rect 375 1430 420 1460
rect 375 1405 385 1430
rect 410 1405 420 1430
rect 375 1385 420 1405
rect 375 1360 385 1385
rect 410 1360 420 1385
rect 375 1330 420 1360
rect 375 1305 385 1330
rect 410 1305 420 1330
rect 375 1285 420 1305
rect 375 1260 385 1285
rect 410 1260 420 1285
rect 375 1230 420 1260
rect 375 1205 385 1230
rect 410 1205 420 1230
rect 375 1185 420 1205
rect 375 1160 385 1185
rect 410 1160 420 1185
rect 375 1130 420 1160
rect 375 1105 385 1130
rect 410 1105 420 1130
rect 375 1085 420 1105
rect 375 1060 385 1085
rect 410 1060 420 1085
rect 375 1030 420 1060
rect 375 1005 385 1030
rect 410 1005 420 1030
rect 375 985 420 1005
rect 375 960 385 985
rect 410 960 420 985
rect 375 930 420 960
rect 375 905 385 930
rect 410 905 420 930
rect 375 885 420 905
rect 375 860 385 885
rect 410 860 420 885
rect 375 830 420 860
rect 375 805 385 830
rect 410 805 420 830
rect 375 785 420 805
rect 375 760 385 785
rect 410 760 420 785
rect 375 730 420 760
rect 375 705 385 730
rect 410 705 420 730
rect 375 685 420 705
rect 375 660 385 685
rect 410 660 420 685
rect 375 630 420 660
rect 375 605 385 630
rect 410 605 420 630
rect 375 585 420 605
rect 375 560 385 585
rect 410 560 420 585
rect 375 530 420 560
rect 375 505 385 530
rect 410 505 420 530
rect 375 485 420 505
rect 375 460 385 485
rect 410 460 420 485
rect 375 430 420 460
rect 375 405 385 430
rect 410 405 420 430
rect 375 385 420 405
rect 375 360 385 385
rect 410 360 420 385
rect 375 330 420 360
rect 375 305 385 330
rect 410 305 420 330
rect 375 285 420 305
rect 375 260 385 285
rect 410 260 420 285
rect 375 230 420 260
rect 375 205 385 230
rect 410 205 420 230
rect 375 185 420 205
rect 375 160 385 185
rect 410 160 420 185
rect 305 100 355 110
rect 305 70 315 100
rect 345 70 355 100
rect 305 60 355 70
rect 195 5 205 30
rect 230 5 240 30
rect 195 -20 240 5
rect 195 -45 205 -20
rect 230 -45 240 -20
rect 195 -70 240 -45
rect 195 -95 205 -70
rect 230 -95 240 -70
rect 195 -120 240 -95
rect 195 -145 205 -120
rect 230 -145 240 -120
rect 195 -155 240 -145
rect 305 30 350 40
rect 305 5 315 30
rect 340 5 350 30
rect 305 -20 350 5
rect 305 -45 315 -20
rect 340 -45 350 -20
rect 305 -70 350 -45
rect 305 -95 315 -70
rect 340 -95 350 -70
rect 305 -120 350 -95
rect 305 -145 315 -120
rect 340 -145 350 -120
rect 305 -1170 350 -145
rect 375 30 420 160
rect 375 5 385 30
rect 410 5 420 30
rect 375 -20 420 5
rect 375 -45 385 -20
rect 410 -45 420 -20
rect 375 -70 420 -45
rect 375 -95 385 -70
rect 410 -95 420 -70
rect 375 -120 420 -95
rect 375 -145 385 -120
rect 410 -145 420 -120
rect 375 -155 420 -145
rect -60 -1180 10 -1170
rect -60 -1230 -50 -1180
rect 0 -1230 10 -1180
rect -60 -1240 10 -1230
rect 115 -1180 185 -1170
rect 115 -1230 125 -1180
rect 175 -1230 185 -1180
rect 115 -1240 185 -1230
rect 295 -1180 365 -1170
rect 295 -1230 305 -1180
rect 355 -1230 365 -1180
rect 295 -1240 365 -1230
<< viali >>
rect -50 1885 0 1935
rect 125 1885 175 1935
rect 305 1885 355 1935
rect -50 -1230 0 -1180
rect 125 -1230 175 -1180
rect 305 -1230 355 -1180
<< metal1 >>
rect -60 1935 10 1945
rect -60 1885 -50 1935
rect 0 1885 10 1935
rect -60 1875 10 1885
rect 115 1935 185 1945
rect 115 1885 125 1935
rect 175 1885 185 1935
rect 115 1875 185 1885
rect 295 1935 365 1945
rect 295 1885 305 1935
rect 355 1885 365 1935
rect 295 1875 365 1885
rect -60 -1180 10 -1170
rect -60 -1230 -50 -1180
rect 0 -1230 10 -1180
rect -60 -1240 10 -1230
rect 115 -1180 185 -1170
rect 115 -1230 125 -1180
rect 175 -1230 185 -1180
rect 115 -1240 185 -1230
rect 295 -1180 365 -1170
rect 295 -1230 305 -1180
rect 355 -1230 365 -1180
rect 295 -1240 365 -1230
<< via1 >>
rect -50 1885 0 1935
rect 125 1885 175 1935
rect 305 1885 355 1935
rect -50 -1230 0 -1180
rect 125 -1230 175 -1180
rect 305 -1230 355 -1180
<< metal2 >>
rect -60 1935 10 1945
rect -60 1885 -50 1935
rect 0 1885 10 1935
rect -60 1875 10 1885
rect 115 1935 185 1945
rect 115 1885 125 1935
rect 175 1885 185 1935
rect 115 1875 185 1885
rect 295 1935 365 1945
rect 295 1885 305 1935
rect 355 1885 365 1935
rect 295 1875 365 1885
rect -60 -1180 10 -1170
rect -60 -1230 -50 -1180
rect 0 -1230 10 -1180
rect -60 -1240 10 -1230
rect 115 -1180 185 -1170
rect 115 -1230 125 -1180
rect 175 -1230 185 -1180
rect 115 -1240 185 -1230
rect 295 -1180 365 -1170
rect 295 -1230 305 -1180
rect 355 -1230 365 -1180
rect 295 -1240 365 -1230
<< via2 >>
rect -50 1885 0 1935
rect 125 1885 175 1935
rect 305 1885 355 1935
rect -50 -1230 0 -1180
rect 125 -1230 175 -1180
rect 305 -1230 355 -1180
<< metal3 >>
rect -60 1935 10 1945
rect -60 1885 -50 1935
rect 0 1885 10 1935
rect -60 1875 10 1885
rect 115 1935 185 1945
rect 115 1885 125 1935
rect 175 1885 185 1935
rect 115 1875 185 1885
rect 295 1935 365 1945
rect 295 1885 305 1935
rect 355 1885 365 1935
rect 295 1875 365 1885
rect -60 -1180 10 -1170
rect -60 -1230 -50 -1180
rect 0 -1230 10 -1180
rect -60 -1240 10 -1230
rect 115 -1180 185 -1170
rect 115 -1230 125 -1180
rect 175 -1230 185 -1180
rect 115 -1240 185 -1230
rect 295 -1180 365 -1170
rect 295 -1230 305 -1180
rect 355 -1230 365 -1180
rect 295 -1240 365 -1230
<< via3 >>
rect -50 1885 0 1935
rect 125 1885 175 1935
rect 305 1885 355 1935
rect -50 -1230 0 -1180
rect 125 -1230 175 -1180
rect 305 -1230 355 -1180
<< metal4 >>
rect -80 1935 450 1955
rect -80 1885 -50 1935
rect 0 1885 125 1935
rect 175 1885 305 1935
rect 355 1885 450 1935
rect -80 1865 450 1885
rect -80 -1180 450 -1160
rect -80 -1230 -50 -1180
rect 0 -1230 125 -1180
rect 175 -1230 305 -1180
rect 355 -1230 450 -1180
rect -80 -1250 450 -1230
<< end >>
