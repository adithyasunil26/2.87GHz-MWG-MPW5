magic
tech sky130A
timestamp 1647865536
<< locali >>
rect -665 8178 -464 8216
rect -665 8047 -635 8178
rect -504 8047 -464 8178
rect -665 8017 -464 8047
rect 457 6820 560 6992
rect 4516 6611 5896 6828
rect 10650 5456 10773 5464
rect 10650 5356 10660 5456
rect 10764 5356 10773 5456
rect 10650 5341 10773 5356
rect -22 444 161 613
rect 1446 -30 1498 1375
rect 1931 0 1983 1359
rect 2426 93 2478 1401
rect 1440 -111 1500 -30
rect 1386 -119 1500 -111
rect -2173 -245 1500 -119
rect -2173 -249 1495 -245
rect -2173 -9118 -2064 -249
rect 1386 -250 1495 -249
rect 1927 -335 1983 0
rect 2421 -58 2478 93
rect -1869 -336 1987 -335
rect -1926 -431 1987 -336
rect -1926 -1977 -1839 -431
rect -1702 -512 -1576 -502
rect 2421 -512 2474 -58
rect 2901 -62 2953 1365
rect 3396 -34 3448 1370
rect 3999 190 4051 1437
rect -1702 -596 2479 -512
rect -1934 -8213 -1830 -1977
rect -1702 -6898 -1576 -596
rect -1450 -665 -1239 -661
rect 2895 -665 2953 -62
rect -1450 -675 2963 -665
rect -1452 -770 2963 -675
rect -1452 -772 1200 -770
rect -1452 -781 -1239 -772
rect -1452 -5319 -1336 -781
rect -1206 -880 -1122 -877
rect -1206 -885 2992 -880
rect 3395 -885 3455 -34
rect -1206 -963 3455 -885
rect -1206 -968 3453 -963
rect -1206 -1455 -1122 -968
rect 3998 -1039 4055 190
rect -1213 -1495 -1122 -1455
rect -1012 -1044 -937 -1040
rect -144 -1044 4060 -1039
rect -1012 -1137 4060 -1044
rect -1012 -1147 -113 -1137
rect -1213 -3202 -1124 -1495
rect -1012 -2032 -937 -1147
rect -1012 -2058 -732 -2032
rect -1012 -2162 -872 -2058
rect -750 -2162 -732 -2058
rect -1012 -2180 -732 -2162
rect -1213 -3648 -1125 -3202
rect -1213 -3663 -718 -3648
rect -1213 -3778 -880 -3663
rect -766 -3778 -718 -3663
rect -1213 -3796 -718 -3778
rect -898 -3802 -749 -3796
rect -1458 -5343 -862 -5319
rect -1458 -5462 -1206 -5343
rect -1081 -5462 -862 -5343
rect -1458 -5483 -862 -5462
rect -1702 -6935 -757 -6898
rect -1702 -7065 -1136 -6935
rect -994 -7065 -757 -6935
rect -1702 -7093 -757 -7065
rect -1934 -8708 -1824 -8213
rect -1934 -8735 -877 -8708
rect -1934 -8842 -1301 -8735
rect -1183 -8842 -877 -8735
rect -1934 -8870 -877 -8842
rect -2178 -9225 -2064 -9118
rect -2178 -10307 -2068 -9225
rect -1455 -10307 -1236 -10296
rect -2183 -10323 -1083 -10307
rect -2183 -10493 -1433 -10323
rect -1263 -10493 -1083 -10323
rect -2183 -10509 -1083 -10493
rect -1455 -10515 -1236 -10509
<< viali >>
rect -635 8047 -504 8178
rect 724 6790 789 6850
rect 3834 6790 3903 6858
rect 10660 5356 10764 5456
rect 33 3154 137 3250
rect -872 -2162 -750 -2058
rect -880 -3778 -766 -3663
rect -1206 -5462 -1081 -5343
rect -1136 -7065 -994 -6935
rect -1301 -8842 -1183 -8735
rect -1433 -10493 -1263 -10323
<< metal1 >>
rect -665 8178 -464 8216
rect -665 8047 -635 8178
rect -504 8047 -464 8178
rect -665 8017 -464 8047
rect -628 6149 -528 8017
rect 5408 7360 11141 7361
rect 232 7343 11141 7360
rect 232 7236 244 7343
rect 343 7236 11141 7343
rect 232 7228 11141 7236
rect 232 7227 5694 7228
rect -167 6902 5 6921
rect -167 6764 -149 6902
rect -11 6868 5 6902
rect -11 6850 816 6868
rect -11 6790 724 6850
rect 789 6790 816 6850
rect -11 6778 816 6790
rect 3826 6858 3913 6867
rect 3826 6790 3834 6858
rect 3903 6790 3913 6858
rect 3826 6779 3913 6790
rect -11 6776 318 6778
rect -11 6764 5 6776
rect -167 6748 5 6764
rect -628 6114 -504 6149
rect 183 6114 956 6116
rect -628 6022 956 6114
rect -628 6016 239 6022
rect -628 6015 128 6016
rect 10650 5458 10773 5464
rect 11028 5458 11140 7228
rect 10650 5456 11140 5458
rect 10650 5356 10660 5456
rect 10764 5356 11140 5456
rect 10650 5344 11140 5356
rect 10650 5341 10773 5344
rect 14 3250 156 3280
rect 14 3154 33 3250
rect 137 3154 156 3250
rect 14 3122 156 3154
rect -890 -2058 -719 -2030
rect -890 -2162 -872 -2058
rect -750 -2162 -719 -2058
rect -890 -2186 -719 -2162
rect -898 -3663 -749 -3648
rect -898 -3778 -880 -3663
rect -766 -3778 -749 -3663
rect -898 -3802 -749 -3778
rect -1234 -5343 -1050 -5322
rect -1234 -5462 -1206 -5343
rect -1081 -5462 -1050 -5343
rect -1234 -5480 -1050 -5462
rect -1157 -6935 -973 -6910
rect -1157 -7065 -1136 -6935
rect -994 -7065 -973 -6935
rect -1157 -7086 -973 -7065
rect -1320 -8735 -1161 -8712
rect -1320 -8842 -1301 -8735
rect -1183 -8842 -1161 -8735
rect -1320 -8866 -1161 -8842
rect -1455 -10323 -1236 -10296
rect -1455 -10493 -1433 -10323
rect -1263 -10493 -1236 -10323
rect -1455 -10515 -1236 -10493
<< via1 >>
rect -635 8047 -504 8178
rect 244 7236 343 7343
rect -149 6764 -11 6902
rect 3834 6790 3903 6858
rect 33 3154 137 3250
rect -872 -2162 -750 -2058
rect -880 -3778 -766 -3663
rect -1206 -5462 -1081 -5343
rect -1136 -7065 -994 -6935
rect -1301 -8842 -1183 -8735
rect -1433 -10493 -1263 -10323
<< metal2 >>
rect -1834 11459 -1332 11501
rect -1834 11357 -1476 11459
rect -1371 11357 -1332 11459
rect -1834 11318 -1332 11357
rect -1834 7371 -1632 11318
rect -980 9793 -515 9830
rect -980 9683 -664 9793
rect -551 9683 -515 9793
rect -980 9656 -515 9683
rect -978 9609 -864 9656
rect -979 9587 -864 9609
rect -979 7563 -866 9587
rect -665 8178 -464 8216
rect -665 8047 -635 8178
rect -504 8047 -464 8178
rect -665 8017 -464 8047
rect 366 7563 3517 7568
rect -979 7473 5712 7563
rect -979 7466 437 7473
rect 3464 7472 5712 7473
rect 5621 7455 5712 7472
rect 5621 7429 5713 7455
rect -984 7371 372 7373
rect -1834 7343 372 7371
rect -1834 7236 244 7343
rect 343 7236 372 7343
rect -1834 7218 372 7236
rect -1834 7216 -478 7218
rect -167 6902 5 6921
rect -167 6764 -149 6902
rect -11 6764 5 6902
rect 3826 6858 3913 6867
rect 3826 6790 3834 6858
rect 3903 6790 3913 6858
rect 3826 6779 3913 6790
rect 5628 6808 5713 7429
rect -167 6748 5 6764
rect 5628 6710 6272 6808
rect 5355 5956 5571 5958
rect 4434 5842 5571 5956
rect 5355 5841 5571 5842
rect 5475 5450 5571 5841
rect 5475 5431 6151 5450
rect 5475 5376 6152 5431
rect 14 3250 156 3280
rect 14 3154 33 3250
rect 137 3154 156 3250
rect 14 3122 156 3154
rect -890 -2058 -719 -2030
rect -890 -2162 -872 -2058
rect -750 -2162 -719 -2058
rect -890 -2186 -719 -2162
rect -898 -3663 -749 -3648
rect -898 -3778 -880 -3663
rect -766 -3778 -749 -3663
rect -898 -3802 -749 -3778
rect -1234 -5343 -1050 -5322
rect -1234 -5462 -1206 -5343
rect -1081 -5462 -1050 -5343
rect -1234 -5480 -1050 -5462
rect -1157 -6935 -973 -6910
rect -1157 -7065 -1136 -6935
rect -994 -7065 -973 -6935
rect -1157 -7086 -973 -7065
rect -1320 -8735 -1161 -8712
rect -1320 -8842 -1301 -8735
rect -1183 -8842 -1161 -8735
rect -1320 -8866 -1161 -8842
rect -1455 -10323 -1236 -10296
rect -1455 -10493 -1433 -10323
rect -1263 -10493 -1236 -10323
rect -1455 -10515 -1236 -10493
<< via2 >>
rect -1476 11357 -1371 11459
rect -664 9683 -551 9793
rect -635 8047 -504 8178
rect -149 6764 -11 6902
rect 3834 6790 3903 6858
rect 33 3154 137 3250
rect -872 -2162 -750 -2058
rect -880 -3778 -766 -3663
rect -1206 -5462 -1081 -5343
rect -1136 -7065 -994 -6935
rect -1301 -8842 -1183 -8735
rect -1433 -10493 -1263 -10323
<< metal3 >>
rect -1504 11459 -1346 11479
rect -1504 11357 -1476 11459
rect -1371 11357 -1346 11459
rect -1504 11335 -1346 11357
rect -676 9793 -542 9805
rect -676 9683 -664 9793
rect -551 9683 -542 9793
rect -676 9674 -542 9683
rect -665 8178 -464 8216
rect -665 8047 -635 8178
rect -504 8047 -464 8178
rect -665 8017 -464 8047
rect -167 6902 5 6921
rect -167 6764 -149 6902
rect -11 6764 5 6902
rect 3826 6858 3913 6867
rect 3826 6790 3834 6858
rect 3903 6790 3913 6858
rect 3826 6779 3913 6790
rect -167 6748 5 6764
rect 14 3250 156 3280
rect 14 3154 33 3250
rect 137 3154 156 3250
rect 14 3122 156 3154
rect -890 -2058 -719 -2030
rect -890 -2162 -872 -2058
rect -750 -2162 -719 -2058
rect -890 -2186 -719 -2162
rect -898 -3663 -749 -3648
rect -898 -3778 -880 -3663
rect -766 -3778 -749 -3663
rect -898 -3802 -749 -3778
rect -1234 -5343 -1050 -5322
rect -1234 -5462 -1206 -5343
rect -1081 -5462 -1050 -5343
rect -1234 -5480 -1050 -5462
rect -1157 -6935 -973 -6910
rect -1157 -7065 -1136 -6935
rect -994 -7065 -973 -6935
rect -1157 -7086 -973 -7065
rect -1320 -8735 -1161 -8712
rect -1320 -8842 -1301 -8735
rect -1183 -8842 -1161 -8735
rect -1320 -8866 -1161 -8842
rect -1455 -10323 -1236 -10296
rect -1455 -10493 -1433 -10323
rect -1263 -10493 -1236 -10323
rect -1455 -10515 -1236 -10493
<< via3 >>
rect -1476 11357 -1371 11459
rect -664 9683 -551 9793
rect -635 8047 -504 8178
rect -149 6764 -11 6902
rect 3834 6790 3903 6858
rect 33 3154 137 3250
rect -872 -2162 -750 -2058
rect -880 -3778 -766 -3663
rect -1206 -5462 -1081 -5343
rect -1136 -7065 -994 -6935
rect -1301 -8842 -1183 -8735
rect -1433 -10493 -1263 -10323
<< metal4 >>
rect -2967 11789 -2640 11800
rect -2967 11637 25 11789
rect -2967 11315 -2640 11637
rect -1428 11479 -293 11487
rect -1504 11459 -293 11479
rect -1504 11357 -1476 11459
rect -1371 11357 -293 11459
rect -1504 11335 -293 11357
rect -2957 10935 -2647 11315
rect -2972 10826 -2647 10935
rect -2972 10118 -2652 10826
rect -2972 10041 -69 10118
rect -2962 9978 -69 10041
rect -2962 8476 -2652 9978
rect -687 9793 -408 9825
rect -687 9683 -664 9793
rect -551 9683 -408 9793
rect -687 9661 -408 9683
rect -702 8476 -417 8479
rect -2962 8336 -64 8476
rect -2962 3370 -2652 8336
rect -702 8330 -417 8336
rect -665 8186 -464 8216
rect -665 8178 -324 8186
rect -665 8047 -635 8178
rect -504 8055 -324 8178
rect -504 8047 -464 8055
rect -665 8017 -464 8047
rect -167 6902 5 6921
rect -167 6764 -149 6902
rect -11 6764 5 6902
rect 3826 6858 5200 6876
rect 3826 6790 3834 6858
rect 3903 6790 5200 6858
rect 3826 6779 5200 6790
rect -167 6748 5 6764
rect 5108 6205 5200 6779
rect 5108 6094 6540 6205
rect 5108 6091 5200 6094
rect -2962 3250 167 3370
rect -2962 3154 33 3250
rect 137 3154 167 3250
rect -2962 3037 167 3154
rect -2962 -1749 -2652 3037
rect -2962 -1880 -364 -1749
rect -2962 -3367 -2652 -1880
rect -937 -2058 -654 -2014
rect -937 -2162 -872 -2058
rect -750 -2162 -654 -2058
rect -937 -2188 -654 -2162
rect -1305 -3367 -1213 -3361
rect -2962 -3498 -1213 -3367
rect -2962 -5020 -2652 -3498
rect -1305 -3502 -1213 -3498
rect -1125 -3367 -1002 -3361
rect -1125 -3498 -340 -3367
rect -1125 -3502 -1002 -3498
rect -950 -3663 -643 -3645
rect -950 -3778 -880 -3663
rect -766 -3778 -643 -3663
rect -950 -3799 -643 -3778
rect -898 -3802 -749 -3799
rect -2962 -5151 -450 -5020
rect -2962 -6646 -2652 -5151
rect -1338 -5343 -713 -5319
rect -1338 -5462 -1206 -5343
rect -1081 -5462 -713 -5343
rect -1338 -5483 -713 -5462
rect -2962 -6777 -412 -6646
rect -2962 -8426 -2652 -6777
rect -1383 -6935 -672 -6888
rect -1383 -7065 -1136 -6935
rect -994 -7065 -672 -6935
rect -1383 -7103 -672 -7065
rect -2962 -8557 -485 -8426
rect -2962 -10044 -2652 -8557
rect -1663 -8735 -844 -8692
rect -1663 -8842 -1301 -8735
rect -1183 -8842 -844 -8735
rect -1663 -8880 -844 -8842
rect -2962 -10174 -471 -10044
rect -2527 -10175 -471 -10174
rect -1576 -10323 -771 -10296
rect -1576 -10493 -1433 -10323
rect -1263 -10493 -771 -10323
rect -1576 -10504 -771 -10493
rect -1455 -10515 -1236 -10504
<< via4 >>
rect -149 6764 -11 6902
<< metal5 >>
rect -217 10904 28 11003
rect -227 10562 31 10904
rect -222 8956 23 9326
rect -186 7374 30 7801
rect -186 7274 29 7374
rect -1362 7270 29 7274
rect -1384 7206 29 7270
rect -1384 7019 31 7206
rect -1384 388 -1163 7019
rect -190 7006 30 7019
rect -190 6902 28 7006
rect -190 6764 -149 6902
rect -11 6764 28 6902
rect -190 6721 28 6764
rect -1387 382 -365 388
rect -1387 165 -360 382
rect -576 -1273 -360 165
rect -606 -2520 -363 -2506
rect -606 -2877 -318 -2520
rect -606 -3116 -496 -2877
rect -611 -4103 -519 -4023
rect -642 -4552 -338 -4103
rect -655 -5993 -360 -5805
rect -685 -6161 -360 -5993
rect -685 -6395 -575 -6161
rect -703 -7680 -381 -7419
rect -737 -7941 -381 -7680
rect -737 -8082 -627 -7941
rect -716 -9196 -596 -9189
rect -716 -9424 -449 -9196
rect -711 -9559 -449 -9424
rect -711 -9700 -601 -9559
use tapered_buf  tapered_buf_7
timestamp 1647818295
transform 1 0 -374 0 1 -9948
box -470 -910 43675 401
use tapered_buf  tapered_buf_6
timestamp 1647818295
transform 1 0 -414 0 1 -8329
box -470 -910 43675 401
use tapered_buf  tapered_buf_5
timestamp 1647818295
transform 1 0 -335 0 1 -6548
box -470 -910 43675 401
use tapered_buf  tapered_buf_4
timestamp 1647818295
transform 1 0 -375 0 1 -4929
box -470 -910 43675 401
use tapered_buf  tapered_buf_3
timestamp 1647818295
transform 1 0 -256 0 1 -3271
box -470 -910 43675 401
use tapered_buf  tapered_buf_2
timestamp 1647818295
transform 1 0 -296 0 1 -1652
box -470 -910 43675 401
use ro_complete  ro_complete_0
timestamp 1647865156
transform 1 0 348 0 1 5690
box -348 -5690 4661 1440
use tapered_buf  tapered_buf_0
timestamp 1647818295
transform 1 0 100 0 1 8579
box -470 -910 43675 401
use divider  divider_0
timestamp 1647865156
transform 1 0 6289 0 1 4964
box -490 -235 4690 2150
use tapered_buf  tapered_buf_1
timestamp 1647818295
transform 1 0 60 0 1 10198
box -470 -910 43675 401
use tapered_buf  tapered_buf_8
timestamp 1647818295
transform 1 0 65 0 1 11875
box -470 -910 43675 401
<< labels >>
rlabel metal4 -2844 3190 -2844 3190 1 gnd!
rlabel space -819 -9903 -819 -9903 1 a0
rlabel space -854 -8280 -854 -8280 1 a1
rlabel space -779 -6505 -779 -6505 1 a2
rlabel space -798 -4893 -798 -4893 1 a3
rlabel space -701 -3231 -701 -3231 1 a4
rlabel space -728 -1606 -728 -1606 1 a5
rlabel space -107 11937 -107 11937 1 vdd!
rlabel metal5 -112 10587 -112 10587 1 vdd!
rlabel space -324 8611 -324 8611 1 vcont
rlabel space -338 9736 -338 9736 1 out
rlabel space -395 10231 -395 10231 1 mc2
rlabel space -390 11890 -390 11890 1 out
<< end >>
