magic
tech sky130A
magscale 1 2
timestamp 1640799896
<< nwell >>
rect -250 320 1600 1010
rect -116 -750 186 -397
rect 534 -752 836 -399
rect 1202 -756 1504 -403
<< nmos >>
rect -110 -20 -50 180
rect 640 -20 700 180
rect 1400 -20 1460 180
<< pmos >>
rect -110 360 -50 760
rect 640 360 700 760
rect 1400 360 1460 760
<< varactor >>
rect 17 -688 53 -488
rect 667 -690 703 -490
rect 1335 -694 1371 -494
<< ndiff >>
rect -210 150 -110 180
rect -210 10 -180 150
rect -140 10 -110 150
rect -210 -20 -110 10
rect -50 150 50 180
rect -50 10 -20 150
rect 20 10 50 150
rect -50 -20 50 10
rect 540 150 640 180
rect 540 10 570 150
rect 610 10 640 150
rect 540 -20 640 10
rect 700 150 800 180
rect 700 10 730 150
rect 770 10 800 150
rect 700 -20 800 10
rect 1300 150 1400 180
rect 1300 10 1330 150
rect 1370 10 1400 150
rect 1300 -20 1400 10
rect 1460 150 1560 180
rect 1460 10 1490 150
rect 1530 10 1560 150
rect 1460 -20 1560 10
<< pdiff >>
rect -210 730 -110 760
rect -210 390 -180 730
rect -140 390 -110 730
rect -210 360 -110 390
rect -50 730 50 760
rect -50 390 -20 730
rect 20 390 50 730
rect -50 360 50 390
rect 540 730 640 760
rect 540 390 570 730
rect 610 390 640 730
rect 540 360 640 390
rect 700 730 800 760
rect 700 390 730 730
rect 770 390 800 730
rect 700 360 800 390
rect 1300 730 1400 760
rect 1300 390 1330 730
rect 1370 390 1400 730
rect 1300 360 1400 390
rect 1460 730 1560 760
rect 1460 390 1490 730
rect 1530 390 1560 730
rect 1460 360 1560 390
<< ndiffc >>
rect -180 10 -140 150
rect -20 10 20 150
rect 570 10 610 150
rect 730 10 770 150
rect 1330 10 1370 150
rect 1490 10 1530 150
<< pdiffc >>
rect -180 390 -140 730
rect -20 390 20 730
rect 570 390 610 730
rect 730 390 770 730
rect 1330 390 1370 730
rect 1490 390 1530 730
<< psubdiff >>
rect 0 -120 230 -90
rect 0 -170 30 -120
rect 200 -170 230 -120
rect 0 -200 230 -170
rect 500 -120 800 -90
rect 500 -180 530 -120
rect 770 -180 800 -120
rect 500 -200 800 -180
rect 1050 -120 1280 -90
rect 1050 -170 1080 -120
rect 1250 -170 1280 -120
rect 1050 -200 1280 -170
rect 300 -270 430 -240
rect 300 -340 330 -270
rect 400 -340 430 -270
rect 300 -370 430 -340
rect 300 -650 430 -620
rect 300 -720 330 -650
rect 400 -720 430 -650
rect 300 -750 430 -720
<< nsubdiff >>
rect 510 950 830 970
rect 510 880 540 950
rect 800 880 830 950
rect 510 860 830 880
rect -80 -512 17 -488
rect -80 -664 -68 -512
rect -34 -664 17 -512
rect -80 -688 17 -664
rect 53 -512 150 -488
rect 53 -664 104 -512
rect 138 -664 150 -512
rect 570 -514 667 -490
rect 53 -688 150 -664
rect 570 -666 582 -514
rect 616 -666 667 -514
rect 570 -690 667 -666
rect 703 -514 800 -490
rect 703 -666 754 -514
rect 788 -666 800 -514
rect 703 -690 800 -666
rect 1238 -518 1335 -494
rect 1238 -670 1250 -518
rect 1284 -670 1335 -518
rect 1238 -694 1335 -670
rect 1371 -518 1468 -494
rect 1371 -670 1422 -518
rect 1456 -670 1468 -518
rect 1371 -694 1468 -670
<< psubdiffcont >>
rect 30 -170 200 -120
rect 530 -180 770 -120
rect 1080 -170 1250 -120
rect 330 -340 400 -270
rect 330 -720 400 -650
<< nsubdiffcont >>
rect 540 880 800 950
rect -68 -664 -34 -512
rect 104 -664 138 -512
rect 582 -666 616 -514
rect 754 -666 788 -514
rect 1250 -670 1284 -518
rect 1422 -670 1456 -518
<< poly >>
rect -110 760 -50 790
rect 640 760 700 790
rect 1400 760 1460 790
rect -110 300 -50 360
rect 640 300 700 360
rect 1400 300 1460 360
rect -190 280 -50 300
rect -190 240 -170 280
rect -130 240 -50 280
rect -190 220 -50 240
rect 560 280 700 300
rect 560 240 580 280
rect 620 240 700 280
rect 560 220 700 240
rect 1320 280 1460 300
rect 1320 240 1340 280
rect 1380 240 1460 280
rect 1320 220 1460 240
rect -110 180 -50 220
rect 640 180 700 220
rect 1400 180 1460 220
rect -110 -50 -50 -20
rect 640 -50 700 -20
rect 1400 -50 1460 -20
rect 2 -416 68 -400
rect 2 -450 18 -416
rect 52 -450 68 -416
rect 2 -466 68 -450
rect 652 -418 718 -402
rect 652 -452 668 -418
rect 702 -452 718 -418
rect 17 -488 53 -466
rect 652 -468 718 -452
rect 1320 -422 1386 -406
rect 1320 -456 1336 -422
rect 1370 -456 1386 -422
rect 667 -490 703 -468
rect 1320 -472 1386 -456
rect 17 -714 53 -688
rect 1335 -494 1371 -472
rect 667 -716 703 -690
rect 1335 -720 1371 -694
<< polycont >>
rect -170 240 -130 280
rect 580 240 620 280
rect 1340 240 1380 280
rect 18 -450 52 -416
rect 668 -452 702 -418
rect 1336 -456 1370 -422
<< locali >>
rect -250 950 1600 1010
rect -250 880 540 950
rect 800 880 1600 950
rect -250 830 1600 880
rect -200 730 -120 830
rect -200 390 -180 730
rect -140 390 -120 730
rect -200 370 -120 390
rect -40 730 40 750
rect -40 390 -20 730
rect 20 390 40 730
rect -190 290 -110 300
rect -190 230 -180 290
rect -120 230 -110 290
rect -190 220 -110 230
rect -40 290 40 390
rect 550 730 630 830
rect 550 390 570 730
rect 610 390 630 730
rect 550 370 630 390
rect 710 730 790 750
rect 710 390 730 730
rect 770 390 790 730
rect -40 230 560 290
rect -200 150 -120 170
rect -200 10 -180 150
rect -140 10 -120 150
rect -200 -80 -120 10
rect -40 150 40 230
rect 710 290 790 390
rect 1310 730 1390 830
rect 1310 390 1330 730
rect 1370 390 1390 730
rect 1310 370 1390 390
rect 1470 730 1550 750
rect 1470 390 1490 730
rect 1530 390 1550 730
rect 1470 310 1550 390
rect 710 230 1320 290
rect -40 10 -20 150
rect 20 10 40 150
rect -40 -10 40 10
rect 550 150 630 170
rect 550 10 570 150
rect 610 10 630 150
rect 550 -80 630 10
rect 710 150 790 230
rect 1470 210 1570 310
rect 710 10 730 150
rect 770 10 790 150
rect 710 -10 790 10
rect 1310 150 1390 170
rect 1310 10 1330 150
rect 1370 10 1390 150
rect 1310 -80 1390 10
rect 1470 150 1550 210
rect 1470 10 1490 150
rect 1530 10 1550 150
rect 1470 -10 1550 10
rect -230 -120 1600 -80
rect -230 -170 30 -120
rect 200 -170 530 -120
rect -230 -180 530 -170
rect 770 -170 1080 -120
rect 1250 -170 1600 -120
rect 770 -180 1600 -170
rect -230 -220 1600 -180
rect 290 -270 440 -220
rect 290 -340 330 -270
rect 400 -340 440 -270
rect 2 -450 18 -416
rect 52 -450 68 -416
rect -68 -512 -34 -496
rect -68 -680 -34 -664
rect 104 -512 138 -496
rect 104 -680 138 -664
rect 290 -650 440 -340
rect 652 -452 668 -418
rect 702 -452 718 -418
rect 1320 -456 1336 -422
rect 1370 -456 1386 -422
rect 290 -720 330 -650
rect 400 -720 440 -650
rect 582 -514 616 -498
rect 582 -682 616 -666
rect 754 -514 788 -498
rect 754 -682 788 -666
rect 1250 -518 1284 -502
rect 1250 -686 1284 -670
rect 1422 -518 1456 -502
rect 1422 -686 1456 -670
rect 1636 -680 1670 -510
rect 290 -800 440 -720
<< viali >>
rect -180 280 -120 290
rect -180 240 -170 280
rect -170 240 -130 280
rect -130 240 -120 280
rect -180 230 -120 240
rect 560 280 640 300
rect 560 240 580 280
rect 580 240 620 280
rect 620 240 640 280
rect 560 220 640 240
rect 1320 280 1400 300
rect 1320 240 1340 280
rect 1340 240 1380 280
rect 1380 240 1400 280
rect 1320 220 1400 240
rect 1570 230 1630 290
rect 18 -450 52 -416
rect -68 -664 -34 -512
rect 104 -664 138 -512
rect 668 -452 702 -418
rect 1336 -456 1370 -422
rect 582 -666 616 -514
rect 754 -666 788 -514
rect 1250 -670 1284 -518
rect 1422 -670 1456 -518
<< metal1 >>
rect -200 290 -110 310
rect -200 230 -180 290
rect -120 230 -110 290
rect -200 210 -110 230
rect 270 300 660 310
rect 270 220 560 300
rect 640 220 660 300
rect 270 210 660 220
rect 950 300 1420 310
rect 950 220 1320 300
rect 1400 220 1420 300
rect 950 210 1420 220
rect 1550 290 1650 310
rect 1550 230 1570 290
rect 1630 230 1650 290
rect 270 -100 370 210
rect -10 -200 370 -100
rect -10 -416 90 -200
rect 950 -260 1050 210
rect 1550 -100 1650 230
rect -10 -450 18 -416
rect 52 -450 90 -416
rect -10 -470 90 -450
rect 640 -308 1050 -260
rect 1300 -200 1650 -100
rect 640 -418 740 -308
rect 640 -452 668 -418
rect 702 -452 740 -418
rect 640 -470 740 -452
rect 1300 -422 1400 -200
rect 1300 -456 1336 -422
rect 1370 -456 1400 -422
rect 1300 -470 1400 -456
rect -130 -512 1656 -500
rect -130 -664 -68 -512
rect -34 -664 104 -512
rect 138 -514 1656 -512
rect 138 -664 582 -514
rect -130 -666 582 -664
rect 616 -666 754 -514
rect 788 -518 1656 -514
rect 788 -666 1250 -518
rect -130 -670 1250 -666
rect 1284 -670 1422 -518
rect 1456 -670 1656 -518
rect -130 -680 1656 -670
rect 1244 -682 1290 -680
rect 1416 -682 1462 -680
<< via1 >>
rect -180 230 -120 290
rect 1570 230 1630 290
<< metal2 >>
rect -200 290 1650 310
rect -200 230 -180 290
rect -120 230 1570 290
rect 1630 230 1650 290
rect -200 210 1650 230
<< labels >>
rlabel locali 1400 900 1400 900 1 vdd
rlabel locali 1360 -160 1360 -160 1 gnd
rlabel viali 1600 260 1600 260 1 out3
rlabel locali 10 200 10 200 1 out1
rlabel locali 750 190 750 190 1 out2
rlabel locali 1510 190 1510 190 1 out3
rlabel locali 1666 -610 1666 -610 1 vcont
<< end >>
