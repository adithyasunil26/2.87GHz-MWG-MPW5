magic
tech sky130A
timestamp 1647810727
<< locali >>
rect 5076 1340 5818 1489
rect 4847 790 4958 799
rect -384 575 55 722
rect 4847 698 4859 790
rect 4949 698 4958 790
rect 4847 689 4958 698
rect 5109 81 5851 230
<< viali >>
rect 4859 698 4949 790
<< metal1 >>
rect 7867 1139 7942 1144
rect 7476 1114 7942 1139
rect 7519 996 7545 997
rect 7466 977 7545 996
rect 4847 793 4958 799
rect 4847 791 5351 793
rect 4847 790 5493 791
rect -480 730 -295 750
rect -480 568 -467 730
rect -308 568 -295 730
rect 4847 698 4859 790
rect 4949 702 5493 790
rect 4949 698 5497 702
rect 4847 689 4958 698
rect 5316 697 5497 698
rect 5425 583 5497 697
rect 7519 653 7545 977
rect -480 552 -295 568
rect 5424 566 5497 583
rect 5389 550 5534 566
rect 5389 454 5403 550
rect 5518 454 5534 550
rect 5389 438 5534 454
rect 7488 59 7560 653
rect 2050 -94 4971 -84
rect -520 -96 4971 -94
rect 7485 -96 7565 59
rect 7867 5 7942 1114
rect -520 -100 7565 -96
rect -525 -171 7565 -100
rect 7865 -163 7945 5
rect -525 -172 7557 -171
rect -525 -188 32 -172
rect 2050 -174 7557 -172
rect 2050 -175 4971 -174
rect -525 -2102 -380 -188
rect -60 -316 29 -314
rect -60 -318 4956 -316
rect 7862 -318 7951 -163
rect -60 -399 7951 -318
rect -60 -402 7940 -399
rect -60 -707 29 -402
rect 2035 -404 7940 -402
rect 2035 -407 4956 -404
rect -143 -742 50 -707
rect -143 -873 -108 -742
rect 13 -873 50 -742
rect -143 -897 50 -873
rect -542 -2128 -354 -2102
rect -542 -2252 -518 -2128
rect -384 -2252 -354 -2128
rect -542 -2273 -354 -2252
<< via1 >>
rect -467 568 -308 730
rect 5403 454 5518 550
rect -108 -873 13 -742
rect -518 -2252 -384 -2128
<< metal2 >>
rect -590 6498 -406 6516
rect -590 6365 -571 6498
rect -425 6365 -406 6498
rect -590 6349 -406 6365
rect -552 1658 -444 6349
rect -275 5109 -121 5121
rect -275 4994 -259 5109
rect -133 4994 -121 5109
rect -275 4980 -121 4994
rect -244 3039 -161 4980
rect -42 3574 90 3586
rect -42 3473 -30 3574
rect 77 3473 90 3574
rect -42 3463 90 3473
rect 3 3188 48 3463
rect 2229 3189 3802 3191
rect 213 3188 5364 3189
rect 3 3187 5364 3188
rect 5594 3187 5648 3188
rect 3 3138 5648 3187
rect 3 3136 5364 3138
rect 3 3134 259 3136
rect 3791 3134 5364 3136
rect -244 3037 252 3039
rect -244 2978 361 3037
rect -135 2976 361 2978
rect 300 2099 358 2976
rect -552 1568 7 1658
rect -86 794 4 1568
rect 5594 1220 5648 3138
rect 5594 1145 5915 1220
rect -86 791 258 794
rect -480 730 -295 750
rect -480 568 -467 730
rect -308 568 -295 730
rect -86 736 312 791
rect -86 725 258 736
rect -86 724 4 725
rect -480 552 -295 568
rect 5389 550 5534 566
rect 5389 454 5403 550
rect 5518 454 5534 550
rect 5389 438 5534 454
rect 5432 378 5502 438
rect 5432 375 5616 378
rect 5432 301 5918 375
rect -143 -742 50 -707
rect -143 -873 -108 -742
rect 13 -873 50 -742
rect -143 -897 50 -873
rect -542 -2128 -354 -2102
rect -542 -2252 -518 -2128
rect -384 -2150 -354 -2128
rect -384 -2244 56 -2150
rect -384 -2252 -354 -2244
rect -542 -2273 -354 -2252
<< via2 >>
rect -571 6365 -425 6498
rect -259 4994 -133 5109
rect -30 3473 77 3574
rect -467 568 -308 730
<< metal3 >>
rect -590 6498 -406 6516
rect -590 6365 -571 6498
rect -425 6365 -406 6498
rect -590 6349 -406 6365
rect -275 5109 -121 5121
rect -275 4994 -259 5109
rect -133 4994 -121 5109
rect -275 4980 -121 4994
rect -42 3574 90 3586
rect -42 3473 -30 3574
rect 77 3473 90 3574
rect -42 3463 90 3473
rect -480 730 -295 750
rect -480 568 -467 730
rect -308 568 -295 730
rect -480 552 -295 568
<< via3 >>
rect -571 6365 -425 6498
rect -259 4994 -133 5109
rect -30 3473 77 3574
rect -467 568 -308 730
<< metal4 >>
rect -926 6659 308 6794
rect -924 6016 -768 6659
rect -590 6498 61 6532
rect -590 6365 -571 6498
rect -425 6365 61 6498
rect -590 6349 61 6365
rect -929 5424 -768 6016
rect -929 5415 308 5424
rect -926 5289 308 5415
rect -924 4075 -768 5289
rect -275 5109 63 5137
rect -275 4994 -259 5109
rect -133 4994 63 5109
rect -275 4980 63 4994
rect -570 4075 67 4078
rect -924 3936 354 4075
rect -924 3931 -287 3936
rect -105 3931 354 3936
rect -924 713 -768 3931
rect -37 3586 86 3777
rect -42 3574 90 3586
rect -42 3473 -30 3574
rect 77 3473 90 3574
rect -42 3463 90 3473
rect 4174 1459 5867 1465
rect 4174 1414 5983 1459
rect 8466 1421 8575 3429
rect 4174 1403 5867 1414
rect 7463 1369 8575 1421
rect -480 730 -295 750
rect -480 714 -467 730
rect -559 713 -467 714
rect -924 577 -467 713
rect -924 -959 -768 577
rect -559 573 -467 577
rect -480 568 -467 573
rect -308 568 -295 730
rect -480 552 -295 568
rect 8466 -612 8575 1369
rect -924 -1134 329 -959
rect -924 -2333 -768 -1134
rect -947 -2508 293 -2333
<< metal5 >>
rect 186 6072 404 6077
rect 179 5655 414 6072
rect 186 4503 404 4707
rect 145 -1871 363 -1667
use tapered_buf  tapered_buf_4
timestamp 1647784636
transform 1 0 473 0 1 6893
box -470 -910 43675 400
use pd  pd_1
timestamp 1647810585
transform 1 0 6015 0 1 779
box -215 -855 1685 810
use divider  divider_0
timestamp 1647769399
transform 1 0 489 0 1 316
box -490 -235 4690 2150
use tapered_buf  tapered_buf_1
timestamp 1647784636
transform 1 0 473 0 1 5523
box -470 -910 43675 400
use tapered_buf  tapered_buf_0
timestamp 1647784636
transform 1 0 468 0 1 4170
box -470 -910 43675 400
use tapered_buf  tapered_buf_3
timestamp 1647784636
transform 1 0 429 0 1 -2234
box -470 -910 43675 400
use tapered_buf  tapered_buf_2
timestamp 1647784636
transform 1 0 434 0 1 -881
box -470 -910 43675 400
<< labels >>
rlabel space 40 -1345 40 -1345 1 up
rlabel space -14 -2692 -14 -2692 1 down
rlabel space 48 4207 48 4207 1 ref
rlabel space 64 5553 64 5553 1 div
rlabel space 64 6923 64 6923 1 div
rlabel space 18 6944 18 6944 1 clk
rlabel space 32 5564 32 5564 1 mc2
rlabel space 13 4217 13 4217 1 ref
rlabel metal4 8501 2091 8501 2091 1 vdd!
rlabel metal4 -877 1968 -877 1968 1 gnd!
<< end >>
