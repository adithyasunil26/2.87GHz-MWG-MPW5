magic
tech sky130A
timestamp 1640958486
<< nwell >>
rect 0 680 1530 690
rect 0 580 1555 680
rect 1430 360 1555 580
rect 995 -615 1155 -410
rect 0 -730 1155 -615
<< psubdiff >>
rect -210 790 -130 805
rect -210 740 -195 790
rect -145 740 -130 790
rect -210 725 -130 740
rect -65 790 15 805
rect -65 740 -50 790
rect 0 740 15 790
rect -65 725 15 740
rect 295 790 375 805
rect 295 740 310 790
rect 360 740 375 790
rect 295 725 375 740
rect 655 790 735 805
rect 655 740 670 790
rect 720 740 735 790
rect 655 725 735 740
rect 1015 790 1095 805
rect 1015 740 1030 790
rect 1080 740 1095 790
rect 1015 725 1095 740
rect 1375 790 1455 805
rect 1375 740 1390 790
rect 1440 740 1455 790
rect 1375 725 1455 740
rect 1600 710 1680 725
rect 1600 660 1615 710
rect 1665 660 1680 710
rect 1600 645 1680 660
rect -210 430 -130 445
rect -210 380 -195 430
rect -145 380 -130 430
rect -210 365 -130 380
rect 1600 350 1680 365
rect 1600 300 1615 350
rect 1665 300 1680 350
rect 1600 285 1680 300
rect -210 70 -130 85
rect -210 20 -195 70
rect -145 20 -130 70
rect -210 5 -130 20
rect 1365 -40 1445 -25
rect 1365 -90 1380 -40
rect 1430 -90 1445 -40
rect 1365 -105 1445 -90
rect 1230 -210 1310 -195
rect 1230 -260 1245 -210
rect 1295 -260 1310 -210
rect 1230 -275 1310 -260
rect -210 -290 -130 -275
rect -210 -340 -195 -290
rect -145 -340 -130 -290
rect -210 -355 -130 -340
rect 1230 -570 1310 -555
rect 1230 -620 1245 -570
rect 1295 -620 1310 -570
rect 1230 -635 1310 -620
rect -210 -650 -130 -635
rect -210 -700 -195 -650
rect -145 -700 -130 -650
rect -210 -715 -130 -700
rect -65 -785 15 -770
rect -65 -835 -50 -785
rect 0 -835 15 -785
rect -65 -850 15 -835
rect 295 -785 375 -770
rect 295 -835 310 -785
rect 360 -835 375 -785
rect 295 -850 375 -835
rect 655 -785 735 -770
rect 655 -835 670 -785
rect 720 -835 735 -785
rect 655 -850 735 -835
rect 1015 -785 1095 -770
rect 1015 -835 1030 -785
rect 1080 -835 1095 -785
rect 1015 -850 1095 -835
<< nsubdiff >>
rect 1445 525 1515 540
rect 1445 485 1460 525
rect 1500 485 1515 525
rect 1445 470 1515 485
rect 1050 -515 1120 -500
rect 1050 -555 1065 -515
rect 1105 -555 1120 -515
rect 1050 -570 1120 -555
<< psubdiffcont >>
rect -195 740 -145 790
rect -50 740 0 790
rect 310 740 360 790
rect 670 740 720 790
rect 1030 740 1080 790
rect 1390 740 1440 790
rect 1615 660 1665 710
rect -195 380 -145 430
rect 1615 300 1665 350
rect -195 20 -145 70
rect 1380 -90 1430 -40
rect 1245 -260 1295 -210
rect -195 -340 -145 -290
rect 1245 -620 1295 -570
rect -195 -700 -145 -650
rect -50 -835 0 -785
rect 310 -835 360 -785
rect 670 -835 720 -785
rect 1030 -835 1080 -785
<< nsubdiffcont >>
rect 1460 485 1500 525
rect 1065 -555 1105 -515
<< locali >>
rect -215 790 1685 810
rect -215 740 -195 790
rect -145 740 -50 790
rect 0 740 310 790
rect 360 740 670 790
rect 720 740 1030 790
rect 1080 740 1390 790
rect 1440 740 1685 790
rect -215 720 1685 740
rect -215 430 -125 720
rect 1595 710 1685 720
rect 1595 660 1615 710
rect 1665 660 1685 710
rect 1450 525 1510 535
rect 1450 485 1460 525
rect 1500 485 1510 525
rect 1450 475 1510 485
rect -215 380 -195 430
rect -145 380 -125 430
rect -215 70 -125 380
rect 1595 350 1685 660
rect 1595 300 1615 350
rect 1665 300 1685 350
rect -215 20 -195 70
rect -145 50 -125 70
rect -145 20 60 50
rect -215 15 60 20
rect -215 -290 -125 15
rect 1595 -20 1685 300
rect -215 -340 -195 -290
rect -145 -340 -125 -290
rect -215 -650 -125 -340
rect 1225 -40 1685 -20
rect 1225 -90 1380 -40
rect 1430 -90 1685 -40
rect 1225 -110 1685 -90
rect 1225 -210 1315 -110
rect 1225 -260 1245 -210
rect 1295 -260 1315 -210
rect 1055 -515 1115 -505
rect 1055 -555 1065 -515
rect 1105 -555 1115 -515
rect 1055 -565 1115 -555
rect -215 -700 -195 -650
rect -145 -700 -125 -650
rect -215 -765 -125 -700
rect 1225 -570 1315 -260
rect 1225 -620 1245 -570
rect 1295 -620 1315 -570
rect 1225 -765 1315 -620
rect -215 -785 1315 -765
rect -215 -835 -50 -785
rect 0 -835 310 -785
rect 360 -835 670 -785
rect 720 -835 1030 -785
rect 1080 -835 1315 -785
rect -215 -855 1315 -835
<< viali >>
rect 1460 485 1500 525
rect 30 320 50 340
rect 1080 280 1100 300
rect 1435 280 1455 300
rect 30 -385 50 -365
rect 1065 -555 1105 -515
<< metal1 >>
rect 1450 525 1510 535
rect 1450 485 1460 525
rect 1500 485 1510 525
rect 1450 475 1510 485
rect 20 345 60 350
rect 20 315 25 345
rect 55 315 60 345
rect 20 310 60 315
rect 1005 335 1050 350
rect 1200 335 1470 350
rect 1005 300 1020 335
rect 1070 300 1110 310
rect 1070 285 1080 300
rect 1020 280 1080 285
rect 1100 280 1110 300
rect 1020 270 1110 280
rect 1425 305 1465 310
rect 1425 275 1430 305
rect 1460 275 1465 305
rect 1425 270 1465 275
rect 1020 215 1035 270
rect 1020 200 1470 215
rect 20 -360 60 -355
rect 1020 -360 1035 200
rect 20 -390 25 -360
rect 55 -390 60 -360
rect 20 -395 60 -390
rect 1055 -515 1115 -505
rect 1055 -555 1065 -515
rect 1105 -555 1115 -515
rect 1055 -565 1115 -555
<< via1 >>
rect 1460 485 1500 525
rect 25 340 55 345
rect 25 320 30 340
rect 30 320 50 340
rect 50 320 55 340
rect 25 315 55 320
rect 1430 300 1460 305
rect 1430 280 1435 300
rect 1435 280 1455 300
rect 1455 280 1460 300
rect 1430 275 1460 280
rect 25 -365 55 -360
rect 25 -385 30 -365
rect 30 -385 50 -365
rect 50 -385 55 -365
rect 25 -390 55 -385
rect 1065 -555 1105 -515
<< metal2 >>
rect 1450 525 1510 535
rect 1450 485 1460 525
rect 1500 485 1510 525
rect 1450 475 1510 485
rect -115 395 0 410
rect 20 345 60 350
rect 20 315 25 345
rect 55 315 60 345
rect 20 310 60 315
rect 1420 305 1470 315
rect 1420 295 1430 305
rect 415 280 1430 295
rect 420 265 505 280
rect 1420 275 1430 280
rect 1460 275 1470 305
rect 1420 265 1470 275
rect 490 -310 505 265
rect 425 -325 505 -310
rect 15 -360 65 -350
rect 15 -390 25 -360
rect 55 -390 65 -360
rect 15 -400 65 -390
rect -115 -455 0 -440
rect 1055 -515 1115 -505
rect 1055 -555 1065 -515
rect 1105 -555 1115 -515
rect 1055 -565 1115 -555
<< via2 >>
rect 1460 485 1500 525
rect 25 315 55 345
rect 25 -390 55 -360
rect 1065 -555 1105 -515
<< metal3 >>
rect 1450 525 1510 535
rect 1450 485 1460 525
rect 1500 485 1510 525
rect 1450 475 1510 485
rect 15 350 65 355
rect 15 310 20 350
rect 60 310 65 350
rect 15 305 65 310
rect 15 -355 65 -350
rect 15 -395 20 -355
rect 60 -395 65 -355
rect 15 -400 65 -395
rect 1055 -515 1115 -505
rect 1055 -555 1065 -515
rect 1105 -555 1115 -515
rect 1055 -565 1115 -555
<< via3 >>
rect 1460 485 1500 525
rect 20 345 60 350
rect 20 315 25 345
rect 25 315 55 345
rect 55 315 60 345
rect 20 310 60 315
rect 20 -360 60 -355
rect 20 -390 25 -360
rect 25 -390 55 -360
rect 55 -390 60 -360
rect 20 -395 60 -390
rect 1065 -555 1105 -515
<< metal4 >>
rect -70 640 20 670
rect 720 640 925 670
rect -70 350 -40 640
rect 1405 600 1490 630
rect 1445 535 1490 600
rect 1445 525 1510 535
rect 1445 485 1460 525
rect 1500 485 1510 525
rect 1445 480 1510 485
rect 1450 475 1510 480
rect 15 350 65 355
rect -70 320 20 350
rect -70 -360 -40 320
rect 15 310 20 320
rect 60 310 65 350
rect 15 305 65 310
rect 10 -65 1020 20
rect 15 -355 65 -350
rect 15 -360 20 -355
rect -70 -390 20 -360
rect -70 -685 -40 -390
rect 15 -395 20 -390
rect 60 -395 65 -355
rect 15 -400 65 -395
rect 1050 -505 1095 -500
rect 1050 -515 1115 -505
rect 1050 -555 1065 -515
rect 1105 -555 1115 -515
rect 1050 -560 1115 -555
rect 1055 -565 1115 -560
rect 1065 -685 1105 -565
rect -70 -715 20 -685
rect 1020 -715 1105 -685
use tspc_r  tspc_r_0
timestamp 1640958486
transform 1 0 145 0 1 380
box -145 -380 875 305
use tspc_r  tspc_r_1
timestamp 1640958486
transform 1 0 145 0 -1 -425
box -145 -380 875 305
use and_pd  and_pd_0
timestamp 1640958486
transform 1 0 1100 0 1 395
box -120 -375 335 275
<< labels >>
rlabel nwell 980 600 1050 630 1 VDD
rlabel nwell 980 630 1020 640 1 VDD
rlabel space 985 50 1020 120 1 GND
rlabel space 985 85 1050 120 1 GND
rlabel metal4 10 -65 1020 20 1 GND
rlabel metal4 -70 -715 -40 670 1 VDD
rlabel metal2 -115 395 -70 410 1 REF
rlabel metal2 -115 -455 -70 -440 1 DIV
rlabel metal1 1415 335 1470 350 1 UP
rlabel metal1 1415 200 1470 215 1 DOWN
rlabel metal2 1435 280 1460 305 1 R
rlabel metal2 1140 280 1185 295 1 R
<< end >>
