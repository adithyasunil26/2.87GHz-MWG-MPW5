magic
tech sky130A
timestamp 1647883901
<< psubdiff >>
rect 83392 340047 84757 340157
rect 83392 338865 83511 340047
rect 84635 338865 84757 340047
rect 83392 338762 84757 338865
rect 90350 340048 91715 340158
rect 90350 338866 90469 340048
rect 91593 338866 91715 340048
rect 90350 338763 91715 338866
rect 97168 340027 98533 340137
rect 97168 338845 97287 340027
rect 98411 338845 98533 340027
rect 97168 338742 98533 338845
rect 104133 340028 105498 340138
rect 104133 338846 104252 340028
rect 105376 338846 105498 340028
rect 104133 338743 105498 338846
rect 111091 340029 112456 340139
rect 111091 338847 111210 340029
rect 112334 338847 112456 340029
rect 111091 338744 112456 338847
rect 118011 340028 119376 340138
rect 118011 338846 118130 340028
rect 119254 338846 119376 340028
rect 118011 338743 119376 338846
rect 124976 340029 126341 340139
rect 124976 338847 125095 340029
rect 126219 338847 126341 340029
rect 124976 338744 126341 338847
rect 131934 340030 133299 340140
rect 131934 338848 132053 340030
rect 133177 338848 133299 340030
rect 131934 338745 133299 338848
rect 138851 340034 140216 340144
rect 138851 338852 138970 340034
rect 140094 338852 140216 340034
rect 138851 338749 140216 338852
rect 145816 340035 147181 340145
rect 145816 338853 145935 340035
rect 147059 338853 147181 340035
rect 145816 338750 147181 338853
rect 152774 340036 154139 340146
rect 152774 338854 152893 340036
rect 154017 338854 154139 340036
rect 152774 338751 154139 338854
rect 159691 340034 161056 340144
rect 159691 338852 159810 340034
rect 160934 338852 161056 340034
rect 159691 338749 161056 338852
rect 166656 340035 168021 340145
rect 166656 338853 166775 340035
rect 167899 338853 168021 340035
rect 166656 338750 168021 338853
rect 173614 340036 174979 340146
rect 173614 338854 173733 340036
rect 174857 338854 174979 340036
rect 173614 338751 174979 338854
rect 180419 340029 181784 340139
rect 180419 338847 180538 340029
rect 181662 338847 181784 340029
rect 180419 338744 181784 338847
rect 187384 340030 188749 340140
rect 187384 338848 187503 340030
rect 188627 338848 188749 340030
rect 187384 338745 188749 338848
rect 194342 340031 195707 340141
rect 194342 338849 194461 340031
rect 195585 338849 195707 340031
rect 194342 338746 195707 338849
rect 201262 340030 202627 340140
rect 201262 338848 201381 340030
rect 202505 338848 202627 340030
rect 201262 338745 202627 338848
rect 208227 340031 209592 340141
rect 208227 338849 208346 340031
rect 209470 338849 209592 340031
rect 208227 338746 209592 338849
rect 215185 340032 216550 340142
rect 215185 338850 215304 340032
rect 216428 338850 216550 340032
rect 215185 338747 216550 338850
rect 96894 332897 98259 333007
rect 96894 331715 97013 332897
rect 98137 331715 98259 332897
rect 96894 331612 98259 331715
rect 103859 332898 105224 333008
rect 103859 331716 103978 332898
rect 105102 331716 105224 332898
rect 103859 331613 105224 331716
rect 138577 332904 139942 333014
rect 138577 331722 138696 332904
rect 139820 331722 139942 332904
rect 138577 331619 139942 331722
rect 145542 332905 146907 333015
rect 145542 331723 145661 332905
rect 146785 331723 146907 332905
rect 145542 331620 146907 331723
rect 152500 332906 153865 333016
rect 152500 331724 152619 332906
rect 153743 331724 153865 332906
rect 152500 331621 153865 331724
rect 159417 332904 160782 333014
rect 159417 331722 159536 332904
rect 160660 331722 160782 332904
rect 159417 331619 160782 331722
rect 166382 332905 167747 333015
rect 166382 331723 166501 332905
rect 167625 331723 167747 332905
rect 166382 331620 167747 331723
rect 173340 332906 174705 333016
rect 173340 331724 173459 332906
rect 174583 331724 174705 332906
rect 173340 331621 174705 331724
rect 180145 332899 181510 333009
rect 180145 331717 180264 332899
rect 181388 331717 181510 332899
rect 180145 331614 181510 331717
rect 187110 332900 188475 333010
rect 187110 331718 187229 332900
rect 188353 331718 188475 332900
rect 187110 331615 188475 331718
rect 194068 332901 195433 333011
rect 194068 331719 194187 332901
rect 195311 331719 195433 332901
rect 194068 331616 195433 331719
rect 200988 332900 202353 333010
rect 200988 331718 201107 332900
rect 202231 331718 202353 332900
rect 200988 331615 202353 331718
rect 207953 332901 209318 333011
rect 207953 331719 208072 332901
rect 209196 331719 209318 332901
rect 207953 331616 209318 331719
rect 214911 332902 216276 333012
rect 214911 331720 215030 332902
rect 216154 331720 216276 332902
rect 214911 331617 216276 331720
rect 97168 326569 98533 326679
rect 97168 325387 97287 326569
rect 98411 325387 98533 326569
rect 97168 325284 98533 325387
rect 104133 326570 105498 326680
rect 104133 325388 104252 326570
rect 105376 325388 105498 326570
rect 104133 325285 105498 325388
rect 138851 326576 140216 326686
rect 138851 325394 138970 326576
rect 140094 325394 140216 326576
rect 138851 325291 140216 325394
rect 145816 326577 147181 326687
rect 145816 325395 145935 326577
rect 147059 325395 147181 326577
rect 145816 325292 147181 325395
rect 152774 326578 154139 326688
rect 152774 325396 152893 326578
rect 154017 325396 154139 326578
rect 152774 325293 154139 325396
rect 159691 326576 161056 326686
rect 159691 325394 159810 326576
rect 160934 325394 161056 326576
rect 159691 325291 161056 325394
rect 166656 326577 168021 326687
rect 166656 325395 166775 326577
rect 167899 325395 168021 326577
rect 166656 325292 168021 325395
rect 173614 326578 174979 326688
rect 173614 325396 173733 326578
rect 174857 325396 174979 326578
rect 173614 325293 174979 325396
rect 180419 326571 181784 326681
rect 180419 325389 180538 326571
rect 181662 325389 181784 326571
rect 180419 325286 181784 325389
rect 187384 326572 188749 326682
rect 187384 325390 187503 326572
rect 188627 325390 188749 326572
rect 187384 325287 188749 325390
rect 194342 326573 195707 326683
rect 194342 325391 194461 326573
rect 195585 325391 195707 326573
rect 194342 325288 195707 325391
rect 201262 326572 202627 326682
rect 201262 325390 201381 326572
rect 202505 325390 202627 326572
rect 201262 325287 202627 325390
rect 208227 326573 209592 326683
rect 208227 325391 208346 326573
rect 209470 325391 209592 326573
rect 208227 325288 209592 325391
rect 215185 326574 216550 326684
rect 215185 325392 215304 326574
rect 216428 325392 216550 326574
rect 215185 325289 216550 325392
rect 96894 319439 98259 319549
rect 96894 318257 97013 319439
rect 98137 318257 98259 319439
rect 96894 318154 98259 318257
rect 103859 319440 105224 319550
rect 103859 318258 103978 319440
rect 105102 318258 105224 319440
rect 103859 318155 105224 318258
rect 138577 319446 139942 319556
rect 138577 318264 138696 319446
rect 139820 318264 139942 319446
rect 138577 318161 139942 318264
rect 145542 319447 146907 319557
rect 145542 318265 145661 319447
rect 146785 318265 146907 319447
rect 145542 318162 146907 318265
rect 152500 319448 153865 319558
rect 152500 318266 152619 319448
rect 153743 318266 153865 319448
rect 152500 318163 153865 318266
rect 159417 319446 160782 319556
rect 159417 318264 159536 319446
rect 160660 318264 160782 319446
rect 159417 318161 160782 318264
rect 166382 319447 167747 319557
rect 166382 318265 166501 319447
rect 167625 318265 167747 319447
rect 166382 318162 167747 318265
rect 173340 319448 174705 319558
rect 173340 318266 173459 319448
rect 174583 318266 174705 319448
rect 173340 318163 174705 318266
rect 180145 319441 181510 319551
rect 180145 318259 180264 319441
rect 181388 318259 181510 319441
rect 180145 318156 181510 318259
rect 187110 319442 188475 319552
rect 187110 318260 187229 319442
rect 188353 318260 188475 319442
rect 187110 318157 188475 318260
rect 194068 319443 195433 319553
rect 194068 318261 194187 319443
rect 195311 318261 195433 319443
rect 194068 318158 195433 318261
rect 200988 319442 202353 319552
rect 200988 318260 201107 319442
rect 202231 318260 202353 319442
rect 200988 318157 202353 318260
rect 207953 319443 209318 319553
rect 207953 318261 208072 319443
rect 209196 318261 209318 319443
rect 207953 318158 209318 318261
rect 214911 319444 216276 319554
rect 214911 318262 215030 319444
rect 216154 318262 216276 319444
rect 214911 318159 216276 318262
rect 97174 312308 98539 312418
rect 97174 311126 97293 312308
rect 98417 311126 98539 312308
rect 97174 311023 98539 311126
rect 104139 312309 105504 312419
rect 104139 311127 104258 312309
rect 105382 311127 105504 312309
rect 104139 311024 105504 311127
rect 138857 312315 140222 312425
rect 138857 311133 138976 312315
rect 140100 311133 140222 312315
rect 138857 311030 140222 311133
rect 145822 312316 147187 312426
rect 145822 311134 145941 312316
rect 147065 311134 147187 312316
rect 145822 311031 147187 311134
rect 152780 312317 154145 312427
rect 152780 311135 152899 312317
rect 154023 311135 154145 312317
rect 152780 311032 154145 311135
rect 159697 312315 161062 312425
rect 159697 311133 159816 312315
rect 160940 311133 161062 312315
rect 159697 311030 161062 311133
rect 166662 312316 168027 312426
rect 166662 311134 166781 312316
rect 167905 311134 168027 312316
rect 166662 311031 168027 311134
rect 173620 312317 174985 312427
rect 173620 311135 173739 312317
rect 174863 311135 174985 312317
rect 173620 311032 174985 311135
rect 180425 312310 181790 312420
rect 180425 311128 180544 312310
rect 181668 311128 181790 312310
rect 180425 311025 181790 311128
rect 187390 312311 188755 312421
rect 187390 311129 187509 312311
rect 188633 311129 188755 312311
rect 187390 311026 188755 311129
rect 194348 312312 195713 312422
rect 194348 311130 194467 312312
rect 195591 311130 195713 312312
rect 194348 311027 195713 311130
rect 201268 312311 202633 312421
rect 201268 311129 201387 312311
rect 202511 311129 202633 312311
rect 201268 311026 202633 311129
rect 208233 312312 209598 312422
rect 208233 311130 208352 312312
rect 209476 311130 209598 312312
rect 208233 311027 209598 311130
rect 215191 312313 216556 312423
rect 215191 311131 215310 312313
rect 216434 311131 216556 312313
rect 215191 311028 216556 311131
rect 83124 305198 84489 305308
rect 83124 304016 83243 305198
rect 84367 304016 84489 305198
rect 83124 303913 84489 304016
rect 90082 305199 91447 305309
rect 90082 304017 90201 305199
rect 91325 304017 91447 305199
rect 90082 303914 91447 304017
rect 96900 305178 98265 305288
rect 96900 303996 97019 305178
rect 98143 303996 98265 305178
rect 96900 303893 98265 303996
rect 103865 305179 105230 305289
rect 103865 303997 103984 305179
rect 105108 303997 105230 305179
rect 103865 303894 105230 303997
rect 110823 305180 112188 305290
rect 110823 303998 110942 305180
rect 112066 303998 112188 305180
rect 110823 303895 112188 303998
rect 117743 305179 119108 305289
rect 117743 303997 117862 305179
rect 118986 303997 119108 305179
rect 117743 303894 119108 303997
rect 124708 305180 126073 305290
rect 124708 303998 124827 305180
rect 125951 303998 126073 305180
rect 124708 303895 126073 303998
rect 131666 305181 133031 305291
rect 131666 303999 131785 305181
rect 132909 303999 133031 305181
rect 131666 303896 133031 303999
rect 138583 305185 139948 305295
rect 138583 304003 138702 305185
rect 139826 304003 139948 305185
rect 138583 303900 139948 304003
rect 145548 305186 146913 305296
rect 145548 304004 145667 305186
rect 146791 304004 146913 305186
rect 145548 303901 146913 304004
rect 152506 305187 153871 305297
rect 152506 304005 152625 305187
rect 153749 304005 153871 305187
rect 152506 303902 153871 304005
rect 159423 305185 160788 305295
rect 159423 304003 159542 305185
rect 160666 304003 160788 305185
rect 159423 303900 160788 304003
rect 166388 305186 167753 305296
rect 166388 304004 166507 305186
rect 167631 304004 167753 305186
rect 166388 303901 167753 304004
rect 173346 305187 174711 305297
rect 173346 304005 173465 305187
rect 174589 304005 174711 305187
rect 173346 303902 174711 304005
rect 180151 305180 181516 305290
rect 180151 303998 180270 305180
rect 181394 303998 181516 305180
rect 180151 303895 181516 303998
rect 187116 305181 188481 305291
rect 187116 303999 187235 305181
rect 188359 303999 188481 305181
rect 187116 303896 188481 303999
rect 194074 305182 195439 305292
rect 194074 304000 194193 305182
rect 195317 304000 195439 305182
rect 194074 303897 195439 304000
rect 200994 305181 202359 305291
rect 200994 303999 201113 305181
rect 202237 303999 202359 305181
rect 200994 303896 202359 303999
rect 207959 305182 209324 305292
rect 207959 304000 208078 305182
rect 209202 304000 209324 305182
rect 207959 303897 209324 304000
rect 214917 305183 216282 305293
rect 214917 304001 215036 305183
rect 216160 304001 216282 305183
rect 214917 303898 216282 304001
rect 97263 295949 98628 296059
rect 97263 294767 97382 295949
rect 98506 294767 98628 295949
rect 97263 294664 98628 294767
rect 104228 295950 105593 296060
rect 104228 294768 104347 295950
rect 105471 294768 105593 295950
rect 104228 294665 105593 294768
rect 138946 295956 140311 296066
rect 138946 294774 139065 295956
rect 140189 294774 140311 295956
rect 138946 294671 140311 294774
rect 145911 295957 147276 296067
rect 145911 294775 146030 295957
rect 147154 294775 147276 295957
rect 145911 294672 147276 294775
rect 152869 295958 154234 296068
rect 152869 294776 152988 295958
rect 154112 294776 154234 295958
rect 152869 294673 154234 294776
rect 159786 295956 161151 296066
rect 159786 294774 159905 295956
rect 161029 294774 161151 295956
rect 159786 294671 161151 294774
rect 166751 295957 168116 296067
rect 166751 294775 166870 295957
rect 167994 294775 168116 295957
rect 166751 294672 168116 294775
rect 187479 295952 188844 296062
rect 187479 294770 187598 295952
rect 188722 294770 188844 295952
rect 187479 294667 188844 294770
rect 194437 295953 195802 296063
rect 194437 294771 194556 295953
rect 195680 294771 195802 295953
rect 194437 294668 195802 294771
rect 96989 288819 98354 288929
rect 96989 287637 97108 288819
rect 98232 287637 98354 288819
rect 96989 287534 98354 287637
rect 103954 288820 105319 288930
rect 103954 287638 104073 288820
rect 105197 287638 105319 288820
rect 103954 287535 105319 287638
rect 138672 288826 140037 288936
rect 138672 287644 138791 288826
rect 139915 287644 140037 288826
rect 138672 287541 140037 287644
rect 145637 288827 147002 288937
rect 145637 287645 145756 288827
rect 146880 287645 147002 288827
rect 145637 287542 147002 287645
rect 152595 288828 153960 288938
rect 152595 287646 152714 288828
rect 153838 287646 153960 288828
rect 152595 287543 153960 287646
rect 159512 288826 160877 288936
rect 159512 287644 159631 288826
rect 160755 287644 160877 288826
rect 159512 287541 160877 287644
rect 166477 288827 167842 288937
rect 166477 287645 166596 288827
rect 167720 287645 167842 288827
rect 166477 287542 167842 287645
rect 187205 288822 188570 288932
rect 187205 287640 187324 288822
rect 188448 287640 188570 288822
rect 187205 287537 188570 287640
rect 194163 288823 195528 288933
rect 194163 287641 194282 288823
rect 195406 287641 195528 288823
rect 194163 287538 195528 287641
rect 97097 282406 98462 282516
rect 97097 281224 97216 282406
rect 98340 281224 98462 282406
rect 97097 281121 98462 281224
rect 104062 282407 105427 282517
rect 104062 281225 104181 282407
rect 105305 281225 105427 282407
rect 104062 281122 105427 281225
rect 138780 282413 140145 282523
rect 138780 281231 138899 282413
rect 140023 281231 140145 282413
rect 138780 281128 140145 281231
rect 145745 282414 147110 282524
rect 145745 281232 145864 282414
rect 146988 281232 147110 282414
rect 145745 281129 147110 281232
rect 152703 282415 154068 282525
rect 152703 281233 152822 282415
rect 153946 281233 154068 282415
rect 152703 281130 154068 281233
rect 159620 282413 160985 282523
rect 159620 281231 159739 282413
rect 160863 281231 160985 282413
rect 159620 281128 160985 281231
rect 166585 282414 167950 282524
rect 166585 281232 166704 282414
rect 167828 281232 167950 282414
rect 166585 281129 167950 281232
rect 187313 282409 188678 282519
rect 187313 281227 187432 282409
rect 188556 281227 188678 282409
rect 187313 281124 188678 281227
rect 194271 282410 195636 282520
rect 194271 281228 194390 282410
rect 195514 281228 195636 282410
rect 194271 281125 195636 281228
rect 69656 273562 71021 273672
rect 69656 272380 69775 273562
rect 70899 272380 71021 273562
rect 69656 272277 71021 272380
rect 76573 273560 77938 273670
rect 76573 272378 76692 273560
rect 77816 272378 77938 273560
rect 76573 272275 77938 272378
rect 83538 273561 84903 273671
rect 83538 272379 83657 273561
rect 84781 272379 84903 273561
rect 83538 272276 84903 272379
rect 90496 273562 91861 273672
rect 90496 272380 90615 273562
rect 91739 272380 91861 273562
rect 90496 272277 91861 272380
rect 97314 273541 98679 273651
rect 97314 272359 97433 273541
rect 98557 272359 98679 273541
rect 97314 272256 98679 272359
rect 104279 273542 105644 273652
rect 104279 272360 104398 273542
rect 105522 272360 105644 273542
rect 104279 272257 105644 272360
rect 111237 273543 112602 273653
rect 111237 272361 111356 273543
rect 112480 272361 112602 273543
rect 111237 272258 112602 272361
rect 118157 273542 119522 273652
rect 118157 272360 118276 273542
rect 119400 272360 119522 273542
rect 118157 272257 119522 272360
rect 125122 273543 126487 273653
rect 125122 272361 125241 273543
rect 126365 272361 126487 273543
rect 125122 272258 126487 272361
rect 132080 273544 133445 273654
rect 132080 272362 132199 273544
rect 133323 272362 133445 273544
rect 132080 272259 133445 272362
rect 138997 273548 140362 273658
rect 138997 272366 139116 273548
rect 140240 272366 140362 273548
rect 138997 272263 140362 272366
rect 145962 273549 147327 273659
rect 145962 272367 146081 273549
rect 147205 272367 147327 273549
rect 145962 272264 147327 272367
rect 152920 273550 154285 273660
rect 152920 272368 153039 273550
rect 154163 272368 154285 273550
rect 152920 272265 154285 272368
rect 159837 273548 161202 273658
rect 159837 272366 159956 273548
rect 161080 272366 161202 273548
rect 159837 272263 161202 272366
rect 166802 273549 168167 273659
rect 166802 272367 166921 273549
rect 168045 272367 168167 273549
rect 166802 272264 168167 272367
rect 173760 273550 175125 273660
rect 173760 272368 173879 273550
rect 175003 272368 175125 273550
rect 173760 272265 175125 272368
rect 180565 273543 181930 273653
rect 180565 272361 180684 273543
rect 181808 272361 181930 273543
rect 180565 272258 181930 272361
rect 187530 273544 188895 273654
rect 187530 272362 187649 273544
rect 188773 272362 188895 273544
rect 187530 272259 188895 272362
rect 194488 273545 195853 273655
rect 194488 272363 194607 273545
rect 195731 272363 195853 273545
rect 194488 272260 195853 272363
rect 201408 273544 202773 273654
rect 201408 272362 201527 273544
rect 202651 272362 202773 273544
rect 201408 272259 202773 272362
rect 208373 273545 209738 273655
rect 208373 272363 208492 273545
rect 209616 272363 209738 273545
rect 208373 272260 209738 272363
rect 215331 273546 216696 273656
rect 215331 272364 215450 273546
rect 216574 272364 216696 273546
rect 215331 272261 216696 272364
rect 222248 273550 223613 273660
rect 222248 272368 222367 273550
rect 223491 272368 223613 273550
rect 222248 272265 223613 272368
rect 69382 266432 70747 266542
rect 69382 265250 69501 266432
rect 70625 265250 70747 266432
rect 69382 265147 70747 265250
rect 76299 266430 77664 266540
rect 76299 265248 76418 266430
rect 77542 265248 77664 266430
rect 76299 265145 77664 265248
rect 83264 266431 84629 266541
rect 83264 265249 83383 266431
rect 84507 265249 84629 266431
rect 83264 265146 84629 265249
rect 90222 266432 91587 266542
rect 90222 265250 90341 266432
rect 91465 265250 91587 266432
rect 90222 265147 91587 265250
rect 97040 266411 98405 266521
rect 97040 265229 97159 266411
rect 98283 265229 98405 266411
rect 97040 265126 98405 265229
rect 104005 266412 105370 266522
rect 104005 265230 104124 266412
rect 105248 265230 105370 266412
rect 104005 265127 105370 265230
rect 110963 266413 112328 266523
rect 110963 265231 111082 266413
rect 112206 265231 112328 266413
rect 110963 265128 112328 265231
rect 117883 266412 119248 266522
rect 117883 265230 118002 266412
rect 119126 265230 119248 266412
rect 117883 265127 119248 265230
rect 124848 266413 126213 266523
rect 124848 265231 124967 266413
rect 126091 265231 126213 266413
rect 124848 265128 126213 265231
rect 131806 266414 133171 266524
rect 131806 265232 131925 266414
rect 133049 265232 133171 266414
rect 131806 265129 133171 265232
rect 138723 266418 140088 266528
rect 138723 265236 138842 266418
rect 139966 265236 140088 266418
rect 138723 265133 140088 265236
rect 145688 266419 147053 266529
rect 145688 265237 145807 266419
rect 146931 265237 147053 266419
rect 145688 265134 147053 265237
rect 152646 266420 154011 266530
rect 152646 265238 152765 266420
rect 153889 265238 154011 266420
rect 152646 265135 154011 265238
rect 159563 266418 160928 266528
rect 159563 265236 159682 266418
rect 160806 265236 160928 266418
rect 159563 265133 160928 265236
rect 166528 266419 167893 266529
rect 166528 265237 166647 266419
rect 167771 265237 167893 266419
rect 166528 265134 167893 265237
rect 173486 266420 174851 266530
rect 173486 265238 173605 266420
rect 174729 265238 174851 266420
rect 173486 265135 174851 265238
rect 180291 266413 181656 266523
rect 180291 265231 180410 266413
rect 181534 265231 181656 266413
rect 180291 265128 181656 265231
rect 187256 266414 188621 266524
rect 187256 265232 187375 266414
rect 188499 265232 188621 266414
rect 187256 265129 188621 265232
rect 194214 266415 195579 266525
rect 194214 265233 194333 266415
rect 195457 265233 195579 266415
rect 194214 265130 195579 265233
rect 201134 266414 202499 266524
rect 201134 265232 201253 266414
rect 202377 265232 202499 266414
rect 201134 265129 202499 265232
rect 208099 266415 209464 266525
rect 208099 265233 208218 266415
rect 209342 265233 209464 266415
rect 208099 265130 209464 265233
rect 215057 266416 216422 266526
rect 215057 265234 215176 266416
rect 216300 265234 216422 266416
rect 215057 265131 216422 265234
rect 221974 266420 223339 266530
rect 221974 265238 222093 266420
rect 223217 265238 223339 266420
rect 221974 265135 223339 265238
rect 69490 260019 70855 260129
rect 69490 258837 69609 260019
rect 70733 258837 70855 260019
rect 69490 258734 70855 258837
rect 76407 260017 77772 260127
rect 76407 258835 76526 260017
rect 77650 258835 77772 260017
rect 76407 258732 77772 258835
rect 83372 260018 84737 260128
rect 83372 258836 83491 260018
rect 84615 258836 84737 260018
rect 83372 258733 84737 258836
rect 90330 260019 91695 260129
rect 90330 258837 90449 260019
rect 91573 258837 91695 260019
rect 90330 258734 91695 258837
rect 97148 259998 98513 260108
rect 97148 258816 97267 259998
rect 98391 258816 98513 259998
rect 97148 258713 98513 258816
rect 104113 259999 105478 260109
rect 104113 258817 104232 259999
rect 105356 258817 105478 259999
rect 104113 258714 105478 258817
rect 111071 260000 112436 260110
rect 111071 258818 111190 260000
rect 112314 258818 112436 260000
rect 111071 258715 112436 258818
rect 117991 259999 119356 260109
rect 117991 258817 118110 259999
rect 119234 258817 119356 259999
rect 117991 258714 119356 258817
rect 124956 260000 126321 260110
rect 124956 258818 125075 260000
rect 126199 258818 126321 260000
rect 124956 258715 126321 258818
rect 131914 260001 133279 260111
rect 131914 258819 132033 260001
rect 133157 258819 133279 260001
rect 131914 258716 133279 258819
rect 138831 260005 140196 260115
rect 138831 258823 138950 260005
rect 140074 258823 140196 260005
rect 138831 258720 140196 258823
rect 145796 260006 147161 260116
rect 145796 258824 145915 260006
rect 147039 258824 147161 260006
rect 145796 258721 147161 258824
rect 152754 260007 154119 260117
rect 152754 258825 152873 260007
rect 153997 258825 154119 260007
rect 152754 258722 154119 258825
rect 159671 260005 161036 260115
rect 159671 258823 159790 260005
rect 160914 258823 161036 260005
rect 159671 258720 161036 258823
rect 166636 260006 168001 260116
rect 166636 258824 166755 260006
rect 167879 258824 168001 260006
rect 166636 258721 168001 258824
rect 173594 260007 174959 260117
rect 173594 258825 173713 260007
rect 174837 258825 174959 260007
rect 173594 258722 174959 258825
rect 180399 260000 181764 260110
rect 180399 258818 180518 260000
rect 181642 258818 181764 260000
rect 180399 258715 181764 258818
rect 187364 260001 188729 260111
rect 187364 258819 187483 260001
rect 188607 258819 188729 260001
rect 187364 258716 188729 258819
rect 194322 260002 195687 260112
rect 194322 258820 194441 260002
rect 195565 258820 195687 260002
rect 194322 258717 195687 258820
rect 201242 260001 202607 260111
rect 201242 258819 201361 260001
rect 202485 258819 202607 260001
rect 201242 258716 202607 258819
rect 208207 260002 209572 260112
rect 208207 258820 208326 260002
rect 209450 258820 209572 260002
rect 208207 258717 209572 258820
rect 215165 260003 216530 260113
rect 215165 258821 215284 260003
rect 216408 258821 216530 260003
rect 215165 258718 216530 258821
rect 222082 260007 223447 260117
rect 222082 258825 222201 260007
rect 223325 258825 223447 260007
rect 222082 258722 223447 258825
rect 83569 249307 84934 249417
rect 83569 248125 83688 249307
rect 84812 248125 84934 249307
rect 83569 248022 84934 248125
rect 90527 249308 91892 249418
rect 90527 248126 90646 249308
rect 91770 248126 91892 249308
rect 90527 248023 91892 248126
rect 97345 249287 98710 249397
rect 97345 248105 97464 249287
rect 98588 248105 98710 249287
rect 97345 248002 98710 248105
rect 104310 249288 105675 249398
rect 104310 248106 104429 249288
rect 105553 248106 105675 249288
rect 104310 248003 105675 248106
rect 111268 249289 112633 249399
rect 111268 248107 111387 249289
rect 112511 248107 112633 249289
rect 111268 248004 112633 248107
rect 118188 249288 119553 249398
rect 118188 248106 118307 249288
rect 119431 248106 119553 249288
rect 118188 248003 119553 248106
rect 125153 249289 126518 249399
rect 125153 248107 125272 249289
rect 126396 248107 126518 249289
rect 125153 248004 126518 248107
rect 132111 249290 133476 249400
rect 132111 248108 132230 249290
rect 133354 248108 133476 249290
rect 132111 248005 133476 248108
rect 139028 249294 140393 249404
rect 139028 248112 139147 249294
rect 140271 248112 140393 249294
rect 139028 248009 140393 248112
rect 145993 249295 147358 249405
rect 145993 248113 146112 249295
rect 147236 248113 147358 249295
rect 145993 248010 147358 248113
rect 152951 249296 154316 249406
rect 152951 248114 153070 249296
rect 154194 248114 154316 249296
rect 152951 248011 154316 248114
rect 159868 249294 161233 249404
rect 159868 248112 159987 249294
rect 161111 248112 161233 249294
rect 159868 248009 161233 248112
rect 166833 249295 168198 249405
rect 166833 248113 166952 249295
rect 168076 248113 168198 249295
rect 166833 248010 168198 248113
rect 173791 249296 175156 249406
rect 173791 248114 173910 249296
rect 175034 248114 175156 249296
rect 173791 248011 175156 248114
rect 180596 249289 181961 249399
rect 180596 248107 180715 249289
rect 181839 248107 181961 249289
rect 180596 248004 181961 248107
rect 187561 249290 188926 249400
rect 187561 248108 187680 249290
rect 188804 248108 188926 249290
rect 187561 248005 188926 248108
rect 194519 249291 195884 249401
rect 194519 248109 194638 249291
rect 195762 248109 195884 249291
rect 194519 248006 195884 248109
rect 201439 249290 202804 249400
rect 201439 248108 201558 249290
rect 202682 248108 202804 249290
rect 201439 248005 202804 248108
rect 208404 249291 209769 249401
rect 208404 248109 208523 249291
rect 209647 248109 209769 249291
rect 208404 248006 209769 248109
rect 215362 249292 216727 249402
rect 215362 248110 215481 249292
rect 216605 248110 216727 249292
rect 215362 248007 216727 248110
rect 222279 249296 223644 249406
rect 222279 248114 222398 249296
rect 223522 248114 223644 249296
rect 222279 248011 223644 248114
rect 83295 242177 84660 242287
rect 83295 240995 83414 242177
rect 84538 240995 84660 242177
rect 83295 240892 84660 240995
rect 90253 242178 91618 242288
rect 90253 240996 90372 242178
rect 91496 240996 91618 242178
rect 90253 240893 91618 240996
rect 97071 242157 98436 242267
rect 97071 240975 97190 242157
rect 98314 240975 98436 242157
rect 97071 240872 98436 240975
rect 104036 242158 105401 242268
rect 104036 240976 104155 242158
rect 105279 240976 105401 242158
rect 104036 240873 105401 240976
rect 110994 242159 112359 242269
rect 110994 240977 111113 242159
rect 112237 240977 112359 242159
rect 110994 240874 112359 240977
rect 117914 242158 119279 242268
rect 117914 240976 118033 242158
rect 119157 240976 119279 242158
rect 117914 240873 119279 240976
rect 124879 242159 126244 242269
rect 124879 240977 124998 242159
rect 126122 240977 126244 242159
rect 124879 240874 126244 240977
rect 131837 242160 133202 242270
rect 131837 240978 131956 242160
rect 133080 240978 133202 242160
rect 131837 240875 133202 240978
rect 138754 242164 140119 242274
rect 138754 240982 138873 242164
rect 139997 240982 140119 242164
rect 138754 240879 140119 240982
rect 145719 242165 147084 242275
rect 145719 240983 145838 242165
rect 146962 240983 147084 242165
rect 145719 240880 147084 240983
rect 152677 242166 154042 242276
rect 152677 240984 152796 242166
rect 153920 240984 154042 242166
rect 152677 240881 154042 240984
rect 159594 242164 160959 242274
rect 159594 240982 159713 242164
rect 160837 240982 160959 242164
rect 159594 240879 160959 240982
rect 166559 242165 167924 242275
rect 166559 240983 166678 242165
rect 167802 240983 167924 242165
rect 166559 240880 167924 240983
rect 173517 242166 174882 242276
rect 173517 240984 173636 242166
rect 174760 240984 174882 242166
rect 173517 240881 174882 240984
rect 180322 242159 181687 242269
rect 180322 240977 180441 242159
rect 181565 240977 181687 242159
rect 180322 240874 181687 240977
rect 187287 242160 188652 242270
rect 187287 240978 187406 242160
rect 188530 240978 188652 242160
rect 187287 240875 188652 240978
rect 194245 242161 195610 242271
rect 194245 240979 194364 242161
rect 195488 240979 195610 242161
rect 194245 240876 195610 240979
rect 201165 242160 202530 242270
rect 201165 240978 201284 242160
rect 202408 240978 202530 242160
rect 201165 240875 202530 240978
rect 208130 242161 209495 242271
rect 208130 240979 208249 242161
rect 209373 240979 209495 242161
rect 208130 240876 209495 240979
rect 215088 242162 216453 242272
rect 215088 240980 215207 242162
rect 216331 240980 216453 242162
rect 215088 240877 216453 240980
rect 222005 242166 223370 242276
rect 222005 240984 222124 242166
rect 223248 240984 223370 242166
rect 222005 240881 223370 240984
rect 83403 235764 84768 235874
rect 83403 234582 83522 235764
rect 84646 234582 84768 235764
rect 83403 234479 84768 234582
rect 90361 235765 91726 235875
rect 90361 234583 90480 235765
rect 91604 234583 91726 235765
rect 90361 234480 91726 234583
rect 97179 235744 98544 235854
rect 97179 234562 97298 235744
rect 98422 234562 98544 235744
rect 97179 234459 98544 234562
rect 104144 235745 105509 235855
rect 104144 234563 104263 235745
rect 105387 234563 105509 235745
rect 104144 234460 105509 234563
rect 111102 235746 112467 235856
rect 111102 234564 111221 235746
rect 112345 234564 112467 235746
rect 111102 234461 112467 234564
rect 118022 235745 119387 235855
rect 118022 234563 118141 235745
rect 119265 234563 119387 235745
rect 118022 234460 119387 234563
rect 124987 235746 126352 235856
rect 124987 234564 125106 235746
rect 126230 234564 126352 235746
rect 124987 234461 126352 234564
rect 131945 235747 133310 235857
rect 131945 234565 132064 235747
rect 133188 234565 133310 235747
rect 131945 234462 133310 234565
rect 138862 235751 140227 235861
rect 138862 234569 138981 235751
rect 140105 234569 140227 235751
rect 138862 234466 140227 234569
rect 145827 235752 147192 235862
rect 145827 234570 145946 235752
rect 147070 234570 147192 235752
rect 145827 234467 147192 234570
rect 152785 235753 154150 235863
rect 152785 234571 152904 235753
rect 154028 234571 154150 235753
rect 152785 234468 154150 234571
rect 159702 235751 161067 235861
rect 159702 234569 159821 235751
rect 160945 234569 161067 235751
rect 159702 234466 161067 234569
rect 166667 235752 168032 235862
rect 166667 234570 166786 235752
rect 167910 234570 168032 235752
rect 166667 234467 168032 234570
rect 173625 235753 174990 235863
rect 173625 234571 173744 235753
rect 174868 234571 174990 235753
rect 173625 234468 174990 234571
rect 180430 235746 181795 235856
rect 180430 234564 180549 235746
rect 181673 234564 181795 235746
rect 180430 234461 181795 234564
rect 187395 235747 188760 235857
rect 187395 234565 187514 235747
rect 188638 234565 188760 235747
rect 187395 234462 188760 234565
rect 194353 235748 195718 235858
rect 194353 234566 194472 235748
rect 195596 234566 195718 235748
rect 194353 234463 195718 234566
rect 201273 235747 202638 235857
rect 201273 234565 201392 235747
rect 202516 234565 202638 235747
rect 201273 234462 202638 234565
rect 208238 235748 209603 235858
rect 208238 234566 208357 235748
rect 209481 234566 209603 235748
rect 208238 234463 209603 234566
rect 215196 235749 216561 235859
rect 215196 234567 215315 235749
rect 216439 234567 216561 235749
rect 215196 234464 216561 234567
rect 222113 235753 223478 235863
rect 222113 234571 222232 235753
rect 223356 234571 223478 235753
rect 222113 234468 223478 234571
rect 69811 229042 71176 229152
rect 69811 227860 69930 229042
rect 71054 227860 71176 229042
rect 69811 227757 71176 227860
rect 76728 229040 78093 229150
rect 76728 227858 76847 229040
rect 77971 227858 78093 229040
rect 76728 227755 78093 227858
rect 83693 229041 85058 229151
rect 83693 227859 83812 229041
rect 84936 227859 85058 229041
rect 83693 227756 85058 227859
rect 90651 229042 92016 229152
rect 90651 227860 90770 229042
rect 91894 227860 92016 229042
rect 90651 227757 92016 227860
rect 97469 229021 98834 229131
rect 97469 227839 97588 229021
rect 98712 227839 98834 229021
rect 97469 227736 98834 227839
rect 104434 229022 105799 229132
rect 104434 227840 104553 229022
rect 105677 227840 105799 229022
rect 104434 227737 105799 227840
rect 111392 229023 112757 229133
rect 111392 227841 111511 229023
rect 112635 227841 112757 229023
rect 111392 227738 112757 227841
rect 118312 229022 119677 229132
rect 118312 227840 118431 229022
rect 119555 227840 119677 229022
rect 118312 227737 119677 227840
rect 125277 229023 126642 229133
rect 125277 227841 125396 229023
rect 126520 227841 126642 229023
rect 125277 227738 126642 227841
rect 132235 229024 133600 229134
rect 132235 227842 132354 229024
rect 133478 227842 133600 229024
rect 132235 227739 133600 227842
rect 139152 229028 140517 229138
rect 139152 227846 139271 229028
rect 140395 227846 140517 229028
rect 139152 227743 140517 227846
rect 146117 229029 147482 229139
rect 146117 227847 146236 229029
rect 147360 227847 147482 229029
rect 146117 227744 147482 227847
rect 153075 229030 154440 229140
rect 153075 227848 153194 229030
rect 154318 227848 154440 229030
rect 153075 227745 154440 227848
rect 159992 229028 161357 229138
rect 159992 227846 160111 229028
rect 161235 227846 161357 229028
rect 159992 227743 161357 227846
rect 166957 229029 168322 229139
rect 166957 227847 167076 229029
rect 168200 227847 168322 229029
rect 166957 227744 168322 227847
rect 173915 229030 175280 229140
rect 173915 227848 174034 229030
rect 175158 227848 175280 229030
rect 173915 227745 175280 227848
rect 180720 229023 182085 229133
rect 180720 227841 180839 229023
rect 181963 227841 182085 229023
rect 180720 227738 182085 227841
rect 187685 229024 189050 229134
rect 187685 227842 187804 229024
rect 188928 227842 189050 229024
rect 187685 227739 189050 227842
rect 194643 229025 196008 229135
rect 194643 227843 194762 229025
rect 195886 227843 196008 229025
rect 194643 227740 196008 227843
rect 201563 229024 202928 229134
rect 201563 227842 201682 229024
rect 202806 227842 202928 229024
rect 201563 227739 202928 227842
rect 208528 229025 209893 229135
rect 208528 227843 208647 229025
rect 209771 227843 209893 229025
rect 208528 227740 209893 227843
rect 215486 229026 216851 229136
rect 215486 227844 215605 229026
rect 216729 227844 216851 229026
rect 215486 227741 216851 227844
rect 222403 229030 223768 229140
rect 222403 227848 222522 229030
rect 223646 227848 223768 229030
rect 222403 227745 223768 227848
rect 69791 223180 71156 223290
rect 69791 221998 69910 223180
rect 71034 221998 71156 223180
rect 69791 221895 71156 221998
rect 76708 223178 78073 223288
rect 76708 221996 76827 223178
rect 77951 221996 78073 223178
rect 76708 221893 78073 221996
rect 83673 223179 85038 223289
rect 83673 221997 83792 223179
rect 84916 221997 85038 223179
rect 83673 221894 85038 221997
rect 90631 223180 91996 223290
rect 90631 221998 90750 223180
rect 91874 221998 91996 223180
rect 90631 221895 91996 221998
rect 97449 223159 98814 223269
rect 97449 221977 97568 223159
rect 98692 221977 98814 223159
rect 97449 221874 98814 221977
rect 104414 223160 105779 223270
rect 104414 221978 104533 223160
rect 105657 221978 105779 223160
rect 104414 221875 105779 221978
rect 111372 223161 112737 223271
rect 111372 221979 111491 223161
rect 112615 221979 112737 223161
rect 111372 221876 112737 221979
rect 118292 223160 119657 223270
rect 118292 221978 118411 223160
rect 119535 221978 119657 223160
rect 118292 221875 119657 221978
rect 125257 223161 126622 223271
rect 125257 221979 125376 223161
rect 126500 221979 126622 223161
rect 125257 221876 126622 221979
rect 132215 223162 133580 223272
rect 132215 221980 132334 223162
rect 133458 221980 133580 223162
rect 132215 221877 133580 221980
rect 139132 223166 140497 223276
rect 139132 221984 139251 223166
rect 140375 221984 140497 223166
rect 139132 221881 140497 221984
rect 146097 223167 147462 223277
rect 146097 221985 146216 223167
rect 147340 221985 147462 223167
rect 146097 221882 147462 221985
rect 153055 223168 154420 223278
rect 153055 221986 153174 223168
rect 154298 221986 154420 223168
rect 153055 221883 154420 221986
rect 159972 223166 161337 223276
rect 159972 221984 160091 223166
rect 161215 221984 161337 223166
rect 159972 221881 161337 221984
rect 166937 223167 168302 223277
rect 166937 221985 167056 223167
rect 168180 221985 168302 223167
rect 166937 221882 168302 221985
rect 173895 223168 175260 223278
rect 173895 221986 174014 223168
rect 175138 221986 175260 223168
rect 173895 221883 175260 221986
rect 180700 223161 182065 223271
rect 180700 221979 180819 223161
rect 181943 221979 182065 223161
rect 180700 221876 182065 221979
rect 187665 223162 189030 223272
rect 187665 221980 187784 223162
rect 188908 221980 189030 223162
rect 187665 221877 189030 221980
rect 194623 223163 195988 223273
rect 194623 221981 194742 223163
rect 195866 221981 195988 223163
rect 194623 221878 195988 221981
rect 201543 223162 202908 223272
rect 201543 221980 201662 223162
rect 202786 221980 202908 223162
rect 201543 221877 202908 221980
rect 208508 223163 209873 223273
rect 208508 221981 208627 223163
rect 209751 221981 209873 223163
rect 208508 221878 209873 221981
rect 215466 223164 216831 223274
rect 215466 221982 215585 223164
rect 216709 221982 216831 223164
rect 215466 221879 216831 221982
rect 222383 223168 223748 223278
rect 222383 221986 222502 223168
rect 223626 221986 223748 223168
rect 222383 221883 223748 221986
rect 21190 211109 22555 211219
rect 21190 209927 21309 211109
rect 22433 209927 22555 211109
rect 21190 209824 22555 209927
rect 28148 211110 29513 211220
rect 28148 209928 28267 211110
rect 29391 209928 29513 211110
rect 28148 209825 29513 209928
rect 35068 211109 36433 211219
rect 35068 209927 35187 211109
rect 36311 209927 36433 211109
rect 35068 209824 36433 209927
rect 42033 211110 43398 211220
rect 42033 209928 42152 211110
rect 43276 209928 43398 211110
rect 42033 209825 43398 209928
rect 48991 211111 50356 211221
rect 48991 209929 49110 211111
rect 50234 209929 50356 211111
rect 48991 209826 50356 209929
rect 55908 211115 57273 211225
rect 55908 209933 56027 211115
rect 57151 209933 57273 211115
rect 55908 209830 57273 209933
rect 62873 211116 64238 211226
rect 62873 209934 62992 211116
rect 64116 209934 64238 211116
rect 62873 209831 64238 209934
rect 97489 211096 98854 211206
rect 97489 209914 97608 211096
rect 98732 209914 98854 211096
rect 97489 209811 98854 209914
rect 104454 211097 105819 211207
rect 104454 209915 104573 211097
rect 105697 209915 105819 211097
rect 104454 209812 105819 209915
rect 139172 211103 140537 211213
rect 139172 209921 139291 211103
rect 140415 209921 140537 211103
rect 139172 209818 140537 209921
rect 146137 211104 147502 211214
rect 146137 209922 146256 211104
rect 147380 209922 147502 211104
rect 146137 209819 147502 209922
rect 153095 211105 154460 211215
rect 153095 209923 153214 211105
rect 154338 209923 154460 211105
rect 153095 209820 154460 209923
rect 160012 211103 161377 211213
rect 160012 209921 160131 211103
rect 161255 209921 161377 211103
rect 160012 209818 161377 209921
rect 166977 211104 168342 211214
rect 166977 209922 167096 211104
rect 168220 209922 168342 211104
rect 166977 209819 168342 209922
rect 264326 211107 265691 211217
rect 264326 209925 264445 211107
rect 265569 209925 265691 211107
rect 264326 209822 265691 209925
rect 271284 211108 272649 211218
rect 271284 209926 271403 211108
rect 272527 209926 272649 211108
rect 271284 209823 272649 209926
rect 20916 203979 22281 204089
rect 20916 202797 21035 203979
rect 22159 202797 22281 203979
rect 20916 202694 22281 202797
rect 27874 203980 29239 204090
rect 27874 202798 27993 203980
rect 29117 202798 29239 203980
rect 27874 202695 29239 202798
rect 34794 203979 36159 204089
rect 34794 202797 34913 203979
rect 36037 202797 36159 203979
rect 34794 202694 36159 202797
rect 41759 203980 43124 204090
rect 41759 202798 41878 203980
rect 43002 202798 43124 203980
rect 41759 202695 43124 202798
rect 48717 203981 50082 204091
rect 48717 202799 48836 203981
rect 49960 202799 50082 203981
rect 48717 202696 50082 202799
rect 55634 203985 56999 204095
rect 55634 202803 55753 203985
rect 56877 202803 56999 203985
rect 55634 202700 56999 202803
rect 62599 203986 63964 204096
rect 62599 202804 62718 203986
rect 63842 202804 63964 203986
rect 62599 202701 63964 202804
rect 97215 203966 98580 204076
rect 97215 202784 97334 203966
rect 98458 202784 98580 203966
rect 97215 202681 98580 202784
rect 104180 203967 105545 204077
rect 104180 202785 104299 203967
rect 105423 202785 105545 203967
rect 104180 202682 105545 202785
rect 138898 203973 140263 204083
rect 138898 202791 139017 203973
rect 140141 202791 140263 203973
rect 138898 202688 140263 202791
rect 145863 203974 147228 204084
rect 145863 202792 145982 203974
rect 147106 202792 147228 203974
rect 145863 202689 147228 202792
rect 152821 203975 154186 204085
rect 152821 202793 152940 203975
rect 154064 202793 154186 203975
rect 152821 202690 154186 202793
rect 159738 203973 161103 204083
rect 159738 202791 159857 203973
rect 160981 202791 161103 203973
rect 159738 202688 161103 202791
rect 166703 203974 168068 204084
rect 166703 202792 166822 203974
rect 167946 202792 168068 203974
rect 166703 202689 168068 202792
rect 264052 203977 265417 204087
rect 264052 202795 264171 203977
rect 265295 202795 265417 203977
rect 264052 202692 265417 202795
rect 271010 203978 272375 204088
rect 271010 202796 271129 203978
rect 272253 202796 272375 203978
rect 271010 202693 272375 202796
rect 21024 197566 22389 197676
rect 21024 196384 21143 197566
rect 22267 196384 22389 197566
rect 21024 196281 22389 196384
rect 27982 197567 29347 197677
rect 27982 196385 28101 197567
rect 29225 196385 29347 197567
rect 27982 196282 29347 196385
rect 34902 197566 36267 197676
rect 34902 196384 35021 197566
rect 36145 196384 36267 197566
rect 34902 196281 36267 196384
rect 41867 197567 43232 197677
rect 41867 196385 41986 197567
rect 43110 196385 43232 197567
rect 41867 196282 43232 196385
rect 48825 197568 50190 197678
rect 48825 196386 48944 197568
rect 50068 196386 50190 197568
rect 48825 196283 50190 196386
rect 55742 197572 57107 197682
rect 55742 196390 55861 197572
rect 56985 196390 57107 197572
rect 55742 196287 57107 196390
rect 62707 197573 64072 197683
rect 62707 196391 62826 197573
rect 63950 196391 64072 197573
rect 62707 196288 64072 196391
rect 97323 197553 98688 197663
rect 97323 196371 97442 197553
rect 98566 196371 98688 197553
rect 97323 196268 98688 196371
rect 104288 197554 105653 197664
rect 104288 196372 104407 197554
rect 105531 196372 105653 197554
rect 104288 196269 105653 196372
rect 139006 197560 140371 197670
rect 139006 196378 139125 197560
rect 140249 196378 140371 197560
rect 139006 196275 140371 196378
rect 145971 197561 147336 197671
rect 145971 196379 146090 197561
rect 147214 196379 147336 197561
rect 145971 196276 147336 196379
rect 152929 197562 154294 197672
rect 152929 196380 153048 197562
rect 154172 196380 154294 197562
rect 152929 196277 154294 196380
rect 159846 197560 161211 197670
rect 159846 196378 159965 197560
rect 161089 196378 161211 197560
rect 159846 196275 161211 196378
rect 166811 197561 168176 197671
rect 166811 196379 166930 197561
rect 168054 196379 168176 197561
rect 166811 196276 168176 196379
rect 264160 197564 265525 197674
rect 264160 196382 264279 197564
rect 265403 196382 265525 197564
rect 264160 196279 265525 196382
rect 271118 197565 272483 197675
rect 271118 196383 271237 197565
rect 272361 196383 272483 197565
rect 271118 196280 272483 196383
rect 97476 193203 98841 193313
rect 97476 192021 97595 193203
rect 98719 192021 98841 193203
rect 97476 191918 98841 192021
rect 104441 193204 105806 193314
rect 104441 192022 104560 193204
rect 105684 192022 105806 193204
rect 104441 191919 105806 192022
rect 139159 193210 140524 193320
rect 139159 192028 139278 193210
rect 140402 192028 140524 193210
rect 139159 191925 140524 192028
rect 146124 193211 147489 193321
rect 146124 192029 146243 193211
rect 147367 192029 147489 193211
rect 146124 191926 147489 192029
rect 153082 193212 154447 193322
rect 153082 192030 153201 193212
rect 154325 192030 154447 193212
rect 153082 191927 154447 192030
rect 159999 193210 161364 193320
rect 159999 192028 160118 193210
rect 161242 192028 161364 193210
rect 159999 191925 161364 192028
rect 166964 193211 168329 193321
rect 166964 192029 167083 193211
rect 168207 192029 168329 193211
rect 166964 191926 168329 192029
rect 264313 193214 265678 193324
rect 264313 192032 264432 193214
rect 265556 192032 265678 193214
rect 264313 191929 265678 192032
rect 271271 193215 272636 193325
rect 271271 192033 271390 193215
rect 272514 192033 272636 193215
rect 271271 191930 272636 192033
rect 76461 186092 77826 186202
rect 76461 184910 76580 186092
rect 77704 184910 77826 186092
rect 76461 184807 77826 184910
rect 83426 186093 84791 186203
rect 83426 184911 83545 186093
rect 84669 184911 84791 186093
rect 83426 184808 84791 184911
rect 90384 186094 91749 186204
rect 90384 184912 90503 186094
rect 91627 184912 91749 186094
rect 90384 184809 91749 184912
rect 97202 186073 98567 186183
rect 97202 184891 97321 186073
rect 98445 184891 98567 186073
rect 97202 184788 98567 184891
rect 104167 186074 105532 186184
rect 104167 184892 104286 186074
rect 105410 184892 105532 186074
rect 104167 184789 105532 184892
rect 138885 186080 140250 186190
rect 138885 184898 139004 186080
rect 140128 184898 140250 186080
rect 138885 184795 140250 184898
rect 145850 186081 147215 186191
rect 145850 184899 145969 186081
rect 147093 184899 147215 186081
rect 145850 184796 147215 184899
rect 152808 186082 154173 186192
rect 152808 184900 152927 186082
rect 154051 184900 154173 186082
rect 152808 184797 154173 184900
rect 159725 186080 161090 186190
rect 159725 184898 159844 186080
rect 160968 184898 161090 186080
rect 159725 184795 161090 184898
rect 166690 186081 168055 186191
rect 166690 184899 166809 186081
rect 167933 184899 168055 186081
rect 166690 184796 168055 184899
rect 173648 186082 175013 186192
rect 173648 184900 173767 186082
rect 174891 184900 175013 186082
rect 173648 184797 175013 184900
rect 180453 186075 181818 186185
rect 180453 184893 180572 186075
rect 181696 184893 181818 186075
rect 180453 184790 181818 184893
rect 187418 186076 188783 186186
rect 187418 184894 187537 186076
rect 188661 184894 188783 186076
rect 187418 184791 188783 184894
rect 194376 186077 195741 186187
rect 194376 184895 194495 186077
rect 195619 184895 195741 186077
rect 194376 184792 195741 184895
rect 201296 186076 202661 186186
rect 201296 184894 201415 186076
rect 202539 184894 202661 186076
rect 201296 184791 202661 184894
rect 208261 186077 209626 186187
rect 208261 184895 208380 186077
rect 209504 184895 209626 186077
rect 208261 184792 209626 184895
rect 215219 186078 216584 186188
rect 215219 184896 215338 186078
rect 216462 184896 216584 186078
rect 215219 184793 216584 184896
rect 222136 186082 223501 186192
rect 222136 184900 222255 186082
rect 223379 184900 223501 186082
rect 222136 184797 223501 184900
rect 229101 186083 230466 186193
rect 229101 184901 229220 186083
rect 230344 184901 230466 186083
rect 229101 184798 230466 184901
rect 236059 186084 237424 186194
rect 236059 184902 236178 186084
rect 237302 184902 237424 186084
rect 236059 184799 237424 184902
rect 242976 186082 244341 186192
rect 242976 184900 243095 186082
rect 244219 184900 244341 186082
rect 242976 184797 244341 184900
rect 249941 186083 251306 186193
rect 249941 184901 250060 186083
rect 251184 184901 251306 186083
rect 249941 184798 251306 184901
rect 256899 186084 258264 186194
rect 256899 184902 257018 186084
rect 258142 184902 258264 186084
rect 256899 184799 258264 184902
rect 264039 186084 265404 186194
rect 264039 184902 264158 186084
rect 265282 184902 265404 186084
rect 264039 184799 265404 184902
rect 270997 186085 272362 186195
rect 270997 184903 271116 186085
rect 272240 184903 272362 186085
rect 270997 184800 272362 184903
rect 278133 186075 279498 186185
rect 278133 184893 278252 186075
rect 279376 184893 279498 186075
rect 278133 184790 279498 184893
rect 76569 179679 77934 179789
rect 76569 178497 76688 179679
rect 77812 178497 77934 179679
rect 76569 178394 77934 178497
rect 83534 179680 84899 179790
rect 83534 178498 83653 179680
rect 84777 178498 84899 179680
rect 83534 178395 84899 178498
rect 90492 179681 91857 179791
rect 90492 178499 90611 179681
rect 91735 178499 91857 179681
rect 90492 178396 91857 178499
rect 97310 179660 98675 179770
rect 97310 178478 97429 179660
rect 98553 178478 98675 179660
rect 97310 178375 98675 178478
rect 104275 179661 105640 179771
rect 104275 178479 104394 179661
rect 105518 178479 105640 179661
rect 104275 178376 105640 178479
rect 111233 179662 112598 179772
rect 111233 178480 111352 179662
rect 112476 178480 112598 179662
rect 111233 178377 112598 178480
rect 118153 179661 119518 179771
rect 118153 178479 118272 179661
rect 119396 178479 119518 179661
rect 118153 178376 119518 178479
rect 125118 179662 126483 179772
rect 125118 178480 125237 179662
rect 126361 178480 126483 179662
rect 125118 178377 126483 178480
rect 132076 179663 133441 179773
rect 132076 178481 132195 179663
rect 133319 178481 133441 179663
rect 132076 178378 133441 178481
rect 138993 179667 140358 179777
rect 138993 178485 139112 179667
rect 140236 178485 140358 179667
rect 138993 178382 140358 178485
rect 145958 179668 147323 179778
rect 145958 178486 146077 179668
rect 147201 178486 147323 179668
rect 145958 178383 147323 178486
rect 152916 179669 154281 179779
rect 152916 178487 153035 179669
rect 154159 178487 154281 179669
rect 152916 178384 154281 178487
rect 159833 179667 161198 179777
rect 159833 178485 159952 179667
rect 161076 178485 161198 179667
rect 159833 178382 161198 178485
rect 166798 179668 168163 179778
rect 166798 178486 166917 179668
rect 168041 178486 168163 179668
rect 166798 178383 168163 178486
rect 173756 179669 175121 179779
rect 173756 178487 173875 179669
rect 174999 178487 175121 179669
rect 173756 178384 175121 178487
rect 180561 179662 181926 179772
rect 180561 178480 180680 179662
rect 181804 178480 181926 179662
rect 180561 178377 181926 178480
rect 187526 179663 188891 179773
rect 187526 178481 187645 179663
rect 188769 178481 188891 179663
rect 187526 178378 188891 178481
rect 194484 179664 195849 179774
rect 194484 178482 194603 179664
rect 195727 178482 195849 179664
rect 194484 178379 195849 178482
rect 201404 179663 202769 179773
rect 201404 178481 201523 179663
rect 202647 178481 202769 179663
rect 201404 178378 202769 178481
rect 208369 179664 209734 179774
rect 208369 178482 208488 179664
rect 209612 178482 209734 179664
rect 208369 178379 209734 178482
rect 215327 179665 216692 179775
rect 215327 178483 215446 179665
rect 216570 178483 216692 179665
rect 215327 178380 216692 178483
rect 222244 179669 223609 179779
rect 222244 178487 222363 179669
rect 223487 178487 223609 179669
rect 222244 178384 223609 178487
rect 229209 179670 230574 179780
rect 229209 178488 229328 179670
rect 230452 178488 230574 179670
rect 229209 178385 230574 178488
rect 236167 179671 237532 179781
rect 236167 178489 236286 179671
rect 237410 178489 237532 179671
rect 236167 178386 237532 178489
rect 243084 179669 244449 179779
rect 243084 178487 243203 179669
rect 244327 178487 244449 179669
rect 243084 178384 244449 178487
rect 250049 179670 251414 179780
rect 250049 178488 250168 179670
rect 251292 178488 251414 179670
rect 250049 178385 251414 178488
rect 257007 179671 258372 179781
rect 257007 178489 257126 179671
rect 258250 178489 258372 179671
rect 257007 178386 258372 178489
rect 264147 179671 265512 179781
rect 264147 178489 264266 179671
rect 265390 178489 265512 179671
rect 264147 178386 265512 178489
rect 271105 179672 272470 179782
rect 271105 178490 271224 179672
rect 272348 178490 272470 179672
rect 271105 178387 272470 178490
rect 278241 179662 279606 179772
rect 278241 178480 278360 179662
rect 279484 178480 279606 179662
rect 278241 178377 279606 178480
rect 69367 173767 70732 173877
rect 69367 172585 69486 173767
rect 70610 172585 70732 173767
rect 69367 172482 70732 172585
rect 76284 173765 77649 173875
rect 76284 172583 76403 173765
rect 77527 172583 77649 173765
rect 76284 172480 77649 172583
rect 83249 173766 84614 173876
rect 83249 172584 83368 173766
rect 84492 172584 84614 173766
rect 83249 172481 84614 172584
rect 90207 173767 91572 173877
rect 90207 172585 90326 173767
rect 91450 172585 91572 173767
rect 90207 172482 91572 172585
rect 97025 173746 98390 173856
rect 97025 172564 97144 173746
rect 98268 172564 98390 173746
rect 97025 172461 98390 172564
rect 103990 173747 105355 173857
rect 103990 172565 104109 173747
rect 105233 172565 105355 173747
rect 103990 172462 105355 172565
rect 110948 173748 112313 173858
rect 110948 172566 111067 173748
rect 112191 172566 112313 173748
rect 110948 172463 112313 172566
rect 117868 173747 119233 173857
rect 117868 172565 117987 173747
rect 119111 172565 119233 173747
rect 117868 172462 119233 172565
rect 124833 173748 126198 173858
rect 124833 172566 124952 173748
rect 126076 172566 126198 173748
rect 124833 172463 126198 172566
rect 131791 173749 133156 173859
rect 131791 172567 131910 173749
rect 133034 172567 133156 173749
rect 131791 172464 133156 172567
rect 138708 173753 140073 173863
rect 138708 172571 138827 173753
rect 139951 172571 140073 173753
rect 138708 172468 140073 172571
rect 145673 173754 147038 173864
rect 145673 172572 145792 173754
rect 146916 172572 147038 173754
rect 145673 172469 147038 172572
rect 152631 173755 153996 173865
rect 152631 172573 152750 173755
rect 153874 172573 153996 173755
rect 152631 172470 153996 172573
rect 159548 173753 160913 173863
rect 159548 172571 159667 173753
rect 160791 172571 160913 173753
rect 159548 172468 160913 172571
rect 166513 173754 167878 173864
rect 166513 172572 166632 173754
rect 167756 172572 167878 173754
rect 166513 172469 167878 172572
rect 173471 173755 174836 173865
rect 173471 172573 173590 173755
rect 174714 172573 174836 173755
rect 173471 172470 174836 172573
rect 180276 173748 181641 173858
rect 180276 172566 180395 173748
rect 181519 172566 181641 173748
rect 180276 172463 181641 172566
rect 187241 173749 188606 173859
rect 187241 172567 187360 173749
rect 188484 172567 188606 173749
rect 187241 172464 188606 172567
rect 194199 173750 195564 173860
rect 194199 172568 194318 173750
rect 195442 172568 195564 173750
rect 194199 172465 195564 172568
rect 201119 173749 202484 173859
rect 201119 172567 201238 173749
rect 202362 172567 202484 173749
rect 201119 172464 202484 172567
rect 208084 173750 209449 173860
rect 208084 172568 208203 173750
rect 209327 172568 209449 173750
rect 208084 172465 209449 172568
rect 215042 173751 216407 173861
rect 215042 172569 215161 173751
rect 216285 172569 216407 173751
rect 215042 172466 216407 172569
rect 221959 173755 223324 173865
rect 221959 172573 222078 173755
rect 223202 172573 223324 173755
rect 221959 172470 223324 172573
rect 228924 173756 230289 173866
rect 228924 172574 229043 173756
rect 230167 172574 230289 173756
rect 228924 172471 230289 172574
rect 235882 173757 237247 173867
rect 235882 172575 236001 173757
rect 237125 172575 237247 173757
rect 235882 172472 237247 172575
rect 242799 173755 244164 173865
rect 242799 172573 242918 173755
rect 244042 172573 244164 173755
rect 242799 172470 244164 172573
rect 249764 173756 251129 173866
rect 249764 172574 249883 173756
rect 251007 172574 251129 173756
rect 249764 172471 251129 172574
rect 256722 173757 258087 173867
rect 256722 172575 256841 173757
rect 257965 172575 258087 173757
rect 256722 172472 258087 172575
rect 263862 173757 265227 173867
rect 263862 172575 263981 173757
rect 265105 172575 265227 173757
rect 263862 172472 265227 172575
rect 270820 173758 272185 173868
rect 270820 172576 270939 173758
rect 272063 172576 272185 173758
rect 270820 172473 272185 172576
rect 277956 173748 279321 173858
rect 277956 172566 278075 173748
rect 279199 172566 279321 173748
rect 277956 172463 279321 172566
rect 69475 167354 70840 167464
rect 69475 166172 69594 167354
rect 70718 166172 70840 167354
rect 69475 166069 70840 166172
rect 76392 167352 77757 167462
rect 76392 166170 76511 167352
rect 77635 166170 77757 167352
rect 76392 166067 77757 166170
rect 83357 167353 84722 167463
rect 83357 166171 83476 167353
rect 84600 166171 84722 167353
rect 83357 166068 84722 166171
rect 90315 167354 91680 167464
rect 90315 166172 90434 167354
rect 91558 166172 91680 167354
rect 90315 166069 91680 166172
rect 97133 167333 98498 167443
rect 97133 166151 97252 167333
rect 98376 166151 98498 167333
rect 97133 166048 98498 166151
rect 104098 167334 105463 167444
rect 104098 166152 104217 167334
rect 105341 166152 105463 167334
rect 104098 166049 105463 166152
rect 111056 167335 112421 167445
rect 111056 166153 111175 167335
rect 112299 166153 112421 167335
rect 111056 166050 112421 166153
rect 117976 167334 119341 167444
rect 117976 166152 118095 167334
rect 119219 166152 119341 167334
rect 117976 166049 119341 166152
rect 124941 167335 126306 167445
rect 124941 166153 125060 167335
rect 126184 166153 126306 167335
rect 124941 166050 126306 166153
rect 131899 167336 133264 167446
rect 131899 166154 132018 167336
rect 133142 166154 133264 167336
rect 131899 166051 133264 166154
rect 138816 167340 140181 167450
rect 138816 166158 138935 167340
rect 140059 166158 140181 167340
rect 138816 166055 140181 166158
rect 145781 167341 147146 167451
rect 145781 166159 145900 167341
rect 147024 166159 147146 167341
rect 145781 166056 147146 166159
rect 152739 167342 154104 167452
rect 152739 166160 152858 167342
rect 153982 166160 154104 167342
rect 152739 166057 154104 166160
rect 159656 167340 161021 167450
rect 159656 166158 159775 167340
rect 160899 166158 161021 167340
rect 159656 166055 161021 166158
rect 166621 167341 167986 167451
rect 166621 166159 166740 167341
rect 167864 166159 167986 167341
rect 166621 166056 167986 166159
rect 173579 167342 174944 167452
rect 173579 166160 173698 167342
rect 174822 166160 174944 167342
rect 173579 166057 174944 166160
rect 180384 167335 181749 167445
rect 180384 166153 180503 167335
rect 181627 166153 181749 167335
rect 180384 166050 181749 166153
rect 187349 167336 188714 167446
rect 187349 166154 187468 167336
rect 188592 166154 188714 167336
rect 187349 166051 188714 166154
rect 194307 167337 195672 167447
rect 194307 166155 194426 167337
rect 195550 166155 195672 167337
rect 194307 166052 195672 166155
rect 201227 167336 202592 167446
rect 201227 166154 201346 167336
rect 202470 166154 202592 167336
rect 201227 166051 202592 166154
rect 208192 167337 209557 167447
rect 208192 166155 208311 167337
rect 209435 166155 209557 167337
rect 208192 166052 209557 166155
rect 215150 167338 216515 167448
rect 215150 166156 215269 167338
rect 216393 166156 216515 167338
rect 215150 166053 216515 166156
rect 222067 167342 223432 167452
rect 222067 166160 222186 167342
rect 223310 166160 223432 167342
rect 222067 166057 223432 166160
rect 229032 167343 230397 167453
rect 229032 166161 229151 167343
rect 230275 166161 230397 167343
rect 229032 166058 230397 166161
rect 235990 167344 237355 167454
rect 235990 166162 236109 167344
rect 237233 166162 237355 167344
rect 235990 166059 237355 166162
rect 242907 167342 244272 167452
rect 242907 166160 243026 167342
rect 244150 166160 244272 167342
rect 242907 166057 244272 166160
rect 249872 167343 251237 167453
rect 249872 166161 249991 167343
rect 251115 166161 251237 167343
rect 249872 166058 251237 166161
rect 256830 167344 258195 167454
rect 256830 166162 256949 167344
rect 258073 166162 258195 167344
rect 256830 166059 258195 166162
rect 263970 167344 265335 167454
rect 263970 166162 264089 167344
rect 265213 166162 265335 167344
rect 263970 166059 265335 166162
rect 270928 167345 272293 167455
rect 270928 166163 271047 167345
rect 272171 166163 272293 167345
rect 270928 166060 272293 166163
rect 278064 167335 279429 167445
rect 278064 166153 278183 167335
rect 279307 166153 279429 167335
rect 278064 166050 279429 166153
rect 21601 160007 22966 160117
rect 21601 158825 21720 160007
rect 22844 158825 22966 160007
rect 21601 158722 22966 158825
rect 28559 160008 29924 160118
rect 28559 158826 28678 160008
rect 29802 158826 29924 160008
rect 28559 158723 29924 158826
rect 35479 160007 36844 160117
rect 35479 158825 35598 160007
rect 36722 158825 36844 160007
rect 35479 158722 36844 158825
rect 56319 160013 57684 160123
rect 56319 158831 56438 160013
rect 57562 158831 57684 160013
rect 56319 158728 57684 158831
rect 63284 160014 64649 160124
rect 63284 158832 63403 160014
rect 64527 158832 64649 160014
rect 63284 158729 64649 158832
rect 97900 159994 99265 160104
rect 97900 158812 98019 159994
rect 99143 158812 99265 159994
rect 97900 158709 99265 158812
rect 104865 159995 106230 160105
rect 104865 158813 104984 159995
rect 106108 158813 106230 159995
rect 104865 158710 106230 158813
rect 139583 160001 140948 160111
rect 139583 158819 139702 160001
rect 140826 158819 140948 160001
rect 139583 158716 140948 158819
rect 146548 160002 147913 160112
rect 146548 158820 146667 160002
rect 147791 158820 147913 160002
rect 146548 158717 147913 158820
rect 153506 160003 154871 160113
rect 153506 158821 153625 160003
rect 154749 158821 154871 160003
rect 153506 158718 154871 158821
rect 160423 160001 161788 160111
rect 160423 158819 160542 160001
rect 161666 158819 161788 160001
rect 160423 158716 161788 158819
rect 167388 160002 168753 160112
rect 167388 158820 167507 160002
rect 168631 158820 168753 160002
rect 167388 158717 168753 158820
rect 188116 159997 189481 160107
rect 188116 158815 188235 159997
rect 189359 158815 189481 159997
rect 188116 158712 189481 158815
rect 195074 159998 196439 160108
rect 195074 158816 195193 159998
rect 196317 158816 196439 159998
rect 195074 158713 196439 158816
rect 229673 159998 231038 160108
rect 229673 158816 229792 159998
rect 230916 158816 231038 159998
rect 229673 158713 231038 158816
rect 236638 159999 238003 160109
rect 236638 158817 236757 159999
rect 237881 158817 238003 159999
rect 236638 158714 238003 158817
rect 243596 160000 244961 160110
rect 243596 158818 243715 160000
rect 244839 158818 244961 160000
rect 243596 158715 244961 158818
rect 250513 160004 251878 160114
rect 250513 158822 250632 160004
rect 251756 158822 251878 160004
rect 250513 158719 251878 158822
rect 257405 159987 258770 160097
rect 257405 158805 257524 159987
rect 258648 158805 258770 159987
rect 257405 158702 258770 158805
rect 264370 159988 265735 160098
rect 264370 158806 264489 159988
rect 265613 158806 265735 159988
rect 264370 158703 265735 158806
rect 271328 159989 272693 160099
rect 271328 158807 271447 159989
rect 272571 158807 272693 159989
rect 271328 158704 272693 158807
rect 278245 159993 279610 160103
rect 278245 158811 278364 159993
rect 279488 158811 279610 159993
rect 278245 158708 279610 158811
rect 21886 155174 23251 155284
rect 21886 153992 22005 155174
rect 23129 153992 23251 155174
rect 21886 153889 23251 153992
rect 28844 155175 30209 155285
rect 28844 153993 28963 155175
rect 30087 153993 30209 155175
rect 28844 153890 30209 153993
rect 35764 155174 37129 155284
rect 35764 153992 35883 155174
rect 37007 153992 37129 155174
rect 35764 153889 37129 153992
rect 56604 155180 57969 155290
rect 56604 153998 56723 155180
rect 57847 153998 57969 155180
rect 56604 153895 57969 153998
rect 63569 155181 64934 155291
rect 63569 153999 63688 155181
rect 64812 153999 64934 155181
rect 63569 153896 64934 153999
rect 98185 155161 99550 155271
rect 98185 153979 98304 155161
rect 99428 153979 99550 155161
rect 98185 153876 99550 153979
rect 105150 155162 106515 155272
rect 105150 153980 105269 155162
rect 106393 153980 106515 155162
rect 105150 153877 106515 153980
rect 139868 155168 141233 155278
rect 139868 153986 139987 155168
rect 141111 153986 141233 155168
rect 139868 153883 141233 153986
rect 146833 155169 148198 155279
rect 146833 153987 146952 155169
rect 148076 153987 148198 155169
rect 146833 153884 148198 153987
rect 153791 155170 155156 155280
rect 153791 153988 153910 155170
rect 155034 153988 155156 155170
rect 153791 153885 155156 153988
rect 160708 155168 162073 155278
rect 160708 153986 160827 155168
rect 161951 153986 162073 155168
rect 160708 153883 162073 153986
rect 167673 155169 169038 155279
rect 167673 153987 167792 155169
rect 168916 153987 169038 155169
rect 167673 153884 169038 153987
rect 188401 155164 189766 155274
rect 188401 153982 188520 155164
rect 189644 153982 189766 155164
rect 188401 153879 189766 153982
rect 195359 155165 196724 155275
rect 195359 153983 195478 155165
rect 196602 153983 196724 155165
rect 195359 153880 196724 153983
rect 229958 155165 231323 155275
rect 229958 153983 230077 155165
rect 231201 153983 231323 155165
rect 229958 153880 231323 153983
rect 236923 155166 238288 155276
rect 236923 153984 237042 155166
rect 238166 153984 238288 155166
rect 236923 153881 238288 153984
rect 243881 155167 245246 155277
rect 243881 153985 244000 155167
rect 245124 153985 245246 155167
rect 243881 153882 245246 153985
rect 250798 155171 252163 155281
rect 250798 153989 250917 155171
rect 252041 153989 252163 155171
rect 250798 153886 252163 153989
rect 257690 155154 259055 155264
rect 257690 153972 257809 155154
rect 258933 153972 259055 155154
rect 257690 153869 259055 153972
rect 264655 155155 266020 155265
rect 264655 153973 264774 155155
rect 265898 153973 266020 155155
rect 264655 153870 266020 153973
rect 271613 155156 272978 155266
rect 271613 153974 271732 155156
rect 272856 153974 272978 155156
rect 271613 153871 272978 153974
rect 278530 155160 279895 155270
rect 278530 153978 278649 155160
rect 279773 153978 279895 155160
rect 278530 153875 279895 153978
rect 21957 149914 23322 150024
rect 21957 148732 22076 149914
rect 23200 148732 23322 149914
rect 21957 148629 23322 148732
rect 28915 149915 30280 150025
rect 28915 148733 29034 149915
rect 30158 148733 30280 149915
rect 28915 148630 30280 148733
rect 35835 149914 37200 150024
rect 35835 148732 35954 149914
rect 37078 148732 37200 149914
rect 35835 148629 37200 148732
rect 56675 149920 58040 150030
rect 56675 148738 56794 149920
rect 57918 148738 58040 149920
rect 56675 148635 58040 148738
rect 63640 149921 65005 150031
rect 63640 148739 63759 149921
rect 64883 148739 65005 149921
rect 63640 148636 65005 148739
rect 98256 149901 99621 150011
rect 98256 148719 98375 149901
rect 99499 148719 99621 149901
rect 98256 148616 99621 148719
rect 105221 149902 106586 150012
rect 105221 148720 105340 149902
rect 106464 148720 106586 149902
rect 105221 148617 106586 148720
rect 139939 149908 141304 150018
rect 139939 148726 140058 149908
rect 141182 148726 141304 149908
rect 139939 148623 141304 148726
rect 146904 149909 148269 150019
rect 146904 148727 147023 149909
rect 148147 148727 148269 149909
rect 146904 148624 148269 148727
rect 153862 149910 155227 150020
rect 153862 148728 153981 149910
rect 155105 148728 155227 149910
rect 153862 148625 155227 148728
rect 160779 149908 162144 150018
rect 160779 148726 160898 149908
rect 162022 148726 162144 149908
rect 160779 148623 162144 148726
rect 167744 149909 169109 150019
rect 167744 148727 167863 149909
rect 168987 148727 169109 149909
rect 167744 148624 169109 148727
rect 188472 149904 189837 150014
rect 188472 148722 188591 149904
rect 189715 148722 189837 149904
rect 188472 148619 189837 148722
rect 195430 149905 196795 150015
rect 195430 148723 195549 149905
rect 196673 148723 196795 149905
rect 195430 148620 196795 148723
rect 230029 149905 231394 150015
rect 230029 148723 230148 149905
rect 231272 148723 231394 149905
rect 230029 148620 231394 148723
rect 236994 149906 238359 150016
rect 236994 148724 237113 149906
rect 238237 148724 238359 149906
rect 236994 148621 238359 148724
rect 243952 149907 245317 150017
rect 243952 148725 244071 149907
rect 245195 148725 245317 149907
rect 243952 148622 245317 148725
rect 250869 149911 252234 150021
rect 250869 148729 250988 149911
rect 252112 148729 252234 149911
rect 250869 148626 252234 148729
rect 257761 149894 259126 150004
rect 257761 148712 257880 149894
rect 259004 148712 259126 149894
rect 257761 148609 259126 148712
rect 264726 149895 266091 150005
rect 264726 148713 264845 149895
rect 265969 148713 266091 149895
rect 264726 148610 266091 148713
rect 271684 149896 273049 150006
rect 271684 148714 271803 149896
rect 272927 148714 273049 149896
rect 271684 148611 273049 148714
rect 278601 149900 279966 150010
rect 278601 148718 278720 149900
rect 279844 148718 279966 149900
rect 278601 148615 279966 148718
rect 21886 144440 23251 144550
rect 21886 143258 22005 144440
rect 23129 143258 23251 144440
rect 21886 143155 23251 143258
rect 28844 144441 30209 144551
rect 28844 143259 28963 144441
rect 30087 143259 30209 144441
rect 28844 143156 30209 143259
rect 35764 144440 37129 144550
rect 35764 143258 35883 144440
rect 37007 143258 37129 144440
rect 35764 143155 37129 143258
rect 56604 144446 57969 144556
rect 56604 143264 56723 144446
rect 57847 143264 57969 144446
rect 56604 143161 57969 143264
rect 63569 144447 64934 144557
rect 63569 143265 63688 144447
rect 64812 143265 64934 144447
rect 63569 143162 64934 143265
rect 98185 144427 99550 144537
rect 98185 143245 98304 144427
rect 99428 143245 99550 144427
rect 98185 143142 99550 143245
rect 105150 144428 106515 144538
rect 105150 143246 105269 144428
rect 106393 143246 106515 144428
rect 105150 143143 106515 143246
rect 139868 144434 141233 144544
rect 139868 143252 139987 144434
rect 141111 143252 141233 144434
rect 139868 143149 141233 143252
rect 146833 144435 148198 144545
rect 146833 143253 146952 144435
rect 148076 143253 148198 144435
rect 146833 143150 148198 143253
rect 153791 144436 155156 144546
rect 153791 143254 153910 144436
rect 155034 143254 155156 144436
rect 153791 143151 155156 143254
rect 160708 144434 162073 144544
rect 160708 143252 160827 144434
rect 161951 143252 162073 144434
rect 160708 143149 162073 143252
rect 167673 144435 169038 144545
rect 167673 143253 167792 144435
rect 168916 143253 169038 144435
rect 167673 143150 169038 143253
rect 188401 144430 189766 144540
rect 188401 143248 188520 144430
rect 189644 143248 189766 144430
rect 188401 143145 189766 143248
rect 195359 144431 196724 144541
rect 195359 143249 195478 144431
rect 196602 143249 196724 144431
rect 195359 143146 196724 143249
rect 22028 138328 23393 138438
rect 22028 137146 22147 138328
rect 23271 137146 23393 138328
rect 22028 137043 23393 137146
rect 28986 138329 30351 138439
rect 28986 137147 29105 138329
rect 30229 137147 30351 138329
rect 28986 137044 30351 137147
rect 35906 138328 37271 138438
rect 35906 137146 36025 138328
rect 37149 137146 37271 138328
rect 35906 137043 37271 137146
rect 56746 138334 58111 138444
rect 56746 137152 56865 138334
rect 57989 137152 58111 138334
rect 56746 137049 58111 137152
rect 63711 138335 65076 138445
rect 63711 137153 63830 138335
rect 64954 137153 65076 138335
rect 63711 137050 65076 137153
rect 98327 138315 99692 138425
rect 98327 137133 98446 138315
rect 99570 137133 99692 138315
rect 98327 137030 99692 137133
rect 105292 138316 106657 138426
rect 105292 137134 105411 138316
rect 106535 137134 106657 138316
rect 105292 137031 106657 137134
rect 140010 138322 141375 138432
rect 140010 137140 140129 138322
rect 141253 137140 141375 138322
rect 140010 137037 141375 137140
rect 146975 138323 148340 138433
rect 146975 137141 147094 138323
rect 148218 137141 148340 138323
rect 146975 137038 148340 137141
rect 153933 138324 155298 138434
rect 153933 137142 154052 138324
rect 155176 137142 155298 138324
rect 153933 137039 155298 137142
rect 160850 138322 162215 138432
rect 160850 137140 160969 138322
rect 162093 137140 162215 138322
rect 160850 137037 162215 137140
rect 167815 138323 169180 138433
rect 167815 137141 167934 138323
rect 169058 137141 169180 138323
rect 167815 137038 169180 137141
rect 188543 138318 189908 138428
rect 188543 137136 188662 138318
rect 189786 137136 189908 138318
rect 188543 137033 189908 137136
rect 195501 138319 196866 138429
rect 195501 137137 195620 138319
rect 196744 137137 196866 138319
rect 195501 137034 196866 137137
rect 21818 130454 23183 130564
rect 21818 129272 21937 130454
rect 23061 129272 23183 130454
rect 21818 129169 23183 129272
rect 28776 130455 30141 130565
rect 28776 129273 28895 130455
rect 30019 129273 30141 130455
rect 28776 129170 30141 129273
rect 35696 130454 37061 130564
rect 35696 129272 35815 130454
rect 36939 129272 37061 130454
rect 35696 129169 37061 129272
rect 42661 130455 44026 130565
rect 42661 129273 42780 130455
rect 43904 129273 44026 130455
rect 42661 129170 44026 129273
rect 49619 130456 50984 130566
rect 49619 129274 49738 130456
rect 50862 129274 50984 130456
rect 49619 129171 50984 129274
rect 56536 130460 57901 130570
rect 56536 129278 56655 130460
rect 57779 129278 57901 130460
rect 56536 129175 57901 129278
rect 63501 130461 64866 130571
rect 63501 129279 63620 130461
rect 64744 129279 64866 130461
rect 63501 129176 64866 129279
rect 70459 130462 71824 130572
rect 70459 129280 70578 130462
rect 71702 129280 71824 130462
rect 70459 129177 71824 129280
rect 77376 130460 78741 130570
rect 77376 129278 77495 130460
rect 78619 129278 78741 130460
rect 77376 129175 78741 129278
rect 84341 130461 85706 130571
rect 84341 129279 84460 130461
rect 85584 129279 85706 130461
rect 84341 129176 85706 129279
rect 91299 130462 92664 130572
rect 91299 129280 91418 130462
rect 92542 129280 92664 130462
rect 91299 129177 92664 129280
rect 98117 130441 99482 130551
rect 98117 129259 98236 130441
rect 99360 129259 99482 130441
rect 98117 129156 99482 129259
rect 105082 130442 106447 130552
rect 105082 129260 105201 130442
rect 106325 129260 106447 130442
rect 105082 129157 106447 129260
rect 112040 130443 113405 130553
rect 112040 129261 112159 130443
rect 113283 129261 113405 130443
rect 112040 129158 113405 129261
rect 118960 130442 120325 130552
rect 118960 129260 119079 130442
rect 120203 129260 120325 130442
rect 118960 129157 120325 129260
rect 125925 130443 127290 130553
rect 125925 129261 126044 130443
rect 127168 129261 127290 130443
rect 125925 129158 127290 129261
rect 132883 130444 134248 130554
rect 132883 129262 133002 130444
rect 134126 129262 134248 130444
rect 132883 129159 134248 129262
rect 139800 130448 141165 130558
rect 139800 129266 139919 130448
rect 141043 129266 141165 130448
rect 139800 129163 141165 129266
rect 146765 130449 148130 130559
rect 146765 129267 146884 130449
rect 148008 129267 148130 130449
rect 146765 129164 148130 129267
rect 153723 130450 155088 130560
rect 153723 129268 153842 130450
rect 154966 129268 155088 130450
rect 153723 129165 155088 129268
rect 160640 130448 162005 130558
rect 160640 129266 160759 130448
rect 161883 129266 162005 130448
rect 160640 129163 162005 129266
rect 167605 130449 168970 130559
rect 167605 129267 167724 130449
rect 168848 129267 168970 130449
rect 167605 129164 168970 129267
rect 174563 130450 175928 130560
rect 174563 129268 174682 130450
rect 175806 129268 175928 130450
rect 174563 129165 175928 129268
rect 181368 130443 182733 130553
rect 181368 129261 181487 130443
rect 182611 129261 182733 130443
rect 181368 129158 182733 129261
rect 188333 130444 189698 130554
rect 188333 129262 188452 130444
rect 189576 129262 189698 130444
rect 188333 129159 189698 129262
rect 195291 130445 196656 130555
rect 195291 129263 195410 130445
rect 196534 129263 196656 130445
rect 195291 129160 196656 129263
rect 97634 119125 98999 119235
rect 97634 117943 97753 119125
rect 98877 117943 98999 119125
rect 97634 117840 98999 117943
rect 104599 119126 105964 119236
rect 104599 117944 104718 119126
rect 105842 117944 105964 119126
rect 104599 117841 105964 117944
rect 139317 119132 140682 119242
rect 139317 117950 139436 119132
rect 140560 117950 140682 119132
rect 139317 117847 140682 117950
rect 146282 119133 147647 119243
rect 146282 117951 146401 119133
rect 147525 117951 147647 119133
rect 146282 117848 147647 117951
rect 153240 119134 154605 119244
rect 153240 117952 153359 119134
rect 154483 117952 154605 119134
rect 153240 117849 154605 117952
rect 160157 119132 161522 119242
rect 160157 117950 160276 119132
rect 161400 117950 161522 119132
rect 160157 117847 161522 117950
rect 167122 119133 168487 119243
rect 167122 117951 167241 119133
rect 168365 117951 168487 119133
rect 167122 117848 168487 117951
rect 97839 111173 99204 111283
rect 97839 109991 97958 111173
rect 99082 109991 99204 111173
rect 97839 109888 99204 109991
rect 104804 111174 106169 111284
rect 104804 109992 104923 111174
rect 106047 109992 106169 111174
rect 104804 109889 106169 109992
rect 139522 111180 140887 111290
rect 139522 109998 139641 111180
rect 140765 109998 140887 111180
rect 139522 109895 140887 109998
rect 146487 111181 147852 111291
rect 146487 109999 146606 111181
rect 147730 109999 147852 111181
rect 146487 109896 147852 109999
rect 153445 111182 154810 111292
rect 153445 110000 153564 111182
rect 154688 110000 154810 111182
rect 153445 109897 154810 110000
rect 160362 111180 161727 111290
rect 160362 109998 160481 111180
rect 161605 109998 161727 111180
rect 160362 109895 161727 109998
rect 167327 111181 168692 111291
rect 167327 109999 167446 111181
rect 168570 109999 168692 111181
rect 167327 109896 168692 109999
rect 97839 102947 99204 103057
rect 97839 101765 97958 102947
rect 99082 101765 99204 102947
rect 97839 101662 99204 101765
rect 104804 102948 106169 103058
rect 104804 101766 104923 102948
rect 106047 101766 106169 102948
rect 104804 101663 106169 101766
rect 139522 102954 140887 103064
rect 139522 101772 139641 102954
rect 140765 101772 140887 102954
rect 139522 101669 140887 101772
rect 146487 102955 147852 103065
rect 146487 101773 146606 102955
rect 147730 101773 147852 102955
rect 146487 101670 147852 101773
rect 153445 102956 154810 103066
rect 153445 101774 153564 102956
rect 154688 101774 154810 102956
rect 153445 101671 154810 101774
rect 160362 102954 161727 103064
rect 160362 101772 160481 102954
rect 161605 101772 161727 102954
rect 160362 101669 161727 101772
rect 167327 102955 168692 103065
rect 167327 101773 167446 102955
rect 168570 101773 168692 102955
rect 167327 101670 168692 101773
rect 97634 95543 98999 95653
rect 97634 94361 97753 95543
rect 98877 94361 98999 95543
rect 97634 94258 98999 94361
rect 104599 95544 105964 95654
rect 104599 94362 104718 95544
rect 105842 94362 105964 95544
rect 104599 94259 105964 94362
rect 139317 95550 140682 95660
rect 139317 94368 139436 95550
rect 140560 94368 140682 95550
rect 139317 94265 140682 94368
rect 146282 95551 147647 95661
rect 146282 94369 146401 95551
rect 147525 94369 147647 95551
rect 146282 94266 147647 94369
rect 153240 95552 154605 95662
rect 153240 94370 153359 95552
rect 154483 94370 154605 95552
rect 153240 94267 154605 94370
rect 160157 95550 161522 95660
rect 160157 94368 160276 95550
rect 161400 94368 161522 95550
rect 160157 94265 161522 94368
rect 167122 95551 168487 95661
rect 167122 94369 167241 95551
rect 168365 94369 168487 95551
rect 167122 94266 168487 94369
rect 97360 88413 98725 88523
rect 97360 87231 97479 88413
rect 98603 87231 98725 88413
rect 97360 87128 98725 87231
rect 104325 88414 105690 88524
rect 104325 87232 104444 88414
rect 105568 87232 105690 88414
rect 104325 87129 105690 87232
rect 111283 88415 112648 88525
rect 111283 87233 111402 88415
rect 112526 87233 112648 88415
rect 111283 87130 112648 87233
rect 118203 88414 119568 88524
rect 118203 87232 118322 88414
rect 119446 87232 119568 88414
rect 118203 87129 119568 87232
rect 125168 88415 126533 88525
rect 125168 87233 125287 88415
rect 126411 87233 126533 88415
rect 125168 87130 126533 87233
rect 132126 88416 133491 88526
rect 132126 87234 132245 88416
rect 133369 87234 133491 88416
rect 132126 87131 133491 87234
rect 139043 88420 140408 88530
rect 139043 87238 139162 88420
rect 140286 87238 140408 88420
rect 139043 87135 140408 87238
rect 146008 88421 147373 88531
rect 146008 87239 146127 88421
rect 147251 87239 147373 88421
rect 146008 87136 147373 87239
rect 152966 88422 154331 88532
rect 152966 87240 153085 88422
rect 154209 87240 154331 88422
rect 152966 87137 154331 87240
rect 159883 88420 161248 88530
rect 159883 87238 160002 88420
rect 161126 87238 161248 88420
rect 159883 87135 161248 87238
rect 166848 88421 168213 88531
rect 166848 87239 166967 88421
rect 168091 87239 168213 88421
rect 166848 87136 168213 87239
rect 97468 82000 98833 82110
rect 97468 80818 97587 82000
rect 98711 80818 98833 82000
rect 97468 80715 98833 80818
rect 104433 82001 105798 82111
rect 104433 80819 104552 82001
rect 105676 80819 105798 82001
rect 104433 80716 105798 80819
rect 111391 82002 112756 82112
rect 111391 80820 111510 82002
rect 112634 80820 112756 82002
rect 111391 80717 112756 80820
rect 118311 82001 119676 82111
rect 118311 80819 118430 82001
rect 119554 80819 119676 82001
rect 118311 80716 119676 80819
rect 125276 82002 126641 82112
rect 125276 80820 125395 82002
rect 126519 80820 126641 82002
rect 125276 80717 126641 80820
rect 132234 82003 133599 82113
rect 132234 80821 132353 82003
rect 133477 80821 133599 82003
rect 132234 80718 133599 80821
rect 139151 82007 140516 82117
rect 139151 80825 139270 82007
rect 140394 80825 140516 82007
rect 139151 80722 140516 80825
rect 146116 82008 147481 82118
rect 146116 80826 146235 82008
rect 147359 80826 147481 82008
rect 146116 80723 147481 80826
rect 153074 82009 154439 82119
rect 153074 80827 153193 82009
rect 154317 80827 154439 82009
rect 153074 80724 154439 80827
rect 159991 82007 161356 82117
rect 159991 80825 160110 82007
rect 161234 80825 161356 82007
rect 159991 80722 161356 80825
rect 166956 82008 168321 82118
rect 166956 80826 167075 82008
rect 168199 80826 168321 82008
rect 166956 80723 168321 80826
rect 21035 70833 22400 70943
rect 21035 69651 21154 70833
rect 22278 69651 22400 70833
rect 21035 69548 22400 69651
rect 27993 70834 29358 70944
rect 27993 69652 28112 70834
rect 29236 69652 29358 70834
rect 27993 69549 29358 69652
rect 34913 70833 36278 70943
rect 34913 69651 35032 70833
rect 36156 69651 36278 70833
rect 34913 69548 36278 69651
rect 41878 70834 43243 70944
rect 41878 69652 41997 70834
rect 43121 69652 43243 70834
rect 41878 69549 43243 69652
rect 48836 70835 50201 70945
rect 48836 69653 48955 70835
rect 50079 69653 50201 70835
rect 48836 69550 50201 69653
rect 55753 70839 57118 70949
rect 55753 69657 55872 70839
rect 56996 69657 57118 70839
rect 55753 69554 57118 69657
rect 62718 70840 64083 70950
rect 62718 69658 62837 70840
rect 63961 69658 64083 70840
rect 62718 69555 64083 69658
rect 69676 70841 71041 70951
rect 69676 69659 69795 70841
rect 70919 69659 71041 70841
rect 69676 69556 71041 69659
rect 76593 70839 77958 70949
rect 76593 69657 76712 70839
rect 77836 69657 77958 70839
rect 76593 69554 77958 69657
rect 83558 70840 84923 70950
rect 83558 69658 83677 70840
rect 84801 69658 84923 70840
rect 83558 69555 84923 69658
rect 90516 70841 91881 70951
rect 90516 69659 90635 70841
rect 91759 69659 91881 70841
rect 90516 69556 91881 69659
rect 97334 70820 98699 70930
rect 97334 69638 97453 70820
rect 98577 69638 98699 70820
rect 97334 69535 98699 69638
rect 104299 70821 105664 70931
rect 104299 69639 104418 70821
rect 105542 69639 105664 70821
rect 104299 69536 105664 69639
rect 111257 70822 112622 70932
rect 111257 69640 111376 70822
rect 112500 69640 112622 70822
rect 111257 69537 112622 69640
rect 118177 70821 119542 70931
rect 118177 69639 118296 70821
rect 119420 69639 119542 70821
rect 118177 69536 119542 69639
rect 125142 70822 126507 70932
rect 125142 69640 125261 70822
rect 126385 69640 126507 70822
rect 125142 69537 126507 69640
rect 132100 70823 133465 70933
rect 132100 69641 132219 70823
rect 133343 69641 133465 70823
rect 132100 69538 133465 69641
rect 139017 70827 140382 70937
rect 139017 69645 139136 70827
rect 140260 69645 140382 70827
rect 139017 69542 140382 69645
rect 145982 70828 147347 70938
rect 145982 69646 146101 70828
rect 147225 69646 147347 70828
rect 145982 69543 147347 69646
rect 152940 70829 154305 70939
rect 152940 69647 153059 70829
rect 154183 69647 154305 70829
rect 152940 69544 154305 69647
rect 159857 70827 161222 70937
rect 159857 69645 159976 70827
rect 161100 69645 161222 70827
rect 159857 69542 161222 69645
rect 166822 70828 168187 70938
rect 166822 69646 166941 70828
rect 168065 69646 168187 70828
rect 166822 69543 168187 69646
rect 173780 70829 175145 70939
rect 173780 69647 173899 70829
rect 175023 69647 175145 70829
rect 173780 69544 175145 69647
rect 21000 64593 22365 64703
rect 21000 63411 21119 64593
rect 22243 63411 22365 64593
rect 21000 63308 22365 63411
rect 27958 64594 29323 64704
rect 27958 63412 28077 64594
rect 29201 63412 29323 64594
rect 27958 63309 29323 63412
rect 34878 64593 36243 64703
rect 34878 63411 34997 64593
rect 36121 63411 36243 64593
rect 34878 63308 36243 63411
rect 41843 64594 43208 64704
rect 41843 63412 41962 64594
rect 43086 63412 43208 64594
rect 41843 63309 43208 63412
rect 48801 64595 50166 64705
rect 48801 63413 48920 64595
rect 50044 63413 50166 64595
rect 48801 63310 50166 63413
rect 55718 64599 57083 64709
rect 55718 63417 55837 64599
rect 56961 63417 57083 64599
rect 55718 63314 57083 63417
rect 62683 64600 64048 64710
rect 62683 63418 62802 64600
rect 63926 63418 64048 64600
rect 62683 63315 64048 63418
rect 69641 64601 71006 64711
rect 69641 63419 69760 64601
rect 70884 63419 71006 64601
rect 69641 63316 71006 63419
rect 76558 64599 77923 64709
rect 76558 63417 76677 64599
rect 77801 63417 77923 64599
rect 76558 63314 77923 63417
rect 83523 64600 84888 64710
rect 83523 63418 83642 64600
rect 84766 63418 84888 64600
rect 83523 63315 84888 63418
rect 90481 64601 91846 64711
rect 90481 63419 90600 64601
rect 91724 63419 91846 64601
rect 90481 63316 91846 63419
rect 97299 64580 98664 64690
rect 97299 63398 97418 64580
rect 98542 63398 98664 64580
rect 97299 63295 98664 63398
rect 104264 64581 105629 64691
rect 104264 63399 104383 64581
rect 105507 63399 105629 64581
rect 104264 63296 105629 63399
rect 111222 64582 112587 64692
rect 111222 63400 111341 64582
rect 112465 63400 112587 64582
rect 111222 63297 112587 63400
rect 118142 64581 119507 64691
rect 118142 63399 118261 64581
rect 119385 63399 119507 64581
rect 118142 63296 119507 63399
rect 125107 64582 126472 64692
rect 125107 63400 125226 64582
rect 126350 63400 126472 64582
rect 125107 63297 126472 63400
rect 132065 64583 133430 64693
rect 132065 63401 132184 64583
rect 133308 63401 133430 64583
rect 132065 63298 133430 63401
rect 138982 64587 140347 64697
rect 138982 63405 139101 64587
rect 140225 63405 140347 64587
rect 138982 63302 140347 63405
rect 145947 64588 147312 64698
rect 145947 63406 146066 64588
rect 147190 63406 147312 64588
rect 145947 63303 147312 63406
rect 152905 64589 154270 64699
rect 152905 63407 153024 64589
rect 154148 63407 154270 64589
rect 152905 63304 154270 63407
rect 159822 64587 161187 64697
rect 159822 63405 159941 64587
rect 161065 63405 161187 64587
rect 159822 63302 161187 63405
rect 166787 64588 168152 64698
rect 166787 63406 166906 64588
rect 168030 63406 168152 64588
rect 166787 63303 168152 63406
rect 173745 64589 175110 64699
rect 173745 63407 173864 64589
rect 174988 63407 175110 64589
rect 173745 63304 175110 63407
rect 20965 58876 22330 58986
rect 20965 57694 21084 58876
rect 22208 57694 22330 58876
rect 20965 57591 22330 57694
rect 27923 58877 29288 58987
rect 27923 57695 28042 58877
rect 29166 57695 29288 58877
rect 27923 57592 29288 57695
rect 34843 58876 36208 58986
rect 34843 57694 34962 58876
rect 36086 57694 36208 58876
rect 34843 57591 36208 57694
rect 41808 58877 43173 58987
rect 41808 57695 41927 58877
rect 43051 57695 43173 58877
rect 41808 57592 43173 57695
rect 48766 58878 50131 58988
rect 48766 57696 48885 58878
rect 50009 57696 50131 58878
rect 48766 57593 50131 57696
rect 55683 58882 57048 58992
rect 55683 57700 55802 58882
rect 56926 57700 57048 58882
rect 55683 57597 57048 57700
rect 62648 58883 64013 58993
rect 62648 57701 62767 58883
rect 63891 57701 64013 58883
rect 62648 57598 64013 57701
rect 69606 58884 70971 58994
rect 69606 57702 69725 58884
rect 70849 57702 70971 58884
rect 69606 57599 70971 57702
rect 76523 58882 77888 58992
rect 76523 57700 76642 58882
rect 77766 57700 77888 58882
rect 76523 57597 77888 57700
rect 83488 58883 84853 58993
rect 83488 57701 83607 58883
rect 84731 57701 84853 58883
rect 83488 57598 84853 57701
rect 90446 58884 91811 58994
rect 90446 57702 90565 58884
rect 91689 57702 91811 58884
rect 90446 57599 91811 57702
rect 97264 58863 98629 58973
rect 97264 57681 97383 58863
rect 98507 57681 98629 58863
rect 97264 57578 98629 57681
rect 104229 58864 105594 58974
rect 104229 57682 104348 58864
rect 105472 57682 105594 58864
rect 104229 57579 105594 57682
rect 111187 58865 112552 58975
rect 111187 57683 111306 58865
rect 112430 57683 112552 58865
rect 111187 57580 112552 57683
rect 118107 58864 119472 58974
rect 118107 57682 118226 58864
rect 119350 57682 119472 58864
rect 118107 57579 119472 57682
rect 125072 58865 126437 58975
rect 125072 57683 125191 58865
rect 126315 57683 126437 58865
rect 125072 57580 126437 57683
rect 132030 58866 133395 58976
rect 132030 57684 132149 58866
rect 133273 57684 133395 58866
rect 132030 57581 133395 57684
rect 138947 58870 140312 58980
rect 138947 57688 139066 58870
rect 140190 57688 140312 58870
rect 138947 57585 140312 57688
rect 145912 58871 147277 58981
rect 145912 57689 146031 58871
rect 147155 57689 147277 58871
rect 145912 57586 147277 57689
rect 152870 58872 154235 58982
rect 152870 57690 152989 58872
rect 154113 57690 154235 58872
rect 152870 57587 154235 57690
rect 159787 58870 161152 58980
rect 159787 57688 159906 58870
rect 161030 57688 161152 58870
rect 159787 57585 161152 57688
rect 166752 58871 168117 58981
rect 166752 57689 166871 58871
rect 167995 57689 168117 58871
rect 166752 57586 168117 57689
rect 173710 58872 175075 58982
rect 173710 57690 173829 58872
rect 174953 57690 175075 58872
rect 173710 57587 175075 57690
rect 20896 52671 22261 52781
rect 20896 51489 21015 52671
rect 22139 51489 22261 52671
rect 20896 51386 22261 51489
rect 27854 52672 29219 52782
rect 27854 51490 27973 52672
rect 29097 51490 29219 52672
rect 27854 51387 29219 51490
rect 34774 52671 36139 52781
rect 34774 51489 34893 52671
rect 36017 51489 36139 52671
rect 34774 51386 36139 51489
rect 41739 52672 43104 52782
rect 41739 51490 41858 52672
rect 42982 51490 43104 52672
rect 41739 51387 43104 51490
rect 48697 52673 50062 52783
rect 48697 51491 48816 52673
rect 49940 51491 50062 52673
rect 48697 51388 50062 51491
rect 55614 52677 56979 52787
rect 55614 51495 55733 52677
rect 56857 51495 56979 52677
rect 55614 51392 56979 51495
rect 62579 52678 63944 52788
rect 62579 51496 62698 52678
rect 63822 51496 63944 52678
rect 62579 51393 63944 51496
rect 69537 52679 70902 52789
rect 69537 51497 69656 52679
rect 70780 51497 70902 52679
rect 69537 51394 70902 51497
rect 76454 52677 77819 52787
rect 76454 51495 76573 52677
rect 77697 51495 77819 52677
rect 76454 51392 77819 51495
rect 83419 52678 84784 52788
rect 83419 51496 83538 52678
rect 84662 51496 84784 52678
rect 83419 51393 84784 51496
rect 90377 52679 91742 52789
rect 90377 51497 90496 52679
rect 91620 51497 91742 52679
rect 90377 51394 91742 51497
rect 97195 52658 98560 52768
rect 97195 51476 97314 52658
rect 98438 51476 98560 52658
rect 97195 51373 98560 51476
rect 104160 52659 105525 52769
rect 104160 51477 104279 52659
rect 105403 51477 105525 52659
rect 104160 51374 105525 51477
rect 111118 52660 112483 52770
rect 111118 51478 111237 52660
rect 112361 51478 112483 52660
rect 111118 51375 112483 51478
rect 118038 52659 119403 52769
rect 118038 51477 118157 52659
rect 119281 51477 119403 52659
rect 118038 51374 119403 51477
rect 125003 52660 126368 52770
rect 125003 51478 125122 52660
rect 126246 51478 126368 52660
rect 125003 51375 126368 51478
rect 131961 52661 133326 52771
rect 131961 51479 132080 52661
rect 133204 51479 133326 52661
rect 131961 51376 133326 51479
rect 138878 52665 140243 52775
rect 138878 51483 138997 52665
rect 140121 51483 140243 52665
rect 138878 51380 140243 51483
rect 145843 52666 147208 52776
rect 145843 51484 145962 52666
rect 147086 51484 147208 52666
rect 145843 51381 147208 51484
rect 152801 52667 154166 52777
rect 152801 51485 152920 52667
rect 154044 51485 154166 52667
rect 152801 51382 154166 51485
rect 159718 52665 161083 52775
rect 159718 51483 159837 52665
rect 160961 51483 161083 52665
rect 159718 51380 161083 51483
rect 166683 52666 168048 52776
rect 166683 51484 166802 52666
rect 167926 51484 168048 52666
rect 166683 51381 168048 51484
rect 173641 52667 175006 52777
rect 173641 51485 173760 52667
rect 174884 51485 175006 52667
rect 173641 51382 175006 51485
rect 138590 44807 139955 44917
rect 138590 43625 138709 44807
rect 139833 43625 139955 44807
rect 138590 43522 139955 43625
rect 145555 44808 146920 44918
rect 145555 43626 145674 44808
rect 146798 43626 146920 44808
rect 145555 43523 146920 43626
rect 152513 44809 153878 44919
rect 152513 43627 152632 44809
rect 153756 43627 153878 44809
rect 152513 43524 153878 43627
rect 159430 44807 160795 44917
rect 159430 43625 159549 44807
rect 160673 43625 160795 44807
rect 159430 43522 160795 43625
rect 166395 44808 167760 44918
rect 166395 43626 166514 44808
rect 167638 43626 167760 44808
rect 166395 43523 167760 43626
rect 173353 44809 174718 44919
rect 173353 43627 173472 44809
rect 174596 43627 174718 44809
rect 173353 43524 174718 43627
rect 138590 38513 139955 38623
rect 138590 37331 138709 38513
rect 139833 37331 139955 38513
rect 138590 37228 139955 37331
rect 145555 38514 146920 38624
rect 145555 37332 145674 38514
rect 146798 37332 146920 38514
rect 145555 37229 146920 37332
rect 152513 38515 153878 38625
rect 152513 37333 152632 38515
rect 153756 37333 153878 38515
rect 152513 37230 153878 37333
rect 159430 38513 160795 38623
rect 159430 37331 159549 38513
rect 160673 37331 160795 38513
rect 159430 37228 160795 37331
rect 166395 38514 167760 38624
rect 166395 37332 166514 38514
rect 167638 37332 167760 38514
rect 166395 37229 167760 37332
rect 173353 38515 174718 38625
rect 173353 37333 173472 38515
rect 174596 37333 174718 38515
rect 173353 37230 174718 37333
rect 138590 32219 139955 32329
rect 138590 31037 138709 32219
rect 139833 31037 139955 32219
rect 138590 30934 139955 31037
rect 145555 32220 146920 32330
rect 145555 31038 145674 32220
rect 146798 31038 146920 32220
rect 145555 30935 146920 31038
rect 152513 32221 153878 32331
rect 152513 31039 152632 32221
rect 153756 31039 153878 32221
rect 152513 30936 153878 31039
rect 159430 32219 160795 32329
rect 159430 31037 159549 32219
rect 160673 31037 160795 32219
rect 159430 30934 160795 31037
rect 166395 32220 167760 32330
rect 166395 31038 166514 32220
rect 167638 31038 167760 32220
rect 166395 30935 167760 31038
rect 173353 32221 174718 32331
rect 173353 31039 173472 32221
rect 174596 31039 174718 32221
rect 173353 30936 174718 31039
<< psubdiffcont >>
rect 83511 338865 84635 340047
rect 90469 338866 91593 340048
rect 97287 338845 98411 340027
rect 104252 338846 105376 340028
rect 111210 338847 112334 340029
rect 118130 338846 119254 340028
rect 125095 338847 126219 340029
rect 132053 338848 133177 340030
rect 138970 338852 140094 340034
rect 145935 338853 147059 340035
rect 152893 338854 154017 340036
rect 159810 338852 160934 340034
rect 166775 338853 167899 340035
rect 173733 338854 174857 340036
rect 180538 338847 181662 340029
rect 187503 338848 188627 340030
rect 194461 338849 195585 340031
rect 201381 338848 202505 340030
rect 208346 338849 209470 340031
rect 215304 338850 216428 340032
rect 97013 331715 98137 332897
rect 103978 331716 105102 332898
rect 138696 331722 139820 332904
rect 145661 331723 146785 332905
rect 152619 331724 153743 332906
rect 159536 331722 160660 332904
rect 166501 331723 167625 332905
rect 173459 331724 174583 332906
rect 180264 331717 181388 332899
rect 187229 331718 188353 332900
rect 194187 331719 195311 332901
rect 201107 331718 202231 332900
rect 208072 331719 209196 332901
rect 215030 331720 216154 332902
rect 97287 325387 98411 326569
rect 104252 325388 105376 326570
rect 138970 325394 140094 326576
rect 145935 325395 147059 326577
rect 152893 325396 154017 326578
rect 159810 325394 160934 326576
rect 166775 325395 167899 326577
rect 173733 325396 174857 326578
rect 180538 325389 181662 326571
rect 187503 325390 188627 326572
rect 194461 325391 195585 326573
rect 201381 325390 202505 326572
rect 208346 325391 209470 326573
rect 215304 325392 216428 326574
rect 97013 318257 98137 319439
rect 103978 318258 105102 319440
rect 138696 318264 139820 319446
rect 145661 318265 146785 319447
rect 152619 318266 153743 319448
rect 159536 318264 160660 319446
rect 166501 318265 167625 319447
rect 173459 318266 174583 319448
rect 180264 318259 181388 319441
rect 187229 318260 188353 319442
rect 194187 318261 195311 319443
rect 201107 318260 202231 319442
rect 208072 318261 209196 319443
rect 215030 318262 216154 319444
rect 97293 311126 98417 312308
rect 104258 311127 105382 312309
rect 138976 311133 140100 312315
rect 145941 311134 147065 312316
rect 152899 311135 154023 312317
rect 159816 311133 160940 312315
rect 166781 311134 167905 312316
rect 173739 311135 174863 312317
rect 180544 311128 181668 312310
rect 187509 311129 188633 312311
rect 194467 311130 195591 312312
rect 201387 311129 202511 312311
rect 208352 311130 209476 312312
rect 215310 311131 216434 312313
rect 83243 304016 84367 305198
rect 90201 304017 91325 305199
rect 97019 303996 98143 305178
rect 103984 303997 105108 305179
rect 110942 303998 112066 305180
rect 117862 303997 118986 305179
rect 124827 303998 125951 305180
rect 131785 303999 132909 305181
rect 138702 304003 139826 305185
rect 145667 304004 146791 305186
rect 152625 304005 153749 305187
rect 159542 304003 160666 305185
rect 166507 304004 167631 305186
rect 173465 304005 174589 305187
rect 180270 303998 181394 305180
rect 187235 303999 188359 305181
rect 194193 304000 195317 305182
rect 201113 303999 202237 305181
rect 208078 304000 209202 305182
rect 215036 304001 216160 305183
rect 97382 294767 98506 295949
rect 104347 294768 105471 295950
rect 139065 294774 140189 295956
rect 146030 294775 147154 295957
rect 152988 294776 154112 295958
rect 159905 294774 161029 295956
rect 166870 294775 167994 295957
rect 187598 294770 188722 295952
rect 194556 294771 195680 295953
rect 97108 287637 98232 288819
rect 104073 287638 105197 288820
rect 138791 287644 139915 288826
rect 145756 287645 146880 288827
rect 152714 287646 153838 288828
rect 159631 287644 160755 288826
rect 166596 287645 167720 288827
rect 187324 287640 188448 288822
rect 194282 287641 195406 288823
rect 97216 281224 98340 282406
rect 104181 281225 105305 282407
rect 138899 281231 140023 282413
rect 145864 281232 146988 282414
rect 152822 281233 153946 282415
rect 159739 281231 160863 282413
rect 166704 281232 167828 282414
rect 187432 281227 188556 282409
rect 194390 281228 195514 282410
rect 69775 272380 70899 273562
rect 76692 272378 77816 273560
rect 83657 272379 84781 273561
rect 90615 272380 91739 273562
rect 97433 272359 98557 273541
rect 104398 272360 105522 273542
rect 111356 272361 112480 273543
rect 118276 272360 119400 273542
rect 125241 272361 126365 273543
rect 132199 272362 133323 273544
rect 139116 272366 140240 273548
rect 146081 272367 147205 273549
rect 153039 272368 154163 273550
rect 159956 272366 161080 273548
rect 166921 272367 168045 273549
rect 173879 272368 175003 273550
rect 180684 272361 181808 273543
rect 187649 272362 188773 273544
rect 194607 272363 195731 273545
rect 201527 272362 202651 273544
rect 208492 272363 209616 273545
rect 215450 272364 216574 273546
rect 222367 272368 223491 273550
rect 69501 265250 70625 266432
rect 76418 265248 77542 266430
rect 83383 265249 84507 266431
rect 90341 265250 91465 266432
rect 97159 265229 98283 266411
rect 104124 265230 105248 266412
rect 111082 265231 112206 266413
rect 118002 265230 119126 266412
rect 124967 265231 126091 266413
rect 131925 265232 133049 266414
rect 138842 265236 139966 266418
rect 145807 265237 146931 266419
rect 152765 265238 153889 266420
rect 159682 265236 160806 266418
rect 166647 265237 167771 266419
rect 173605 265238 174729 266420
rect 180410 265231 181534 266413
rect 187375 265232 188499 266414
rect 194333 265233 195457 266415
rect 201253 265232 202377 266414
rect 208218 265233 209342 266415
rect 215176 265234 216300 266416
rect 222093 265238 223217 266420
rect 69609 258837 70733 260019
rect 76526 258835 77650 260017
rect 83491 258836 84615 260018
rect 90449 258837 91573 260019
rect 97267 258816 98391 259998
rect 104232 258817 105356 259999
rect 111190 258818 112314 260000
rect 118110 258817 119234 259999
rect 125075 258818 126199 260000
rect 132033 258819 133157 260001
rect 138950 258823 140074 260005
rect 145915 258824 147039 260006
rect 152873 258825 153997 260007
rect 159790 258823 160914 260005
rect 166755 258824 167879 260006
rect 173713 258825 174837 260007
rect 180518 258818 181642 260000
rect 187483 258819 188607 260001
rect 194441 258820 195565 260002
rect 201361 258819 202485 260001
rect 208326 258820 209450 260002
rect 215284 258821 216408 260003
rect 222201 258825 223325 260007
rect 83688 248125 84812 249307
rect 90646 248126 91770 249308
rect 97464 248105 98588 249287
rect 104429 248106 105553 249288
rect 111387 248107 112511 249289
rect 118307 248106 119431 249288
rect 125272 248107 126396 249289
rect 132230 248108 133354 249290
rect 139147 248112 140271 249294
rect 146112 248113 147236 249295
rect 153070 248114 154194 249296
rect 159987 248112 161111 249294
rect 166952 248113 168076 249295
rect 173910 248114 175034 249296
rect 180715 248107 181839 249289
rect 187680 248108 188804 249290
rect 194638 248109 195762 249291
rect 201558 248108 202682 249290
rect 208523 248109 209647 249291
rect 215481 248110 216605 249292
rect 222398 248114 223522 249296
rect 83414 240995 84538 242177
rect 90372 240996 91496 242178
rect 97190 240975 98314 242157
rect 104155 240976 105279 242158
rect 111113 240977 112237 242159
rect 118033 240976 119157 242158
rect 124998 240977 126122 242159
rect 131956 240978 133080 242160
rect 138873 240982 139997 242164
rect 145838 240983 146962 242165
rect 152796 240984 153920 242166
rect 159713 240982 160837 242164
rect 166678 240983 167802 242165
rect 173636 240984 174760 242166
rect 180441 240977 181565 242159
rect 187406 240978 188530 242160
rect 194364 240979 195488 242161
rect 201284 240978 202408 242160
rect 208249 240979 209373 242161
rect 215207 240980 216331 242162
rect 222124 240984 223248 242166
rect 83522 234582 84646 235764
rect 90480 234583 91604 235765
rect 97298 234562 98422 235744
rect 104263 234563 105387 235745
rect 111221 234564 112345 235746
rect 118141 234563 119265 235745
rect 125106 234564 126230 235746
rect 132064 234565 133188 235747
rect 138981 234569 140105 235751
rect 145946 234570 147070 235752
rect 152904 234571 154028 235753
rect 159821 234569 160945 235751
rect 166786 234570 167910 235752
rect 173744 234571 174868 235753
rect 180549 234564 181673 235746
rect 187514 234565 188638 235747
rect 194472 234566 195596 235748
rect 201392 234565 202516 235747
rect 208357 234566 209481 235748
rect 215315 234567 216439 235749
rect 222232 234571 223356 235753
rect 69930 227860 71054 229042
rect 76847 227858 77971 229040
rect 83812 227859 84936 229041
rect 90770 227860 91894 229042
rect 97588 227839 98712 229021
rect 104553 227840 105677 229022
rect 111511 227841 112635 229023
rect 118431 227840 119555 229022
rect 125396 227841 126520 229023
rect 132354 227842 133478 229024
rect 139271 227846 140395 229028
rect 146236 227847 147360 229029
rect 153194 227848 154318 229030
rect 160111 227846 161235 229028
rect 167076 227847 168200 229029
rect 174034 227848 175158 229030
rect 180839 227841 181963 229023
rect 187804 227842 188928 229024
rect 194762 227843 195886 229025
rect 201682 227842 202806 229024
rect 208647 227843 209771 229025
rect 215605 227844 216729 229026
rect 222522 227848 223646 229030
rect 69910 221998 71034 223180
rect 76827 221996 77951 223178
rect 83792 221997 84916 223179
rect 90750 221998 91874 223180
rect 97568 221977 98692 223159
rect 104533 221978 105657 223160
rect 111491 221979 112615 223161
rect 118411 221978 119535 223160
rect 125376 221979 126500 223161
rect 132334 221980 133458 223162
rect 139251 221984 140375 223166
rect 146216 221985 147340 223167
rect 153174 221986 154298 223168
rect 160091 221984 161215 223166
rect 167056 221985 168180 223167
rect 174014 221986 175138 223168
rect 180819 221979 181943 223161
rect 187784 221980 188908 223162
rect 194742 221981 195866 223163
rect 201662 221980 202786 223162
rect 208627 221981 209751 223163
rect 215585 221982 216709 223164
rect 222502 221986 223626 223168
rect 21309 209927 22433 211109
rect 28267 209928 29391 211110
rect 35187 209927 36311 211109
rect 42152 209928 43276 211110
rect 49110 209929 50234 211111
rect 56027 209933 57151 211115
rect 62992 209934 64116 211116
rect 97608 209914 98732 211096
rect 104573 209915 105697 211097
rect 139291 209921 140415 211103
rect 146256 209922 147380 211104
rect 153214 209923 154338 211105
rect 160131 209921 161255 211103
rect 167096 209922 168220 211104
rect 264445 209925 265569 211107
rect 271403 209926 272527 211108
rect 21035 202797 22159 203979
rect 27993 202798 29117 203980
rect 34913 202797 36037 203979
rect 41878 202798 43002 203980
rect 48836 202799 49960 203981
rect 55753 202803 56877 203985
rect 62718 202804 63842 203986
rect 97334 202784 98458 203966
rect 104299 202785 105423 203967
rect 139017 202791 140141 203973
rect 145982 202792 147106 203974
rect 152940 202793 154064 203975
rect 159857 202791 160981 203973
rect 166822 202792 167946 203974
rect 264171 202795 265295 203977
rect 271129 202796 272253 203978
rect 21143 196384 22267 197566
rect 28101 196385 29225 197567
rect 35021 196384 36145 197566
rect 41986 196385 43110 197567
rect 48944 196386 50068 197568
rect 55861 196390 56985 197572
rect 62826 196391 63950 197573
rect 97442 196371 98566 197553
rect 104407 196372 105531 197554
rect 139125 196378 140249 197560
rect 146090 196379 147214 197561
rect 153048 196380 154172 197562
rect 159965 196378 161089 197560
rect 166930 196379 168054 197561
rect 264279 196382 265403 197564
rect 271237 196383 272361 197565
rect 97595 192021 98719 193203
rect 104560 192022 105684 193204
rect 139278 192028 140402 193210
rect 146243 192029 147367 193211
rect 153201 192030 154325 193212
rect 160118 192028 161242 193210
rect 167083 192029 168207 193211
rect 264432 192032 265556 193214
rect 271390 192033 272514 193215
rect 76580 184910 77704 186092
rect 83545 184911 84669 186093
rect 90503 184912 91627 186094
rect 97321 184891 98445 186073
rect 104286 184892 105410 186074
rect 139004 184898 140128 186080
rect 145969 184899 147093 186081
rect 152927 184900 154051 186082
rect 159844 184898 160968 186080
rect 166809 184899 167933 186081
rect 173767 184900 174891 186082
rect 180572 184893 181696 186075
rect 187537 184894 188661 186076
rect 194495 184895 195619 186077
rect 201415 184894 202539 186076
rect 208380 184895 209504 186077
rect 215338 184896 216462 186078
rect 222255 184900 223379 186082
rect 229220 184901 230344 186083
rect 236178 184902 237302 186084
rect 243095 184900 244219 186082
rect 250060 184901 251184 186083
rect 257018 184902 258142 186084
rect 264158 184902 265282 186084
rect 271116 184903 272240 186085
rect 278252 184893 279376 186075
rect 76688 178497 77812 179679
rect 83653 178498 84777 179680
rect 90611 178499 91735 179681
rect 97429 178478 98553 179660
rect 104394 178479 105518 179661
rect 111352 178480 112476 179662
rect 118272 178479 119396 179661
rect 125237 178480 126361 179662
rect 132195 178481 133319 179663
rect 139112 178485 140236 179667
rect 146077 178486 147201 179668
rect 153035 178487 154159 179669
rect 159952 178485 161076 179667
rect 166917 178486 168041 179668
rect 173875 178487 174999 179669
rect 180680 178480 181804 179662
rect 187645 178481 188769 179663
rect 194603 178482 195727 179664
rect 201523 178481 202647 179663
rect 208488 178482 209612 179664
rect 215446 178483 216570 179665
rect 222363 178487 223487 179669
rect 229328 178488 230452 179670
rect 236286 178489 237410 179671
rect 243203 178487 244327 179669
rect 250168 178488 251292 179670
rect 257126 178489 258250 179671
rect 264266 178489 265390 179671
rect 271224 178490 272348 179672
rect 278360 178480 279484 179662
rect 69486 172585 70610 173767
rect 76403 172583 77527 173765
rect 83368 172584 84492 173766
rect 90326 172585 91450 173767
rect 97144 172564 98268 173746
rect 104109 172565 105233 173747
rect 111067 172566 112191 173748
rect 117987 172565 119111 173747
rect 124952 172566 126076 173748
rect 131910 172567 133034 173749
rect 138827 172571 139951 173753
rect 145792 172572 146916 173754
rect 152750 172573 153874 173755
rect 159667 172571 160791 173753
rect 166632 172572 167756 173754
rect 173590 172573 174714 173755
rect 180395 172566 181519 173748
rect 187360 172567 188484 173749
rect 194318 172568 195442 173750
rect 201238 172567 202362 173749
rect 208203 172568 209327 173750
rect 215161 172569 216285 173751
rect 222078 172573 223202 173755
rect 229043 172574 230167 173756
rect 236001 172575 237125 173757
rect 242918 172573 244042 173755
rect 249883 172574 251007 173756
rect 256841 172575 257965 173757
rect 263981 172575 265105 173757
rect 270939 172576 272063 173758
rect 278075 172566 279199 173748
rect 69594 166172 70718 167354
rect 76511 166170 77635 167352
rect 83476 166171 84600 167353
rect 90434 166172 91558 167354
rect 97252 166151 98376 167333
rect 104217 166152 105341 167334
rect 111175 166153 112299 167335
rect 118095 166152 119219 167334
rect 125060 166153 126184 167335
rect 132018 166154 133142 167336
rect 138935 166158 140059 167340
rect 145900 166159 147024 167341
rect 152858 166160 153982 167342
rect 159775 166158 160899 167340
rect 166740 166159 167864 167341
rect 173698 166160 174822 167342
rect 180503 166153 181627 167335
rect 187468 166154 188592 167336
rect 194426 166155 195550 167337
rect 201346 166154 202470 167336
rect 208311 166155 209435 167337
rect 215269 166156 216393 167338
rect 222186 166160 223310 167342
rect 229151 166161 230275 167343
rect 236109 166162 237233 167344
rect 243026 166160 244150 167342
rect 249991 166161 251115 167343
rect 256949 166162 258073 167344
rect 264089 166162 265213 167344
rect 271047 166163 272171 167345
rect 278183 166153 279307 167335
rect 21720 158825 22844 160007
rect 28678 158826 29802 160008
rect 35598 158825 36722 160007
rect 56438 158831 57562 160013
rect 63403 158832 64527 160014
rect 98019 158812 99143 159994
rect 104984 158813 106108 159995
rect 139702 158819 140826 160001
rect 146667 158820 147791 160002
rect 153625 158821 154749 160003
rect 160542 158819 161666 160001
rect 167507 158820 168631 160002
rect 188235 158815 189359 159997
rect 195193 158816 196317 159998
rect 229792 158816 230916 159998
rect 236757 158817 237881 159999
rect 243715 158818 244839 160000
rect 250632 158822 251756 160004
rect 257524 158805 258648 159987
rect 264489 158806 265613 159988
rect 271447 158807 272571 159989
rect 278364 158811 279488 159993
rect 22005 153992 23129 155174
rect 28963 153993 30087 155175
rect 35883 153992 37007 155174
rect 56723 153998 57847 155180
rect 63688 153999 64812 155181
rect 98304 153979 99428 155161
rect 105269 153980 106393 155162
rect 139987 153986 141111 155168
rect 146952 153987 148076 155169
rect 153910 153988 155034 155170
rect 160827 153986 161951 155168
rect 167792 153987 168916 155169
rect 188520 153982 189644 155164
rect 195478 153983 196602 155165
rect 230077 153983 231201 155165
rect 237042 153984 238166 155166
rect 244000 153985 245124 155167
rect 250917 153989 252041 155171
rect 257809 153972 258933 155154
rect 264774 153973 265898 155155
rect 271732 153974 272856 155156
rect 278649 153978 279773 155160
rect 22076 148732 23200 149914
rect 29034 148733 30158 149915
rect 35954 148732 37078 149914
rect 56794 148738 57918 149920
rect 63759 148739 64883 149921
rect 98375 148719 99499 149901
rect 105340 148720 106464 149902
rect 140058 148726 141182 149908
rect 147023 148727 148147 149909
rect 153981 148728 155105 149910
rect 160898 148726 162022 149908
rect 167863 148727 168987 149909
rect 188591 148722 189715 149904
rect 195549 148723 196673 149905
rect 230148 148723 231272 149905
rect 237113 148724 238237 149906
rect 244071 148725 245195 149907
rect 250988 148729 252112 149911
rect 257880 148712 259004 149894
rect 264845 148713 265969 149895
rect 271803 148714 272927 149896
rect 278720 148718 279844 149900
rect 22005 143258 23129 144440
rect 28963 143259 30087 144441
rect 35883 143258 37007 144440
rect 56723 143264 57847 144446
rect 63688 143265 64812 144447
rect 98304 143245 99428 144427
rect 105269 143246 106393 144428
rect 139987 143252 141111 144434
rect 146952 143253 148076 144435
rect 153910 143254 155034 144436
rect 160827 143252 161951 144434
rect 167792 143253 168916 144435
rect 188520 143248 189644 144430
rect 195478 143249 196602 144431
rect 22147 137146 23271 138328
rect 29105 137147 30229 138329
rect 36025 137146 37149 138328
rect 56865 137152 57989 138334
rect 63830 137153 64954 138335
rect 98446 137133 99570 138315
rect 105411 137134 106535 138316
rect 140129 137140 141253 138322
rect 147094 137141 148218 138323
rect 154052 137142 155176 138324
rect 160969 137140 162093 138322
rect 167934 137141 169058 138323
rect 188662 137136 189786 138318
rect 195620 137137 196744 138319
rect 21937 129272 23061 130454
rect 28895 129273 30019 130455
rect 35815 129272 36939 130454
rect 42780 129273 43904 130455
rect 49738 129274 50862 130456
rect 56655 129278 57779 130460
rect 63620 129279 64744 130461
rect 70578 129280 71702 130462
rect 77495 129278 78619 130460
rect 84460 129279 85584 130461
rect 91418 129280 92542 130462
rect 98236 129259 99360 130441
rect 105201 129260 106325 130442
rect 112159 129261 113283 130443
rect 119079 129260 120203 130442
rect 126044 129261 127168 130443
rect 133002 129262 134126 130444
rect 139919 129266 141043 130448
rect 146884 129267 148008 130449
rect 153842 129268 154966 130450
rect 160759 129266 161883 130448
rect 167724 129267 168848 130449
rect 174682 129268 175806 130450
rect 181487 129261 182611 130443
rect 188452 129262 189576 130444
rect 195410 129263 196534 130445
rect 97753 117943 98877 119125
rect 104718 117944 105842 119126
rect 139436 117950 140560 119132
rect 146401 117951 147525 119133
rect 153359 117952 154483 119134
rect 160276 117950 161400 119132
rect 167241 117951 168365 119133
rect 97958 109991 99082 111173
rect 104923 109992 106047 111174
rect 139641 109998 140765 111180
rect 146606 109999 147730 111181
rect 153564 110000 154688 111182
rect 160481 109998 161605 111180
rect 167446 109999 168570 111181
rect 97958 101765 99082 102947
rect 104923 101766 106047 102948
rect 139641 101772 140765 102954
rect 146606 101773 147730 102955
rect 153564 101774 154688 102956
rect 160481 101772 161605 102954
rect 167446 101773 168570 102955
rect 97753 94361 98877 95543
rect 104718 94362 105842 95544
rect 139436 94368 140560 95550
rect 146401 94369 147525 95551
rect 153359 94370 154483 95552
rect 160276 94368 161400 95550
rect 167241 94369 168365 95551
rect 97479 87231 98603 88413
rect 104444 87232 105568 88414
rect 111402 87233 112526 88415
rect 118322 87232 119446 88414
rect 125287 87233 126411 88415
rect 132245 87234 133369 88416
rect 139162 87238 140286 88420
rect 146127 87239 147251 88421
rect 153085 87240 154209 88422
rect 160002 87238 161126 88420
rect 166967 87239 168091 88421
rect 97587 80818 98711 82000
rect 104552 80819 105676 82001
rect 111510 80820 112634 82002
rect 118430 80819 119554 82001
rect 125395 80820 126519 82002
rect 132353 80821 133477 82003
rect 139270 80825 140394 82007
rect 146235 80826 147359 82008
rect 153193 80827 154317 82009
rect 160110 80825 161234 82007
rect 167075 80826 168199 82008
rect 21154 69651 22278 70833
rect 28112 69652 29236 70834
rect 35032 69651 36156 70833
rect 41997 69652 43121 70834
rect 48955 69653 50079 70835
rect 55872 69657 56996 70839
rect 62837 69658 63961 70840
rect 69795 69659 70919 70841
rect 76712 69657 77836 70839
rect 83677 69658 84801 70840
rect 90635 69659 91759 70841
rect 97453 69638 98577 70820
rect 104418 69639 105542 70821
rect 111376 69640 112500 70822
rect 118296 69639 119420 70821
rect 125261 69640 126385 70822
rect 132219 69641 133343 70823
rect 139136 69645 140260 70827
rect 146101 69646 147225 70828
rect 153059 69647 154183 70829
rect 159976 69645 161100 70827
rect 166941 69646 168065 70828
rect 173899 69647 175023 70829
rect 21119 63411 22243 64593
rect 28077 63412 29201 64594
rect 34997 63411 36121 64593
rect 41962 63412 43086 64594
rect 48920 63413 50044 64595
rect 55837 63417 56961 64599
rect 62802 63418 63926 64600
rect 69760 63419 70884 64601
rect 76677 63417 77801 64599
rect 83642 63418 84766 64600
rect 90600 63419 91724 64601
rect 97418 63398 98542 64580
rect 104383 63399 105507 64581
rect 111341 63400 112465 64582
rect 118261 63399 119385 64581
rect 125226 63400 126350 64582
rect 132184 63401 133308 64583
rect 139101 63405 140225 64587
rect 146066 63406 147190 64588
rect 153024 63407 154148 64589
rect 159941 63405 161065 64587
rect 166906 63406 168030 64588
rect 173864 63407 174988 64589
rect 21084 57694 22208 58876
rect 28042 57695 29166 58877
rect 34962 57694 36086 58876
rect 41927 57695 43051 58877
rect 48885 57696 50009 58878
rect 55802 57700 56926 58882
rect 62767 57701 63891 58883
rect 69725 57702 70849 58884
rect 76642 57700 77766 58882
rect 83607 57701 84731 58883
rect 90565 57702 91689 58884
rect 97383 57681 98507 58863
rect 104348 57682 105472 58864
rect 111306 57683 112430 58865
rect 118226 57682 119350 58864
rect 125191 57683 126315 58865
rect 132149 57684 133273 58866
rect 139066 57688 140190 58870
rect 146031 57689 147155 58871
rect 152989 57690 154113 58872
rect 159906 57688 161030 58870
rect 166871 57689 167995 58871
rect 173829 57690 174953 58872
rect 21015 51489 22139 52671
rect 27973 51490 29097 52672
rect 34893 51489 36017 52671
rect 41858 51490 42982 52672
rect 48816 51491 49940 52673
rect 55733 51495 56857 52677
rect 62698 51496 63822 52678
rect 69656 51497 70780 52679
rect 76573 51495 77697 52677
rect 83538 51496 84662 52678
rect 90496 51497 91620 52679
rect 97314 51476 98438 52658
rect 104279 51477 105403 52659
rect 111237 51478 112361 52660
rect 118157 51477 119281 52659
rect 125122 51478 126246 52660
rect 132080 51479 133204 52661
rect 138997 51483 140121 52665
rect 145962 51484 147086 52666
rect 152920 51485 154044 52667
rect 159837 51483 160961 52665
rect 166802 51484 167926 52666
rect 173760 51485 174884 52667
rect 138709 43625 139833 44807
rect 145674 43626 146798 44808
rect 152632 43627 153756 44809
rect 159549 43625 160673 44807
rect 166514 43626 167638 44808
rect 173472 43627 174596 44809
rect 138709 37331 139833 38513
rect 145674 37332 146798 38514
rect 152632 37333 153756 38515
rect 159549 37331 160673 38513
rect 166514 37332 167638 38514
rect 173472 37333 174596 38515
rect 138709 31037 139833 32219
rect 145674 31038 146798 32220
rect 152632 31039 153756 32221
rect 159549 31037 160673 32219
rect 166514 31038 167638 32220
rect 173472 31039 174596 32221
<< locali >>
rect 79696 340492 100486 340530
rect 102753 340517 141064 340530
rect 143513 340517 189653 340530
rect 102753 340495 189653 340517
rect 192003 340495 220030 340530
rect 102753 340492 220030 340495
rect 79696 340048 220030 340492
rect 79696 340047 90469 340048
rect 79696 338865 83511 340047
rect 84635 338866 90469 340047
rect 91593 340036 220030 340048
rect 91593 340035 152893 340036
rect 91593 340034 145935 340035
rect 91593 340030 138970 340034
rect 91593 340029 132053 340030
rect 91593 340028 111210 340029
rect 91593 340027 104252 340028
rect 91593 338866 97287 340027
rect 84635 338865 97287 338866
rect 79696 338845 97287 338865
rect 98411 338846 104252 340027
rect 105376 338847 111210 340028
rect 112334 340028 125095 340029
rect 112334 338847 118130 340028
rect 105376 338846 118130 338847
rect 119254 338847 125095 340028
rect 126219 338848 132053 340029
rect 133177 338852 138970 340030
rect 140094 338853 145935 340034
rect 147059 338854 152893 340035
rect 154017 340035 173733 340036
rect 154017 340034 166775 340035
rect 154017 338854 159810 340034
rect 147059 338853 159810 338854
rect 140094 338852 159810 338853
rect 160934 339949 166775 340034
rect 160934 338852 164500 339949
rect 133177 338848 164500 338852
rect 126219 338847 164500 338848
rect 119254 338846 164500 338847
rect 98411 338845 164500 338846
rect 79696 338774 164500 338845
rect 165766 338853 166775 339949
rect 167899 338854 173733 340035
rect 174857 340032 220030 340036
rect 174857 340031 215304 340032
rect 174857 340030 194461 340031
rect 174857 340029 187503 340030
rect 174857 338854 180538 340029
rect 167899 338853 180538 338854
rect 165766 338847 180538 338853
rect 181662 338848 187503 340029
rect 188627 338849 194461 340030
rect 195585 340030 208346 340031
rect 195585 338849 201381 340030
rect 188627 338848 201381 338849
rect 202505 338849 208346 340030
rect 209470 338850 215304 340031
rect 216428 338850 220030 340032
rect 209470 338849 220030 338850
rect 202505 338848 220030 338849
rect 181662 338847 220030 338848
rect 165766 338774 220030 338847
rect 79696 338423 220030 338774
rect 100639 333400 102538 338423
rect 141388 333400 143287 338423
rect 189962 333400 191861 338423
rect 94867 332898 107106 333400
rect 94867 332897 103978 332898
rect 94867 331715 97013 332897
rect 98137 331716 103978 332897
rect 105102 331716 107106 332898
rect 98137 331715 107106 331716
rect 94867 331293 107106 331715
rect 136177 332906 220030 333400
rect 136177 332905 152619 332906
rect 136177 332904 145661 332905
rect 136177 331722 138696 332904
rect 139820 331723 145661 332904
rect 146785 331724 152619 332905
rect 153743 332905 173459 332906
rect 153743 332904 166501 332905
rect 153743 331724 159536 332904
rect 146785 331723 159536 331724
rect 139820 331722 159536 331723
rect 160660 332863 166501 332904
rect 160660 331722 164481 332863
rect 136177 331688 164481 331722
rect 165747 331723 166501 332863
rect 167625 331724 173459 332905
rect 174583 332902 220030 332906
rect 174583 332901 215030 332902
rect 174583 332900 194187 332901
rect 174583 332899 187229 332900
rect 174583 331724 180264 332899
rect 167625 331723 180264 331724
rect 165747 331717 180264 331723
rect 181388 331718 187229 332899
rect 188353 331719 194187 332900
rect 195311 332900 208072 332901
rect 195311 331719 201107 332900
rect 188353 331718 201107 331719
rect 202231 331719 208072 332900
rect 209196 331720 215030 332901
rect 216154 331720 220030 332902
rect 209196 331719 220030 331720
rect 202231 331718 220030 331719
rect 181388 331717 220030 331718
rect 165747 331688 220030 331717
rect 136177 331293 220030 331688
rect 100593 330649 102644 331293
rect 141388 330649 143422 331293
rect 100593 327072 102621 330649
rect 141394 327719 143422 330649
rect 141388 327072 143422 327719
rect 189886 330649 191921 331293
rect 189886 327072 191914 330649
rect 94867 326570 107106 327072
rect 94867 326569 104252 326570
rect 94867 325387 97287 326569
rect 98411 325388 104252 326569
rect 105376 325388 107106 326570
rect 98411 325387 107106 325388
rect 94867 324965 107106 325387
rect 136177 326578 220030 327072
rect 136177 326577 152893 326578
rect 136177 326576 145935 326577
rect 136177 325394 138970 326576
rect 140094 325395 145935 326576
rect 147059 325396 152893 326577
rect 154017 326577 173733 326578
rect 154017 326576 166775 326577
rect 154017 325396 159810 326576
rect 147059 325395 159810 325396
rect 140094 325394 159810 325395
rect 160934 326491 166775 326576
rect 160934 325394 164500 326491
rect 136177 325316 164500 325394
rect 165766 325395 166775 326491
rect 167899 325396 173733 326577
rect 174857 326574 220030 326578
rect 174857 326573 215304 326574
rect 174857 326572 194461 326573
rect 174857 326571 187503 326572
rect 174857 325396 180538 326571
rect 167899 325395 180538 325396
rect 165766 325389 180538 325395
rect 181662 325390 187503 326571
rect 188627 325391 194461 326572
rect 195585 326572 208346 326573
rect 195585 325391 201381 326572
rect 188627 325390 201381 325391
rect 202505 325391 208346 326572
rect 209470 325392 215304 326573
rect 216428 325392 220030 326574
rect 209470 325391 220030 325392
rect 202505 325390 220030 325391
rect 181662 325389 220030 325390
rect 165766 325316 220030 325389
rect 136177 324965 220030 325316
rect 100593 319942 102621 324965
rect 141388 319942 143422 324965
rect 189886 319942 191914 324965
rect 94867 319440 107106 319942
rect 94867 319439 103978 319440
rect 94867 318257 97013 319439
rect 98137 318258 103978 319439
rect 105102 318258 107106 319440
rect 98137 318257 107106 318258
rect 94867 317835 107106 318257
rect 136177 319448 220030 319942
rect 136177 319447 152619 319448
rect 136177 319446 145661 319447
rect 136177 318264 138696 319446
rect 139820 318265 145661 319446
rect 146785 318266 152619 319447
rect 153743 319447 173459 319448
rect 153743 319446 166501 319447
rect 153743 318266 159536 319446
rect 146785 318265 159536 318266
rect 139820 318264 159536 318265
rect 160660 319405 166501 319446
rect 160660 318264 164481 319405
rect 136177 318230 164481 318264
rect 165747 318265 166501 319405
rect 167625 318266 173459 319447
rect 174583 319444 220030 319448
rect 174583 319443 215030 319444
rect 174583 319442 194187 319443
rect 174583 319441 187229 319442
rect 174583 318266 180264 319441
rect 167625 318265 180264 318266
rect 165747 318259 180264 318265
rect 181388 318260 187229 319441
rect 188353 318261 194187 319442
rect 195311 319442 208072 319443
rect 195311 318261 201107 319442
rect 188353 318260 201107 318261
rect 202231 318261 208072 319442
rect 209196 318262 215030 319443
rect 216154 318262 220030 319444
rect 209196 318261 220030 318262
rect 202231 318260 220030 318261
rect 181388 318259 220030 318260
rect 165747 318230 220030 318259
rect 136177 317835 220030 318230
rect 100593 317191 102644 317835
rect 141388 317191 143422 317835
rect 100593 313001 102621 317191
rect 141394 313182 143422 317191
rect 189886 317191 191921 317835
rect 100645 312811 102544 313001
rect 141394 312811 143293 313182
rect 189886 313114 191914 317191
rect 189968 312811 191867 313114
rect 94867 312309 107106 312811
rect 94867 312308 104258 312309
rect 94867 311126 97293 312308
rect 98417 311127 104258 312308
rect 105382 311127 107106 312309
rect 98417 311126 107106 311127
rect 94867 310704 107106 311126
rect 136177 312317 220036 312811
rect 136177 312316 152899 312317
rect 136177 312315 145941 312316
rect 136177 311133 138976 312315
rect 140100 311134 145941 312315
rect 147065 311135 152899 312316
rect 154023 312316 173739 312317
rect 154023 312315 166781 312316
rect 154023 311135 159816 312315
rect 147065 311134 159816 311135
rect 140100 311133 159816 311134
rect 160940 312230 166781 312315
rect 160940 311133 164506 312230
rect 136177 311055 164506 311133
rect 165772 311134 166781 312230
rect 167905 311135 173739 312316
rect 174863 312313 220036 312317
rect 174863 312312 215310 312313
rect 174863 312311 194467 312312
rect 174863 312310 187509 312311
rect 174863 311135 180544 312310
rect 167905 311134 180544 311135
rect 165772 311128 180544 311134
rect 181668 311129 187509 312310
rect 188633 311130 194467 312311
rect 195591 312311 208352 312312
rect 195591 311130 201387 312311
rect 188633 311129 201387 311130
rect 202511 311130 208352 312311
rect 209476 311131 215310 312312
rect 216434 311131 220036 312313
rect 209476 311130 220036 311131
rect 202511 311129 220036 311130
rect 181668 311128 220036 311129
rect 165772 311055 220036 311128
rect 136177 310704 220036 311055
rect 100645 305681 102544 310704
rect 141394 305681 143293 310704
rect 189968 305681 191867 310704
rect 78600 305199 220036 305681
rect 78600 305198 90201 305199
rect 78600 304016 83243 305198
rect 84367 304017 90201 305198
rect 91325 305187 220036 305199
rect 91325 305186 152625 305187
rect 91325 305185 145667 305186
rect 91325 305181 138702 305185
rect 91325 305180 131785 305181
rect 91325 305179 110942 305180
rect 91325 305178 103984 305179
rect 91325 304017 97019 305178
rect 84367 304016 97019 304017
rect 78600 303996 97019 304016
rect 98143 303997 103984 305178
rect 105108 303998 110942 305179
rect 112066 305179 124827 305180
rect 112066 303998 117862 305179
rect 105108 303997 117862 303998
rect 118986 303998 124827 305179
rect 125951 303999 131785 305180
rect 132909 304003 138702 305181
rect 139826 304004 145667 305185
rect 146791 304005 152625 305186
rect 153749 305186 173465 305187
rect 153749 305185 166507 305186
rect 153749 304005 159542 305185
rect 146791 304004 159542 304005
rect 139826 304003 159542 304004
rect 160666 305144 166507 305185
rect 160666 304003 164487 305144
rect 132909 303999 164487 304003
rect 125951 303998 164487 303999
rect 118986 303997 164487 303998
rect 98143 303996 164487 303997
rect 78600 303969 164487 303996
rect 165753 304004 166507 305144
rect 167631 304005 173465 305186
rect 174589 305183 220036 305187
rect 174589 305182 215036 305183
rect 174589 305181 194193 305182
rect 174589 305180 187235 305181
rect 174589 304005 180270 305180
rect 167631 304004 180270 304005
rect 165753 303998 180270 304004
rect 181394 303999 187235 305180
rect 188359 304000 194193 305181
rect 195317 305181 208078 305182
rect 195317 304000 201113 305181
rect 188359 303999 201113 304000
rect 202237 304000 208078 305181
rect 209202 304001 215036 305182
rect 216160 304001 220036 305183
rect 209202 304000 220036 304001
rect 202237 303999 220036 304000
rect 181394 303998 220036 303999
rect 165753 303969 220036 303998
rect 78600 303574 220036 303969
rect 100645 302753 102650 303574
rect 141394 302753 143412 303574
rect 100686 296667 102650 302753
rect 141448 296736 143412 302753
rect 189963 297099 191927 303574
rect 189963 296770 191956 297099
rect 100734 296452 102633 296667
rect 141483 296452 143382 296736
rect 190057 296452 191956 296770
rect 94994 295950 107999 296452
rect 94994 295949 104347 295950
rect 94994 294767 97382 295949
rect 98506 294768 104347 295949
rect 105471 294768 107999 295950
rect 98506 294767 107999 294768
rect 94994 294345 107999 294767
rect 136177 295958 170475 296452
rect 136177 295957 152988 295958
rect 136177 295956 146030 295957
rect 136177 294774 139065 295956
rect 140189 294775 146030 295956
rect 147154 294776 152988 295957
rect 154112 295957 170475 295958
rect 154112 295956 166870 295957
rect 154112 294776 159905 295956
rect 147154 294775 159905 294776
rect 140189 294774 159905 294775
rect 161029 295871 166870 295956
rect 161029 294774 164595 295871
rect 136177 294696 164595 294774
rect 165861 294775 166870 295871
rect 167994 294775 170475 295957
rect 165861 294696 170475 294775
rect 136177 294345 170475 294696
rect 183225 295953 197760 296452
rect 183225 295952 194556 295953
rect 183225 294770 187598 295952
rect 188722 294771 194556 295952
rect 195680 294771 197760 295953
rect 188722 294770 197760 294771
rect 183225 294345 197760 294770
rect 100734 289322 102633 294345
rect 141483 289322 143382 294345
rect 190057 289322 191956 294345
rect 94994 288820 107999 289322
rect 94994 288819 104073 288820
rect 94994 287637 97108 288819
rect 98232 287638 104073 288819
rect 105197 287638 107999 288820
rect 98232 287637 107999 287638
rect 94994 287215 107999 287637
rect 136177 288828 170475 289322
rect 136177 288827 152714 288828
rect 136177 288826 145756 288827
rect 136177 287644 138791 288826
rect 139915 287645 145756 288826
rect 146880 287646 152714 288827
rect 153838 288827 170475 288828
rect 153838 288826 166596 288827
rect 153838 287646 159631 288826
rect 146880 287645 159631 287646
rect 139915 287644 159631 287645
rect 160755 288785 166596 288826
rect 160755 287644 164576 288785
rect 136177 287610 164576 287644
rect 165842 287645 166596 288785
rect 167720 287645 170475 288827
rect 165842 287610 170475 287645
rect 136177 287215 170475 287610
rect 183225 288823 197760 289322
rect 183225 288822 194282 288823
rect 183225 287640 187324 288822
rect 188448 287641 194282 288822
rect 195406 287641 197760 288823
rect 188448 287640 197760 287641
rect 183225 287215 197760 287640
rect 100734 282909 102633 287215
rect 141483 282909 143382 287215
rect 190057 282909 191956 287215
rect 94994 282407 107999 282909
rect 94994 282406 104181 282407
rect 94994 281224 97216 282406
rect 98340 281225 104181 282406
rect 105305 281225 107999 282407
rect 98340 281224 107999 281225
rect 94994 280802 107999 281224
rect 136177 282415 170475 282909
rect 136177 282414 152822 282415
rect 136177 282413 145864 282414
rect 136177 281231 138899 282413
rect 140023 281232 145864 282413
rect 146988 281233 152822 282414
rect 153946 282414 170475 282415
rect 153946 282413 166704 282414
rect 153946 281233 159739 282413
rect 146988 281232 159739 281233
rect 140023 281231 159739 281232
rect 160863 282383 166704 282413
rect 160863 281231 164539 282383
rect 136177 281208 164539 281231
rect 165805 281232 166704 282383
rect 167828 281232 170475 282414
rect 165805 281208 170475 281232
rect 136177 280802 170475 281208
rect 183225 282410 197760 282909
rect 183225 282409 194390 282410
rect 183225 281227 187432 282409
rect 188556 281228 194390 282409
rect 195514 281228 197760 282410
rect 188556 281227 197760 281228
rect 183225 280802 197760 281227
rect 100327 274044 102704 280802
rect 141089 274044 143466 280802
rect 189461 274691 191838 280802
rect 189461 274044 192007 274691
rect 66323 273562 226094 274044
rect 66323 272380 69775 273562
rect 70899 273561 90615 273562
rect 70899 273560 83657 273561
rect 70899 272380 76692 273560
rect 66323 272378 76692 272380
rect 77816 272379 83657 273560
rect 84781 272380 90615 273561
rect 91739 273550 226094 273562
rect 91739 273549 153039 273550
rect 91739 273548 146081 273549
rect 91739 273544 139116 273548
rect 91739 273543 132199 273544
rect 91739 273542 111356 273543
rect 91739 273541 104398 273542
rect 91739 272380 97433 273541
rect 84781 272379 97433 272380
rect 77816 272378 97433 272379
rect 66323 272359 97433 272378
rect 98557 272360 104398 273541
rect 105522 272361 111356 273542
rect 112480 273542 125241 273543
rect 112480 272361 118276 273542
rect 105522 272360 118276 272361
rect 119400 272361 125241 273542
rect 126365 272362 132199 273543
rect 133323 272366 139116 273544
rect 140240 272367 146081 273548
rect 147205 272368 153039 273549
rect 154163 273549 173879 273550
rect 154163 273548 166921 273549
rect 154163 272368 159956 273548
rect 147205 272367 159956 272368
rect 140240 272366 159956 272367
rect 161080 273463 166921 273548
rect 161080 272366 164646 273463
rect 133323 272362 164646 272366
rect 126365 272361 164646 272362
rect 119400 272360 164646 272361
rect 98557 272359 164646 272360
rect 66323 272288 164646 272359
rect 165912 272367 166921 273463
rect 168045 272368 173879 273549
rect 175003 273546 222367 273550
rect 175003 273545 215450 273546
rect 175003 273544 194607 273545
rect 175003 273543 187649 273544
rect 175003 272368 180684 273543
rect 168045 272367 180684 272368
rect 165912 272361 180684 272367
rect 181808 272362 187649 273543
rect 188773 272363 194607 273544
rect 195731 273544 208492 273545
rect 195731 272363 201527 273544
rect 188773 272362 201527 272363
rect 202651 272363 208492 273544
rect 209616 272364 215450 273545
rect 216574 272368 222367 273546
rect 223491 272368 226094 273550
rect 216574 272364 226094 272368
rect 209616 272363 226094 272364
rect 202651 272362 226094 272363
rect 181808 272361 226094 272362
rect 165912 272288 226094 272361
rect 66323 271937 226094 272288
rect 100785 266914 102684 271937
rect 141534 266914 143433 271937
rect 190108 266914 192007 271937
rect 66323 266432 226094 266914
rect 66323 265250 69501 266432
rect 70625 266431 90341 266432
rect 70625 266430 83383 266431
rect 70625 265250 76418 266430
rect 66323 265248 76418 265250
rect 77542 265249 83383 266430
rect 84507 265250 90341 266431
rect 91465 266420 226094 266432
rect 91465 266419 152765 266420
rect 91465 266418 145807 266419
rect 91465 266414 138842 266418
rect 91465 266413 131925 266414
rect 91465 266412 111082 266413
rect 91465 266411 104124 266412
rect 91465 265250 97159 266411
rect 84507 265249 97159 265250
rect 77542 265248 97159 265249
rect 66323 265229 97159 265248
rect 98283 265230 104124 266411
rect 105248 265231 111082 266412
rect 112206 266412 124967 266413
rect 112206 265231 118002 266412
rect 105248 265230 118002 265231
rect 119126 265231 124967 266412
rect 126091 265232 131925 266413
rect 133049 265236 138842 266414
rect 139966 265237 145807 266418
rect 146931 265238 152765 266419
rect 153889 266419 173605 266420
rect 153889 266418 166647 266419
rect 153889 265238 159682 266418
rect 146931 265237 159682 265238
rect 139966 265236 159682 265237
rect 160806 266377 166647 266418
rect 160806 265236 164627 266377
rect 133049 265232 164627 265236
rect 126091 265231 164627 265232
rect 119126 265230 164627 265231
rect 98283 265229 164627 265230
rect 66323 265202 164627 265229
rect 165893 265237 166647 266377
rect 167771 265238 173605 266419
rect 174729 266416 222093 266420
rect 174729 266415 215176 266416
rect 174729 266414 194333 266415
rect 174729 266413 187375 266414
rect 174729 265238 180410 266413
rect 167771 265237 180410 265238
rect 165893 265231 180410 265237
rect 181534 265232 187375 266413
rect 188499 265233 194333 266414
rect 195457 266414 208218 266415
rect 195457 265233 201253 266414
rect 188499 265232 201253 265233
rect 202377 265233 208218 266414
rect 209342 265234 215176 266415
rect 216300 265238 222093 266416
rect 223217 265238 226094 266420
rect 216300 265234 226094 265238
rect 209342 265233 226094 265234
rect 202377 265232 226094 265233
rect 181534 265231 226094 265232
rect 165893 265202 226094 265231
rect 66323 264807 226094 265202
rect 100785 260501 102684 264807
rect 141534 260501 143433 264807
rect 190108 260501 192007 264807
rect 66323 260019 226094 260501
rect 66323 258837 69609 260019
rect 70733 260018 90449 260019
rect 70733 260017 83491 260018
rect 70733 258837 76526 260017
rect 66323 258835 76526 258837
rect 77650 258836 83491 260017
rect 84615 258837 90449 260018
rect 91573 260007 226094 260019
rect 91573 260006 152873 260007
rect 91573 260005 145915 260006
rect 91573 260001 138950 260005
rect 91573 260000 132033 260001
rect 91573 259999 111190 260000
rect 91573 259998 104232 259999
rect 91573 258837 97267 259998
rect 84615 258836 97267 258837
rect 77650 258835 97267 258836
rect 66323 258816 97267 258835
rect 98391 258817 104232 259998
rect 105356 258818 111190 259999
rect 112314 259999 125075 260000
rect 112314 258818 118110 259999
rect 105356 258817 118110 258818
rect 119234 258818 125075 259999
rect 126199 258819 132033 260000
rect 133157 258823 138950 260001
rect 140074 258824 145915 260005
rect 147039 258825 152873 260006
rect 153997 260006 173713 260007
rect 153997 260005 166755 260006
rect 153997 258825 159790 260005
rect 147039 258824 159790 258825
rect 140074 258823 159790 258824
rect 160914 259975 166755 260005
rect 160914 258823 164590 259975
rect 133157 258819 164590 258823
rect 126199 258818 164590 258819
rect 119234 258817 164590 258818
rect 98391 258816 164590 258817
rect 66323 258800 164590 258816
rect 165856 258824 166755 259975
rect 167879 258825 173713 260006
rect 174837 260003 222201 260007
rect 174837 260002 215284 260003
rect 174837 260001 194441 260002
rect 174837 260000 187483 260001
rect 174837 258825 180518 260000
rect 167879 258824 180518 258825
rect 165856 258818 180518 258824
rect 181642 258819 187483 260000
rect 188607 258820 194441 260001
rect 195565 260001 208326 260002
rect 195565 258820 201361 260001
rect 188607 258819 201361 258820
rect 202485 258820 208326 260001
rect 209450 258821 215284 260002
rect 216408 258825 222201 260003
rect 223325 258825 226094 260007
rect 216408 258821 226094 258825
rect 209450 258820 226094 258821
rect 202485 258819 226094 258820
rect 181642 258818 226094 258819
rect 165856 258800 226094 258818
rect 66323 258394 226094 258800
rect 100447 257821 102801 258394
rect 141318 257821 143513 258394
rect 100748 250077 102801 257821
rect 141460 250096 143513 257821
rect 189592 250437 191978 258394
rect 100816 249790 102715 250077
rect 141565 249790 143464 250096
rect 189592 249790 192038 250437
rect 80519 249308 226125 249790
rect 80519 249307 90646 249308
rect 80519 248125 83688 249307
rect 84812 248126 90646 249307
rect 91770 249296 226125 249308
rect 91770 249295 153070 249296
rect 91770 249294 146112 249295
rect 91770 249290 139147 249294
rect 91770 249289 132230 249290
rect 91770 249288 111387 249289
rect 91770 249287 104429 249288
rect 91770 248126 97464 249287
rect 84812 248125 97464 248126
rect 80519 248105 97464 248125
rect 98588 248106 104429 249287
rect 105553 248107 111387 249288
rect 112511 249288 125272 249289
rect 112511 248107 118307 249288
rect 105553 248106 118307 248107
rect 119431 248107 125272 249288
rect 126396 248108 132230 249289
rect 133354 248112 139147 249290
rect 140271 248113 146112 249294
rect 147236 248114 153070 249295
rect 154194 249295 173910 249296
rect 154194 249294 166952 249295
rect 154194 248114 159987 249294
rect 147236 248113 159987 248114
rect 140271 248112 159987 248113
rect 161111 249209 166952 249294
rect 161111 248112 164677 249209
rect 133354 248108 164677 248112
rect 126396 248107 164677 248108
rect 119431 248106 164677 248107
rect 98588 248105 164677 248106
rect 80519 248034 164677 248105
rect 165943 248113 166952 249209
rect 168076 248114 173910 249295
rect 175034 249292 222398 249296
rect 175034 249291 215481 249292
rect 175034 249290 194638 249291
rect 175034 249289 187680 249290
rect 175034 248114 180715 249289
rect 168076 248113 180715 248114
rect 165943 248107 180715 248113
rect 181839 248108 187680 249289
rect 188804 248109 194638 249290
rect 195762 249290 208523 249291
rect 195762 248109 201558 249290
rect 188804 248108 201558 248109
rect 202682 248109 208523 249290
rect 209647 248110 215481 249291
rect 216605 248114 222398 249292
rect 223522 248114 226125 249296
rect 216605 248110 226125 248114
rect 209647 248109 226125 248110
rect 202682 248108 226125 248109
rect 181839 248107 226125 248108
rect 165943 248034 226125 248107
rect 80519 247683 226125 248034
rect 100816 242660 102715 247683
rect 141565 242660 143464 247683
rect 190139 242660 192038 247683
rect 80519 242178 226125 242660
rect 80519 242177 90372 242178
rect 80519 240995 83414 242177
rect 84538 240996 90372 242177
rect 91496 242166 226125 242178
rect 91496 242165 152796 242166
rect 91496 242164 145838 242165
rect 91496 242160 138873 242164
rect 91496 242159 131956 242160
rect 91496 242158 111113 242159
rect 91496 242157 104155 242158
rect 91496 240996 97190 242157
rect 84538 240995 97190 240996
rect 80519 240975 97190 240995
rect 98314 240976 104155 242157
rect 105279 240977 111113 242158
rect 112237 242158 124998 242159
rect 112237 240977 118033 242158
rect 105279 240976 118033 240977
rect 119157 240977 124998 242158
rect 126122 240978 131956 242159
rect 133080 240982 138873 242160
rect 139997 240983 145838 242164
rect 146962 240984 152796 242165
rect 153920 242165 173636 242166
rect 153920 242164 166678 242165
rect 153920 240984 159713 242164
rect 146962 240983 159713 240984
rect 139997 240982 159713 240983
rect 160837 242123 166678 242164
rect 160837 240982 164658 242123
rect 133080 240978 164658 240982
rect 126122 240977 164658 240978
rect 119157 240976 164658 240977
rect 98314 240975 164658 240976
rect 80519 240948 164658 240975
rect 165924 240983 166678 242123
rect 167802 240984 173636 242165
rect 174760 242162 222124 242166
rect 174760 242161 215207 242162
rect 174760 242160 194364 242161
rect 174760 242159 187406 242160
rect 174760 240984 180441 242159
rect 167802 240983 180441 240984
rect 165924 240977 180441 240983
rect 181565 240978 187406 242159
rect 188530 240979 194364 242160
rect 195488 242160 208249 242161
rect 195488 240979 201284 242160
rect 188530 240978 201284 240979
rect 202408 240979 208249 242160
rect 209373 240980 215207 242161
rect 216331 240984 222124 242162
rect 223248 240984 226125 242166
rect 216331 240980 226125 240984
rect 209373 240979 226125 240980
rect 202408 240978 226125 240979
rect 181565 240977 226125 240978
rect 165924 240948 226125 240977
rect 80519 240553 226125 240948
rect 100816 236247 102715 240553
rect 141565 236247 143464 240553
rect 190139 236247 192038 240553
rect 80519 235765 226125 236247
rect 80519 235764 90480 235765
rect 80519 234582 83522 235764
rect 84646 234583 90480 235764
rect 91604 235753 226125 235765
rect 91604 235752 152904 235753
rect 91604 235751 145946 235752
rect 91604 235747 138981 235751
rect 91604 235746 132064 235747
rect 91604 235745 111221 235746
rect 91604 235744 104263 235745
rect 91604 234583 97298 235744
rect 84646 234582 97298 234583
rect 80519 234562 97298 234582
rect 98422 234563 104263 235744
rect 105387 234564 111221 235745
rect 112345 235745 125106 235746
rect 112345 234564 118141 235745
rect 105387 234563 118141 234564
rect 119265 234564 125106 235745
rect 126230 234565 132064 235746
rect 133188 234569 138981 235747
rect 140105 234570 145946 235751
rect 147070 234571 152904 235752
rect 154028 235752 173744 235753
rect 154028 235751 166786 235752
rect 154028 234571 159821 235751
rect 147070 234570 159821 234571
rect 140105 234569 159821 234570
rect 160945 235721 166786 235751
rect 160945 234569 164621 235721
rect 133188 234565 164621 234569
rect 126230 234564 164621 234565
rect 119265 234563 164621 234564
rect 98422 234562 164621 234563
rect 80519 234546 164621 234562
rect 165887 234570 166786 235721
rect 167910 234571 173744 235752
rect 174868 235749 222232 235753
rect 174868 235748 215315 235749
rect 174868 235747 194472 235748
rect 174868 235746 187514 235747
rect 174868 234571 180549 235746
rect 167910 234570 180549 234571
rect 165887 234564 180549 234570
rect 181673 234565 187514 235746
rect 188638 234566 194472 235747
rect 195596 235747 208357 235748
rect 195596 234566 201392 235747
rect 188638 234565 201392 234566
rect 202516 234566 208357 235747
rect 209481 234567 215315 235748
rect 216439 234571 222232 235749
rect 223356 234571 226125 235753
rect 216439 234567 226125 234571
rect 209481 234566 226125 234567
rect 202516 234565 226125 234566
rect 181673 234564 226125 234565
rect 165887 234546 226125 234564
rect 80519 234140 226125 234546
rect 100478 233567 102850 234140
rect 141349 233567 143486 234140
rect 100933 230190 102850 233567
rect 100940 229524 102839 230190
rect 141413 229545 143486 233567
rect 189617 233567 191774 234140
rect 141413 229524 143588 229545
rect 189617 229524 191690 233567
rect 69559 229503 191690 229524
rect 192275 229503 226544 229524
rect 69559 229042 226544 229503
rect 69559 227860 69930 229042
rect 71054 229041 90770 229042
rect 71054 229040 83812 229041
rect 71054 227860 76847 229040
rect 69559 227858 76847 227860
rect 77971 227859 83812 229040
rect 84936 227860 90770 229041
rect 91894 229030 226544 229042
rect 91894 229029 153194 229030
rect 91894 229028 146236 229029
rect 91894 229024 139271 229028
rect 91894 229023 132354 229024
rect 91894 229022 111511 229023
rect 91894 229021 104553 229022
rect 91894 227860 97588 229021
rect 84936 227859 97588 227860
rect 77971 227858 97588 227859
rect 69559 227839 97588 227858
rect 98712 227840 104553 229021
rect 105677 227841 111511 229022
rect 112635 229022 125396 229023
rect 112635 227841 118431 229022
rect 105677 227840 118431 227841
rect 119555 227841 125396 229022
rect 126520 227842 132354 229023
rect 133478 227846 139271 229024
rect 140395 227847 146236 229028
rect 147360 227848 153194 229029
rect 154318 229029 174034 229030
rect 154318 229028 167076 229029
rect 154318 227848 160111 229028
rect 147360 227847 160111 227848
rect 140395 227846 160111 227847
rect 161235 228943 167076 229028
rect 161235 227846 164801 228943
rect 133478 227842 164801 227846
rect 126520 227841 164801 227842
rect 119555 227840 164801 227841
rect 98712 227839 164801 227840
rect 69559 227768 164801 227839
rect 166067 227847 167076 228943
rect 168200 227848 174034 229029
rect 175158 229026 222522 229030
rect 175158 229025 215605 229026
rect 175158 229024 194762 229025
rect 175158 229023 187804 229024
rect 175158 227848 180839 229023
rect 168200 227847 180839 227848
rect 166067 227841 180839 227847
rect 181963 227842 187804 229023
rect 188928 227843 194762 229024
rect 195886 229024 208647 229025
rect 195886 227843 201682 229024
rect 188928 227842 201682 227843
rect 202806 227843 208647 229024
rect 209771 227844 215605 229025
rect 216729 227848 222522 229026
rect 223646 227848 226544 229030
rect 216729 227844 226544 227848
rect 209771 227843 226544 227844
rect 202806 227842 226544 227843
rect 181963 227841 226544 227842
rect 166067 227768 226544 227841
rect 69559 227417 226544 227768
rect 100884 226887 102839 227417
rect 141689 226887 143654 227417
rect 100884 223662 102836 226887
rect 141702 224776 143654 226887
rect 141669 223662 143654 224776
rect 190179 226887 192162 227417
rect 190179 224776 192131 226887
rect 190179 223662 192142 224776
rect 69559 223180 226544 223662
rect 69559 221998 69910 223180
rect 71034 223179 90750 223180
rect 71034 223178 83792 223179
rect 71034 221998 76827 223178
rect 69559 221996 76827 221998
rect 77951 221997 83792 223178
rect 84916 221998 90750 223179
rect 91874 223168 226544 223180
rect 91874 223167 153174 223168
rect 91874 223166 146216 223167
rect 91874 223162 139251 223166
rect 91874 223161 132334 223162
rect 91874 223160 111491 223161
rect 91874 223159 104533 223160
rect 91874 221998 97568 223159
rect 84916 221997 97568 221998
rect 77951 221996 97568 221997
rect 69559 221977 97568 221996
rect 98692 221978 104533 223159
rect 105657 221979 111491 223160
rect 112615 223160 125376 223161
rect 112615 221979 118411 223160
rect 105657 221978 118411 221979
rect 119535 221979 125376 223160
rect 126500 221980 132334 223161
rect 133458 221984 139251 223162
rect 140375 221985 146216 223166
rect 147340 221986 153174 223167
rect 154298 223167 174014 223168
rect 154298 223166 167056 223167
rect 154298 221986 160091 223166
rect 147340 221985 160091 221986
rect 140375 221984 160091 221985
rect 161215 223081 167056 223166
rect 161215 221984 164781 223081
rect 133458 221980 164781 221984
rect 126500 221979 164781 221980
rect 119535 221978 164781 221979
rect 98692 221977 164781 221978
rect 69559 221906 164781 221977
rect 166047 221985 167056 223081
rect 168180 221986 174014 223167
rect 175138 223164 222502 223168
rect 175138 223163 215585 223164
rect 175138 223162 194742 223163
rect 175138 223161 187784 223162
rect 175138 221986 180819 223161
rect 168180 221985 180819 221986
rect 166047 221979 180819 221985
rect 181943 221980 187784 223161
rect 188908 221981 194742 223162
rect 195866 223162 208627 223163
rect 195866 221981 201662 223162
rect 188908 221980 201662 221981
rect 202786 221981 208627 223162
rect 209751 221982 215585 223163
rect 216709 221986 222502 223164
rect 223626 221986 226544 223168
rect 216709 221982 226544 221986
rect 209751 221981 226544 221982
rect 202786 221980 226544 221981
rect 181943 221979 226544 221980
rect 166047 221906 226544 221979
rect 69559 221555 226544 221906
rect 59047 212180 60999 220696
rect 100884 213295 102836 221555
rect 141669 221025 143654 221555
rect 100884 212669 102859 213295
rect 59084 211599 60983 212180
rect 66008 211599 96677 211657
rect 100960 211599 102859 212669
rect 141702 212477 143654 221025
rect 190179 221025 192142 221555
rect 190179 216801 192131 221025
rect 141709 211599 143608 212477
rect 18223 211578 31024 211599
rect 33596 211578 108521 211599
rect 18223 211116 108521 211578
rect 18223 211115 62992 211116
rect 18223 211111 56027 211115
rect 18223 211110 49110 211111
rect 18223 211109 28267 211110
rect 18223 209927 21309 211109
rect 22433 209928 28267 211109
rect 29391 211109 42152 211110
rect 29391 209928 35187 211109
rect 22433 209927 35187 209928
rect 36311 209928 42152 211109
rect 43276 209929 49110 211110
rect 50234 209933 56027 211111
rect 57151 209934 62992 211115
rect 64116 211097 108521 211116
rect 64116 211096 104573 211097
rect 64116 209934 97608 211096
rect 57151 209933 97608 209934
rect 50234 209929 97608 209933
rect 43276 209928 97608 209929
rect 36311 209927 97608 209928
rect 18223 209914 97608 209927
rect 98732 209915 104573 211096
rect 105697 209915 108521 211097
rect 98732 209914 108521 209915
rect 18223 209558 108521 209914
rect 18223 209492 67183 209558
rect 94909 209492 108521 209558
rect 136248 211105 170528 211599
rect 136248 211104 153214 211105
rect 136248 211103 146256 211104
rect 136248 209921 139291 211103
rect 140415 209922 146256 211103
rect 147380 209923 153214 211104
rect 154338 211104 170528 211105
rect 154338 211103 167096 211104
rect 154338 209923 160131 211103
rect 147380 209922 160131 209923
rect 140415 209921 160131 209922
rect 161255 211018 167096 211103
rect 161255 209921 164821 211018
rect 136248 209843 164821 209921
rect 166087 209922 167096 211018
rect 168220 209922 170528 211104
rect 166087 209843 170528 209922
rect 136248 209492 170528 209843
rect 31238 204469 33137 209492
rect 59084 204469 60983 209492
rect 100960 204469 102859 209492
rect 141709 204469 143608 209492
rect 18223 203986 67183 204469
rect 18223 203985 62718 203986
rect 18223 203981 55753 203985
rect 18223 203980 48836 203981
rect 18223 203979 27993 203980
rect 18223 202797 21035 203979
rect 22159 202798 27993 203979
rect 29117 203979 41878 203980
rect 29117 202798 34913 203979
rect 22159 202797 34913 202798
rect 36037 202798 41878 203979
rect 43002 202799 48836 203980
rect 49960 202803 55753 203981
rect 56877 202804 62718 203985
rect 63842 202804 67183 203986
rect 56877 202803 67183 202804
rect 49960 202799 67183 202803
rect 43002 202798 67183 202799
rect 36037 202797 67183 202798
rect 18223 202362 67183 202797
rect 94909 203967 108521 204469
rect 94909 203966 104299 203967
rect 94909 202784 97334 203966
rect 98458 202785 104299 203966
rect 105423 202785 108521 203967
rect 98458 202784 108521 202785
rect 94909 202362 108521 202784
rect 136248 203975 170528 204469
rect 136248 203974 152940 203975
rect 136248 203973 145982 203974
rect 136248 202791 139017 203973
rect 140141 202792 145982 203973
rect 147106 202793 152940 203974
rect 154064 203974 170528 203975
rect 154064 203973 166822 203974
rect 154064 202793 159857 203973
rect 147106 202792 159857 202793
rect 140141 202791 159857 202792
rect 160981 203932 166822 203973
rect 160981 202791 164802 203932
rect 136248 202757 164802 202791
rect 166068 202792 166822 203932
rect 167946 202792 170528 203974
rect 166068 202757 170528 202792
rect 136248 202362 170528 202757
rect 31238 198056 33137 202362
rect 59084 198056 60983 202362
rect 100960 198056 102859 202362
rect 141709 198056 143608 202362
rect 18223 197573 67183 198056
rect 18223 197572 62826 197573
rect 18223 197568 55861 197572
rect 18223 197567 48944 197568
rect 18223 197566 28101 197567
rect 18223 196384 21143 197566
rect 22267 196385 28101 197566
rect 29225 197566 41986 197567
rect 29225 196385 35021 197566
rect 22267 196384 35021 196385
rect 36145 196385 41986 197566
rect 43110 196386 48944 197567
rect 50068 196390 55861 197568
rect 56985 196391 62826 197572
rect 63950 196391 67183 197573
rect 56985 196390 67183 196391
rect 50068 196386 67183 196390
rect 43110 196385 67183 196386
rect 36145 196384 67183 196385
rect 18223 195949 67183 196384
rect 94909 197554 108521 198056
rect 94909 197553 104407 197554
rect 94909 196371 97442 197553
rect 98566 196372 104407 197553
rect 105531 196372 108521 197554
rect 98566 196371 108521 196372
rect 94909 195949 108521 196371
rect 136248 197562 170528 198056
rect 136248 197561 153048 197562
rect 136248 197560 146090 197561
rect 136248 196378 139125 197560
rect 140249 196379 146090 197560
rect 147214 196380 153048 197561
rect 154172 197561 170528 197562
rect 154172 197560 166930 197561
rect 154172 196380 159965 197560
rect 147214 196379 159965 196380
rect 140249 196378 159965 196379
rect 161089 197530 166930 197560
rect 161089 196378 164765 197530
rect 136248 196355 164765 196378
rect 166031 196379 166930 197530
rect 168054 196379 170528 197561
rect 166031 196355 170528 196379
rect 136248 195949 170528 196355
rect 30914 195886 33004 195949
rect 58685 195928 60775 195949
rect 100622 194676 102712 195949
rect 141493 194676 143583 195949
rect 100622 193706 102846 194676
rect 141493 193706 143595 194676
rect 94909 193204 108521 193706
rect 94909 193203 104560 193204
rect 94909 192021 97595 193203
rect 98719 192022 104560 193203
rect 105684 192022 108521 193204
rect 98719 192021 108521 192022
rect 94909 191599 108521 192021
rect 136248 193212 170528 193706
rect 136248 193211 153201 193212
rect 136248 193210 146243 193211
rect 136248 192028 139278 193210
rect 140402 192029 146243 193210
rect 147367 192030 153201 193211
rect 154325 193211 170528 193212
rect 154325 193210 167083 193211
rect 154325 192030 160118 193210
rect 147367 192029 160118 192030
rect 140402 192028 160118 192029
rect 161242 193125 167083 193210
rect 161242 192028 164808 193125
rect 136248 191950 164808 192028
rect 166074 192029 167083 193125
rect 168207 192029 170528 193211
rect 166074 191950 170528 192029
rect 136248 191599 170528 191950
rect 100947 186576 102846 191599
rect 141696 186576 143595 191599
rect 190120 189863 192151 216801
rect 267372 212458 269324 215436
rect 267418 211599 269317 212458
rect 260514 211108 275385 211599
rect 260514 211107 271403 211108
rect 260514 209925 264445 211107
rect 265569 209926 271403 211107
rect 272527 209926 275385 211108
rect 265569 209925 275385 209926
rect 260514 209492 275385 209925
rect 267418 204469 269317 209492
rect 260514 203978 275385 204469
rect 260514 203977 271129 203978
rect 260514 202795 264171 203977
rect 265295 202796 271129 203977
rect 272253 202796 275385 203978
rect 265295 202795 275385 202796
rect 260514 202362 275385 202795
rect 267418 198056 269317 202362
rect 260514 197565 275385 198056
rect 260514 197564 271237 197565
rect 260514 196382 264279 197564
rect 265403 196383 271237 197564
rect 272361 196383 275385 197565
rect 265403 196382 275385 196383
rect 260514 195949 275385 196382
rect 267305 193706 269395 195949
rect 260514 193215 275385 193706
rect 260514 193214 271390 193215
rect 260514 192032 264432 193214
rect 265556 192033 271390 193214
rect 272514 192033 275385 193215
rect 265556 192032 275385 192033
rect 260514 191599 275385 192032
rect 190120 188908 192169 189863
rect 190270 186576 192169 188908
rect 232553 186576 234452 189863
rect 267405 186576 269304 191599
rect 73528 186094 108521 186576
rect 73528 186093 90503 186094
rect 73528 186092 83545 186093
rect 73528 184910 76580 186092
rect 77704 184911 83545 186092
rect 84669 184912 90503 186093
rect 91627 186074 108521 186094
rect 91627 186073 104286 186074
rect 91627 184912 97321 186073
rect 84669 184911 97321 184912
rect 77704 184910 97321 184911
rect 73528 184891 97321 184910
rect 98445 184892 104286 186073
rect 105410 184892 108521 186074
rect 98445 184891 108521 184892
rect 73528 184469 108521 184891
rect 136248 186538 279909 186576
rect 136248 186085 280952 186538
rect 136248 186084 271116 186085
rect 136248 186083 236178 186084
rect 136248 186082 229220 186083
rect 136248 186081 152927 186082
rect 136248 186080 145969 186081
rect 136248 184898 139004 186080
rect 140128 184899 145969 186080
rect 147093 184900 152927 186081
rect 154051 186081 173767 186082
rect 154051 186080 166809 186081
rect 154051 184900 159844 186080
rect 147093 184899 159844 184900
rect 140128 184898 159844 184899
rect 160968 186039 166809 186080
rect 160968 184898 164789 186039
rect 136248 184864 164789 184898
rect 166055 184899 166809 186039
rect 167933 184900 173767 186081
rect 174891 186078 222255 186082
rect 174891 186077 215338 186078
rect 174891 186076 194495 186077
rect 174891 186075 187537 186076
rect 174891 184900 180572 186075
rect 167933 184899 180572 184900
rect 166055 184893 180572 184899
rect 181696 184894 187537 186075
rect 188661 184895 194495 186076
rect 195619 186076 208380 186077
rect 195619 184895 201415 186076
rect 188661 184894 201415 184895
rect 202539 184895 208380 186076
rect 209504 184896 215338 186077
rect 216462 184900 222255 186078
rect 223379 184901 229220 186082
rect 230344 184902 236178 186083
rect 237302 186083 257018 186084
rect 237302 186082 250060 186083
rect 237302 184902 243095 186082
rect 230344 184901 243095 184902
rect 223379 184900 243095 184901
rect 244219 184901 250060 186082
rect 251184 184902 257018 186083
rect 258142 184902 264158 186084
rect 265282 184903 271116 186084
rect 272240 186075 280952 186085
rect 272240 184903 278252 186075
rect 265282 184902 278252 184903
rect 251184 184901 278252 184902
rect 244219 184900 278252 184901
rect 216462 184896 278252 184900
rect 209504 184895 278252 184896
rect 202539 184894 278252 184895
rect 181696 184893 278252 184894
rect 279376 184893 280952 186075
rect 166055 184864 280952 184893
rect 136248 184488 280952 184864
rect 136248 184469 279909 184488
rect 100947 180163 102846 184469
rect 141696 180163 143595 184469
rect 190270 180163 192169 184469
rect 232553 180163 234452 184469
rect 267405 180163 269304 184469
rect 73528 180125 280017 180163
rect 73528 179681 281060 180125
rect 73528 179680 90611 179681
rect 73528 179679 83653 179680
rect 73528 178497 76688 179679
rect 77812 178498 83653 179679
rect 84777 178499 90611 179680
rect 91735 179672 281060 179681
rect 91735 179671 271224 179672
rect 91735 179670 236286 179671
rect 91735 179669 229328 179670
rect 91735 179668 153035 179669
rect 91735 179667 146077 179668
rect 91735 179663 139112 179667
rect 91735 179662 132195 179663
rect 91735 179661 111352 179662
rect 91735 179660 104394 179661
rect 91735 178499 97429 179660
rect 84777 178498 97429 178499
rect 77812 178497 97429 178498
rect 73528 178478 97429 178497
rect 98553 178479 104394 179660
rect 105518 178480 111352 179661
rect 112476 179661 125237 179662
rect 112476 178480 118272 179661
rect 105518 178479 118272 178480
rect 119396 178480 125237 179661
rect 126361 178481 132195 179662
rect 133319 178485 139112 179663
rect 140236 178486 146077 179667
rect 147201 178487 153035 179668
rect 154159 179668 173875 179669
rect 154159 179667 166917 179668
rect 154159 178487 159952 179667
rect 147201 178486 159952 178487
rect 140236 178485 159952 178486
rect 161076 179637 166917 179667
rect 161076 178485 164752 179637
rect 133319 178481 164752 178485
rect 126361 178480 164752 178481
rect 119396 178479 164752 178480
rect 98553 178478 164752 178479
rect 73528 178462 164752 178478
rect 166018 178486 166917 179637
rect 168041 178487 173875 179668
rect 174999 179665 222363 179669
rect 174999 179664 215446 179665
rect 174999 179663 194603 179664
rect 174999 179662 187645 179663
rect 174999 178487 180680 179662
rect 168041 178486 180680 178487
rect 166018 178480 180680 178486
rect 181804 178481 187645 179662
rect 188769 178482 194603 179663
rect 195727 179663 208488 179664
rect 195727 178482 201523 179663
rect 188769 178481 201523 178482
rect 202647 178482 208488 179663
rect 209612 178483 215446 179664
rect 216570 178487 222363 179665
rect 223487 178488 229328 179669
rect 230452 178489 236286 179670
rect 237410 179670 257126 179671
rect 237410 179669 250168 179670
rect 237410 178489 243203 179669
rect 230452 178488 243203 178489
rect 223487 178487 243203 178488
rect 244327 178488 250168 179669
rect 251292 178489 257126 179670
rect 258250 178489 264266 179671
rect 265390 178490 271224 179671
rect 272348 179662 281060 179672
rect 272348 178490 278360 179662
rect 265390 178489 278360 178490
rect 251292 178488 278360 178489
rect 244327 178487 278360 178488
rect 216570 178483 278360 178487
rect 209612 178482 278360 178483
rect 202647 178481 278360 178482
rect 181804 178480 278360 178481
rect 279484 178480 281060 179662
rect 166018 178462 281060 178480
rect 73528 178075 281060 178462
rect 73528 178056 280017 178075
rect 100609 176358 102830 178056
rect 100674 174249 102830 176358
rect 141462 174249 143618 178056
rect 189815 176358 192042 178056
rect 189886 174249 192042 176358
rect 232171 176358 234269 178056
rect 267266 176358 269382 178056
rect 232171 175011 234265 176358
rect 267266 175011 269360 176358
rect 232171 174249 234275 175011
rect 267228 174249 269360 175011
rect 65177 174211 279732 174249
rect 65177 173767 280775 174211
rect 65177 172585 69486 173767
rect 70610 173766 90326 173767
rect 70610 173765 83368 173766
rect 70610 172585 76403 173765
rect 65177 172583 76403 172585
rect 77527 172584 83368 173765
rect 84492 172585 90326 173766
rect 91450 173758 280775 173767
rect 91450 173757 270939 173758
rect 91450 173756 236001 173757
rect 91450 173755 229043 173756
rect 91450 173754 152750 173755
rect 91450 173753 145792 173754
rect 91450 173749 138827 173753
rect 91450 173748 131910 173749
rect 91450 173747 111067 173748
rect 91450 173746 104109 173747
rect 91450 172585 97144 173746
rect 84492 172584 97144 172585
rect 77527 172583 97144 172584
rect 65177 172564 97144 172583
rect 98268 172565 104109 173746
rect 105233 172566 111067 173747
rect 112191 173747 124952 173748
rect 112191 172566 117987 173747
rect 105233 172565 117987 172566
rect 119111 172566 124952 173747
rect 126076 172567 131910 173748
rect 133034 172571 138827 173749
rect 139951 172572 145792 173753
rect 146916 172573 152750 173754
rect 153874 173754 173590 173755
rect 153874 173753 166632 173754
rect 153874 172573 159667 173753
rect 146916 172572 159667 172573
rect 139951 172571 159667 172572
rect 160791 173712 166632 173753
rect 160791 172571 164612 173712
rect 133034 172567 164612 172571
rect 126076 172566 164612 172567
rect 119111 172565 164612 172566
rect 98268 172564 164612 172565
rect 65177 172537 164612 172564
rect 165878 172572 166632 173712
rect 167756 172573 173590 173754
rect 174714 173751 222078 173755
rect 174714 173750 215161 173751
rect 174714 173749 194318 173750
rect 174714 173748 187360 173749
rect 174714 172573 180395 173748
rect 167756 172572 180395 172573
rect 165878 172566 180395 172572
rect 181519 172567 187360 173748
rect 188484 172568 194318 173749
rect 195442 173749 208203 173750
rect 195442 172568 201238 173749
rect 188484 172567 201238 172568
rect 202362 172568 208203 173749
rect 209327 172569 215161 173750
rect 216285 172573 222078 173751
rect 223202 172574 229043 173755
rect 230167 172575 236001 173756
rect 237125 173756 256841 173757
rect 237125 173755 249883 173756
rect 237125 172575 242918 173755
rect 230167 172574 242918 172575
rect 223202 172573 242918 172574
rect 244042 172574 249883 173755
rect 251007 172575 256841 173756
rect 257965 172575 263981 173757
rect 265105 172576 270939 173757
rect 272063 173748 280775 173758
rect 272063 172576 278075 173748
rect 265105 172575 278075 172576
rect 251007 172574 278075 172575
rect 244042 172573 278075 172574
rect 216285 172569 278075 172573
rect 209327 172568 278075 172569
rect 202362 172567 278075 172568
rect 181519 172566 278075 172567
rect 279199 172566 280775 173748
rect 165878 172537 280775 172566
rect 65177 172161 280775 172537
rect 65177 172142 279732 172161
rect 100674 167836 102830 172142
rect 141462 167836 143618 172142
rect 189886 167836 192042 172142
rect 232171 167836 234275 172142
rect 267228 167836 269360 172142
rect 65177 167798 279840 167836
rect 65177 167354 280883 167798
rect 65177 166172 69594 167354
rect 70718 167353 90434 167354
rect 70718 167352 83476 167353
rect 70718 166172 76511 167352
rect 65177 166170 76511 166172
rect 77635 166171 83476 167352
rect 84600 166172 90434 167353
rect 91558 167345 280883 167354
rect 91558 167344 271047 167345
rect 91558 167343 236109 167344
rect 91558 167342 229151 167343
rect 91558 167341 152858 167342
rect 91558 167340 145900 167341
rect 91558 167336 138935 167340
rect 91558 167335 132018 167336
rect 91558 167334 111175 167335
rect 91558 167333 104217 167334
rect 91558 166172 97252 167333
rect 84600 166171 97252 166172
rect 77635 166170 97252 166171
rect 65177 166151 97252 166170
rect 98376 166152 104217 167333
rect 105341 166153 111175 167334
rect 112299 167334 125060 167335
rect 112299 166153 118095 167334
rect 105341 166152 118095 166153
rect 119219 166153 125060 167334
rect 126184 166154 132018 167335
rect 133142 166158 138935 167336
rect 140059 166159 145900 167340
rect 147024 166160 152858 167341
rect 153982 167341 173698 167342
rect 153982 167340 166740 167341
rect 153982 166160 159775 167340
rect 147024 166159 159775 166160
rect 140059 166158 159775 166159
rect 160899 167310 166740 167340
rect 160899 166158 164575 167310
rect 133142 166154 164575 166158
rect 126184 166153 164575 166154
rect 119219 166152 164575 166153
rect 98376 166151 164575 166152
rect 65177 166135 164575 166151
rect 165841 166159 166740 167310
rect 167864 166160 173698 167341
rect 174822 167338 222186 167342
rect 174822 167337 215269 167338
rect 174822 167336 194426 167337
rect 174822 167335 187468 167336
rect 174822 166160 180503 167335
rect 167864 166159 180503 166160
rect 165841 166153 180503 166159
rect 181627 166154 187468 167335
rect 188592 166155 194426 167336
rect 195550 167336 208311 167337
rect 195550 166155 201346 167336
rect 188592 166154 201346 166155
rect 202470 166155 208311 167336
rect 209435 166156 215269 167337
rect 216393 166160 222186 167338
rect 223310 166161 229151 167342
rect 230275 166162 236109 167343
rect 237233 167343 256949 167344
rect 237233 167342 249991 167343
rect 237233 166162 243026 167342
rect 230275 166161 243026 166162
rect 223310 166160 243026 166161
rect 244150 166161 249991 167342
rect 251115 166162 256949 167343
rect 258073 166162 264089 167344
rect 265213 166163 271047 167344
rect 272171 167335 280883 167345
rect 272171 166163 278183 167335
rect 265213 166162 278183 166163
rect 251115 166161 278183 166162
rect 244150 166160 278183 166161
rect 216393 166156 278183 166160
rect 209435 166155 278183 166156
rect 202470 166154 278183 166155
rect 181627 166153 278183 166154
rect 279307 166153 280883 167335
rect 165841 166135 280883 166153
rect 65177 165748 280883 166135
rect 65177 165729 279840 165748
rect 100432 164985 102830 165729
rect 141303 164985 143618 165729
rect 189638 164985 192042 165729
rect 232002 164985 234265 165729
rect 267115 164985 269360 165729
rect 100674 160497 102830 164985
rect 141462 160497 143618 164985
rect 189886 160497 192042 164985
rect 232171 160498 234265 164985
rect 18634 160008 38196 160497
rect 18634 160007 28678 160008
rect 18634 158825 21720 160007
rect 22844 158826 28678 160007
rect 29802 160007 38196 160008
rect 29802 158826 35598 160007
rect 22844 158825 35598 158826
rect 36722 158825 38196 160007
rect 18634 158394 38196 158825
rect 18634 158390 31100 158394
rect 31314 155664 33327 158394
rect 34165 158390 38196 158394
rect 54328 160014 66931 160497
rect 54328 160013 63403 160014
rect 54328 158831 56438 160013
rect 57562 158832 63403 160013
rect 64527 158832 66931 160014
rect 57562 158831 66931 158832
rect 54328 158390 66931 158831
rect 95161 159995 108521 160497
rect 95161 159994 104984 159995
rect 95161 158812 98019 159994
rect 99143 158813 104984 159994
rect 106108 158813 108521 159995
rect 99143 158812 108521 158813
rect 95161 158390 108521 158812
rect 136751 160488 143618 160497
rect 144252 160488 171536 160497
rect 136751 160049 171536 160488
rect 136751 160003 164841 160049
rect 136751 160002 153625 160003
rect 136751 160001 146667 160002
rect 136751 158819 139702 160001
rect 140826 158820 146667 160001
rect 147791 158821 153625 160002
rect 154749 160001 164841 160003
rect 154749 158821 160542 160001
rect 147791 158820 160542 158821
rect 140826 158819 160542 158820
rect 161666 158874 164841 160001
rect 166107 160002 171536 160049
rect 166107 158874 167507 160002
rect 161666 158820 167507 158874
rect 168631 158820 171536 160002
rect 161666 158819 171536 158820
rect 136751 158390 171536 158819
rect 185400 159998 197751 160497
rect 185400 159997 195193 159998
rect 185400 158815 188235 159997
rect 189359 158816 195193 159997
rect 196317 158816 197751 159998
rect 189359 158815 197751 158816
rect 185400 158390 197751 158815
rect 227494 160004 253730 160498
rect 267266 160487 269360 164985
rect 227494 160000 250632 160004
rect 227494 159999 243715 160000
rect 227494 159998 236757 159999
rect 227494 158816 229792 159998
rect 230916 158817 236757 159998
rect 237881 158818 243715 159999
rect 244839 158822 250632 160000
rect 251756 158822 253730 160004
rect 244839 158818 253730 158822
rect 237881 158817 253730 158818
rect 230916 158816 253730 158817
rect 227494 158391 253730 158816
rect 253787 159993 281462 160487
rect 253787 159989 278364 159993
rect 253787 159988 271447 159989
rect 253787 159987 264489 159988
rect 253787 158805 257524 159987
rect 258648 158806 264489 159987
rect 265613 158807 271447 159988
rect 272571 158811 278364 159989
rect 279488 158811 281462 159993
rect 272571 158807 281462 158811
rect 265613 158806 281462 158807
rect 258648 158805 281462 158806
rect 59124 158325 61394 158390
rect 101090 158325 103270 158390
rect 141462 158376 144019 158390
rect 141763 158325 144019 158376
rect 190340 158360 192593 158390
rect 59124 155664 61137 158325
rect 101090 155664 103103 158325
rect 141763 155664 143776 158325
rect 190340 155664 192353 158360
rect 232171 155665 234265 158391
rect 253787 158380 281462 158805
rect 18919 155175 38196 155664
rect 18919 155174 28963 155175
rect 18919 153992 22005 155174
rect 23129 153993 28963 155174
rect 30087 155174 38196 155175
rect 30087 153993 35883 155174
rect 23129 153992 35883 153993
rect 37007 153992 38196 155174
rect 18919 153561 38196 153992
rect 18919 153557 33327 153561
rect 34450 153557 38196 153561
rect 54328 155181 66931 155664
rect 54328 155180 63688 155181
rect 54328 153998 56723 155180
rect 57847 153999 63688 155180
rect 64812 153999 66931 155181
rect 57847 153998 66931 153999
rect 54328 153557 66931 153998
rect 95161 155162 108521 155664
rect 95161 155161 105269 155162
rect 95161 153979 98304 155161
rect 99428 153980 105269 155161
rect 106393 153980 108521 155162
rect 99428 153979 108521 153980
rect 95161 153557 108521 153979
rect 136751 155209 171536 155664
rect 136751 155170 164822 155209
rect 136751 155169 153910 155170
rect 136751 155168 146952 155169
rect 136751 153986 139987 155168
rect 141111 153987 146952 155168
rect 148076 153988 153910 155169
rect 155034 155168 164822 155170
rect 155034 153988 160827 155168
rect 148076 153987 160827 153988
rect 141111 153986 160827 153987
rect 161951 154034 164822 155168
rect 166088 155169 171536 155209
rect 166088 154034 167792 155169
rect 161951 153987 167792 154034
rect 168916 153987 171536 155169
rect 161951 153986 171536 153987
rect 136751 153557 171536 153986
rect 185400 155165 197751 155664
rect 185400 155164 195478 155165
rect 185400 153982 188520 155164
rect 189644 153983 195478 155164
rect 196602 153983 197751 155165
rect 189644 153982 197751 153983
rect 185400 153557 197751 153982
rect 227494 155654 254015 155665
rect 267266 155654 269360 158380
rect 227494 155171 281747 155654
rect 227494 155167 250917 155171
rect 227494 155166 244000 155167
rect 227494 155165 237042 155166
rect 227494 153983 230077 155165
rect 231201 153984 237042 155165
rect 238166 153985 244000 155166
rect 245124 153989 250917 155167
rect 252041 155160 281747 155171
rect 252041 155156 278649 155160
rect 252041 155155 271732 155156
rect 252041 155154 264774 155155
rect 252041 153989 257809 155154
rect 245124 153985 257809 153989
rect 238166 153984 257809 153985
rect 231201 153983 257809 153984
rect 227494 153972 257809 153983
rect 258933 153973 264774 155154
rect 265898 153974 271732 155155
rect 272856 153978 278649 155156
rect 279773 153978 281747 155160
rect 272856 153974 281747 153978
rect 265898 153973 281747 153974
rect 258933 153972 281747 153973
rect 227494 153558 281747 153972
rect 31314 150404 33327 153557
rect 59124 153492 61679 153557
rect 101090 153492 103555 153557
rect 141763 153492 144304 153557
rect 190340 153527 192878 153557
rect 59124 150404 61137 153492
rect 101090 150404 103103 153492
rect 141763 150404 143776 153492
rect 190340 150404 192353 153527
rect 232171 150405 234265 153558
rect 253787 153547 281747 153558
rect 18990 149915 38196 150404
rect 18990 149914 29034 149915
rect 18990 148732 22076 149914
rect 23200 148733 29034 149914
rect 30158 149914 38196 149915
rect 30158 148733 35954 149914
rect 23200 148732 35954 148733
rect 37078 148732 38196 149914
rect 18990 148301 38196 148732
rect 18990 148297 33327 148301
rect 34521 148297 38196 148301
rect 54328 149921 66931 150404
rect 54328 149920 63759 149921
rect 54328 148738 56794 149920
rect 57918 148739 63759 149920
rect 64883 148739 66931 149921
rect 57918 148738 66931 148739
rect 54328 148297 66931 148738
rect 95161 149902 108521 150404
rect 95161 149901 105340 149902
rect 95161 148719 98375 149901
rect 99499 148720 105340 149901
rect 106464 148720 108521 149902
rect 99499 148719 108521 148720
rect 95161 148297 108521 148719
rect 136751 149939 171536 150404
rect 136751 149910 164803 149939
rect 136751 149909 153981 149910
rect 136751 149908 147023 149909
rect 136751 148726 140058 149908
rect 141182 148727 147023 149908
rect 148147 148728 153981 149909
rect 155105 149908 164803 149910
rect 155105 148728 160898 149908
rect 148147 148727 160898 148728
rect 141182 148726 160898 148727
rect 162022 148764 164803 149908
rect 166069 149909 171536 149939
rect 166069 148764 167863 149909
rect 162022 148727 167863 148764
rect 168987 148727 171536 149909
rect 162022 148726 171536 148727
rect 136751 148297 171536 148726
rect 185400 149905 197751 150404
rect 185400 149904 195549 149905
rect 185400 148722 188591 149904
rect 189715 148723 195549 149904
rect 196673 148723 197751 149905
rect 189715 148722 197751 148723
rect 185400 148297 197751 148722
rect 227494 150394 254086 150405
rect 267266 150394 269360 153547
rect 227494 149911 281818 150394
rect 227494 149907 250988 149911
rect 227494 149906 244071 149907
rect 227494 149905 237113 149906
rect 227494 148723 230148 149905
rect 231272 148724 237113 149905
rect 238237 148725 244071 149906
rect 245195 148729 250988 149907
rect 252112 149900 281818 149911
rect 252112 149896 278720 149900
rect 252112 149895 271803 149896
rect 252112 149894 264845 149895
rect 252112 148729 257880 149894
rect 245195 148725 257880 148729
rect 238237 148724 257880 148725
rect 231272 148723 257880 148724
rect 227494 148712 257880 148723
rect 259004 148713 264845 149894
rect 265969 148714 271803 149895
rect 272927 148718 278720 149896
rect 279844 148718 281818 149900
rect 272927 148714 281818 148718
rect 265969 148713 281818 148714
rect 259004 148712 281818 148713
rect 227494 148298 281818 148712
rect 31314 144930 33327 148297
rect 59124 148232 61750 148297
rect 101090 148232 103626 148297
rect 141763 148232 144375 148297
rect 190340 148267 192949 148297
rect 253787 148287 281818 148298
rect 59124 144930 61137 148232
rect 101090 144930 103103 148232
rect 141763 144930 143776 148232
rect 190340 144930 192353 148267
rect 18919 144441 38196 144930
rect 18919 144440 28963 144441
rect 18919 143258 22005 144440
rect 23129 143259 28963 144440
rect 30087 144440 38196 144441
rect 30087 143259 35883 144440
rect 23129 143258 35883 143259
rect 37007 143258 38196 144440
rect 18919 142827 38196 143258
rect 18919 142823 33327 142827
rect 34450 142823 38196 142827
rect 54328 144447 66931 144930
rect 54328 144446 63688 144447
rect 54328 143264 56723 144446
rect 57847 143265 63688 144446
rect 64812 143265 66931 144447
rect 57847 143264 66931 143265
rect 54328 142823 66931 143264
rect 95161 144428 108521 144930
rect 95161 144427 105269 144428
rect 95161 143245 98304 144427
rect 99428 143246 105269 144427
rect 106393 143246 108521 144428
rect 99428 143245 108521 143246
rect 95161 142823 108521 143245
rect 136751 144436 171536 144930
rect 136751 144435 153910 144436
rect 136751 144434 146952 144435
rect 136751 143252 139987 144434
rect 141111 143253 146952 144434
rect 148076 143254 153910 144435
rect 155034 144435 171536 144436
rect 155034 144434 167792 144435
rect 155034 143254 160827 144434
rect 148076 143253 160827 143254
rect 141111 143252 160827 143253
rect 161951 144387 167792 144434
rect 161951 143252 164785 144387
rect 136751 143212 164785 143252
rect 166051 143253 167792 144387
rect 168916 143253 171536 144435
rect 166051 143212 171536 143253
rect 136751 142823 171536 143212
rect 185400 144431 197751 144930
rect 185400 144430 195478 144431
rect 185400 143248 188520 144430
rect 189644 143249 195478 144430
rect 196602 143249 197751 144431
rect 189644 143248 197751 143249
rect 185400 142823 197751 143248
rect 31314 138818 33327 142823
rect 59124 142758 61679 142823
rect 101090 142758 103555 142823
rect 141763 142758 144304 142823
rect 190340 142793 192878 142823
rect 59124 138818 61137 142758
rect 101090 138818 103103 142758
rect 141763 138818 143776 142758
rect 190340 138818 192353 142793
rect 19061 138329 38196 138818
rect 19061 138328 29105 138329
rect 19061 137146 22147 138328
rect 23271 137147 29105 138328
rect 30229 138328 38196 138329
rect 30229 137147 36025 138328
rect 23271 137146 36025 137147
rect 37149 137146 38196 138328
rect 19061 136715 38196 137146
rect 19061 136711 33327 136715
rect 34592 136711 38196 136715
rect 54328 138335 66931 138818
rect 54328 138334 63830 138335
rect 54328 137152 56865 138334
rect 57989 137153 63830 138334
rect 64954 137153 66931 138335
rect 57989 137152 66931 137153
rect 54328 136711 66931 137152
rect 95161 138316 108521 138818
rect 95161 138315 105411 138316
rect 95161 137133 98446 138315
rect 99570 137134 105411 138315
rect 106535 137134 108521 138316
rect 99570 137133 108521 137134
rect 95161 136711 108521 137133
rect 136751 138324 171536 138818
rect 136751 138323 154052 138324
rect 136751 138322 147094 138323
rect 136751 137140 140129 138322
rect 141253 137141 147094 138322
rect 148218 137142 154052 138323
rect 155176 138323 171536 138324
rect 155176 138322 167934 138323
rect 155176 137142 160969 138322
rect 148218 137141 160969 137142
rect 141253 137140 160969 137141
rect 162093 138197 167934 138322
rect 162093 137140 164785 138197
rect 136751 137022 164785 137140
rect 166051 137141 167934 138197
rect 169058 137141 171536 138323
rect 166051 137022 171536 137141
rect 136751 136711 171536 137022
rect 185400 138319 197751 138818
rect 185400 138318 195620 138319
rect 185400 137136 188662 138318
rect 189786 137137 195620 138318
rect 196744 137137 197751 138319
rect 189786 137136 197751 137137
rect 185400 136711 197751 137136
rect 31314 130944 33327 136711
rect 59124 136646 61821 136711
rect 101090 136646 103697 136711
rect 141763 136646 144446 136711
rect 190340 136681 193020 136711
rect 59124 130944 61137 136646
rect 101090 130944 103103 136646
rect 141763 130944 143776 136646
rect 190340 130944 192353 136681
rect 18851 130462 200168 130944
rect 18851 130461 70578 130462
rect 18851 130460 63620 130461
rect 18851 130456 56655 130460
rect 18851 130455 49738 130456
rect 18851 130454 28895 130455
rect 18851 129272 21937 130454
rect 23061 129273 28895 130454
rect 30019 130454 42780 130455
rect 30019 129273 35815 130454
rect 23061 129272 35815 129273
rect 36939 129273 42780 130454
rect 43904 129274 49738 130455
rect 50862 129278 56655 130456
rect 57779 129279 63620 130460
rect 64744 129280 70578 130461
rect 71702 130461 91418 130462
rect 71702 130460 84460 130461
rect 71702 129280 77495 130460
rect 64744 129279 77495 129280
rect 57779 129278 77495 129279
rect 78619 129279 84460 130460
rect 85584 129280 91418 130461
rect 92542 130450 200168 130462
rect 92542 130449 153842 130450
rect 92542 130448 146884 130449
rect 92542 130444 139919 130448
rect 92542 130443 133002 130444
rect 92542 130442 112159 130443
rect 92542 130441 105201 130442
rect 92542 129280 98236 130441
rect 85584 129279 98236 129280
rect 78619 129278 98236 129279
rect 50862 129274 98236 129278
rect 43904 129273 98236 129274
rect 36939 129272 98236 129273
rect 18851 129259 98236 129272
rect 99360 129260 105201 130441
rect 106325 129261 112159 130442
rect 113283 130442 126044 130443
rect 113283 129261 119079 130442
rect 106325 129260 119079 129261
rect 120203 129261 126044 130442
rect 127168 129262 133002 130443
rect 134126 129266 139919 130444
rect 141043 129267 146884 130448
rect 148008 129268 153842 130449
rect 154966 130449 174682 130450
rect 154966 130448 167724 130449
rect 154966 129268 160759 130448
rect 148008 129267 160759 129268
rect 141043 129266 160759 129267
rect 161883 129267 167724 130448
rect 168848 129268 174682 130449
rect 175806 130445 200168 130450
rect 175806 130444 195410 130445
rect 175806 130443 188452 130444
rect 175806 129268 181487 130443
rect 168848 129267 181487 129268
rect 161883 129266 181487 129267
rect 134126 129262 181487 129266
rect 127168 129261 181487 129262
rect 182611 129262 188452 130443
rect 189576 129263 195410 130444
rect 196534 129263 200168 130445
rect 189576 129262 200168 129263
rect 182611 129261 200168 129262
rect 120203 129260 200168 129261
rect 99360 129259 200168 129260
rect 18851 128841 200168 129259
rect 18851 128837 33327 128841
rect 34382 128837 200168 128841
rect 31314 121523 33327 128837
rect 59124 128772 61611 128837
rect 101090 128772 103487 128837
rect 141763 128772 144236 128837
rect 190340 128807 192810 128837
rect 59124 121523 61137 128772
rect 101090 119628 103103 128772
rect 141763 119628 143776 128772
rect 190340 121685 192353 128807
rect 94909 119126 107765 119628
rect 94909 119125 104718 119126
rect 94909 117943 97753 119125
rect 98877 117944 104718 119125
rect 105842 117944 107765 119126
rect 98877 117943 107765 117944
rect 94909 117521 107765 117943
rect 138012 119134 171454 119628
rect 138012 119133 153359 119134
rect 138012 119132 146401 119133
rect 138012 117950 139436 119132
rect 140560 117951 146401 119132
rect 147525 117952 153359 119133
rect 154483 119133 171454 119134
rect 154483 119132 167241 119133
rect 154483 117952 160276 119132
rect 147525 117951 160276 117952
rect 140560 117950 160276 117951
rect 161400 119093 167241 119132
rect 161400 117950 164793 119093
rect 138012 117918 164793 117950
rect 166059 117951 167241 119093
rect 168365 117951 171454 119133
rect 166059 117918 171454 117951
rect 138012 117521 171454 117918
rect 101090 116639 103103 117521
rect 141763 117070 143776 117521
rect 101105 111676 103004 116639
rect 141854 111676 143753 117070
rect 94909 111174 107765 111676
rect 94909 111173 104923 111174
rect 94909 109991 97958 111173
rect 99082 109992 104923 111173
rect 106047 109992 107765 111174
rect 99082 109991 107765 109992
rect 94909 109569 107765 109991
rect 138012 111182 171454 111676
rect 138012 111181 153564 111182
rect 138012 111180 146606 111181
rect 138012 109998 139641 111180
rect 140765 109999 146606 111180
rect 147730 110000 153564 111181
rect 154688 111181 171454 111182
rect 154688 111180 167446 111181
rect 154688 110000 160481 111180
rect 147730 109999 160481 110000
rect 140765 109998 160481 109999
rect 161605 111166 167446 111180
rect 161605 109998 164902 111166
rect 138012 109991 164902 109998
rect 166168 109999 167446 111166
rect 168570 109999 171454 111181
rect 166168 109991 171454 109999
rect 138012 109569 171454 109991
rect 101105 103450 103004 109569
rect 141854 103450 143753 109569
rect 94909 102948 107765 103450
rect 94909 102947 104923 102948
rect 94909 101765 97958 102947
rect 99082 101766 104923 102947
rect 106047 101766 107765 102948
rect 99082 101765 107765 101766
rect 94909 101343 107765 101765
rect 138012 102964 171454 103450
rect 138012 102956 165003 102964
rect 138012 102955 153564 102956
rect 138012 102954 146606 102955
rect 138012 101772 139641 102954
rect 140765 101773 146606 102954
rect 147730 101774 153564 102955
rect 154688 102954 165003 102956
rect 154688 101774 160481 102954
rect 147730 101773 160481 101774
rect 140765 101772 160481 101773
rect 161605 101789 165003 102954
rect 166269 102955 171454 102964
rect 166269 101789 167446 102955
rect 161605 101773 167446 101789
rect 168570 101773 171454 102955
rect 161605 101772 171454 101773
rect 138012 101343 171454 101772
rect 101105 96046 103004 101343
rect 141854 96046 143753 101343
rect 94909 95544 107765 96046
rect 94909 95543 104718 95544
rect 94909 94361 97753 95543
rect 98877 94362 104718 95543
rect 105842 94362 107765 95544
rect 98877 94361 107765 94362
rect 94909 93939 107765 94361
rect 138012 95552 171454 96046
rect 138012 95551 153359 95552
rect 138012 95550 146401 95551
rect 138012 94368 139436 95550
rect 140560 94369 146401 95550
rect 147525 94370 153359 95551
rect 154483 95551 171454 95552
rect 154483 95550 167241 95551
rect 154483 94370 160276 95550
rect 147525 94369 160276 94370
rect 140560 94368 160276 94369
rect 161400 95465 167241 95550
rect 161400 94368 164966 95465
rect 138012 94290 164966 94368
rect 166232 94369 167241 95465
rect 168365 94369 171454 95551
rect 166232 94290 171454 94369
rect 138012 93939 171454 94290
rect 101105 88916 103004 93939
rect 141854 88916 143753 93939
rect 94454 88422 171454 88916
rect 94454 88421 153085 88422
rect 94454 88420 146127 88421
rect 94454 88416 139162 88420
rect 94454 88415 132245 88416
rect 94454 88414 111402 88415
rect 94454 88413 104444 88414
rect 94454 87231 97479 88413
rect 98603 87232 104444 88413
rect 105568 87233 111402 88414
rect 112526 88414 125287 88415
rect 112526 87233 118322 88414
rect 105568 87232 118322 87233
rect 119446 87233 125287 88414
rect 126411 87234 132245 88415
rect 133369 87238 139162 88416
rect 140286 87239 146127 88420
rect 147251 87240 153085 88421
rect 154209 88421 171454 88422
rect 154209 88420 166967 88421
rect 154209 87240 160002 88420
rect 147251 87239 160002 87240
rect 140286 87238 160002 87239
rect 161126 88379 166967 88420
rect 161126 87238 164947 88379
rect 133369 87234 164947 87238
rect 126411 87233 164947 87234
rect 119446 87232 164947 87233
rect 98603 87231 164947 87232
rect 94454 87204 164947 87231
rect 166213 87239 166967 88379
rect 168091 87239 171454 88421
rect 166213 87204 171454 87239
rect 94454 86809 171454 87204
rect 101105 82503 103004 86809
rect 141854 82503 143753 86809
rect 94454 82009 171454 82503
rect 94454 82008 153193 82009
rect 94454 82007 146235 82008
rect 94454 82003 139270 82007
rect 94454 82002 132353 82003
rect 94454 82001 111510 82002
rect 94454 82000 104552 82001
rect 94454 80818 97587 82000
rect 98711 80819 104552 82000
rect 105676 80820 111510 82001
rect 112634 82001 125395 82002
rect 112634 80820 118430 82001
rect 105676 80819 118430 80820
rect 119554 80820 125395 82001
rect 126519 80821 132353 82002
rect 133477 80825 139270 82003
rect 140394 80826 146235 82007
rect 147359 80827 153193 82008
rect 154317 82008 171454 82009
rect 154317 82007 167075 82008
rect 154317 80827 160110 82007
rect 147359 80826 160110 80827
rect 140394 80825 160110 80826
rect 161234 81977 167075 82007
rect 161234 80825 164910 81977
rect 133477 80821 164910 80825
rect 126519 80820 164910 80821
rect 119554 80819 164910 80820
rect 98711 80818 164910 80819
rect 94454 80802 164910 80818
rect 166176 80826 167075 81977
rect 168199 80826 171454 82008
rect 166176 80802 171454 80826
rect 94454 80396 171454 80802
rect 100767 71584 102857 80396
rect 31059 71323 33699 71555
rect 60920 71323 60994 71584
rect 100767 71323 102870 71584
rect 141638 71323 143728 80396
rect 18234 71274 58830 71323
rect 60920 71274 176227 71323
rect 18234 70841 176227 71274
rect 18234 70840 69795 70841
rect 18234 70839 62837 70840
rect 18234 70835 55872 70839
rect 18234 70834 48955 70835
rect 18234 70833 28112 70834
rect 18234 69651 21154 70833
rect 22278 69652 28112 70833
rect 29236 70833 41997 70834
rect 29236 69652 35032 70833
rect 22278 69651 35032 69652
rect 36156 69652 41997 70833
rect 43121 69653 48955 70834
rect 50079 69657 55872 70835
rect 56996 69658 62837 70839
rect 63961 69659 69795 70840
rect 70919 70840 90635 70841
rect 70919 70839 83677 70840
rect 70919 69659 76712 70839
rect 63961 69658 76712 69659
rect 56996 69657 76712 69658
rect 77836 69658 83677 70839
rect 84801 69659 90635 70840
rect 91759 70829 176227 70841
rect 91759 70828 153059 70829
rect 91759 70827 146101 70828
rect 91759 70823 139136 70827
rect 91759 70822 132219 70823
rect 91759 70821 111376 70822
rect 91759 70820 104418 70821
rect 91759 69659 97453 70820
rect 84801 69658 97453 69659
rect 77836 69657 97453 69658
rect 50079 69653 97453 69657
rect 43121 69652 97453 69653
rect 36156 69651 97453 69652
rect 18234 69638 97453 69651
rect 98577 69639 104418 70820
rect 105542 69640 111376 70821
rect 112500 70821 125261 70822
rect 112500 69640 118296 70821
rect 105542 69639 118296 69640
rect 119420 69640 125261 70821
rect 126385 69641 132219 70822
rect 133343 69645 139136 70823
rect 140260 69646 146101 70827
rect 147225 69647 153059 70828
rect 154183 70828 173899 70829
rect 154183 70827 166941 70828
rect 154183 69647 159976 70827
rect 147225 69646 159976 69647
rect 140260 69645 159976 69646
rect 161100 70727 166941 70827
rect 161100 69645 164892 70727
rect 133343 69641 164892 69645
rect 126385 69640 164892 69641
rect 119420 69639 164892 69640
rect 98577 69638 164892 69639
rect 18234 69552 164892 69638
rect 166158 69646 166941 70727
rect 168065 69647 173899 70828
rect 175023 69647 176227 70829
rect 168065 69646 176227 69647
rect 166158 69552 176227 69646
rect 18234 69216 176227 69552
rect 31059 65083 33699 69216
rect 58830 65083 61404 69216
rect 100767 65083 102857 69216
rect 141638 65083 143728 69216
rect 18199 64732 176227 65083
rect 18199 64601 164818 64732
rect 18199 64600 69760 64601
rect 18199 64599 62802 64600
rect 18199 64595 55837 64599
rect 18199 64594 48920 64595
rect 18199 64593 28077 64594
rect 18199 63411 21119 64593
rect 22243 63412 28077 64593
rect 29201 64593 41962 64594
rect 29201 63412 34997 64593
rect 22243 63411 34997 63412
rect 36121 63412 41962 64593
rect 43086 63413 48920 64594
rect 50044 63417 55837 64595
rect 56961 63418 62802 64599
rect 63926 63419 69760 64600
rect 70884 64600 90600 64601
rect 70884 64599 83642 64600
rect 70884 63419 76677 64599
rect 63926 63418 76677 63419
rect 56961 63417 76677 63418
rect 77801 63418 83642 64599
rect 84766 63419 90600 64600
rect 91724 64589 164818 64601
rect 91724 64588 153024 64589
rect 91724 64587 146066 64588
rect 91724 64583 139101 64587
rect 91724 64582 132184 64583
rect 91724 64581 111341 64582
rect 91724 64580 104383 64581
rect 91724 63419 97418 64580
rect 84766 63418 97418 63419
rect 77801 63417 97418 63418
rect 50044 63413 97418 63417
rect 43086 63412 97418 63413
rect 36121 63411 97418 63412
rect 18199 63398 97418 63411
rect 98542 63399 104383 64580
rect 105507 63400 111341 64581
rect 112465 64581 125226 64582
rect 112465 63400 118261 64581
rect 105507 63399 118261 63400
rect 119385 63400 125226 64581
rect 126350 63401 132184 64582
rect 133308 63405 139101 64583
rect 140225 63406 146066 64587
rect 147190 63407 153024 64588
rect 154148 64587 164818 64589
rect 154148 63407 159941 64587
rect 147190 63406 159941 63407
rect 140225 63405 159941 63406
rect 161065 63557 164818 64587
rect 166084 64589 176227 64732
rect 166084 64588 173864 64589
rect 166084 63557 166906 64588
rect 161065 63406 166906 63557
rect 168030 63407 173864 64588
rect 174988 63407 176227 64589
rect 168030 63406 176227 63407
rect 161065 63405 176227 63406
rect 133308 63401 176227 63405
rect 126350 63400 176227 63401
rect 119385 63399 176227 63400
rect 98542 63398 176227 63399
rect 18199 62976 176227 63398
rect 31059 59366 33699 62976
rect 58830 59366 61404 62976
rect 100767 59366 102857 62976
rect 141638 59366 143728 62976
rect 18164 58904 176227 59366
rect 18164 58884 164855 58904
rect 18164 58883 69725 58884
rect 18164 58882 62767 58883
rect 18164 58878 55802 58882
rect 18164 58877 48885 58878
rect 18164 58876 28042 58877
rect 18164 57694 21084 58876
rect 22208 57695 28042 58876
rect 29166 58876 41927 58877
rect 29166 57695 34962 58876
rect 22208 57694 34962 57695
rect 36086 57695 41927 58876
rect 43051 57696 48885 58877
rect 50009 57700 55802 58878
rect 56926 57701 62767 58882
rect 63891 57702 69725 58883
rect 70849 58883 90565 58884
rect 70849 58882 83607 58883
rect 70849 57702 76642 58882
rect 63891 57701 76642 57702
rect 56926 57700 76642 57701
rect 77766 57701 83607 58882
rect 84731 57702 90565 58883
rect 91689 58872 164855 58884
rect 91689 58871 152989 58872
rect 91689 58870 146031 58871
rect 91689 58866 139066 58870
rect 91689 58865 132149 58866
rect 91689 58864 111306 58865
rect 91689 58863 104348 58864
rect 91689 57702 97383 58863
rect 84731 57701 97383 57702
rect 77766 57700 97383 57701
rect 50009 57696 97383 57700
rect 43051 57695 97383 57696
rect 36086 57694 97383 57695
rect 18164 57681 97383 57694
rect 98507 57682 104348 58863
rect 105472 57683 111306 58864
rect 112430 58864 125191 58865
rect 112430 57683 118226 58864
rect 105472 57682 118226 57683
rect 119350 57683 125191 58864
rect 126315 57684 132149 58865
rect 133273 57688 139066 58866
rect 140190 57689 146031 58870
rect 147155 57690 152989 58871
rect 154113 58870 164855 58872
rect 154113 57690 159906 58870
rect 147155 57689 159906 57690
rect 140190 57688 159906 57689
rect 161030 57729 164855 58870
rect 166121 58872 176227 58904
rect 166121 58871 173829 58872
rect 166121 57729 166871 58871
rect 161030 57689 166871 57729
rect 167995 57690 173829 58871
rect 174953 57690 176227 58872
rect 167995 57689 176227 57690
rect 161030 57688 176227 57689
rect 133273 57684 176227 57688
rect 126315 57683 176227 57684
rect 119350 57682 176227 57683
rect 98507 57681 176227 57682
rect 18164 57259 176227 57681
rect 31059 53161 33699 57259
rect 58830 53161 61404 57259
rect 100767 53161 102857 57259
rect 141638 53422 143728 57259
rect 141581 53161 143728 53422
rect 18095 52817 176227 53161
rect 18095 52679 164929 52817
rect 18095 52678 69656 52679
rect 18095 52677 62698 52678
rect 18095 52673 55733 52677
rect 18095 52672 48816 52673
rect 18095 52671 27973 52672
rect 18095 51489 21015 52671
rect 22139 51490 27973 52671
rect 29097 52671 41858 52672
rect 29097 51490 34893 52671
rect 22139 51489 34893 51490
rect 36017 51490 41858 52671
rect 42982 51491 48816 52672
rect 49940 51495 55733 52673
rect 56857 51496 62698 52677
rect 63822 51497 69656 52678
rect 70780 52678 90496 52679
rect 70780 52677 83538 52678
rect 70780 51497 76573 52677
rect 63822 51496 76573 51497
rect 56857 51495 76573 51496
rect 77697 51496 83538 52677
rect 84662 51497 90496 52678
rect 91620 52667 164929 52679
rect 91620 52666 152920 52667
rect 91620 52665 145962 52666
rect 91620 52661 138997 52665
rect 91620 52660 132080 52661
rect 91620 52659 111237 52660
rect 91620 52658 104279 52659
rect 91620 51497 97314 52658
rect 84662 51496 97314 51497
rect 77697 51495 97314 51496
rect 49940 51491 97314 51495
rect 42982 51490 97314 51491
rect 36017 51489 97314 51490
rect 18095 51476 97314 51489
rect 98438 51477 104279 52658
rect 105403 51478 111237 52659
rect 112361 52659 125122 52660
rect 112361 51478 118157 52659
rect 105403 51477 118157 51478
rect 119281 51478 125122 52659
rect 126246 51479 132080 52660
rect 133204 51483 138997 52661
rect 140121 51484 145962 52665
rect 147086 51485 152920 52666
rect 154044 52665 164929 52667
rect 154044 51485 159837 52665
rect 147086 51484 159837 51485
rect 140121 51483 159837 51484
rect 160961 51642 164929 52665
rect 166195 52667 176227 52817
rect 166195 52666 173760 52667
rect 166195 51642 166802 52666
rect 160961 51484 166802 51642
rect 167926 51485 173760 52666
rect 174884 51485 176227 52667
rect 167926 51484 176227 51485
rect 160961 51483 176227 51484
rect 133204 51479 176227 51483
rect 126246 51478 176227 51479
rect 119281 51477 176227 51478
rect 98438 51476 176227 51477
rect 18095 51054 176227 51476
rect 100312 47394 102598 51054
rect 141218 45303 143504 51054
rect 135410 44959 176227 45303
rect 135410 44809 164641 44959
rect 135410 44808 152632 44809
rect 135410 44807 145674 44808
rect 135410 43625 138709 44807
rect 139833 43626 145674 44807
rect 146798 43627 152632 44808
rect 153756 44807 164641 44809
rect 153756 43627 159549 44807
rect 146798 43626 159549 43627
rect 139833 43625 159549 43626
rect 160673 43784 164641 44807
rect 165907 44809 176227 44959
rect 165907 44808 173472 44809
rect 165907 43784 166514 44808
rect 160673 43626 166514 43784
rect 167638 43627 173472 44808
rect 174596 43627 176227 44809
rect 167638 43626 176227 43627
rect 160673 43625 176227 43626
rect 135410 43196 176227 43625
rect 141218 39009 143504 43196
rect 135410 38665 176227 39009
rect 135410 38515 164641 38665
rect 135410 38514 152632 38515
rect 135410 38513 145674 38514
rect 135410 37331 138709 38513
rect 139833 37332 145674 38513
rect 146798 37333 152632 38514
rect 153756 38513 164641 38515
rect 153756 37333 159549 38513
rect 146798 37332 159549 37333
rect 139833 37331 159549 37332
rect 160673 37490 164641 38513
rect 165907 38515 176227 38665
rect 165907 38514 173472 38515
rect 165907 37490 166514 38514
rect 160673 37332 166514 37490
rect 167638 37333 173472 38514
rect 174596 37333 176227 38515
rect 167638 37332 176227 37333
rect 160673 37331 176227 37332
rect 135410 36902 176227 37331
rect 141218 32715 143504 36902
rect 135410 32371 176227 32715
rect 135410 32221 164641 32371
rect 135410 32220 152632 32221
rect 135410 32219 145674 32220
rect 135410 31037 138709 32219
rect 139833 31038 145674 32219
rect 146798 31039 152632 32220
rect 153756 32219 164641 32221
rect 153756 31039 159549 32219
rect 146798 31038 159549 31039
rect 139833 31037 159549 31038
rect 160673 31196 164641 32219
rect 165907 32221 176227 32371
rect 165907 32220 173472 32221
rect 165907 31196 166514 32220
rect 160673 31038 166514 31196
rect 167638 31039 173472 32220
rect 174596 31039 176227 32221
rect 167638 31038 176227 31039
rect 160673 31037 176227 31038
rect 135410 30608 176227 31037
rect 141218 23755 143504 30608
<< viali >>
rect 164500 338774 165766 339949
rect 164481 331688 165747 332863
rect 164500 325316 165766 326491
rect 164481 318230 165747 319405
rect 164506 311055 165772 312230
rect 164487 303969 165753 305144
rect 164595 294696 165861 295871
rect 164576 287610 165842 288785
rect 164539 281208 165805 282383
rect 164646 272288 165912 273463
rect 164627 265202 165893 266377
rect 164590 258800 165856 259975
rect 164677 248034 165943 249209
rect 164658 240948 165924 242123
rect 164621 234546 165887 235721
rect 164801 227768 166067 228943
rect 164781 221906 166047 223081
rect 164821 209843 166087 211018
rect 164802 202757 166068 203932
rect 164765 196355 166031 197530
rect 164808 191950 166074 193125
rect 164789 184864 166055 186039
rect 164752 178462 166018 179637
rect 164612 172537 165878 173712
rect 164575 166135 165841 167310
rect 164841 158874 166107 160049
rect 164822 154034 166088 155209
rect 164803 148764 166069 149939
rect 164785 143212 166051 144387
rect 164785 137022 166051 138197
rect 164793 117918 166059 119093
rect 164902 109991 166168 111166
rect 165003 101789 166269 102964
rect 164966 94290 166232 95465
rect 164947 87204 166213 88379
rect 164910 80802 166176 81977
rect 164892 69552 166158 70727
rect 164818 63557 166084 64732
rect 164855 57729 166121 58904
rect 164929 51642 166195 52817
rect 164641 43784 165907 44959
rect 164641 37490 165907 38665
rect 164641 31196 165907 32371
<< metal1 >>
rect 164427 339949 165848 340032
rect 164427 338774 164500 339949
rect 165766 338774 165848 339949
rect 164427 338683 165848 338774
rect 164408 332863 165829 332946
rect 164408 331688 164481 332863
rect 165747 331688 165829 332863
rect 164408 331597 165829 331688
rect 164427 326491 165848 326574
rect 164427 325316 164500 326491
rect 165766 325316 165848 326491
rect 164427 325225 165848 325316
rect 164408 319405 165829 319488
rect 164408 318230 164481 319405
rect 165747 318230 165829 319405
rect 164408 318139 165829 318230
rect 164433 312230 165854 312313
rect 164433 311055 164506 312230
rect 165772 311055 165854 312230
rect 164433 310964 165854 311055
rect 164414 305144 165835 305227
rect 164414 303969 164487 305144
rect 165753 303969 165835 305144
rect 164414 303878 165835 303969
rect 164522 295871 165943 295954
rect 164522 294696 164595 295871
rect 165861 294696 165943 295871
rect 164522 294605 165943 294696
rect 164503 288785 165924 288868
rect 164503 287610 164576 288785
rect 165842 287610 165924 288785
rect 164503 287519 165924 287610
rect 164466 282383 165887 282466
rect 164466 281208 164539 282383
rect 165805 281208 165887 282383
rect 164466 281117 165887 281208
rect 164573 273463 165994 273546
rect 164573 272288 164646 273463
rect 165912 272288 165994 273463
rect 164573 272197 165994 272288
rect 164554 266377 165975 266460
rect 164554 265202 164627 266377
rect 165893 265202 165975 266377
rect 164554 265111 165975 265202
rect 164517 259975 165938 260058
rect 164517 258800 164590 259975
rect 165856 258800 165938 259975
rect 164517 258709 165938 258800
rect 164604 249209 166025 249292
rect 164604 248034 164677 249209
rect 165943 248034 166025 249209
rect 164604 247943 166025 248034
rect 164585 242123 166006 242206
rect 164585 240948 164658 242123
rect 165924 240948 166006 242123
rect 164585 240857 166006 240948
rect 164548 235721 165969 235804
rect 164548 234546 164621 235721
rect 165887 234546 165969 235721
rect 164548 234455 165969 234546
rect 164728 228943 166149 229026
rect 164728 227768 164801 228943
rect 166067 227768 166149 228943
rect 164728 227677 166149 227768
rect 164708 223081 166129 223164
rect 164708 221906 164781 223081
rect 166047 221906 166129 223081
rect 164708 221815 166129 221906
rect 164748 211018 166169 211101
rect 164748 209843 164821 211018
rect 166087 209843 166169 211018
rect 164748 209752 166169 209843
rect 164729 203932 166150 204015
rect 164729 202757 164802 203932
rect 166068 202757 166150 203932
rect 164729 202666 166150 202757
rect 164692 197530 166113 197613
rect 164692 196355 164765 197530
rect 166031 196355 166113 197530
rect 164692 196264 166113 196355
rect 164735 193125 166156 193208
rect 164735 191950 164808 193125
rect 166074 191950 166156 193125
rect 164735 191859 166156 191950
rect 164716 186039 166137 186122
rect 164716 184864 164789 186039
rect 166055 184864 166137 186039
rect 164716 184773 166137 184864
rect 164679 179637 166100 179720
rect 164679 178462 164752 179637
rect 166018 178462 166100 179637
rect 164679 178371 166100 178462
rect 164539 173712 165960 173795
rect 164539 172537 164612 173712
rect 165878 172537 165960 173712
rect 164539 172446 165960 172537
rect 164502 167310 165923 167393
rect 164502 166135 164575 167310
rect 165841 166135 165923 167310
rect 164502 166044 165923 166135
rect 164768 160049 166189 160132
rect 164768 158874 164841 160049
rect 166107 158874 166189 160049
rect 164768 158783 166189 158874
rect 164749 155209 166170 155292
rect 164749 154034 164822 155209
rect 166088 154034 166170 155209
rect 164749 153943 166170 154034
rect 164730 149939 166151 150022
rect 164730 148764 164803 149939
rect 166069 148764 166151 149939
rect 164730 148673 166151 148764
rect 164712 144387 166133 144470
rect 164712 143212 164785 144387
rect 166051 143212 166133 144387
rect 164712 143121 166133 143212
rect 164712 138197 166133 138280
rect 164712 137022 164785 138197
rect 166051 137022 166133 138197
rect 164712 136931 166133 137022
rect 164720 119093 166141 119176
rect 164720 117918 164793 119093
rect 166059 117918 166141 119093
rect 164720 117827 166141 117918
rect 164829 111166 166250 111249
rect 164829 109991 164902 111166
rect 166168 109991 166250 111166
rect 164829 109900 166250 109991
rect 164930 102964 166351 103047
rect 164930 101789 165003 102964
rect 166269 101789 166351 102964
rect 164930 101698 166351 101789
rect 164893 95465 166314 95548
rect 164893 94290 164966 95465
rect 166232 94290 166314 95465
rect 164893 94199 166314 94290
rect 164874 88379 166295 88462
rect 164874 87204 164947 88379
rect 166213 87204 166295 88379
rect 164874 87113 166295 87204
rect 164837 81977 166258 82060
rect 164837 80802 164910 81977
rect 166176 80802 166258 81977
rect 164837 80711 166258 80802
rect 164819 70727 166240 70810
rect 164819 69552 164892 70727
rect 166158 69552 166240 70727
rect 164819 69461 166240 69552
rect 164745 64732 166166 64815
rect 164745 63557 164818 64732
rect 166084 63557 166166 64732
rect 164745 63466 166166 63557
rect 164782 58904 166203 58987
rect 164782 57729 164855 58904
rect 166121 57729 166203 58904
rect 164782 57638 166203 57729
rect 164856 52817 166277 52900
rect 164856 51642 164929 52817
rect 166195 51642 166277 52817
rect 164856 51551 166277 51642
rect 164568 44959 165989 45042
rect 164568 43784 164641 44959
rect 165907 43784 165989 44959
rect 164568 43693 165989 43784
rect 164568 38665 165989 38748
rect 164568 37490 164641 38665
rect 165907 37490 165989 38665
rect 164568 37399 165989 37490
rect 164568 32371 165989 32454
rect 164568 31196 164641 32371
rect 165907 31196 165989 32371
rect 164568 31105 165989 31196
<< via1 >>
rect 164500 338774 165766 339949
rect 164481 331688 165747 332863
rect 164500 325316 165766 326491
rect 164481 318230 165747 319405
rect 164506 311055 165772 312230
rect 164487 303969 165753 305144
rect 164595 294696 165861 295871
rect 164576 287610 165842 288785
rect 164539 281208 165805 282383
rect 164646 272288 165912 273463
rect 164627 265202 165893 266377
rect 164590 258800 165856 259975
rect 164677 248034 165943 249209
rect 164658 240948 165924 242123
rect 164621 234546 165887 235721
rect 164801 227768 166067 228943
rect 164781 221906 166047 223081
rect 164821 209843 166087 211018
rect 164802 202757 166068 203932
rect 164765 196355 166031 197530
rect 164808 191950 166074 193125
rect 164789 184864 166055 186039
rect 164752 178462 166018 179637
rect 164612 172537 165878 173712
rect 164575 166135 165841 167310
rect 164841 158874 166107 160049
rect 164822 154034 166088 155209
rect 164803 148764 166069 149939
rect 164785 143212 166051 144387
rect 164785 137022 166051 138197
rect 164793 117918 166059 119093
rect 164902 109991 166168 111166
rect 165003 101789 166269 102964
rect 164966 94290 166232 95465
rect 164947 87204 166213 88379
rect 164910 80802 166176 81977
rect 164892 69552 166158 70727
rect 164818 63557 166084 64732
rect 164855 57729 166121 58904
rect 164929 51642 166195 52817
rect 164641 43784 165907 44959
rect 164641 37490 165907 38665
rect 164641 31196 165907 32371
<< metal2 >>
rect 164427 339949 165848 340032
rect 164427 338774 164500 339949
rect 165766 338774 165848 339949
rect 164427 338683 165848 338774
rect 164408 332863 165829 332946
rect 164408 331688 164481 332863
rect 165747 331688 165829 332863
rect 164408 331597 165829 331688
rect 164427 326491 165848 326574
rect 164427 325316 164500 326491
rect 165766 325316 165848 326491
rect 164427 325225 165848 325316
rect 164408 319405 165829 319488
rect 164408 318230 164481 319405
rect 165747 318230 165829 319405
rect 164408 318139 165829 318230
rect 164433 312230 165854 312313
rect 164433 311055 164506 312230
rect 165772 311055 165854 312230
rect 164433 310964 165854 311055
rect 164414 305144 165835 305227
rect 164414 303969 164487 305144
rect 165753 303969 165835 305144
rect 164414 303878 165835 303969
rect 164522 295871 165943 295954
rect 164522 294696 164595 295871
rect 165861 294696 165943 295871
rect 164522 294605 165943 294696
rect 164503 288785 165924 288868
rect 164503 287610 164576 288785
rect 165842 287610 165924 288785
rect 164503 287519 165924 287610
rect 164466 282383 165887 282466
rect 164466 281208 164539 282383
rect 165805 281208 165887 282383
rect 164466 281117 165887 281208
rect 164573 273463 165994 273546
rect 164573 272288 164646 273463
rect 165912 272288 165994 273463
rect 164573 272197 165994 272288
rect 164554 266377 165975 266460
rect 164554 265202 164627 266377
rect 165893 265202 165975 266377
rect 164554 265111 165975 265202
rect 164517 259975 165938 260058
rect 164517 258800 164590 259975
rect 165856 258800 165938 259975
rect 164517 258709 165938 258800
rect 164604 249209 166025 249292
rect 164604 248034 164677 249209
rect 165943 248034 166025 249209
rect 164604 247943 166025 248034
rect 164585 242123 166006 242206
rect 164585 240948 164658 242123
rect 165924 240948 166006 242123
rect 164585 240857 166006 240948
rect 164548 235721 165969 235804
rect 164548 234546 164621 235721
rect 165887 234546 165969 235721
rect 164548 234455 165969 234546
rect 164728 228943 166149 229026
rect 164728 227768 164801 228943
rect 166067 227768 166149 228943
rect 164728 227677 166149 227768
rect 164708 223081 166129 223164
rect 164708 221906 164781 223081
rect 166047 221906 166129 223081
rect 164708 221815 166129 221906
rect 164748 211018 166169 211101
rect 164748 209843 164821 211018
rect 166087 209843 166169 211018
rect 164748 209752 166169 209843
rect 164729 203932 166150 204015
rect 164729 202757 164802 203932
rect 166068 202757 166150 203932
rect 164729 202666 166150 202757
rect 164692 197530 166113 197613
rect 164692 196355 164765 197530
rect 166031 196355 166113 197530
rect 164692 196264 166113 196355
rect 164735 193125 166156 193208
rect 164735 191950 164808 193125
rect 166074 191950 166156 193125
rect 164735 191859 166156 191950
rect 164716 186039 166137 186122
rect 164716 184864 164789 186039
rect 166055 184864 166137 186039
rect 164716 184773 166137 184864
rect 164679 179637 166100 179720
rect 164679 178462 164752 179637
rect 166018 178462 166100 179637
rect 164679 178371 166100 178462
rect 164539 173712 165960 173795
rect 164539 172537 164612 173712
rect 165878 172537 165960 173712
rect 164539 172446 165960 172537
rect 164502 167310 165923 167393
rect 164502 166135 164575 167310
rect 165841 166135 165923 167310
rect 164502 166044 165923 166135
rect 164768 160049 166189 160132
rect 164768 158874 164841 160049
rect 166107 158874 166189 160049
rect 164768 158783 166189 158874
rect 164749 155209 166170 155292
rect 164749 154034 164822 155209
rect 166088 154034 166170 155209
rect 164749 153943 166170 154034
rect 164730 149939 166151 150022
rect 164730 148764 164803 149939
rect 166069 148764 166151 149939
rect 164730 148673 166151 148764
rect 164712 144387 166133 144470
rect 164712 143212 164785 144387
rect 166051 143212 166133 144387
rect 164712 143121 166133 143212
rect 164712 138197 166133 138280
rect 164712 137022 164785 138197
rect 166051 137022 166133 138197
rect 164712 136931 166133 137022
rect 164720 119093 166141 119176
rect 164720 117918 164793 119093
rect 166059 117918 166141 119093
rect 164720 117827 166141 117918
rect 164829 111166 166250 111249
rect 164829 109991 164902 111166
rect 166168 109991 166250 111166
rect 164829 109900 166250 109991
rect 164930 102964 166351 103047
rect 164930 101789 165003 102964
rect 166269 101789 166351 102964
rect 164930 101698 166351 101789
rect 164893 95465 166314 95548
rect 164893 94290 164966 95465
rect 166232 94290 166314 95465
rect 164893 94199 166314 94290
rect 164874 88379 166295 88462
rect 164874 87204 164947 88379
rect 166213 87204 166295 88379
rect 164874 87113 166295 87204
rect 164837 81977 166258 82060
rect 164837 80802 164910 81977
rect 166176 80802 166258 81977
rect 164837 80711 166258 80802
rect 164819 70727 166240 70810
rect 164819 69552 164892 70727
rect 166158 69552 166240 70727
rect 164819 69461 166240 69552
rect 164745 64732 166166 64815
rect 164745 63557 164818 64732
rect 166084 63557 166166 64732
rect 164745 63466 166166 63557
rect 164782 58904 166203 58987
rect 164782 57729 164855 58904
rect 166121 57729 166203 58904
rect 164782 57638 166203 57729
rect 164856 52817 166277 52900
rect 164856 51642 164929 52817
rect 166195 51642 166277 52817
rect 164856 51551 166277 51642
rect 164568 44959 165989 45042
rect 164568 43784 164641 44959
rect 165907 43784 165989 44959
rect 164568 43693 165989 43784
rect 164568 38665 165989 38748
rect 164568 37490 164641 38665
rect 165907 37490 165989 38665
rect 164568 37399 165989 37490
rect 164568 32371 165989 32454
rect 164568 31196 164641 32371
rect 165907 31196 165989 32371
rect 164568 31105 165989 31196
rect 262 -400 318 240
rect 853 -400 909 240
rect 1444 -400 1500 240
rect 2035 -400 2091 240
rect 2626 -400 2682 240
rect 3217 -400 3273 240
rect 3808 -400 3864 240
rect 4399 -400 4455 240
rect 4990 -400 5046 240
rect 5581 -400 5637 240
rect 6172 -400 6228 240
rect 6763 -400 6819 240
rect 7354 -400 7410 240
rect 7945 -400 8001 240
rect 8536 -400 8592 240
rect 9127 -400 9183 240
rect 9718 -400 9774 240
rect 10309 -400 10365 240
rect 10900 -400 10956 240
rect 11491 -400 11547 240
rect 12082 -400 12138 240
rect 12673 -400 12729 240
rect 13264 -400 13320 240
rect 13855 -400 13911 240
rect 14446 -400 14502 240
rect 15037 -400 15093 240
rect 15628 -400 15684 240
rect 16219 -400 16275 240
rect 16810 -400 16866 240
rect 17401 -400 17457 240
rect 17992 -400 18048 240
rect 18583 -400 18639 240
rect 19174 -400 19230 240
rect 19765 -400 19821 240
rect 20356 -400 20412 240
rect 20947 -400 21003 240
rect 21538 -400 21594 240
rect 22129 -400 22185 240
rect 22720 -400 22776 240
rect 23311 -400 23367 240
rect 23902 -400 23958 240
rect 24493 -400 24549 240
rect 25084 -400 25140 240
rect 25675 -400 25731 240
rect 26266 -400 26322 240
rect 26857 -400 26913 240
rect 27448 -400 27504 240
rect 28039 -400 28095 240
rect 28630 -400 28686 240
rect 29221 -400 29277 240
rect 29812 -400 29868 240
rect 30403 -400 30459 240
rect 30994 -400 31050 240
rect 31585 -400 31641 240
rect 32176 -400 32232 240
rect 32767 -400 32823 240
rect 33358 -400 33414 240
rect 33949 -400 34005 240
rect 34540 -400 34596 240
rect 35131 -400 35187 240
rect 35722 -400 35778 240
rect 36313 -400 36369 240
rect 36904 -400 36960 240
rect 37495 -400 37551 240
rect 38086 -400 38142 240
rect 38677 -400 38733 240
rect 39268 -400 39324 240
rect 39859 -400 39915 240
rect 40450 -400 40506 240
rect 41041 -400 41097 240
rect 41632 -400 41688 240
rect 42223 -400 42279 240
rect 42814 -400 42870 240
rect 43405 -400 43461 240
rect 43996 -400 44052 240
rect 44587 -400 44643 240
rect 45178 -400 45234 240
rect 45769 -400 45825 240
rect 46360 -400 46416 240
rect 46951 -400 47007 240
rect 47542 -400 47598 240
rect 48133 -400 48189 240
rect 48724 -400 48780 240
rect 49315 -400 49371 240
rect 49906 -400 49962 240
rect 50497 -400 50553 240
rect 51088 -400 51144 240
rect 51679 -400 51735 240
rect 52270 -400 52326 240
rect 52861 -400 52917 240
rect 53452 -400 53508 240
rect 54043 -400 54099 240
rect 54634 -400 54690 240
rect 55225 -400 55281 240
rect 55816 -400 55872 240
rect 56407 -400 56463 240
rect 56998 -400 57054 240
rect 57589 -400 57645 240
rect 58180 -400 58236 240
rect 58771 -400 58827 240
rect 59362 -400 59418 240
rect 59953 -400 60009 240
rect 60544 -400 60600 240
rect 61135 -400 61191 240
rect 61726 -400 61782 240
rect 62317 -400 62373 240
rect 62908 -400 62964 240
rect 63499 -400 63555 240
rect 64090 -400 64146 240
rect 64681 -400 64737 240
rect 65272 -400 65328 240
rect 65863 -400 65919 240
rect 66454 -400 66510 240
rect 67045 -400 67101 240
rect 67636 -400 67692 240
rect 68227 -400 68283 240
rect 68818 -400 68874 240
rect 69409 -400 69465 240
rect 70000 -400 70056 240
rect 70591 -400 70647 240
rect 71182 -400 71238 240
rect 71773 -400 71829 240
rect 72364 -400 72420 240
rect 72955 -400 73011 240
rect 73546 -400 73602 240
rect 74137 -400 74193 240
rect 74728 -400 74784 240
rect 75319 -400 75375 240
rect 75910 -400 75966 240
rect 76501 -400 76557 240
rect 77092 -400 77148 240
rect 77683 -400 77739 240
rect 78274 -400 78330 240
rect 78865 -400 78921 240
rect 79456 -400 79512 240
rect 80047 -400 80103 240
rect 80638 -400 80694 240
rect 81229 -400 81285 240
rect 81820 -400 81876 240
rect 82411 -400 82467 240
rect 83002 -400 83058 240
rect 83593 -400 83649 240
rect 84184 -400 84240 240
rect 84775 -400 84831 240
rect 85366 -400 85422 240
rect 85957 -400 86013 240
rect 86548 -400 86604 240
rect 87139 -400 87195 240
rect 87730 -400 87786 240
rect 88321 -400 88377 240
rect 88912 -400 88968 240
rect 89503 -400 89559 240
rect 90094 -400 90150 240
rect 90685 -400 90741 240
rect 91276 -400 91332 240
rect 91867 -400 91923 240
rect 92458 -400 92514 240
rect 93049 -400 93105 240
rect 93640 -400 93696 240
rect 94231 -400 94287 240
rect 94822 -400 94878 240
rect 95413 -400 95469 240
rect 96004 -400 96060 240
rect 96595 -400 96651 240
rect 97186 -400 97242 240
rect 97777 -400 97833 240
rect 98368 -400 98424 240
rect 98959 -400 99015 240
rect 99550 -400 99606 240
rect 100141 -400 100197 240
rect 100732 -400 100788 240
rect 101323 -400 101379 240
rect 101914 -400 101970 240
rect 102505 -400 102561 240
rect 103096 -400 103152 240
rect 103687 -400 103743 240
rect 104278 -400 104334 240
rect 104869 -400 104925 240
rect 105460 -400 105516 240
rect 106051 -400 106107 240
rect 106642 -400 106698 240
rect 107233 -400 107289 240
rect 107824 -400 107880 240
rect 108415 -400 108471 240
rect 109006 -400 109062 240
rect 109597 -400 109653 240
rect 110188 -400 110244 240
rect 110779 -400 110835 240
rect 111370 -400 111426 240
rect 111961 -400 112017 240
rect 112552 -400 112608 240
rect 113143 -400 113199 240
rect 113734 -400 113790 240
rect 114325 -400 114381 240
rect 114916 -400 114972 240
rect 115507 -400 115563 240
rect 116098 -400 116154 240
rect 116689 -400 116745 240
rect 117280 -400 117336 240
rect 117871 -400 117927 240
rect 118462 -400 118518 240
rect 119053 -400 119109 240
rect 119644 -400 119700 240
rect 120235 -400 120291 240
rect 120826 -400 120882 240
rect 121417 -400 121473 240
rect 122008 -400 122064 240
rect 122599 -400 122655 240
rect 123190 -400 123246 240
rect 123781 -400 123837 240
rect 124372 -400 124428 240
rect 124963 -400 125019 240
rect 125554 -400 125610 240
rect 126145 -400 126201 240
rect 126736 -400 126792 240
rect 127327 -400 127383 240
rect 127918 -400 127974 240
rect 128509 -400 128565 240
rect 129100 -400 129156 240
rect 129691 -400 129747 240
rect 130282 -400 130338 240
rect 130873 -400 130929 240
rect 131464 -400 131520 240
rect 132055 -400 132111 240
rect 132646 -400 132702 240
rect 133237 -400 133293 240
rect 133828 -400 133884 240
rect 134419 -400 134475 240
rect 135010 -400 135066 240
rect 135601 -400 135657 240
rect 136192 -400 136248 240
rect 136783 -400 136839 240
rect 137374 -400 137430 240
rect 137965 -400 138021 240
rect 138556 -400 138612 240
rect 139147 -400 139203 240
rect 139738 -400 139794 240
rect 140329 -400 140385 240
rect 140920 -400 140976 240
rect 141511 -400 141567 240
rect 142102 -400 142158 240
rect 142693 -400 142749 240
rect 143284 -400 143340 240
rect 143875 -400 143931 240
rect 144466 -400 144522 240
rect 145057 -400 145113 240
rect 145648 -400 145704 240
rect 146239 -400 146295 240
rect 146830 -400 146886 240
rect 147421 -400 147477 240
rect 148012 -400 148068 240
rect 148603 -400 148659 240
rect 149194 -400 149250 240
rect 149785 -400 149841 240
rect 150376 -400 150432 240
rect 150967 -400 151023 240
rect 151558 -400 151614 240
rect 152149 -400 152205 240
rect 152740 -400 152796 240
rect 153331 -400 153387 240
rect 153922 -400 153978 240
rect 154513 -400 154569 240
rect 155104 -400 155160 240
rect 155695 -400 155751 240
rect 156286 -400 156342 240
rect 156877 -400 156933 240
rect 157468 -400 157524 240
rect 158059 -400 158115 240
rect 158650 -400 158706 240
rect 159241 -400 159297 240
rect 159832 -400 159888 240
rect 160423 -400 160479 240
rect 161014 -400 161070 240
rect 161605 -400 161661 240
rect 162196 -400 162252 240
rect 162787 -400 162843 240
rect 163378 -400 163434 240
rect 163969 -400 164025 240
rect 164560 -400 164616 240
rect 165151 -400 165207 240
rect 165742 -400 165798 240
rect 166333 -400 166389 240
rect 166924 -400 166980 240
rect 167515 -400 167571 240
rect 168106 -400 168162 240
rect 168697 -400 168753 240
rect 169288 -400 169344 240
rect 169879 -400 169935 240
rect 170470 -400 170526 240
rect 171061 -400 171117 240
rect 171652 -400 171708 240
rect 172243 -400 172299 240
rect 172834 -400 172890 240
rect 173425 -400 173481 240
rect 174016 -400 174072 240
rect 174607 -400 174663 240
rect 175198 -400 175254 240
rect 175789 -400 175845 240
rect 176380 -400 176436 240
rect 176971 -400 177027 240
rect 177562 -400 177618 240
rect 178153 -400 178209 240
rect 178744 -400 178800 240
rect 179335 -400 179391 240
rect 179926 -400 179982 240
rect 180517 -400 180573 240
rect 181108 -400 181164 240
rect 181699 -400 181755 240
rect 182290 -400 182346 240
rect 182881 -400 182937 240
rect 183472 -400 183528 240
rect 184063 -400 184119 240
rect 184654 -400 184710 240
rect 185245 -400 185301 240
rect 185836 -400 185892 240
rect 186427 -400 186483 240
rect 187018 -400 187074 240
rect 187609 -400 187665 240
rect 188200 -400 188256 240
rect 188791 -400 188847 240
rect 189382 -400 189438 240
rect 189973 -400 190029 240
rect 190564 -400 190620 240
rect 191155 -400 191211 240
rect 191746 -400 191802 240
rect 192337 -400 192393 240
rect 192928 -400 192984 240
rect 193519 -400 193575 240
rect 194110 -400 194166 240
rect 194701 -400 194757 240
rect 195292 -400 195348 240
rect 195883 -400 195939 240
rect 196474 -400 196530 240
rect 197065 -400 197121 240
rect 197656 -400 197712 240
rect 198247 -400 198303 240
rect 198838 -400 198894 240
rect 199429 -400 199485 240
rect 200020 -400 200076 240
rect 200611 -400 200667 240
rect 201202 -400 201258 240
rect 201793 -400 201849 240
rect 202384 -400 202440 240
rect 202975 -400 203031 240
rect 203566 -400 203622 240
rect 204157 -400 204213 240
rect 204748 -400 204804 240
rect 205339 -400 205395 240
rect 205930 -400 205986 240
rect 206521 -400 206577 240
rect 207112 -400 207168 240
rect 207703 -400 207759 240
rect 208294 -400 208350 240
rect 208885 -400 208941 240
rect 209476 -400 209532 240
rect 210067 -400 210123 240
rect 210658 -400 210714 240
rect 211249 -400 211305 240
rect 211840 -400 211896 240
rect 212431 -400 212487 240
rect 213022 -400 213078 240
rect 213613 -400 213669 240
rect 214204 -400 214260 240
rect 214795 -400 214851 240
rect 215386 -400 215442 240
rect 215977 -400 216033 240
rect 216568 -400 216624 240
rect 217159 -400 217215 240
rect 217750 -400 217806 240
rect 218341 -400 218397 240
rect 218932 -400 218988 240
rect 219523 -400 219579 240
rect 220114 -400 220170 240
rect 220705 -400 220761 240
rect 221296 -400 221352 240
rect 221887 -400 221943 240
rect 222478 -400 222534 240
rect 223069 -400 223125 240
rect 223660 -400 223716 240
rect 224251 -400 224307 240
rect 224842 -400 224898 240
rect 225433 -400 225489 240
rect 226024 -400 226080 240
rect 226615 -400 226671 240
rect 227206 -400 227262 240
rect 227797 -400 227853 240
rect 228388 -400 228444 240
rect 228979 -400 229035 240
rect 229570 -400 229626 240
rect 230161 -400 230217 240
rect 230752 -400 230808 240
rect 231343 -400 231399 240
rect 231934 -400 231990 240
rect 232525 -400 232581 240
rect 233116 -400 233172 240
rect 233707 -400 233763 240
rect 234298 -400 234354 240
rect 234889 -400 234945 240
rect 235480 -400 235536 240
rect 236071 -400 236127 240
rect 236662 -400 236718 240
rect 237253 -400 237309 240
rect 237844 -400 237900 240
rect 238435 -400 238491 240
rect 239026 -400 239082 240
rect 239617 -400 239673 240
rect 240208 -400 240264 240
rect 240799 -400 240855 240
rect 241390 -400 241446 240
rect 241981 -400 242037 240
rect 242572 -400 242628 240
rect 243163 -400 243219 240
rect 243754 -400 243810 240
rect 244345 -400 244401 240
rect 244936 -400 244992 240
rect 245527 -400 245583 240
rect 246118 -400 246174 240
rect 246709 -400 246765 240
rect 247300 -400 247356 240
rect 247891 -400 247947 240
rect 248482 -400 248538 240
rect 249073 -400 249129 240
rect 249664 -400 249720 240
rect 250255 -400 250311 240
rect 250846 -400 250902 240
rect 251437 -400 251493 240
rect 252028 -400 252084 240
rect 252619 -400 252675 240
rect 253210 -400 253266 240
rect 253801 -400 253857 240
rect 254392 -400 254448 240
rect 254983 -400 255039 240
rect 255574 -400 255630 240
rect 256165 -400 256221 240
rect 256756 -400 256812 240
rect 257347 -400 257403 240
rect 257938 -400 257994 240
rect 258529 -400 258585 240
rect 259120 -400 259176 240
rect 259711 -400 259767 240
rect 260302 -400 260358 240
rect 260893 -400 260949 240
rect 261484 -400 261540 240
rect 262075 -400 262131 240
rect 262666 -400 262722 240
rect 263257 -400 263313 240
rect 263848 -400 263904 240
rect 264439 -400 264495 240
rect 265030 -400 265086 240
rect 265621 -400 265677 240
rect 266212 -400 266268 240
rect 266803 -400 266859 240
rect 267394 -400 267450 240
rect 267985 -400 268041 240
rect 268576 -400 268632 240
rect 269167 -400 269223 240
rect 269758 -400 269814 240
rect 270349 -400 270405 240
rect 270940 -400 270996 240
rect 271531 -400 271587 240
rect 272122 -400 272178 240
rect 272713 -400 272769 240
rect 273304 -400 273360 240
rect 273895 -400 273951 240
rect 274486 -400 274542 240
rect 275077 -400 275133 240
rect 275668 -400 275724 240
rect 276259 -400 276315 240
rect 276850 -400 276906 240
rect 277441 -400 277497 240
rect 278032 -400 278088 240
rect 278623 -400 278679 240
rect 279214 -400 279270 240
rect 279805 -400 279861 240
rect 280396 -400 280452 240
rect 280987 -400 281043 240
rect 281578 -400 281634 240
rect 282169 -400 282225 240
rect 282760 -400 282816 240
rect 283351 -400 283407 240
rect 283942 -400 283998 240
rect 284533 -400 284589 240
rect 285124 -400 285180 240
rect 285715 -400 285771 240
rect 286306 -400 286362 240
rect 286897 -400 286953 240
rect 287488 -400 287544 240
rect 288079 -400 288135 240
rect 288670 -400 288726 240
rect 289261 -400 289317 240
rect 289852 -400 289908 240
rect 290443 -400 290499 240
rect 291034 -400 291090 240
rect 291625 -400 291681 240
<< via2 >>
rect 164500 338774 165766 339949
rect 164481 331688 165747 332863
rect 164500 325316 165766 326491
rect 164481 318230 165747 319405
rect 164506 311055 165772 312230
rect 164487 303969 165753 305144
rect 164595 294696 165861 295871
rect 164576 287610 165842 288785
rect 164539 281208 165805 282383
rect 164646 272288 165912 273463
rect 164627 265202 165893 266377
rect 164590 258800 165856 259975
rect 164677 248034 165943 249209
rect 164658 240948 165924 242123
rect 164621 234546 165887 235721
rect 164801 227768 166067 228943
rect 164781 221906 166047 223081
rect 164821 209843 166087 211018
rect 164802 202757 166068 203932
rect 164765 196355 166031 197530
rect 164808 191950 166074 193125
rect 164789 184864 166055 186039
rect 164752 178462 166018 179637
rect 164612 172537 165878 173712
rect 164575 166135 165841 167310
rect 164841 158874 166107 160049
rect 164822 154034 166088 155209
rect 164803 148764 166069 149939
rect 164785 143212 166051 144387
rect 164785 137022 166051 138197
rect 164793 117918 166059 119093
rect 164902 109991 166168 111166
rect 165003 101789 166269 102964
rect 164966 94290 166232 95465
rect 164947 87204 166213 88379
rect 164910 80802 166176 81977
rect 164892 69552 166158 70727
rect 164818 63557 166084 64732
rect 164855 57729 166121 58904
rect 164929 51642 166195 52817
rect 164641 43784 165907 44959
rect 164641 37490 165907 38665
rect 164641 31196 165907 32371
<< metal3 >>
rect 8097 351150 10597 352400
rect 34097 351150 36597 352400
rect 60097 351150 62597 352400
rect 82797 351150 85297 352400
rect 85447 351150 86547 352400
rect 86697 351150 87797 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 111297 351150 112397 352400
rect 112547 351150 113647 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 162147 351150 163247 352400
rect 163397 351150 164497 352400
rect 164647 351150 167147 352400
rect 206697 351150 209197 352400
rect 232697 351150 235197 352400
rect 255297 351170 257697 352400
rect 260297 351170 262697 352400
rect 8376 349233 10412 351150
rect 34331 349233 36367 351150
rect 60339 349338 62375 351150
rect 82963 349244 84999 351150
rect 88168 349208 90204 351150
rect 108814 349155 110850 351150
rect 114054 349155 116090 351150
rect 159668 349191 161704 351150
rect 164874 349155 166910 351150
rect 206890 349311 208926 351150
rect 232866 349389 234902 351150
rect 255440 349320 257476 351170
rect 260451 349303 262487 351170
rect 283297 351150 285797 352400
rect 283588 349206 285624 351150
rect -400 342364 850 342621
rect -400 340471 4906 342364
rect 291150 341209 292400 341492
rect -400 340121 850 340471
rect 164427 339949 165848 340032
rect 164427 338774 164500 339949
rect 165766 338774 165848 339949
rect 287117 339172 292400 341209
rect 291150 338992 292400 339172
rect 164427 338683 165848 338774
rect 164408 332863 165829 332946
rect 164408 331688 164481 332863
rect 165747 331688 165829 332863
rect 164408 331597 165829 331688
rect 164427 326491 165848 326574
rect 164427 325316 164500 326491
rect 165766 325316 165848 326491
rect 164427 325225 165848 325316
rect -400 324049 830 324321
rect -400 322156 4976 324049
rect -400 321921 830 322156
rect 291170 322092 292400 322292
rect 287015 320055 292400 322092
rect 291170 319892 292400 320055
rect 164408 319405 165829 319488
rect -400 319125 830 319321
rect -400 317232 4906 319125
rect 164408 318230 164481 319405
rect 165747 318230 165829 319405
rect 164408 318139 165829 318230
rect -400 316921 830 317232
rect 291170 317127 292400 317292
rect 287114 315090 292400 317127
rect 291170 314892 292400 315090
rect 164433 312230 165854 312313
rect 164433 311055 164506 312230
rect 165772 311055 165854 312230
rect 164433 310964 165854 311055
rect 164414 305144 165835 305227
rect 164414 303969 164487 305144
rect 165753 303969 165835 305144
rect 164414 303878 165835 303969
rect 164522 295871 165943 295954
rect 164522 294696 164595 295871
rect 165861 294696 165943 295871
rect 291760 294736 292400 294792
rect 164522 294605 165943 294696
rect 291760 294145 292400 294201
rect 291760 293554 292400 293610
rect 291760 292963 292400 293019
rect 287531 292428 291858 292545
rect 287531 292372 292400 292428
rect 287531 292267 291858 292372
rect 287523 291837 291850 291977
rect 287523 291781 292400 291837
rect 287523 291699 291850 291781
rect 164503 288785 165924 288868
rect 164503 287610 164576 288785
rect 165842 287610 165924 288785
rect 164503 287519 165924 287610
rect 164466 282383 165887 282466
rect -400 281893 830 282121
rect -400 280000 4941 281893
rect 164466 281208 164539 282383
rect 165805 281208 165887 282383
rect 164466 281117 165887 281208
rect -400 279721 830 280000
rect 273285 277424 287287 277475
rect 291170 277424 292400 277681
rect -400 276863 830 277121
rect 273285 276989 292400 277424
rect -400 274970 4906 276863
rect 273285 275847 273813 276989
rect 275123 275847 292400 276989
rect 273285 275531 292400 275847
rect 273285 275503 287287 275531
rect 291170 275281 292400 275531
rect -400 274721 830 274970
rect 164573 273463 165994 273546
rect 164573 272288 164646 273463
rect 165912 272288 165994 273463
rect 291170 272430 292400 272681
rect 164573 272197 165994 272288
rect 286997 270537 292400 272430
rect 291170 270281 292400 270537
rect 164554 266377 165975 266460
rect 164554 265202 164627 266377
rect 165893 265202 165975 266377
rect 164554 265111 165975 265202
rect 164517 259975 165938 260058
rect 164517 258800 164590 259975
rect 165856 258800 165938 259975
rect 164517 258709 165938 258800
rect 176 255821 1564 255918
rect -400 255765 1564 255821
rect 176 255663 1564 255765
rect 190 255230 1578 255336
rect -400 255174 1578 255230
rect 190 255081 1578 255174
rect -400 254583 240 254639
rect -400 253992 240 254048
rect -400 253401 240 253457
rect -400 252810 240 252866
rect 291760 250025 292400 250081
rect 291760 249434 292400 249490
rect 164604 249209 166025 249292
rect 164604 248034 164677 249209
rect 165943 248034 166025 249209
rect 291760 248843 292400 248899
rect 291760 248252 292400 248308
rect 164604 247943 166025 248034
rect 291760 247661 292400 247717
rect 291760 247070 292400 247126
rect 164585 242123 166006 242206
rect 164585 240948 164658 242123
rect 165924 240948 166006 242123
rect 164585 240857 166006 240948
rect 164548 235721 165969 235804
rect 164548 234546 164621 235721
rect 165887 234546 165969 235721
rect 164548 234455 165969 234546
rect 153 234210 1541 234292
rect -400 234154 1541 234210
rect 153 234037 1541 234154
rect 176 233619 1564 233734
rect -400 233563 1564 233619
rect 176 233479 1564 233563
rect -400 232972 240 233028
rect -400 232381 240 232437
rect -400 231790 240 231846
rect -400 231199 240 231255
rect 164728 228943 166149 229026
rect 164728 227768 164801 228943
rect 166067 227768 166149 228943
rect 291760 227814 292400 227870
rect 164728 227677 166149 227768
rect 291760 227223 292400 227279
rect 291760 226632 292400 226688
rect 291760 226041 292400 226097
rect 291760 225450 292400 225506
rect 291760 224859 292400 224915
rect 164708 223081 166129 223164
rect 164708 221906 164781 223081
rect 166047 221906 166129 223081
rect 164708 221815 166129 221906
rect 171 212599 1559 212727
rect -400 212543 1559 212599
rect 171 212472 1559 212543
rect 175 212008 1563 212112
rect -400 211952 1563 212008
rect 175 211857 1563 211952
rect -400 211361 240 211417
rect 164748 211018 166169 211101
rect -400 210770 240 210826
rect -400 210179 240 210235
rect 164748 209843 164821 211018
rect 166087 209843 166169 211018
rect 164748 209752 166169 209843
rect -400 209588 240 209644
rect 291760 205603 292400 205659
rect 291760 205012 292400 205068
rect 291760 204421 292400 204477
rect 164729 203932 166150 204015
rect 164729 202757 164802 203932
rect 166068 202757 166150 203932
rect 291760 203830 292400 203886
rect 291760 203239 292400 203295
rect 164729 202666 166150 202757
rect 291760 202648 292400 202704
rect 164692 197530 166113 197613
rect 164692 196355 164765 197530
rect 166031 196355 166113 197530
rect 164692 196264 166113 196355
rect 164735 193125 166156 193208
rect 164735 191950 164808 193125
rect 166074 191950 166156 193125
rect 164735 191859 166156 191950
rect 185 190988 1573 191097
rect -400 190932 1573 190988
rect 185 190842 1573 190932
rect 204 190397 1592 190525
rect -400 190341 1592 190397
rect 204 190270 1592 190341
rect -400 189750 240 189806
rect -400 189159 240 189215
rect -400 188568 240 188624
rect -400 187977 240 188033
rect 164716 186039 166137 186122
rect 164716 184864 164789 186039
rect 166055 184864 166137 186039
rect 164716 184773 166137 184864
rect 291760 182392 292400 182448
rect 291760 181801 292400 181857
rect 291760 181210 292400 181266
rect 291760 180619 292400 180675
rect 291760 180028 292400 180084
rect 164679 179637 166100 179720
rect 164679 178462 164752 179637
rect 166018 178462 166100 179637
rect 291760 179437 292400 179493
rect 164679 178371 166100 178462
rect 164539 173712 165960 173795
rect 164539 172537 164612 173712
rect 165878 172537 165960 173712
rect 164539 172446 165960 172537
rect 181 169377 1569 169509
rect -400 169321 1569 169377
rect 181 169254 1569 169321
rect 199 168786 1587 168886
rect -400 168730 1587 168786
rect 199 168631 1587 168730
rect -400 168139 240 168195
rect -400 167548 240 167604
rect 164502 167310 165923 167393
rect -400 166957 240 167013
rect -400 166366 240 166422
rect 164502 166135 164575 167310
rect 165841 166135 165923 167310
rect 164502 166044 165923 166135
rect 164768 160049 166189 160132
rect 164768 158874 164841 160049
rect 166107 158874 166189 160049
rect 291760 159781 292400 159837
rect 291760 159190 292400 159246
rect 164768 158783 166189 158874
rect 291760 158599 292400 158655
rect 291760 158008 292400 158064
rect 291760 157417 292400 157473
rect 291760 156826 292400 156882
rect 164749 155209 166170 155292
rect 164749 154034 164822 155209
rect 166088 154034 166170 155209
rect 164749 153943 166170 154034
rect 164730 149939 166151 150022
rect 164730 148764 164803 149939
rect 166069 148764 166151 149939
rect 164730 148673 166151 148764
rect 190 147766 1578 147897
rect -400 147710 1578 147766
rect 190 147642 1578 147710
rect 218 147175 1606 147320
rect -400 147119 1606 147175
rect 218 147065 1606 147119
rect -400 146528 240 146584
rect -400 145937 240 145993
rect -400 145346 240 145402
rect -400 144755 240 144811
rect 164712 144387 166133 144470
rect 164712 143212 164785 144387
rect 166051 143212 166133 144387
rect 164712 143121 166133 143212
rect 164712 138197 166133 138280
rect 164712 137022 164785 138197
rect 166051 137022 166133 138197
rect 291760 137570 292400 137626
rect 164712 136931 166133 137022
rect 291760 136979 292400 137035
rect 291760 136388 292400 136444
rect 291760 135797 292400 135853
rect 291760 135206 292400 135262
rect 291760 134615 292400 134671
rect 195 126255 1583 126392
rect -400 126199 1583 126255
rect 195 126137 1583 126199
rect 204 125664 1592 125824
rect -400 125608 1592 125664
rect 204 125569 1592 125608
rect -400 125017 240 125073
rect -400 124426 240 124482
rect -400 123835 240 123891
rect -400 123244 240 123300
rect 164720 119093 166141 119176
rect 164720 117918 164793 119093
rect 166059 117918 166141 119093
rect 164720 117827 166141 117918
rect 291170 117615 292400 120015
rect 291170 112615 292400 115015
rect 164829 111166 166250 111249
rect 164829 109991 164902 111166
rect 166168 109991 166250 111166
rect 164829 109900 166250 109991
rect -400 109532 830 109844
rect -400 107639 4916 109532
rect -400 107444 830 107639
rect -400 104575 830 104844
rect -400 102682 4916 104575
rect 164930 102964 166351 103047
rect -400 102444 830 102682
rect 164930 101789 165003 102964
rect 166269 101789 166351 102964
rect 164930 101698 166351 101789
rect 291170 95715 292400 98115
rect 164893 95465 166314 95548
rect 164893 94290 164966 95465
rect 166232 94290 166314 95465
rect 164893 94199 166314 94290
rect 291170 90715 292400 93115
rect -400 88533 830 88844
rect -400 86640 4920 88533
rect 164874 88379 166295 88462
rect 164874 87204 164947 88379
rect 166213 87204 166295 88379
rect 164874 87113 166295 87204
rect -400 86444 830 86640
rect -400 83589 830 83844
rect -400 81696 4990 83589
rect 164837 81977 166258 82060
rect -400 81444 830 81696
rect 164837 80802 164910 81977
rect 166176 80802 166258 81977
rect 164837 80711 166258 80802
rect 280813 75549 287932 75721
rect 291170 75549 292400 75815
rect 280813 75451 292400 75549
rect 280813 73748 281123 75451
rect 282980 73748 292400 75451
rect 280813 73656 292400 73748
rect 280813 73527 288755 73656
rect 280813 73516 286531 73527
rect 291170 73415 292400 73656
rect 164819 70727 166240 70810
rect 164819 69552 164892 70727
rect 166158 69552 166240 70727
rect 164819 69461 166240 69552
rect 287067 70535 288755 70545
rect 291170 70535 292400 70815
rect 287067 68984 292400 70535
rect 287095 68642 292400 68984
rect 291170 68415 292400 68642
rect 164745 64732 166166 64815
rect 164745 63557 164818 64732
rect 166084 63557 166166 64732
rect 164745 63466 166166 63557
rect 181 62444 1569 62587
rect -400 62388 1569 62444
rect 181 62332 1569 62388
rect 199 61853 1587 62001
rect -400 61797 1587 61853
rect 199 61746 1587 61797
rect -400 61206 240 61262
rect -400 60615 240 60671
rect -400 60024 240 60080
rect -400 59433 240 59489
rect 164782 58904 166203 58987
rect 164782 57729 164855 58904
rect 166121 57729 166203 58904
rect 164782 57638 166203 57729
rect 164856 52817 166277 52900
rect 164856 51642 164929 52817
rect 166195 51642 166277 52817
rect 164856 51551 166277 51642
rect 291760 47559 292400 47615
rect 291760 46968 292400 47024
rect 291760 46377 292400 46433
rect 291760 45786 292400 45842
rect 164568 44959 165989 45042
rect 164568 43784 164641 44959
rect 165907 43784 165989 44959
rect 164568 43693 165989 43784
rect 195 40833 1583 41003
rect -400 40777 1583 40833
rect 195 40748 1583 40777
rect 204 40242 1592 40399
rect -400 40186 1592 40242
rect 204 40144 1592 40186
rect -400 39595 240 39651
rect -400 39004 240 39060
rect 164568 38665 165989 38748
rect -400 38413 240 38469
rect -400 37822 240 37878
rect 164568 37490 164641 38665
rect 165907 37490 165989 38665
rect 164568 37399 165989 37490
rect 164568 32371 165989 32454
rect 164568 31196 164641 32371
rect 165907 31196 165989 32371
rect 164568 31105 165989 31196
rect 291760 25230 292400 25286
rect 291760 24639 292400 24695
rect 291760 24048 292400 24104
rect 291760 23457 292400 23513
rect 199 19222 1587 19359
rect -400 19166 1587 19222
rect 199 19104 1587 19166
rect 195 18631 1583 18746
rect -400 18575 1583 18631
rect 195 18491 1583 18575
rect -400 17984 240 18040
rect -400 17393 240 17449
rect -400 16802 240 16858
rect -400 16211 240 16267
rect 291760 12001 292400 12057
rect 291760 11410 292400 11466
rect 291760 10819 292400 10875
rect 291760 10228 292400 10284
rect 291760 9637 292400 9693
rect 291760 9046 292400 9102
rect 195 8511 1583 8651
rect -400 8455 1583 8511
rect 291760 8455 292400 8511
rect 195 8396 1583 8455
rect 213 7920 1601 8041
rect -400 7864 1601 7920
rect 291760 7864 292400 7920
rect 213 7786 1601 7864
rect -400 7273 240 7329
rect 291760 7273 292400 7329
rect -400 6682 240 6738
rect 291760 6682 292400 6738
rect -400 6091 240 6147
rect 291760 6091 292400 6147
rect -400 5500 240 5556
rect 291760 5500 292400 5556
rect -400 4909 240 4965
rect 291760 4909 292400 4965
rect -400 4318 240 4374
rect 291760 4318 292400 4374
rect -400 3727 240 3783
rect 291760 3727 292400 3783
rect -400 3136 240 3192
rect 291760 3136 292400 3192
rect -400 2545 240 2601
rect 291760 2545 292400 2601
rect -400 1954 240 2010
rect 291760 1954 292400 2010
rect -400 1363 240 1419
rect 291760 1363 292400 1419
rect -400 772 240 828
rect 291760 772 292400 828
<< via3 >>
rect 164500 338774 165766 339949
rect 164481 331688 165747 332863
rect 164500 325316 165766 326491
rect 164481 318230 165747 319405
rect 164506 311055 165772 312230
rect 164487 303969 165753 305144
rect 164595 294696 165861 295871
rect 164576 287610 165842 288785
rect 164539 281208 165805 282383
rect 273813 275847 275123 276989
rect 164646 272288 165912 273463
rect 164627 265202 165893 266377
rect 164590 258800 165856 259975
rect 164677 248034 165943 249209
rect 164658 240948 165924 242123
rect 164621 234546 165887 235721
rect 164801 227768 166067 228943
rect 164781 221906 166047 223081
rect 164821 209843 166087 211018
rect 164802 202757 166068 203932
rect 164765 196355 166031 197530
rect 164808 191950 166074 193125
rect 164789 184864 166055 186039
rect 164752 178462 166018 179637
rect 164612 172537 165878 173712
rect 164575 166135 165841 167310
rect 164841 158874 166107 160049
rect 164822 154034 166088 155209
rect 164803 148764 166069 149939
rect 164785 143212 166051 144387
rect 164785 137022 166051 138197
rect 164793 117918 166059 119093
rect 164902 109991 166168 111166
rect 165003 101789 166269 102964
rect 164966 94290 166232 95465
rect 164947 87204 166213 88379
rect 164910 80802 166176 81977
rect 281123 73748 282980 75451
rect 164892 69552 166158 70727
rect 164818 63557 166084 64732
rect 164855 57729 166121 58904
rect 164929 51642 166195 52817
rect 164641 43784 165907 44959
rect 164641 37490 165907 38665
rect 164641 31196 165907 32371
<< metal4 >>
rect 82797 351150 85297 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 164647 351150 167147 352400
rect 82963 349244 84999 351150
rect 88168 349208 90204 351150
rect 108814 349155 110850 351150
rect 114054 349155 116090 351150
rect 159668 349191 161704 351150
rect 164874 349155 166910 351150
rect 164359 341807 166659 342174
rect 164270 341177 166659 341807
rect 163899 339949 166659 341177
rect 163899 338774 164500 339949
rect 165766 338774 166659 339949
rect 163899 337301 166659 338774
rect 163899 333969 166665 337301
rect 163791 332863 166665 333969
rect 163791 331688 164481 332863
rect 165747 331688 166665 332863
rect 163791 331547 166665 331688
rect 163789 330649 166665 331547
rect 164365 328716 166665 330649
rect 164359 328349 166665 328716
rect 164270 327719 166665 328349
rect 163899 326491 166665 327719
rect 163899 325316 164500 326491
rect 165766 325316 166665 326491
rect 163899 320511 166665 325316
rect 163791 319405 166665 320511
rect 10583 318426 11415 318528
rect 10583 301349 11422 318426
rect 163791 318230 164481 319405
rect 165747 318230 166665 319405
rect 163791 318089 166665 318230
rect 163789 317191 166665 318089
rect 164365 314088 166665 317191
rect 164276 313458 166665 314088
rect 163905 312230 166665 313458
rect 163905 311055 164506 312230
rect 165772 311055 166665 312230
rect 163905 306250 166665 311055
rect 163797 305144 166665 306250
rect 163797 303969 164487 305144
rect 165753 303969 166665 305144
rect 163797 303828 166665 303969
rect 163795 302921 166665 303828
rect 163905 302753 166665 302921
rect 9451 301304 18902 301349
rect 9451 301000 83398 301304
rect 164365 301000 166665 302753
rect 233832 301000 234467 306499
rect 241132 301000 241198 301061
rect 9451 299000 241198 301000
rect 9451 298973 83398 299000
rect 9451 298867 18902 298973
rect 164365 297099 166665 299000
rect 163994 295871 166665 297099
rect 163994 294696 164595 295871
rect 165861 294696 166665 295871
rect 163994 289891 166665 294696
rect 163886 288785 166665 289891
rect 163886 287610 164576 288785
rect 165842 287610 166665 288785
rect 163886 287469 166665 287610
rect 163884 286562 166665 287469
rect 163994 282383 166665 286562
rect 163994 281208 164539 282383
rect 165805 282016 166665 282383
rect 165805 281208 166759 282016
rect 163994 281056 166759 281208
rect 163992 280229 166759 281056
rect 164356 274691 166759 280229
rect 273495 276989 275423 277344
rect 273495 275847 273813 276989
rect 275123 275847 275423 276989
rect 273495 275548 275423 275847
rect 164045 273463 166759 274691
rect 164045 272288 164646 273463
rect 165912 272547 166759 273463
rect 165912 272524 166735 272547
rect 165912 272288 166716 272524
rect 164045 267483 166716 272288
rect 163937 266377 166716 267483
rect 163937 265202 164627 266377
rect 165893 265202 166716 266377
rect 163937 265061 166716 265202
rect 163935 264154 166716 265061
rect 12067 257000 12435 260680
rect 164045 259975 166716 264154
rect 164045 258800 164590 259975
rect 165856 259608 166716 259975
rect 165856 258800 166810 259608
rect 164045 258648 166810 258800
rect 164043 257821 166810 258648
rect 164365 257000 166810 257821
rect 266660 257000 267646 259231
rect 10000 256998 17520 257000
rect 29189 256998 62683 257000
rect 10000 256982 62683 256998
rect 70642 256982 275000 257000
rect 10000 255000 275000 256982
rect 164365 250449 166665 255000
rect 164365 250437 166790 250449
rect 164076 249209 166790 250437
rect 164076 248034 164677 249209
rect 165943 248293 166790 249209
rect 165943 248270 166766 248293
rect 165943 248034 166747 248270
rect 164076 243229 166747 248034
rect 163968 242123 166747 243229
rect 163968 240948 164658 242123
rect 165924 240948 166747 242123
rect 163968 240807 166747 240948
rect 163966 239900 166747 240807
rect 164076 235721 166747 239900
rect 164076 234546 164621 235721
rect 165887 235354 166747 235721
rect 165887 234546 166841 235354
rect 164076 234394 166841 234546
rect 164074 233567 166841 234394
rect 164365 233402 166841 233567
rect 164365 232000 166665 233402
rect 226048 232000 233060 232026
rect 69559 230000 233060 232000
rect 141157 229989 144509 230000
rect 164200 228943 166666 230000
rect 226048 229978 233060 230000
rect 164200 227768 164801 228943
rect 166067 227768 166666 228943
rect 164200 227671 166666 227768
rect 164200 226887 166717 227671
rect 164365 224776 166665 226887
rect 164180 223081 166665 224776
rect 164180 221906 164781 223081
rect 166047 221906 166665 223081
rect 164180 221809 166665 221906
rect 164180 221025 166697 221809
rect 164365 220000 166665 221025
rect 10000 219916 13587 220000
rect 42004 219916 226465 220000
rect 10000 218000 226465 219916
rect 164365 213295 166665 218000
rect 164220 212168 166665 213295
rect 164220 211018 166686 212168
rect 164220 209843 164821 211018
rect 166087 209843 166686 211018
rect 164220 209746 166686 209843
rect 164220 208839 166737 209746
rect 164220 205038 166665 208839
rect 164112 203932 166665 205038
rect 164112 202757 164802 203932
rect 166068 202757 166665 203932
rect 164112 202616 166665 202757
rect 164110 201709 166665 202616
rect 164220 197530 166665 201709
rect 164220 196355 164765 197530
rect 166031 196355 166665 197530
rect 164220 196203 166665 196355
rect 164218 194676 166665 196203
rect 164207 194275 166665 194676
rect 164207 193125 166673 194275
rect 164207 191950 164808 193125
rect 166074 191950 166673 193125
rect 164207 191853 166673 191950
rect 164207 190946 166724 191853
rect 164207 187145 166665 190946
rect 164099 186039 166665 187145
rect 164099 184864 164789 186039
rect 166055 184864 166665 186039
rect 164099 184723 166665 184864
rect 164097 183816 166665 184723
rect 164207 179637 166665 183816
rect 164207 178462 164752 179637
rect 166018 178462 166665 179637
rect 164207 178310 166665 178462
rect 164205 176358 166665 178310
rect 164365 175011 166665 176358
rect 164030 174818 166665 175011
rect 163922 173712 166665 174818
rect 163922 172537 164612 173712
rect 165878 172537 166665 173712
rect 163922 172396 166665 172537
rect 163920 171489 166665 172396
rect 10534 165067 10981 168538
rect 164030 167310 166665 171489
rect 164030 166135 164575 167310
rect 165841 166135 166665 167310
rect 164030 165983 166665 166135
rect 10534 165029 11651 165067
rect 9697 165000 12075 165029
rect 32579 165000 33270 165217
rect 62513 165000 64054 165233
rect 164028 165000 166665 165983
rect 9697 163000 276000 165000
rect 9697 162893 12075 163000
rect 164365 160826 166665 163000
rect 164148 160049 167097 160826
rect 164148 158874 164841 160049
rect 166107 158874 167097 160049
rect 164148 158644 167097 158874
rect 164148 158070 167148 158644
rect 164365 155993 166665 158070
rect 164365 155209 167382 155993
rect 164365 154034 164822 155209
rect 166088 154034 167382 155209
rect 164365 153811 167382 154034
rect 164365 153237 167433 153811
rect 164365 150733 166665 153237
rect 164365 149939 167453 150733
rect 164365 148764 164803 149939
rect 166069 148764 167453 149939
rect 164365 148551 167453 148764
rect 164365 147977 167504 148551
rect 164365 145259 166665 147977
rect 164365 144387 167382 145259
rect 164365 143212 164785 144387
rect 166051 143212 167382 144387
rect 164365 143077 167382 143212
rect 164365 142503 167433 143077
rect 164365 139147 166665 142503
rect 164365 138197 167524 139147
rect 164365 137022 164785 138197
rect 166051 137022 167524 138197
rect 164365 136965 167524 137022
rect 164365 136391 167575 136965
rect 164365 131451 166665 136391
rect 164365 129091 167314 131451
rect 164365 128188 167365 129091
rect 164365 127000 166665 128188
rect 199052 127000 213617 127015
rect 12000 126577 213617 127000
rect 12000 125970 214266 126577
rect 12000 125000 213617 125970
rect 164365 120197 166665 125000
rect 199052 124968 213617 125000
rect 164365 119093 166831 120197
rect 164365 117918 164793 119093
rect 166059 117918 166831 119093
rect 164365 117775 166831 117918
rect 164365 116868 166882 117775
rect 164365 112245 166665 116868
rect 164365 111166 167036 112245
rect 164365 109991 164902 111166
rect 166168 109991 167036 111166
rect 164365 109823 167036 109991
rect 164365 108916 167087 109823
rect 164365 104019 166665 108916
rect 164365 102964 167036 104019
rect 164365 101789 165003 102964
rect 166269 101789 167036 102964
rect 164365 101597 167036 101789
rect 164365 100690 167087 101597
rect 164365 96615 166665 100690
rect 164365 95465 166831 96615
rect 164365 94290 164966 95465
rect 166232 94290 166831 95465
rect 164365 94193 166831 94290
rect 164365 93286 166882 94193
rect 13442 75873 14342 90992
rect 164365 89485 166665 93286
rect 164257 88379 166665 89485
rect 164257 87204 164947 88379
rect 166213 87204 166665 88379
rect 164257 87063 166665 87204
rect 164255 86156 166665 87063
rect 164365 81977 166665 86156
rect 164365 80802 164910 81977
rect 166176 80802 166665 81977
rect 164365 80650 166665 80802
rect 17351 75873 18404 78306
rect 164363 75873 166716 80650
rect 7143 75802 189636 75873
rect 272179 75802 279373 75823
rect 7143 75789 279373 75802
rect 7143 75451 283186 75789
rect 7143 73748 281123 75451
rect 282980 73748 283186 75451
rect 7143 73413 283186 73748
rect 7143 73379 274546 73413
rect 278502 73408 283186 73413
rect 164363 71584 166716 73379
rect 187580 73310 274546 73379
rect 164231 70727 166716 71584
rect 164231 69552 164892 70727
rect 166158 69552 166716 70727
rect 164231 69470 166716 69552
rect 164229 69372 166716 69470
rect 164229 68908 166665 69372
rect 164365 65344 166665 68908
rect 164196 64732 166665 65344
rect 164196 63557 164818 64732
rect 166084 63557 166665 64732
rect 164196 63230 166665 63557
rect 164194 62668 166665 63230
rect 164365 59627 166665 62668
rect 164161 58904 166665 59627
rect 164161 57729 164855 58904
rect 166121 57729 166665 58904
rect 164161 57513 166665 57729
rect 164159 56951 166665 57513
rect 164365 53422 166665 56951
rect 164092 52817 166665 53422
rect 164092 51642 164929 52817
rect 166195 51642 166665 52817
rect 164092 51308 166665 51642
rect 164090 50746 166665 51308
rect 164365 45727 166665 50746
rect 164349 45476 166665 45727
rect 163804 44959 166977 45476
rect 163804 43784 164641 44959
rect 165907 43784 166977 44959
rect 163804 43450 166977 43784
rect 163802 43049 166977 43450
rect 164349 42901 166665 43049
rect 164365 39433 166665 42901
rect 164349 39182 166665 39433
rect 163804 38665 166977 39182
rect 163804 37490 164641 38665
rect 165907 37490 166977 38665
rect 163804 37156 166977 37490
rect 163802 36755 166977 37156
rect 164349 36607 166665 36755
rect 164365 33139 166665 36607
rect 164349 32888 166665 33139
rect 163804 32371 166977 32888
rect 163804 31196 164641 32371
rect 165907 31196 166977 32371
rect 163804 30862 166977 31196
rect 163802 30461 166977 30862
rect 164349 30313 166665 30461
rect 11000 27995 19174 28000
rect 26432 27995 27306 29969
rect 164365 28000 166665 30313
rect 51796 27995 99535 28000
rect 11000 27979 99535 27995
rect 104181 27979 176227 28000
rect 11000 26000 176227 27979
rect 95970 25823 107673 26000
rect 164365 24479 166665 26000
<< via4 >>
rect 273813 275847 275123 276989
<< metal5 >>
rect 82797 351150 85297 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 164647 351150 167147 352400
rect 82963 349244 84999 351150
rect 88168 349208 90204 351150
rect 108814 349155 110850 351150
rect 114054 349155 116090 351150
rect 159668 349191 161704 351150
rect 164874 349155 166910 351150
rect 10000 341000 279000 343000
rect 12130 331056 12441 341000
rect 28333 340927 29338 341000
rect 100337 340994 103311 341000
rect 140522 340966 144447 341000
rect 156586 340685 160000 341000
rect 189353 340946 193169 341000
rect 156557 337000 160000 340685
rect 156557 333969 159446 337000
rect 156478 332036 159446 333969
rect 156419 330649 159446 332036
rect 157052 328716 159393 330649
rect 157046 328349 159393 328716
rect 156957 327719 159393 328349
rect 156586 327227 159393 327719
rect 156557 323816 159393 327227
rect 236749 325976 237463 341000
rect 238022 340997 240372 341000
rect 156557 320511 159446 323816
rect 156478 318578 159446 320511
rect 156419 317191 159446 318578
rect 157052 314088 159393 317191
rect 156963 313458 159393 314088
rect 156592 312966 159393 313458
rect 156563 309555 159393 312966
rect 156563 306250 159452 309555
rect 156484 304317 159452 306250
rect 156425 302921 159452 304317
rect 156592 302753 159452 302921
rect 157052 297099 159393 302753
rect 156681 296607 159393 297099
rect 156652 293196 159393 296607
rect 156652 289891 159541 293196
rect 156573 287958 159541 289891
rect 156514 286562 159541 287958
rect 156681 286108 159541 286562
rect 156681 281545 159393 286108
rect 156622 281056 159393 281545
rect 156622 280229 159389 281056
rect 157010 277890 159389 280229
rect 255736 277912 260234 277918
rect 255736 277906 272994 277912
rect 255736 277890 275442 277906
rect 9908 276989 275442 277890
rect 9908 275847 273813 276989
rect 275123 275847 275442 276989
rect 9908 275136 275442 275847
rect 9908 275109 272994 275136
rect 9908 274978 260234 275109
rect 9908 274941 17520 274978
rect 29189 274976 260234 274978
rect 9908 274937 14729 274941
rect 29189 274937 256191 274976
rect 13656 268363 14065 274937
rect 157010 274691 159444 274937
rect 156732 274199 159444 274691
rect 156703 270788 159444 274199
rect 156703 267483 159592 270788
rect 229206 268940 231073 274937
rect 156624 265550 159592 267483
rect 156565 264154 159592 265550
rect 156732 263700 159592 264154
rect 156732 259137 159444 263700
rect 156673 258648 159444 259137
rect 156673 257821 159440 258648
rect 157052 256386 159440 257821
rect 157052 253620 159393 256386
rect 156887 250449 159424 253620
rect 156887 250437 159475 250449
rect 156763 249945 159475 250437
rect 156734 246534 159475 249945
rect 122960 245000 130971 245011
rect 156734 245000 159623 246534
rect 227159 245000 228235 245043
rect 9000 243072 228235 245000
rect 9000 243000 226843 243072
rect 16926 242759 17233 243000
rect 26157 242759 27614 243000
rect 122960 242990 130971 243000
rect 156655 241296 159623 243000
rect 156596 239900 159623 241296
rect 156763 239446 159623 239900
rect 227159 239767 228235 243072
rect 156763 234883 159475 239446
rect 227159 238586 234587 239767
rect 156704 234394 159475 234883
rect 156704 233567 159471 234394
rect 157052 233402 159471 233567
rect 157052 230638 159393 233402
rect 156887 230093 159393 230638
rect 156887 229679 159394 230093
rect 156858 227000 159445 229679
rect 69559 225000 226544 227000
rect 157052 224776 159393 225000
rect 156867 223817 159393 224776
rect 156838 221025 159425 223817
rect 157052 213295 159393 221025
rect 156907 212168 159393 213295
rect 156907 211754 159414 212168
rect 156878 205038 159465 211754
rect 156799 203105 159465 205038
rect 156740 202843 159465 203105
rect 156740 201709 159393 202843
rect 156907 196692 159393 201709
rect 156848 194275 159393 196692
rect 156848 193861 159401 194275
rect 156848 193531 159452 193861
rect 156865 187145 159452 193531
rect 156786 185212 159452 187145
rect 156727 184950 159452 185212
rect 156727 183816 159393 184950
rect 53308 181650 61449 181788
rect 9572 179580 61449 181650
rect 11699 178165 12054 179580
rect 59103 176959 61380 179580
rect 156894 178799 159393 183816
rect 156835 177000 159393 178799
rect 65177 176959 277000 177000
rect 59103 175000 277000 176959
rect 59103 174889 70417 175000
rect 156688 174818 159393 175000
rect 156609 172885 159393 174818
rect 156550 171489 159393 172885
rect 156717 166472 159393 171489
rect 156658 164985 159393 166472
rect 157052 160826 159393 164985
rect 156835 158070 159825 160826
rect 157052 155993 159393 158070
rect 157052 153237 160110 155993
rect 157052 150733 159393 153237
rect 157052 147977 160181 150733
rect 157052 145259 159393 147977
rect 157052 142503 160110 145259
rect 157052 139147 159393 142503
rect 157052 136391 160252 139147
rect 157052 135000 159393 136391
rect 198378 135000 215898 135038
rect 11000 133000 215898 135000
rect 21168 120516 22352 133000
rect 157052 131451 159393 133000
rect 198378 132984 215898 133000
rect 157052 128209 160042 131451
rect 215060 131248 215306 132984
rect 157052 128188 160040 128209
rect 21057 117981 22422 120516
rect 15740 116741 22422 117981
rect 15740 107632 16148 116741
rect 21057 116705 22422 116741
rect 157052 120197 159393 128188
rect 157052 116893 159559 120197
rect 157052 116868 159557 116893
rect 157052 112245 159393 116868
rect 157052 108941 159764 112245
rect 157052 108916 159762 108941
rect 157052 104019 159393 108916
rect 157052 100715 159764 104019
rect 157052 100690 159762 100715
rect 157052 96615 159393 100690
rect 157052 93311 159559 96615
rect 157052 93286 159557 93311
rect 157052 89485 159393 93286
rect 156944 87552 159393 89485
rect 156885 86156 159393 87552
rect 157052 81139 159393 86156
rect 156993 79768 159393 81139
rect 156993 71584 159391 79768
rect 156918 70211 159391 71584
rect 156918 69959 159393 70211
rect 156859 68908 159393 69959
rect 157052 65344 159393 68908
rect 156883 63719 159393 65344
rect 156824 62668 159393 63719
rect 157052 59627 159393 62668
rect 156848 58002 159393 59627
rect 156789 56951 159393 58002
rect 157052 53422 159393 56951
rect 156779 51797 159393 53422
rect 156720 50746 159393 51797
rect 157052 50000 159393 50746
rect 11000 48000 176227 50000
rect 22603 47963 25872 48000
rect 157052 45727 159393 48000
rect 157036 45476 159393 45727
rect 156491 43939 159705 45476
rect 156432 43049 159705 43939
rect 157036 42901 159393 43049
rect 157052 39433 159393 42901
rect 157036 39182 159393 39433
rect 156491 37645 159705 39182
rect 156432 36755 159705 37645
rect 157036 36607 159393 36755
rect 157052 33139 159393 36607
rect 157036 32888 159393 33139
rect 156491 31351 159705 32888
rect 156432 30461 159705 31351
rect 157036 30313 159393 30461
rect 157052 24479 159393 30313
<< comment >>
rect -50 352000 292050 352050
rect -50 0 0 352000
rect 292000 0 292050 352000
rect -50 -50 292050 0
use pd_buffered  pd_buffered_0
timestamp 1647883824
transform 1 0 13603 0 1 227298
box -947 -3256 44148 4453
use pll_full_buffered2  pll_full_buffered2_0
timestamp 1647878913
transform 1 0 15639 0 1 87306
box -1629 0 44161 20437
use filter_buffered  filter_buffered_0
timestamp 1647861083
transform 1 0 23052 0 1 29678
box -1 0 44805 14450
use cp_buffered  cp_buffered_0
timestamp 1647878778
transform 1 0 13561 0 1 262981
box -1398 -3598 44144 5452
use ro_divider_buffered  ro_divider_buffered_0
timestamp 1647865947
transform 1 0 235839 0 1 234053
box -2972 -10858 43775 12276
use ro_complete_buffered  ro_complete_buffered_0
timestamp 1647861335
transform 1 0 237047 0 1 315756
box -2962 -10858 43775 10272
use div_pd_buffered  div_pd_buffered_0
timestamp 1647861335
transform 1 0 11556 0 1 170913
box -947 -3226 44148 7340
use divider_buffered  divider_buffered_0
timestamp 1647866572
transform 1 0 214902 0 1 126196
box -746 -1568 44148 5163
use pll_full_buffered1  pll_full_buffered1_1
timestamp 1647879069
transform 1 0 11977 0 1 315152
box -1061 0 44159 15955
<< labels >>
flabel metal3 s 291760 134615 292400 134671 0 FreeSans 560 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -400 190932 240 190988 0 FreeSans 560 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -400 169321 240 169377 0 FreeSans 560 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -400 147710 240 147766 0 FreeSans 560 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -400 126199 240 126255 0 FreeSans 560 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -400 62388 240 62444 0 FreeSans 560 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -400 40777 240 40833 0 FreeSans 560 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -400 19166 240 19222 0 FreeSans 560 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -400 8455 240 8511 0 FreeSans 560 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 291760 156826 292400 156882 0 FreeSans 560 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 291760 179437 292400 179493 0 FreeSans 560 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 291760 202648 292400 202704 0 FreeSans 560 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 291760 224859 292400 224915 0 FreeSans 560 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 291760 247070 292400 247126 0 FreeSans 560 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 291760 291781 292400 291837 0 FreeSans 560 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -400 255765 240 255821 0 FreeSans 560 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -400 234154 240 234210 0 FreeSans 560 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -400 212543 240 212599 0 FreeSans 560 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 291760 135206 292400 135262 0 FreeSans 560 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -400 190341 240 190397 0 FreeSans 560 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -400 168730 240 168786 0 FreeSans 560 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -400 147119 240 147175 0 FreeSans 560 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -400 125608 240 125664 0 FreeSans 560 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -400 61797 240 61853 0 FreeSans 560 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -400 40186 240 40242 0 FreeSans 560 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -400 18575 240 18631 0 FreeSans 560 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -400 7864 240 7920 0 FreeSans 560 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 291760 157417 292400 157473 0 FreeSans 560 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 291760 180028 292400 180084 0 FreeSans 560 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 291760 203239 292400 203295 0 FreeSans 560 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 291760 225450 292400 225506 0 FreeSans 560 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 291760 247661 292400 247717 0 FreeSans 560 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 291760 292372 292400 292428 0 FreeSans 560 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -400 255174 240 255230 0 FreeSans 560 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -400 233563 240 233619 0 FreeSans 560 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -400 211952 240 212008 0 FreeSans 560 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 291150 338992 292400 341492 0 FreeSans 560 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 340121 850 342621 0 FreeSans 560 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 283297 351150 285797 352400 0 FreeSans 960 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 232697 351150 235197 352400 0 FreeSans 960 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 206697 351150 209197 352400 0 FreeSans 960 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 8097 351150 10597 352400 0 FreeSans 960 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 163397 351150 164497 352400 0 FreeSans 960 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 162147 351150 163247 352400 0 FreeSans 960 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 291760 1363 292400 1419 0 FreeSans 560 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 291760 204421 292400 204477 0 FreeSans 560 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 291760 226632 292400 226688 0 FreeSans 560 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 291760 248843 292400 248899 0 FreeSans 560 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 291760 293554 292400 293610 0 FreeSans 560 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -400 253992 240 254048 0 FreeSans 560 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -400 232381 240 232437 0 FreeSans 560 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -400 210770 240 210826 0 FreeSans 560 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -400 189159 240 189215 0 FreeSans 560 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -400 167548 240 167604 0 FreeSans 560 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -400 145937 240 145993 0 FreeSans 560 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 291760 3727 292400 3783 0 FreeSans 560 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -400 124426 240 124482 0 FreeSans 560 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -400 60615 240 60671 0 FreeSans 560 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -400 39004 240 39060 0 FreeSans 560 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -400 17393 240 17449 0 FreeSans 560 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -400 6682 240 6738 0 FreeSans 560 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -400 4318 240 4374 0 FreeSans 560 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -400 1954 240 2010 0 FreeSans 560 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 291760 6091 292400 6147 0 FreeSans 560 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 291760 8455 292400 8511 0 FreeSans 560 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 291760 10819 292400 10875 0 FreeSans 560 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 291760 24048 292400 24104 0 FreeSans 560 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 291760 46377 292400 46433 0 FreeSans 560 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 291760 136388 292400 136444 0 FreeSans 560 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 291760 158599 292400 158655 0 FreeSans 560 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 291760 181210 292400 181266 0 FreeSans 560 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 291760 772 292400 828 0 FreeSans 560 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 291760 203830 292400 203886 0 FreeSans 560 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 291760 226041 292400 226097 0 FreeSans 560 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 291760 248252 292400 248308 0 FreeSans 560 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 291760 292963 292400 293019 0 FreeSans 560 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -400 254583 240 254639 0 FreeSans 560 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -400 232972 240 233028 0 FreeSans 560 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -400 211361 240 211417 0 FreeSans 560 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -400 189750 240 189806 0 FreeSans 560 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -400 168139 240 168195 0 FreeSans 560 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -400 146528 240 146584 0 FreeSans 560 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 291760 3136 292400 3192 0 FreeSans 560 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -400 125017 240 125073 0 FreeSans 560 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -400 61206 240 61262 0 FreeSans 560 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -400 39595 240 39651 0 FreeSans 560 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -400 17984 240 18040 0 FreeSans 560 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -400 7273 240 7329 0 FreeSans 560 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -400 4909 240 4965 0 FreeSans 560 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -400 2545 240 2601 0 FreeSans 560 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 291760 5500 292400 5556 0 FreeSans 560 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 291760 7864 292400 7920 0 FreeSans 560 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 291760 10228 292400 10284 0 FreeSans 560 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 291760 23457 292400 23513 0 FreeSans 560 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 291760 45786 292400 45842 0 FreeSans 560 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 291760 135797 292400 135853 0 FreeSans 560 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 291760 158008 292400 158064 0 FreeSans 560 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 291760 180619 292400 180675 0 FreeSans 560 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 291760 2545 292400 2601 0 FreeSans 560 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 291760 205603 292400 205659 0 FreeSans 560 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 291760 227814 292400 227870 0 FreeSans 560 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 291760 250025 292400 250081 0 FreeSans 560 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 291760 294736 292400 294792 0 FreeSans 560 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -400 252810 240 252866 0 FreeSans 560 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -400 231199 240 231255 0 FreeSans 560 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -400 209588 240 209644 0 FreeSans 560 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -400 187977 240 188033 0 FreeSans 560 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -400 166366 240 166422 0 FreeSans 560 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -400 144755 240 144811 0 FreeSans 560 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 291760 4909 292400 4965 0 FreeSans 560 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -400 123244 240 123300 0 FreeSans 560 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -400 59433 240 59489 0 FreeSans 560 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -400 37822 240 37878 0 FreeSans 560 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -400 16211 240 16267 0 FreeSans 560 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -400 5500 240 5556 0 FreeSans 560 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -400 3136 240 3192 0 FreeSans 560 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -400 772 240 828 0 FreeSans 560 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 291760 7273 292400 7329 0 FreeSans 560 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 291760 9637 292400 9693 0 FreeSans 560 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 291760 12001 292400 12057 0 FreeSans 560 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 291760 25230 292400 25286 0 FreeSans 560 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 291760 47559 292400 47615 0 FreeSans 560 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 291760 137570 292400 137626 0 FreeSans 560 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 291760 159781 292400 159837 0 FreeSans 560 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 291760 182392 292400 182448 0 FreeSans 560 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 291760 1954 292400 2010 0 FreeSans 560 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 291760 205012 292400 205068 0 FreeSans 560 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 291760 227223 292400 227279 0 FreeSans 560 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 291760 249434 292400 249490 0 FreeSans 560 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 291760 294145 292400 294201 0 FreeSans 560 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -400 253401 240 253457 0 FreeSans 560 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -400 231790 240 231846 0 FreeSans 560 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -400 210179 240 210235 0 FreeSans 560 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -400 188568 240 188624 0 FreeSans 560 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -400 166957 240 167013 0 FreeSans 560 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -400 145346 240 145402 0 FreeSans 560 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 291760 4318 292400 4374 0 FreeSans 560 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -400 123835 240 123891 0 FreeSans 560 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -400 60024 240 60080 0 FreeSans 560 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -400 38413 240 38469 0 FreeSans 560 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -400 16802 240 16858 0 FreeSans 560 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -400 6091 240 6147 0 FreeSans 560 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -400 3727 240 3783 0 FreeSans 560 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -400 1363 240 1419 0 FreeSans 560 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 291760 6682 292400 6738 0 FreeSans 560 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 291760 9046 292400 9102 0 FreeSans 560 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 291760 11410 292400 11466 0 FreeSans 560 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 291760 24639 292400 24695 0 FreeSans 560 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 291760 46968 292400 47024 0 FreeSans 560 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 291760 136979 292400 137035 0 FreeSans 560 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 291760 159190 292400 159246 0 FreeSans 560 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 291760 181801 292400 181857 0 FreeSans 560 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 62908 -400 62964 240 0 FreeSans 560 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 240208 -400 240264 240 0 FreeSans 560 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 241981 -400 242037 240 0 FreeSans 560 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 243754 -400 243810 240 0 FreeSans 560 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 245527 -400 245583 240 0 FreeSans 560 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 247300 -400 247356 240 0 FreeSans 560 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 249073 -400 249129 240 0 FreeSans 560 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 250846 -400 250902 240 0 FreeSans 560 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 252619 -400 252675 240 0 FreeSans 560 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 254392 -400 254448 240 0 FreeSans 560 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 256165 -400 256221 240 0 FreeSans 560 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 80638 -400 80694 240 0 FreeSans 560 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 257938 -400 257994 240 0 FreeSans 560 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 259711 -400 259767 240 0 FreeSans 560 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 261484 -400 261540 240 0 FreeSans 560 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 263257 -400 263313 240 0 FreeSans 560 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 265030 -400 265086 240 0 FreeSans 560 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 266803 -400 266859 240 0 FreeSans 560 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 268576 -400 268632 240 0 FreeSans 560 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 270349 -400 270405 240 0 FreeSans 560 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 272122 -400 272178 240 0 FreeSans 560 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 273895 -400 273951 240 0 FreeSans 560 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 82411 -400 82467 240 0 FreeSans 560 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 275668 -400 275724 240 0 FreeSans 560 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 277441 -400 277497 240 0 FreeSans 560 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 279214 -400 279270 240 0 FreeSans 560 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 280987 -400 281043 240 0 FreeSans 560 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 282760 -400 282816 240 0 FreeSans 560 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 284533 -400 284589 240 0 FreeSans 560 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 286306 -400 286362 240 0 FreeSans 560 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 288079 -400 288135 240 0 FreeSans 560 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 84184 -400 84240 240 0 FreeSans 560 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 85957 -400 86013 240 0 FreeSans 560 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 87730 -400 87786 240 0 FreeSans 560 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 89503 -400 89559 240 0 FreeSans 560 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 91276 -400 91332 240 0 FreeSans 560 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 93049 -400 93105 240 0 FreeSans 560 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 94822 -400 94878 240 0 FreeSans 560 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 96595 -400 96651 240 0 FreeSans 560 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 64681 -400 64737 240 0 FreeSans 560 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 98368 -400 98424 240 0 FreeSans 560 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 100141 -400 100197 240 0 FreeSans 560 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 101914 -400 101970 240 0 FreeSans 560 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 103687 -400 103743 240 0 FreeSans 560 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 105460 -400 105516 240 0 FreeSans 560 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 107233 -400 107289 240 0 FreeSans 560 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 109006 -400 109062 240 0 FreeSans 560 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 110779 -400 110835 240 0 FreeSans 560 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 112552 -400 112608 240 0 FreeSans 560 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 114325 -400 114381 240 0 FreeSans 560 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 66454 -400 66510 240 0 FreeSans 560 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 116098 -400 116154 240 0 FreeSans 560 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 117871 -400 117927 240 0 FreeSans 560 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 119644 -400 119700 240 0 FreeSans 560 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 121417 -400 121473 240 0 FreeSans 560 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 123190 -400 123246 240 0 FreeSans 560 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 124963 -400 125019 240 0 FreeSans 560 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 126736 -400 126792 240 0 FreeSans 560 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 128509 -400 128565 240 0 FreeSans 560 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 130282 -400 130338 240 0 FreeSans 560 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 132055 -400 132111 240 0 FreeSans 560 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 68227 -400 68283 240 0 FreeSans 560 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 133828 -400 133884 240 0 FreeSans 560 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 135601 -400 135657 240 0 FreeSans 560 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 137374 -400 137430 240 0 FreeSans 560 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 139147 -400 139203 240 0 FreeSans 560 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 140920 -400 140976 240 0 FreeSans 560 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 142693 -400 142749 240 0 FreeSans 560 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 144466 -400 144522 240 0 FreeSans 560 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 146239 -400 146295 240 0 FreeSans 560 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 148012 -400 148068 240 0 FreeSans 560 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 149785 -400 149841 240 0 FreeSans 560 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 70000 -400 70056 240 0 FreeSans 560 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 151558 -400 151614 240 0 FreeSans 560 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 153331 -400 153387 240 0 FreeSans 560 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 155104 -400 155160 240 0 FreeSans 560 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 156877 -400 156933 240 0 FreeSans 560 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 158650 -400 158706 240 0 FreeSans 560 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 160423 -400 160479 240 0 FreeSans 560 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 162196 -400 162252 240 0 FreeSans 560 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 163969 -400 164025 240 0 FreeSans 560 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 165742 -400 165798 240 0 FreeSans 560 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 167515 -400 167571 240 0 FreeSans 560 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 71773 -400 71829 240 0 FreeSans 560 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 169288 -400 169344 240 0 FreeSans 560 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 171061 -400 171117 240 0 FreeSans 560 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 172834 -400 172890 240 0 FreeSans 560 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 174607 -400 174663 240 0 FreeSans 560 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 176380 -400 176436 240 0 FreeSans 560 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 178153 -400 178209 240 0 FreeSans 560 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 179926 -400 179982 240 0 FreeSans 560 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 181699 -400 181755 240 0 FreeSans 560 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 183472 -400 183528 240 0 FreeSans 560 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 185245 -400 185301 240 0 FreeSans 560 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 73546 -400 73602 240 0 FreeSans 560 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 187018 -400 187074 240 0 FreeSans 560 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 188791 -400 188847 240 0 FreeSans 560 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 190564 -400 190620 240 0 FreeSans 560 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 192337 -400 192393 240 0 FreeSans 560 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 194110 -400 194166 240 0 FreeSans 560 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 195883 -400 195939 240 0 FreeSans 560 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 197656 -400 197712 240 0 FreeSans 560 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 199429 -400 199485 240 0 FreeSans 560 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 201202 -400 201258 240 0 FreeSans 560 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 202975 -400 203031 240 0 FreeSans 560 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 75319 -400 75375 240 0 FreeSans 560 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 204748 -400 204804 240 0 FreeSans 560 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 206521 -400 206577 240 0 FreeSans 560 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 208294 -400 208350 240 0 FreeSans 560 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 210067 -400 210123 240 0 FreeSans 560 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 211840 -400 211896 240 0 FreeSans 560 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 213613 -400 213669 240 0 FreeSans 560 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 215386 -400 215442 240 0 FreeSans 560 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 217159 -400 217215 240 0 FreeSans 560 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 218932 -400 218988 240 0 FreeSans 560 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 220705 -400 220761 240 0 FreeSans 560 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 77092 -400 77148 240 0 FreeSans 560 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 222478 -400 222534 240 0 FreeSans 560 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 224251 -400 224307 240 0 FreeSans 560 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 226024 -400 226080 240 0 FreeSans 560 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 227797 -400 227853 240 0 FreeSans 560 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 229570 -400 229626 240 0 FreeSans 560 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 231343 -400 231399 240 0 FreeSans 560 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 233116 -400 233172 240 0 FreeSans 560 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 234889 -400 234945 240 0 FreeSans 560 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 236662 -400 236718 240 0 FreeSans 560 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 238435 -400 238491 240 0 FreeSans 560 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 78865 -400 78921 240 0 FreeSans 560 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 63499 -400 63555 240 0 FreeSans 560 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 240799 -400 240855 240 0 FreeSans 560 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 242572 -400 242628 240 0 FreeSans 560 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 244345 -400 244401 240 0 FreeSans 560 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 246118 -400 246174 240 0 FreeSans 560 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 247891 -400 247947 240 0 FreeSans 560 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 249664 -400 249720 240 0 FreeSans 560 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 251437 -400 251493 240 0 FreeSans 560 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 253210 -400 253266 240 0 FreeSans 560 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 254983 -400 255039 240 0 FreeSans 560 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 256756 -400 256812 240 0 FreeSans 560 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 81229 -400 81285 240 0 FreeSans 560 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 258529 -400 258585 240 0 FreeSans 560 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 260302 -400 260358 240 0 FreeSans 560 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 262075 -400 262131 240 0 FreeSans 560 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 263848 -400 263904 240 0 FreeSans 560 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 265621 -400 265677 240 0 FreeSans 560 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 267394 -400 267450 240 0 FreeSans 560 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 269167 -400 269223 240 0 FreeSans 560 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 270940 -400 270996 240 0 FreeSans 560 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 272713 -400 272769 240 0 FreeSans 560 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 274486 -400 274542 240 0 FreeSans 560 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 83002 -400 83058 240 0 FreeSans 560 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 276259 -400 276315 240 0 FreeSans 560 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 278032 -400 278088 240 0 FreeSans 560 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 279805 -400 279861 240 0 FreeSans 560 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 281578 -400 281634 240 0 FreeSans 560 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 283351 -400 283407 240 0 FreeSans 560 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 285124 -400 285180 240 0 FreeSans 560 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 286897 -400 286953 240 0 FreeSans 560 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 288670 -400 288726 240 0 FreeSans 560 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 84775 -400 84831 240 0 FreeSans 560 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 86548 -400 86604 240 0 FreeSans 560 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 88321 -400 88377 240 0 FreeSans 560 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 90094 -400 90150 240 0 FreeSans 560 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 91867 -400 91923 240 0 FreeSans 560 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 93640 -400 93696 240 0 FreeSans 560 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 95413 -400 95469 240 0 FreeSans 560 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 97186 -400 97242 240 0 FreeSans 560 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 65272 -400 65328 240 0 FreeSans 560 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 98959 -400 99015 240 0 FreeSans 560 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 100732 -400 100788 240 0 FreeSans 560 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 102505 -400 102561 240 0 FreeSans 560 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 104278 -400 104334 240 0 FreeSans 560 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 106051 -400 106107 240 0 FreeSans 560 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 107824 -400 107880 240 0 FreeSans 560 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 109597 -400 109653 240 0 FreeSans 560 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 111370 -400 111426 240 0 FreeSans 560 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 113143 -400 113199 240 0 FreeSans 560 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 114916 -400 114972 240 0 FreeSans 560 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 67045 -400 67101 240 0 FreeSans 560 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 116689 -400 116745 240 0 FreeSans 560 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 118462 -400 118518 240 0 FreeSans 560 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 120235 -400 120291 240 0 FreeSans 560 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 122008 -400 122064 240 0 FreeSans 560 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 123781 -400 123837 240 0 FreeSans 560 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 125554 -400 125610 240 0 FreeSans 560 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 127327 -400 127383 240 0 FreeSans 560 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 129100 -400 129156 240 0 FreeSans 560 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 130873 -400 130929 240 0 FreeSans 560 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 132646 -400 132702 240 0 FreeSans 560 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 68818 -400 68874 240 0 FreeSans 560 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 134419 -400 134475 240 0 FreeSans 560 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 136192 -400 136248 240 0 FreeSans 560 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 137965 -400 138021 240 0 FreeSans 560 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 139738 -400 139794 240 0 FreeSans 560 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 141511 -400 141567 240 0 FreeSans 560 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 143284 -400 143340 240 0 FreeSans 560 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 145057 -400 145113 240 0 FreeSans 560 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 146830 -400 146886 240 0 FreeSans 560 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 148603 -400 148659 240 0 FreeSans 560 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 150376 -400 150432 240 0 FreeSans 560 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 70591 -400 70647 240 0 FreeSans 560 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 152149 -400 152205 240 0 FreeSans 560 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 153922 -400 153978 240 0 FreeSans 560 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 155695 -400 155751 240 0 FreeSans 560 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 157468 -400 157524 240 0 FreeSans 560 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 159241 -400 159297 240 0 FreeSans 560 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 161014 -400 161070 240 0 FreeSans 560 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 162787 -400 162843 240 0 FreeSans 560 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 164560 -400 164616 240 0 FreeSans 560 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 166333 -400 166389 240 0 FreeSans 560 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 168106 -400 168162 240 0 FreeSans 560 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 72364 -400 72420 240 0 FreeSans 560 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 169879 -400 169935 240 0 FreeSans 560 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 171652 -400 171708 240 0 FreeSans 560 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 173425 -400 173481 240 0 FreeSans 560 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 175198 -400 175254 240 0 FreeSans 560 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 176971 -400 177027 240 0 FreeSans 560 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 178744 -400 178800 240 0 FreeSans 560 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 180517 -400 180573 240 0 FreeSans 560 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 182290 -400 182346 240 0 FreeSans 560 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 184063 -400 184119 240 0 FreeSans 560 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 185836 -400 185892 240 0 FreeSans 560 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 74137 -400 74193 240 0 FreeSans 560 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 187609 -400 187665 240 0 FreeSans 560 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 189382 -400 189438 240 0 FreeSans 560 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 191155 -400 191211 240 0 FreeSans 560 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 192928 -400 192984 240 0 FreeSans 560 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 194701 -400 194757 240 0 FreeSans 560 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 196474 -400 196530 240 0 FreeSans 560 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 198247 -400 198303 240 0 FreeSans 560 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 200020 -400 200076 240 0 FreeSans 560 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 201793 -400 201849 240 0 FreeSans 560 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 203566 -400 203622 240 0 FreeSans 560 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 75910 -400 75966 240 0 FreeSans 560 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 205339 -400 205395 240 0 FreeSans 560 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 207112 -400 207168 240 0 FreeSans 560 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 208885 -400 208941 240 0 FreeSans 560 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 210658 -400 210714 240 0 FreeSans 560 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 212431 -400 212487 240 0 FreeSans 560 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 214204 -400 214260 240 0 FreeSans 560 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 215977 -400 216033 240 0 FreeSans 560 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 217750 -400 217806 240 0 FreeSans 560 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 219523 -400 219579 240 0 FreeSans 560 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 221296 -400 221352 240 0 FreeSans 560 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 77683 -400 77739 240 0 FreeSans 560 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 223069 -400 223125 240 0 FreeSans 560 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 224842 -400 224898 240 0 FreeSans 560 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 226615 -400 226671 240 0 FreeSans 560 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 228388 -400 228444 240 0 FreeSans 560 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 230161 -400 230217 240 0 FreeSans 560 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 231934 -400 231990 240 0 FreeSans 560 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 233707 -400 233763 240 0 FreeSans 560 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 235480 -400 235536 240 0 FreeSans 560 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 237253 -400 237309 240 0 FreeSans 560 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 239026 -400 239082 240 0 FreeSans 560 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 79456 -400 79512 240 0 FreeSans 560 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 64090 -400 64146 240 0 FreeSans 560 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 241390 -400 241446 240 0 FreeSans 560 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 243163 -400 243219 240 0 FreeSans 560 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 244936 -400 244992 240 0 FreeSans 560 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 246709 -400 246765 240 0 FreeSans 560 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 248482 -400 248538 240 0 FreeSans 560 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 250255 -400 250311 240 0 FreeSans 560 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 252028 -400 252084 240 0 FreeSans 560 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 253801 -400 253857 240 0 FreeSans 560 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 255574 -400 255630 240 0 FreeSans 560 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 257347 -400 257403 240 0 FreeSans 560 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 81820 -400 81876 240 0 FreeSans 560 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 259120 -400 259176 240 0 FreeSans 560 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 260893 -400 260949 240 0 FreeSans 560 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 262666 -400 262722 240 0 FreeSans 560 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 264439 -400 264495 240 0 FreeSans 560 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 266212 -400 266268 240 0 FreeSans 560 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 267985 -400 268041 240 0 FreeSans 560 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 269758 -400 269814 240 0 FreeSans 560 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 271531 -400 271587 240 0 FreeSans 560 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 273304 -400 273360 240 0 FreeSans 560 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 275077 -400 275133 240 0 FreeSans 560 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 83593 -400 83649 240 0 FreeSans 560 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 276850 -400 276906 240 0 FreeSans 560 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 278623 -400 278679 240 0 FreeSans 560 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 280396 -400 280452 240 0 FreeSans 560 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 282169 -400 282225 240 0 FreeSans 560 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 283942 -400 283998 240 0 FreeSans 560 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 285715 -400 285771 240 0 FreeSans 560 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 287488 -400 287544 240 0 FreeSans 560 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 289261 -400 289317 240 0 FreeSans 560 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 85366 -400 85422 240 0 FreeSans 560 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 87139 -400 87195 240 0 FreeSans 560 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 88912 -400 88968 240 0 FreeSans 560 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 90685 -400 90741 240 0 FreeSans 560 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 92458 -400 92514 240 0 FreeSans 560 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 94231 -400 94287 240 0 FreeSans 560 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 96004 -400 96060 240 0 FreeSans 560 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 97777 -400 97833 240 0 FreeSans 560 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 65863 -400 65919 240 0 FreeSans 560 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 99550 -400 99606 240 0 FreeSans 560 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 101323 -400 101379 240 0 FreeSans 560 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 103096 -400 103152 240 0 FreeSans 560 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 104869 -400 104925 240 0 FreeSans 560 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 106642 -400 106698 240 0 FreeSans 560 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 108415 -400 108471 240 0 FreeSans 560 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 110188 -400 110244 240 0 FreeSans 560 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 111961 -400 112017 240 0 FreeSans 560 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 113734 -400 113790 240 0 FreeSans 560 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 115507 -400 115563 240 0 FreeSans 560 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 67636 -400 67692 240 0 FreeSans 560 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 117280 -400 117336 240 0 FreeSans 560 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 119053 -400 119109 240 0 FreeSans 560 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 120826 -400 120882 240 0 FreeSans 560 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 122599 -400 122655 240 0 FreeSans 560 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 124372 -400 124428 240 0 FreeSans 560 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 126145 -400 126201 240 0 FreeSans 560 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 127918 -400 127974 240 0 FreeSans 560 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 129691 -400 129747 240 0 FreeSans 560 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 131464 -400 131520 240 0 FreeSans 560 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 133237 -400 133293 240 0 FreeSans 560 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 69409 -400 69465 240 0 FreeSans 560 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 135010 -400 135066 240 0 FreeSans 560 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 136783 -400 136839 240 0 FreeSans 560 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 138556 -400 138612 240 0 FreeSans 560 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 140329 -400 140385 240 0 FreeSans 560 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 142102 -400 142158 240 0 FreeSans 560 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 143875 -400 143931 240 0 FreeSans 560 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 145648 -400 145704 240 0 FreeSans 560 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 147421 -400 147477 240 0 FreeSans 560 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 149194 -400 149250 240 0 FreeSans 560 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 150967 -400 151023 240 0 FreeSans 560 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 71182 -400 71238 240 0 FreeSans 560 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 152740 -400 152796 240 0 FreeSans 560 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 154513 -400 154569 240 0 FreeSans 560 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 156286 -400 156342 240 0 FreeSans 560 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 158059 -400 158115 240 0 FreeSans 560 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 159832 -400 159888 240 0 FreeSans 560 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 161605 -400 161661 240 0 FreeSans 560 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 163378 -400 163434 240 0 FreeSans 560 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 165151 -400 165207 240 0 FreeSans 560 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 166924 -400 166980 240 0 FreeSans 560 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 168697 -400 168753 240 0 FreeSans 560 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 72955 -400 73011 240 0 FreeSans 560 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 170470 -400 170526 240 0 FreeSans 560 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 172243 -400 172299 240 0 FreeSans 560 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 174016 -400 174072 240 0 FreeSans 560 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 175789 -400 175845 240 0 FreeSans 560 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 177562 -400 177618 240 0 FreeSans 560 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 179335 -400 179391 240 0 FreeSans 560 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 181108 -400 181164 240 0 FreeSans 560 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 182881 -400 182937 240 0 FreeSans 560 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 184654 -400 184710 240 0 FreeSans 560 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 186427 -400 186483 240 0 FreeSans 560 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 74728 -400 74784 240 0 FreeSans 560 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 188200 -400 188256 240 0 FreeSans 560 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 189973 -400 190029 240 0 FreeSans 560 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 191746 -400 191802 240 0 FreeSans 560 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 193519 -400 193575 240 0 FreeSans 560 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 195292 -400 195348 240 0 FreeSans 560 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 197065 -400 197121 240 0 FreeSans 560 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 198838 -400 198894 240 0 FreeSans 560 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 200611 -400 200667 240 0 FreeSans 560 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 202384 -400 202440 240 0 FreeSans 560 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 204157 -400 204213 240 0 FreeSans 560 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 76501 -400 76557 240 0 FreeSans 560 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 205930 -400 205986 240 0 FreeSans 560 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 207703 -400 207759 240 0 FreeSans 560 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 209476 -400 209532 240 0 FreeSans 560 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 211249 -400 211305 240 0 FreeSans 560 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 213022 -400 213078 240 0 FreeSans 560 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 214795 -400 214851 240 0 FreeSans 560 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 216568 -400 216624 240 0 FreeSans 560 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 218341 -400 218397 240 0 FreeSans 560 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 220114 -400 220170 240 0 FreeSans 560 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 221887 -400 221943 240 0 FreeSans 560 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 78274 -400 78330 240 0 FreeSans 560 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 223660 -400 223716 240 0 FreeSans 560 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 225433 -400 225489 240 0 FreeSans 560 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 227206 -400 227262 240 0 FreeSans 560 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 228979 -400 229035 240 0 FreeSans 560 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 230752 -400 230808 240 0 FreeSans 560 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 232525 -400 232581 240 0 FreeSans 560 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 234298 -400 234354 240 0 FreeSans 560 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 236071 -400 236127 240 0 FreeSans 560 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 237844 -400 237900 240 0 FreeSans 560 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 239617 -400 239673 240 0 FreeSans 560 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 80047 -400 80103 240 0 FreeSans 560 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 289852 -400 289908 240 0 FreeSans 560 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 290443 -400 290499 240 0 FreeSans 560 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 291034 -400 291090 240 0 FreeSans 560 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 291625 -400 291681 240 0 FreeSans 560 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 291170 319892 292400 322292 0 FreeSans 560 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 291170 314892 292400 317292 0 FreeSans 560 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 321921 830 324321 0 FreeSans 560 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 316921 830 319321 0 FreeSans 560 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 291170 270281 292400 272681 0 FreeSans 560 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 291170 275281 292400 277681 0 FreeSans 560 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 291170 117615 292400 120015 0 FreeSans 560 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 291170 112615 292400 115015 0 FreeSans 560 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 102444 830 104844 0 FreeSans 560 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 107444 830 109844 0 FreeSans 560 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 260297 351170 262697 352400 0 FreeSans 960 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 255297 351170 257697 352400 0 FreeSans 960 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 291170 73415 292400 75815 0 FreeSans 560 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 291170 68415 292400 70815 0 FreeSans 560 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 279721 830 282121 0 FreeSans 560 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 274721 830 277121 0 FreeSans 560 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 291170 95715 292400 98115 0 FreeSans 560 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 291170 90715 292400 93115 0 FreeSans 560 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 86444 830 88844 0 FreeSans 560 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 81444 830 83844 0 FreeSans 560 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 262 -400 318 240 0 FreeSans 560 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 853 -400 909 240 0 FreeSans 560 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 1444 -400 1500 240 0 FreeSans 560 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 3808 -400 3864 240 0 FreeSans 560 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 23902 -400 23958 240 0 FreeSans 560 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 25675 -400 25731 240 0 FreeSans 560 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 27448 -400 27504 240 0 FreeSans 560 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 29221 -400 29277 240 0 FreeSans 560 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 30994 -400 31050 240 0 FreeSans 560 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 32767 -400 32823 240 0 FreeSans 560 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 34540 -400 34596 240 0 FreeSans 560 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 36313 -400 36369 240 0 FreeSans 560 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 38086 -400 38142 240 0 FreeSans 560 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 39859 -400 39915 240 0 FreeSans 560 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 6172 -400 6228 240 0 FreeSans 560 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 41632 -400 41688 240 0 FreeSans 560 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 43405 -400 43461 240 0 FreeSans 560 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 45178 -400 45234 240 0 FreeSans 560 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 46951 -400 47007 240 0 FreeSans 560 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 48724 -400 48780 240 0 FreeSans 560 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 50497 -400 50553 240 0 FreeSans 560 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 52270 -400 52326 240 0 FreeSans 560 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 54043 -400 54099 240 0 FreeSans 560 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 55816 -400 55872 240 0 FreeSans 560 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 57589 -400 57645 240 0 FreeSans 560 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 8536 -400 8592 240 0 FreeSans 560 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 59362 -400 59418 240 0 FreeSans 560 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 61135 -400 61191 240 0 FreeSans 560 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 10900 -400 10956 240 0 FreeSans 560 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 13264 -400 13320 240 0 FreeSans 560 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 15037 -400 15093 240 0 FreeSans 560 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 16810 -400 16866 240 0 FreeSans 560 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 18583 -400 18639 240 0 FreeSans 560 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 20356 -400 20412 240 0 FreeSans 560 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 22129 -400 22185 240 0 FreeSans 560 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 2035 -400 2091 240 0 FreeSans 560 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 4399 -400 4455 240 0 FreeSans 560 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 24493 -400 24549 240 0 FreeSans 560 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 26266 -400 26322 240 0 FreeSans 560 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 28039 -400 28095 240 0 FreeSans 560 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 29812 -400 29868 240 0 FreeSans 560 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 31585 -400 31641 240 0 FreeSans 560 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 33358 -400 33414 240 0 FreeSans 560 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 35131 -400 35187 240 0 FreeSans 560 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 36904 -400 36960 240 0 FreeSans 560 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 38677 -400 38733 240 0 FreeSans 560 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 40450 -400 40506 240 0 FreeSans 560 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 6763 -400 6819 240 0 FreeSans 560 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 42223 -400 42279 240 0 FreeSans 560 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 43996 -400 44052 240 0 FreeSans 560 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 45769 -400 45825 240 0 FreeSans 560 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 47542 -400 47598 240 0 FreeSans 560 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 49315 -400 49371 240 0 FreeSans 560 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 51088 -400 51144 240 0 FreeSans 560 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 52861 -400 52917 240 0 FreeSans 560 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 54634 -400 54690 240 0 FreeSans 560 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 56407 -400 56463 240 0 FreeSans 560 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 58180 -400 58236 240 0 FreeSans 560 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 9127 -400 9183 240 0 FreeSans 560 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 59953 -400 60009 240 0 FreeSans 560 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 61726 -400 61782 240 0 FreeSans 560 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 11491 -400 11547 240 0 FreeSans 560 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 13855 -400 13911 240 0 FreeSans 560 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 15628 -400 15684 240 0 FreeSans 560 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 17401 -400 17457 240 0 FreeSans 560 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 19174 -400 19230 240 0 FreeSans 560 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 20947 -400 21003 240 0 FreeSans 560 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 22720 -400 22776 240 0 FreeSans 560 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 4990 -400 5046 240 0 FreeSans 560 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 25084 -400 25140 240 0 FreeSans 560 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 26857 -400 26913 240 0 FreeSans 560 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 28630 -400 28686 240 0 FreeSans 560 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 30403 -400 30459 240 0 FreeSans 560 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 32176 -400 32232 240 0 FreeSans 560 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 33949 -400 34005 240 0 FreeSans 560 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 35722 -400 35778 240 0 FreeSans 560 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 37495 -400 37551 240 0 FreeSans 560 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 39268 -400 39324 240 0 FreeSans 560 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 41041 -400 41097 240 0 FreeSans 560 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 7354 -400 7410 240 0 FreeSans 560 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 42814 -400 42870 240 0 FreeSans 560 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 44587 -400 44643 240 0 FreeSans 560 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 46360 -400 46416 240 0 FreeSans 560 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 48133 -400 48189 240 0 FreeSans 560 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 49906 -400 49962 240 0 FreeSans 560 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 51679 -400 51735 240 0 FreeSans 560 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 53452 -400 53508 240 0 FreeSans 560 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 55225 -400 55281 240 0 FreeSans 560 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 56998 -400 57054 240 0 FreeSans 560 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 58771 -400 58827 240 0 FreeSans 560 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 9718 -400 9774 240 0 FreeSans 560 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 60544 -400 60600 240 0 FreeSans 560 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 62317 -400 62373 240 0 FreeSans 560 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 12082 -400 12138 240 0 FreeSans 560 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 14446 -400 14502 240 0 FreeSans 560 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 16219 -400 16275 240 0 FreeSans 560 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 17992 -400 18048 240 0 FreeSans 560 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 19765 -400 19821 240 0 FreeSans 560 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 21538 -400 21594 240 0 FreeSans 560 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 23311 -400 23367 240 0 FreeSans 560 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 5581 -400 5637 240 0 FreeSans 560 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 7945 -400 8001 240 0 FreeSans 560 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 10309 -400 10365 240 0 FreeSans 560 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 12673 -400 12729 240 0 FreeSans 560 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 2626 -400 2682 240 0 FreeSans 560 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 3217 -400 3273 240 0 FreeSans 560 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 s 85447 351150 86547 352400 0 FreeSans 960 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 111297 351150 112397 352400 0 FreeSans 960 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 86697 351150 87797 352400 0 FreeSans 960 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 112547 351150 113647 352400 0 FreeSans 960 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal5 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 34097 351150 36597 352400 0 FreeSans 960 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 60097 351150 62597 352400 0 FreeSans 960 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal5 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 292000 352000
<< end >>
