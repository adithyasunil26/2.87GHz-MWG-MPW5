magic
tech sky130A
timestamp 1647883824
<< locali >>
rect -458 708 70 709
rect -470 698 70 708
rect -470 594 -458 698
rect -351 594 70 698
rect -470 585 70 594
rect -470 584 -339 585
<< viali >>
rect -458 594 -351 698
<< metal1 >>
rect 2067 1141 2142 1142
rect 1676 1116 2142 1141
rect 1666 981 1768 997
rect -470 698 -339 708
rect -470 594 -458 698
rect -351 594 -339 698
rect 1683 622 1768 981
rect -470 584 -339 594
rect 1684 57 1765 622
rect 1685 -94 1765 57
rect 2067 7 2142 1116
rect -520 -100 1765 -94
rect -525 -169 1765 -100
rect 2065 -161 2145 7
rect -525 -188 1762 -169
rect -525 -2214 -380 -188
rect -60 -316 29 -314
rect 2062 -316 2151 -161
rect -60 -397 2151 -316
rect -60 -402 2140 -397
rect -60 -707 29 -402
rect -143 -742 50 -707
rect -143 -873 -108 -742
rect 13 -873 50 -742
rect -143 -897 50 -873
rect -542 -2240 -354 -2214
rect -542 -2364 -518 -2240
rect -384 -2364 -354 -2240
rect -542 -2385 -354 -2364
<< via1 >>
rect -458 594 -351 698
rect -108 -873 13 -742
rect -518 -2364 -384 -2240
<< metal2 >>
rect -271 3655 -120 3672
rect -271 3535 -260 3655
rect -137 3535 -120 3655
rect -271 3521 -120 3535
rect -470 698 -339 708
rect -470 594 -458 698
rect -351 594 -339 698
rect -470 584 -339 594
rect -231 344 -170 3521
rect -91 2196 22 2210
rect -91 2099 -81 2196
rect 13 2099 22 2196
rect -91 2085 22 2099
rect -65 1192 -18 2085
rect -68 1176 127 1192
rect -68 1175 48 1176
rect -65 1173 -18 1175
rect -231 322 130 344
rect -143 -742 50 -707
rect -143 -873 -108 -742
rect 13 -873 50 -742
rect -143 -897 50 -873
rect -542 -2240 -354 -2214
rect -542 -2364 -518 -2240
rect -384 -2262 -354 -2240
rect -384 -2356 56 -2262
rect -384 -2364 -354 -2356
rect -542 -2385 -354 -2364
<< via2 >>
rect -260 3535 -137 3655
rect -458 594 -351 698
rect -81 2099 13 2196
<< metal3 >>
rect -271 3655 -120 3672
rect -271 3535 -260 3655
rect -137 3535 -120 3655
rect -271 3521 -120 3535
rect -88 2196 22 2205
rect -88 2099 -81 2196
rect 13 2099 22 2196
rect -88 2093 22 2099
rect -470 698 -339 708
rect -470 594 -458 698
rect -351 594 -339 698
rect -470 584 -339 594
<< via3 >>
rect -260 3535 -137 3655
rect -81 2099 13 2196
rect -458 594 -351 698
<< metal4 >>
rect -926 3818 308 3953
rect -924 2510 -768 3818
rect -283 3655 70 3681
rect -283 3535 -260 3655
rect -137 3535 70 3655
rect -283 3519 70 3535
rect -924 2366 354 2510
rect -924 713 -768 2366
rect -91 2196 22 2210
rect -91 2099 -81 2196
rect 13 2099 22 2196
rect -91 2085 22 2099
rect 4178 1401 4456 1818
rect 1681 1257 4456 1401
rect -924 698 -329 713
rect -924 594 -458 698
rect -351 594 -329 698
rect -924 577 -329 594
rect -924 -959 -768 577
rect 4178 -594 4456 1257
rect -924 -1134 329 -959
rect -924 -2445 -768 -1134
rect -947 -2620 293 -2445
<< metal5 >>
rect 186 2938 404 3236
rect 145 -1983 363 -1667
use pd  pd_0
timestamp 1647883824
transform 1 0 215 0 1 781
box -215 -855 1685 810
use tapered_buf  tapered_buf_0
timestamp 1647818295
transform 1 0 468 0 1 2605
box -470 -910 43675 401
use tapered_buf  tapered_buf_2
timestamp 1647818295
transform 1 0 434 0 1 -881
box -470 -910 43675 401
use tapered_buf  tapered_buf_1
timestamp 1647818295
transform 1 0 473 0 1 4052
box -470 -910 43675 401
use tapered_buf  tapered_buf_3
timestamp 1647818295
transform 1 0 429 0 1 -2346
box -470 -910 43675 401
<< labels >>
rlabel space 48 2642 48 2642 1 ref
rlabel space 40 -1345 40 -1345 1 up
rlabel space 64 4082 64 4082 1 div
rlabel space -14 -2804 -14 -2804 1 down
rlabel metal4 4348 686 4348 686 1 vdd!
rlabel metal4 -852 -1043 -852 -1043 1 gnd!
<< end >>
