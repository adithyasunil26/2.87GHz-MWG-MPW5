magic
tech sky130A
magscale 1 2
timestamp 1647892433
<< locali >>
rect -336 6592 1042 6678
rect -336 6328 -312 6592
rect -48 6328 1042 6592
rect -336 6288 1042 6328
<< viali >>
rect -312 6328 -48 6592
<< metal1 >>
rect -718 27414 -200 27420
rect -718 27392 -18 27414
rect -718 27198 -238 27392
rect -30 27198 -18 27392
rect -718 27180 -18 27198
rect -718 27162 -200 27180
rect -706 11656 -512 27162
rect -706 11616 -510 11656
rect -700 8804 -510 11616
rect -366 8804 1658 8828
rect -700 8766 1658 8804
rect -700 8606 1424 8766
rect 1600 8606 1658 8766
rect -700 8552 1658 8606
rect -700 8546 -176 8552
rect -336 6592 -18 6636
rect -336 6328 -312 6592
rect -48 6328 -18 6592
rect -336 6288 -18 6328
<< via1 >>
rect -238 27198 -30 27392
rect 1424 8606 1600 8766
rect -312 6328 -48 6592
<< metal2 >>
rect -676 31268 124 31368
rect -676 31050 -624 31268
rect -392 31050 124 31268
rect -676 31012 124 31050
rect -260 27392 -18 27414
rect -260 27198 -238 27392
rect -30 27198 -18 27392
rect -260 27180 -18 27198
rect -466 24500 -224 24530
rect -466 24310 -440 24500
rect -246 24310 -224 24500
rect -466 24288 -224 24310
rect -422 22994 -268 24288
rect 4280 23388 7430 23396
rect 4280 23282 37142 23388
rect 4280 23066 4392 23282
rect 4610 23066 37142 23282
rect -426 12392 -264 22994
rect 4280 22974 37142 23066
rect 4280 22954 7430 22974
rect 36778 21168 37108 22974
rect 36780 19476 37106 21168
rect -426 12192 1480 12392
rect 1388 8766 1636 8806
rect 1388 8606 1424 8766
rect 1600 8606 1636 8766
rect 1388 8566 1636 8606
rect -336 6592 -18 6636
rect -336 6328 -312 6592
rect -48 6328 -18 6592
rect -336 6288 -18 6328
<< via2 >>
rect -624 31050 -392 31268
rect -238 27198 -30 27392
rect -440 24310 -246 24500
rect 4392 23066 4610 23282
rect -312 6328 -48 6592
<< metal3 >>
rect -1392 31268 -246 31354
rect -1392 31050 -624 31268
rect -392 31050 -246 31268
rect -1392 30980 -246 31050
rect -1386 23434 -1074 30980
rect -260 27392 -18 27414
rect -260 27198 -238 27392
rect -30 27198 -18 27392
rect -260 27180 -18 27198
rect -466 24500 -224 24530
rect -466 24310 -440 24500
rect -246 24310 -224 24500
rect -466 24288 -224 24310
rect -1386 23282 4714 23434
rect -1386 23066 4392 23282
rect 4610 23066 4714 23282
rect -1386 22868 4714 23066
rect -336 6592 -18 6636
rect -336 6328 -312 6592
rect -48 6328 -18 6592
rect -336 6288 -18 6328
<< via3 >>
rect -238 27198 -30 27392
rect -440 24310 -246 24500
rect -312 6328 -48 6592
<< metal4 >>
rect -2086 30590 576 30898
rect -2084 28058 -1694 30590
rect 4252 29396 4668 29624
rect 4224 28758 4692 29396
rect -2084 27750 594 28058
rect -2084 25186 -1694 27750
rect -278 27392 64 27420
rect -278 27198 -238 27392
rect -30 27198 64 27392
rect -278 27156 64 27198
rect 4250 25830 4666 26722
rect -2084 24878 648 25186
rect -2084 6768 -1694 24878
rect -492 24500 40 24548
rect -492 24310 -440 24500
rect -246 24310 40 24500
rect -492 24262 40 24310
rect 1644 22372 2110 23762
rect -2122 6592 128 6768
rect -2122 6328 -312 6592
rect -48 6328 128 6592
rect -2122 6228 128 6328
<< metal5 >>
rect 390 28804 858 29442
rect 402 26070 842 26528
use DIGITAL_BUFFER_v1  DIGITAL_BUFFER_v1_0
timestamp 1647892099
transform 1 0 966 0 1 31078
box -940 -1820 87350 1165
use tapered_buf  tapered_buf_0
timestamp 1647889165
transform 1 0 964 0 1 25320
box -940 -1820 87350 802
use tapered_buf  tapered_buf_1
timestamp 1647889165
transform 1 0 966 0 1 28206
box -940 -1820 87350 802
use pll_full  pll_full_0
timestamp 1647892433
transform 1 0 11586 0 1 1110
box -11588 -1110 26556 21680
<< labels >>
rlabel space 58 25402 58 25402 1 ref
rlabel space 102 28274 102 28274 1 mc2
rlabel space 114 30194 118 30194 1 vco_out
rlabel metal4 -1994 23028 -1994 23028 1 gnd!
rlabel metal4 4428 26200 4428 26200 1 vdd!
<< end >>
