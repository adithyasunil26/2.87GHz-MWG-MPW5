magic
tech sky130A
timestamp 1647885873
<< locali >>
rect -168 3296 521 3339
rect -168 3164 -156 3296
rect -24 3164 521 3296
rect -168 3144 521 3164
<< viali >>
rect -156 3164 -24 3296
<< metal1 >>
rect -359 13707 -100 13710
rect -359 13696 -9 13707
rect -359 13599 -119 13696
rect -15 13599 -9 13696
rect -359 13590 -9 13599
rect -359 13581 -100 13590
rect -353 5828 -256 13581
rect -353 5808 -255 5828
rect -350 4402 -255 5808
rect -183 4402 829 4414
rect -350 4383 829 4402
rect -350 4303 712 4383
rect 800 4303 829 4383
rect -350 4276 829 4303
rect -350 4273 -88 4276
rect -168 3296 -9 3318
rect -168 3164 -156 3296
rect -24 3164 -9 3296
rect -168 3144 -9 3164
<< via1 >>
rect -119 13599 -15 13696
rect 712 4303 800 4383
rect -156 3164 -24 3296
<< metal2 >>
rect -338 15634 62 15684
rect -338 15525 -312 15634
rect -196 15525 62 15634
rect -338 15506 62 15525
rect -130 13696 -9 13707
rect -130 13599 -119 13696
rect -15 13599 -9 13696
rect -130 13590 -9 13599
rect -233 12250 -112 12265
rect -233 12155 -220 12250
rect -123 12155 -112 12250
rect -233 12144 -112 12155
rect -211 11497 -134 12144
rect 2140 11694 3715 11698
rect 2140 11641 18571 11694
rect 2140 11533 2196 11641
rect 2305 11533 18571 11641
rect -213 6196 -132 11497
rect 2140 11487 18571 11533
rect 2140 11477 3715 11487
rect 18389 10584 18554 11487
rect 18390 9738 18553 10584
rect -213 6096 740 6196
rect 694 4383 818 4403
rect 694 4303 712 4383
rect 800 4303 818 4383
rect 694 4283 818 4303
rect -168 3296 -9 3318
rect -168 3164 -156 3296
rect -24 3164 -9 3296
rect -168 3144 -9 3164
<< via2 >>
rect -312 15525 -196 15634
rect -119 13599 -15 13696
rect -220 12155 -123 12250
rect 2196 11533 2305 11641
rect -156 3164 -24 3296
<< metal3 >>
rect -696 15634 -123 15677
rect -696 15525 -312 15634
rect -196 15525 -123 15634
rect -696 15490 -123 15525
rect -693 11717 -537 15490
rect -130 13696 -9 13707
rect -130 13599 -119 13696
rect -15 13599 -9 13696
rect -130 13590 -9 13599
rect -233 12250 -112 12265
rect -233 12155 -220 12250
rect -123 12155 -112 12250
rect -233 12144 -112 12155
rect -693 11641 2357 11717
rect -693 11533 2196 11641
rect 2305 11533 2357 11641
rect -693 11434 2357 11533
rect -168 3296 -9 3318
rect -168 3164 -156 3296
rect -24 3164 -9 3296
rect -168 3144 -9 3164
<< via3 >>
rect -119 13599 -15 13696
rect -220 12155 -123 12250
rect -156 3164 -24 3296
<< metal4 >>
rect -1043 15295 288 15449
rect -1042 14029 -847 15295
rect 2126 14698 2334 14812
rect 2112 14379 2346 14698
rect -1042 13875 297 14029
rect -1042 12593 -847 13875
rect -139 13696 32 13710
rect -139 13599 -119 13696
rect -15 13599 32 13696
rect -139 13578 32 13599
rect 2125 12915 2333 13361
rect -1042 12439 324 12593
rect -1042 3384 -847 12439
rect -246 12250 20 12274
rect -246 12155 -220 12250
rect -123 12155 20 12250
rect -246 12131 20 12155
rect 822 11186 1055 11881
rect -1061 3296 64 3384
rect -1061 3164 -156 3296
rect -24 3164 64 3296
rect -1061 3114 64 3164
<< metal5 >>
rect 195 14402 429 14721
rect 201 13035 421 13264
use tapered_buf  tapered_buf_0
timestamp 1647818295
transform 1 0 482 0 1 12660
box -470 -910 43675 401
use tapered_buf  tapered_buf_1
timestamp 1647818295
transform 1 0 483 0 1 14103
box -470 -910 43675 401
use tapered_buf  tapered_buf_2
timestamp 1647818295
transform 1 0 484 0 1 15554
box -470 -910 43675 401
use pll_full  pll_full_0
timestamp 1647879007
transform 1 0 5793 0 1 555
box -5794 -555 13278 10840
<< labels >>
rlabel space 29 12701 29 12701 1 ref
rlabel space 51 14137 51 14137 1 mc2
rlabel space 57 15097 59 15097 1 vco_out
rlabel metal4 -997 11514 -997 11514 1 gnd!
rlabel metal4 2214 13100 2214 13100 1 vdd!
<< end >>
