magic
tech sky130A
timestamp 1645397998
<< nmos >>
rect -10 0 30 720
<< ndiff >>
rect -100 700 -10 720
rect -100 650 -80 700
rect -30 650 -10 700
rect -100 595 -10 650
rect -100 545 -80 595
rect -30 545 -10 595
rect -100 490 -10 545
rect -100 440 -80 490
rect -30 440 -10 490
rect -100 385 -10 440
rect -100 335 -80 385
rect -30 335 -10 385
rect -100 280 -10 335
rect -100 230 -80 280
rect -30 230 -10 280
rect -100 175 -10 230
rect -100 125 -80 175
rect -30 125 -10 175
rect -100 70 -10 125
rect -100 20 -80 70
rect -30 20 -10 70
rect -100 0 -10 20
rect 30 700 120 720
rect 30 650 50 700
rect 100 650 120 700
rect 30 595 120 650
rect 30 545 50 595
rect 100 545 120 595
rect 30 490 120 545
rect 30 440 50 490
rect 100 440 120 490
rect 30 385 120 440
rect 30 335 50 385
rect 100 335 120 385
rect 30 280 120 335
rect 30 230 50 280
rect 100 230 120 280
rect 30 175 120 230
rect 30 125 50 175
rect 100 125 120 175
rect 30 70 120 125
rect 30 20 50 70
rect 100 20 120 70
rect 30 0 120 20
<< ndiffc >>
rect -80 650 -30 700
rect -80 545 -30 595
rect -80 440 -30 490
rect -80 335 -30 385
rect -80 230 -30 280
rect -80 125 -30 175
rect -80 20 -30 70
rect 50 650 100 700
rect 50 545 100 595
rect 50 440 100 490
rect 50 335 100 385
rect 50 230 100 280
rect 50 125 100 175
rect 50 20 100 70
<< poly >>
rect -20 790 50 800
rect -20 740 -10 790
rect 40 740 50 790
rect -20 730 50 740
rect -10 720 30 730
rect -10 -20 30 0
<< polycont >>
rect -10 740 40 790
<< locali >>
rect -20 790 50 800
rect -20 740 -10 790
rect 40 740 50 790
rect -20 730 50 740
rect -90 700 -20 710
rect -90 650 -80 700
rect -30 650 -20 700
rect -90 595 -20 650
rect -90 545 -80 595
rect -30 545 -20 595
rect -90 490 -20 545
rect -90 440 -80 490
rect -30 440 -20 490
rect -90 385 -20 440
rect -90 335 -80 385
rect -30 335 -20 385
rect -90 280 -20 335
rect -90 230 -80 280
rect -30 230 -20 280
rect -90 175 -20 230
rect -90 125 -80 175
rect -30 125 -20 175
rect -90 70 -20 125
rect -90 20 -80 70
rect -30 20 -20 70
rect -90 10 -20 20
rect 40 700 110 710
rect 40 650 50 700
rect 100 650 110 700
rect 40 595 110 650
rect 40 545 50 595
rect 100 545 110 595
rect 40 490 110 545
rect 40 440 50 490
rect 100 440 110 490
rect 40 385 110 440
rect 40 335 50 385
rect 100 335 110 385
rect 40 280 110 335
rect 40 230 50 280
rect 100 230 110 280
rect 40 175 110 230
rect 40 125 50 175
rect 100 125 110 175
rect 40 70 110 125
rect 40 20 50 70
rect 100 20 110 70
rect 40 10 110 20
<< end >>
