magic
tech sky130A
timestamp 1647784636
<< nwell >>
rect -35 85 29690 260
rect 35 -710 43675 -470
<< nmos >>
rect 275 0 290 50
rect 360 0 375 50
rect 445 0 460 50
rect 530 0 545 50
rect 810 0 825 50
rect 895 0 910 50
rect 980 0 995 50
rect 1065 0 1080 50
rect 1150 0 1165 50
rect 1235 0 1250 50
rect 1320 0 1335 50
rect 1405 0 1420 50
rect 1490 0 1505 50
rect 1575 0 1590 50
rect 1660 0 1675 50
rect 1745 0 1760 50
rect 1830 0 1845 50
rect 1915 0 1930 50
rect 2000 0 2015 50
rect 2085 0 2100 50
rect 2320 0 2335 50
rect 2405 0 2420 50
rect 2490 0 2505 50
rect 2575 0 2590 50
rect 2660 0 2675 50
rect 2745 0 2760 50
rect 2830 0 2845 50
rect 2915 0 2930 50
rect 3000 0 3015 50
rect 3085 0 3100 50
rect 3170 0 3185 50
rect 3255 0 3270 50
rect 3340 0 3355 50
rect 3425 0 3440 50
rect 3510 0 3525 50
rect 3595 0 3610 50
rect 3680 0 3695 50
rect 3765 0 3780 50
rect 3850 0 3865 50
rect 3935 0 3950 50
rect 4020 0 4035 50
rect 4105 0 4120 50
rect 4190 0 4205 50
rect 4275 0 4290 50
rect 4360 0 4375 50
rect 4445 0 4460 50
rect 4530 0 4545 50
rect 4615 0 4630 50
rect 4700 0 4715 50
rect 4785 0 4800 50
rect 4870 0 4885 50
rect 4955 0 4970 50
rect 5040 0 5055 50
rect 5125 0 5140 50
rect 5210 0 5225 50
rect 5295 0 5310 50
rect 5380 0 5395 50
rect 5465 0 5480 50
rect 5550 0 5565 50
rect 5635 0 5650 50
rect 5720 0 5735 50
rect 5805 0 5820 50
rect 5890 0 5905 50
rect 5975 0 5990 50
rect 6060 0 6075 50
rect 6145 0 6160 50
rect 6230 0 6245 50
rect 6315 0 6330 50
rect 6400 0 6415 50
rect 6485 0 6500 50
rect 6570 0 6585 50
rect 6655 0 6670 50
rect 6740 0 6755 50
rect 6825 0 6840 50
rect 6910 0 6925 50
rect 6995 0 7010 50
rect 7080 0 7095 50
rect 7165 0 7180 50
rect 7250 0 7265 50
rect 7335 0 7350 50
rect 7420 0 7435 50
rect 7505 0 7520 50
rect 7590 0 7605 50
rect 7675 0 7690 50
rect 7910 0 7925 50
rect 7995 0 8010 50
rect 8080 0 8095 50
rect 8165 0 8180 50
rect 8250 0 8265 50
rect 8335 0 8350 50
rect 8420 0 8435 50
rect 8505 0 8520 50
rect 8590 0 8605 50
rect 8675 0 8690 50
rect 8760 0 8775 50
rect 8845 0 8860 50
rect 8930 0 8945 50
rect 9015 0 9030 50
rect 9100 0 9115 50
rect 9185 0 9200 50
rect 9270 0 9285 50
rect 9355 0 9370 50
rect 9440 0 9455 50
rect 9525 0 9540 50
rect 9610 0 9625 50
rect 9695 0 9710 50
rect 9780 0 9795 50
rect 9865 0 9880 50
rect 9950 0 9965 50
rect 10035 0 10050 50
rect 10120 0 10135 50
rect 10205 0 10220 50
rect 10290 0 10305 50
rect 10375 0 10390 50
rect 10460 0 10475 50
rect 10545 0 10560 50
rect 10630 0 10645 50
rect 10715 0 10730 50
rect 10800 0 10815 50
rect 10885 0 10900 50
rect 10970 0 10985 50
rect 11055 0 11070 50
rect 11140 0 11155 50
rect 11225 0 11240 50
rect 11310 0 11325 50
rect 11395 0 11410 50
rect 11480 0 11495 50
rect 11565 0 11580 50
rect 11650 0 11665 50
rect 11735 0 11750 50
rect 11820 0 11835 50
rect 11905 0 11920 50
rect 11990 0 12005 50
rect 12075 0 12090 50
rect 12160 0 12175 50
rect 12245 0 12260 50
rect 12330 0 12345 50
rect 12415 0 12430 50
rect 12500 0 12515 50
rect 12585 0 12600 50
rect 12670 0 12685 50
rect 12755 0 12770 50
rect 12840 0 12855 50
rect 12925 0 12940 50
rect 13010 0 13025 50
rect 13095 0 13110 50
rect 13180 0 13195 50
rect 13265 0 13280 50
rect 13350 0 13365 50
rect 13435 0 13450 50
rect 13520 0 13535 50
rect 13605 0 13620 50
rect 13690 0 13705 50
rect 13775 0 13790 50
rect 13860 0 13875 50
rect 13945 0 13960 50
rect 14030 0 14045 50
rect 14115 0 14130 50
rect 14200 0 14215 50
rect 14285 0 14300 50
rect 14370 0 14385 50
rect 14455 0 14470 50
rect 14540 0 14555 50
rect 14625 0 14640 50
rect 14710 0 14725 50
rect 14795 0 14810 50
rect 14880 0 14895 50
rect 14965 0 14980 50
rect 15050 0 15065 50
rect 15135 0 15150 50
rect 15220 0 15235 50
rect 15305 0 15320 50
rect 15390 0 15405 50
rect 15475 0 15490 50
rect 15560 0 15575 50
rect 15645 0 15660 50
rect 15730 0 15745 50
rect 15815 0 15830 50
rect 15900 0 15915 50
rect 15985 0 16000 50
rect 16070 0 16085 50
rect 16155 0 16170 50
rect 16240 0 16255 50
rect 16325 0 16340 50
rect 16410 0 16425 50
rect 16495 0 16510 50
rect 16580 0 16595 50
rect 16665 0 16680 50
rect 16750 0 16765 50
rect 16835 0 16850 50
rect 16920 0 16935 50
rect 17005 0 17020 50
rect 17090 0 17105 50
rect 17175 0 17190 50
rect 17260 0 17275 50
rect 17345 0 17360 50
rect 17430 0 17445 50
rect 17515 0 17530 50
rect 17600 0 17615 50
rect 17685 0 17700 50
rect 17770 0 17785 50
rect 17855 0 17870 50
rect 17940 0 17955 50
rect 18025 0 18040 50
rect 18110 0 18125 50
rect 18195 0 18210 50
rect 18280 0 18295 50
rect 18365 0 18380 50
rect 18450 0 18465 50
rect 18535 0 18550 50
rect 18620 0 18635 50
rect 18705 0 18720 50
rect 18790 0 18805 50
rect 18875 0 18890 50
rect 18960 0 18975 50
rect 19045 0 19060 50
rect 19130 0 19145 50
rect 19215 0 19230 50
rect 19300 0 19315 50
rect 19385 0 19400 50
rect 19470 0 19485 50
rect 19555 0 19570 50
rect 19640 0 19655 50
rect 19725 0 19740 50
rect 19810 0 19825 50
rect 19895 0 19910 50
rect 19980 0 19995 50
rect 20065 0 20080 50
rect 20150 0 20165 50
rect 20235 0 20250 50
rect 20320 0 20335 50
rect 20405 0 20420 50
rect 20490 0 20505 50
rect 20575 0 20590 50
rect 20660 0 20675 50
rect 20745 0 20760 50
rect 20830 0 20845 50
rect 20915 0 20930 50
rect 21000 0 21015 50
rect 21085 0 21100 50
rect 21170 0 21185 50
rect 21255 0 21270 50
rect 21340 0 21355 50
rect 21425 0 21440 50
rect 21510 0 21525 50
rect 21595 0 21610 50
rect 21680 0 21695 50
rect 21765 0 21780 50
rect 21850 0 21865 50
rect 21935 0 21950 50
rect 22020 0 22035 50
rect 22105 0 22120 50
rect 22190 0 22205 50
rect 22275 0 22290 50
rect 22360 0 22375 50
rect 22445 0 22460 50
rect 22530 0 22545 50
rect 22615 0 22630 50
rect 22700 0 22715 50
rect 22785 0 22800 50
rect 22870 0 22885 50
rect 22955 0 22970 50
rect 23040 0 23055 50
rect 23125 0 23140 50
rect 23210 0 23225 50
rect 23295 0 23310 50
rect 23380 0 23395 50
rect 23465 0 23480 50
rect 23550 0 23565 50
rect 23635 0 23650 50
rect 23720 0 23735 50
rect 23805 0 23820 50
rect 23890 0 23905 50
rect 23975 0 23990 50
rect 24060 0 24075 50
rect 24145 0 24160 50
rect 24230 0 24245 50
rect 24315 0 24330 50
rect 24400 0 24415 50
rect 24485 0 24500 50
rect 24570 0 24585 50
rect 24655 0 24670 50
rect 24740 0 24755 50
rect 24825 0 24840 50
rect 24910 0 24925 50
rect 24995 0 25010 50
rect 25080 0 25095 50
rect 25165 0 25180 50
rect 25250 0 25265 50
rect 25335 0 25350 50
rect 25420 0 25435 50
rect 25505 0 25520 50
rect 25590 0 25605 50
rect 25675 0 25690 50
rect 25760 0 25775 50
rect 25845 0 25860 50
rect 25930 0 25945 50
rect 26015 0 26030 50
rect 26100 0 26115 50
rect 26185 0 26200 50
rect 26270 0 26285 50
rect 26355 0 26370 50
rect 26440 0 26455 50
rect 26525 0 26540 50
rect 26610 0 26625 50
rect 26695 0 26710 50
rect 26780 0 26795 50
rect 26865 0 26880 50
rect 26950 0 26965 50
rect 27035 0 27050 50
rect 27120 0 27135 50
rect 27205 0 27220 50
rect 27290 0 27305 50
rect 27375 0 27390 50
rect 27460 0 27475 50
rect 27545 0 27560 50
rect 27630 0 27645 50
rect 27715 0 27730 50
rect 27800 0 27815 50
rect 27885 0 27900 50
rect 27970 0 27985 50
rect 28055 0 28070 50
rect 28140 0 28155 50
rect 28225 0 28240 50
rect 28310 0 28325 50
rect 28395 0 28410 50
rect 28480 0 28495 50
rect 28565 0 28580 50
rect 28650 0 28665 50
rect 28735 0 28750 50
rect 28820 0 28835 50
rect 28905 0 28920 50
rect 28990 0 29005 50
rect 29075 0 29090 50
rect 29160 0 29175 50
rect 29245 0 29260 50
rect 29330 0 29345 50
rect 29415 0 29430 50
rect 29500 0 29515 50
rect 29585 0 29600 50
rect 65 -70 80 -20
rect 125 -425 140 -325
rect 210 -425 225 -325
rect 295 -425 310 -325
rect 380 -425 395 -325
rect 465 -425 480 -325
rect 550 -425 565 -325
rect 635 -425 650 -325
rect 720 -425 735 -325
rect 805 -425 820 -325
rect 890 -425 905 -325
rect 975 -425 990 -325
rect 1060 -425 1075 -325
rect 1145 -425 1160 -325
rect 1230 -425 1245 -325
rect 1315 -425 1330 -325
rect 1400 -425 1415 -325
rect 1485 -425 1500 -325
rect 1570 -425 1585 -325
rect 1655 -425 1670 -325
rect 1740 -425 1755 -325
rect 1825 -425 1840 -325
rect 1910 -425 1925 -325
rect 1995 -425 2010 -325
rect 2080 -425 2095 -325
rect 2165 -425 2180 -325
rect 2250 -425 2265 -325
rect 2335 -425 2350 -325
rect 2420 -425 2435 -325
rect 2505 -425 2520 -325
rect 2590 -425 2605 -325
rect 2675 -425 2690 -325
rect 2760 -425 2775 -325
rect 2845 -425 2860 -325
rect 2930 -425 2945 -325
rect 3015 -425 3030 -325
rect 3100 -425 3115 -325
rect 3185 -425 3200 -325
rect 3270 -425 3285 -325
rect 3355 -425 3370 -325
rect 3440 -425 3455 -325
rect 3525 -425 3540 -325
rect 3610 -425 3625 -325
rect 3695 -425 3710 -325
rect 3780 -425 3795 -325
rect 3865 -425 3880 -325
rect 3950 -425 3965 -325
rect 4035 -425 4050 -325
rect 4120 -425 4135 -325
rect 4205 -425 4220 -325
rect 4290 -425 4305 -325
rect 4375 -425 4390 -325
rect 4460 -425 4475 -325
rect 4545 -425 4560 -325
rect 4630 -425 4645 -325
rect 4715 -425 4730 -325
rect 4800 -425 4815 -325
rect 4885 -425 4900 -325
rect 4970 -425 4985 -325
rect 5055 -425 5070 -325
rect 5140 -425 5155 -325
rect 5225 -425 5240 -325
rect 5310 -425 5325 -325
rect 5395 -425 5410 -325
rect 5480 -425 5495 -325
rect 5565 -425 5580 -325
rect 5650 -425 5665 -325
rect 5735 -425 5750 -325
rect 5820 -425 5835 -325
rect 5905 -425 5920 -325
rect 5990 -425 6005 -325
rect 6075 -425 6090 -325
rect 6160 -425 6175 -325
rect 6245 -425 6260 -325
rect 6330 -425 6345 -325
rect 6415 -425 6430 -325
rect 6500 -425 6515 -325
rect 6585 -425 6600 -325
rect 6670 -425 6685 -325
rect 6755 -425 6770 -325
rect 6840 -425 6855 -325
rect 6925 -425 6940 -325
rect 7010 -425 7025 -325
rect 7095 -425 7110 -325
rect 7180 -425 7195 -325
rect 7265 -425 7280 -325
rect 7350 -425 7365 -325
rect 7435 -425 7450 -325
rect 7520 -425 7535 -325
rect 7605 -425 7620 -325
rect 7690 -425 7705 -325
rect 7775 -425 7790 -325
rect 7860 -425 7875 -325
rect 7945 -425 7960 -325
rect 8030 -425 8045 -325
rect 8115 -425 8130 -325
rect 8200 -425 8215 -325
rect 8285 -425 8300 -325
rect 8370 -425 8385 -325
rect 8455 -425 8470 -325
rect 8540 -425 8555 -325
rect 8625 -425 8640 -325
rect 8710 -425 8725 -325
rect 8795 -425 8810 -325
rect 8880 -425 8895 -325
rect 8965 -425 8980 -325
rect 9050 -425 9065 -325
rect 9135 -425 9150 -325
rect 9220 -425 9235 -325
rect 9305 -425 9320 -325
rect 9390 -425 9405 -325
rect 9475 -425 9490 -325
rect 9560 -425 9575 -325
rect 9645 -425 9660 -325
rect 9730 -425 9745 -325
rect 9815 -425 9830 -325
rect 9900 -425 9915 -325
rect 9985 -425 10000 -325
rect 10070 -425 10085 -325
rect 10155 -425 10170 -325
rect 10240 -425 10255 -325
rect 10325 -425 10340 -325
rect 10410 -425 10425 -325
rect 10495 -425 10510 -325
rect 10580 -425 10595 -325
rect 10665 -425 10680 -325
rect 10750 -425 10765 -325
rect 10835 -425 10850 -325
rect 10920 -425 10935 -325
rect 11005 -425 11020 -325
rect 11090 -425 11105 -325
rect 11175 -425 11190 -325
rect 11260 -425 11275 -325
rect 11345 -425 11360 -325
rect 11430 -425 11445 -325
rect 11515 -425 11530 -325
rect 11600 -425 11615 -325
rect 11685 -425 11700 -325
rect 11770 -425 11785 -325
rect 11855 -425 11870 -325
rect 11940 -425 11955 -325
rect 12025 -425 12040 -325
rect 12110 -425 12125 -325
rect 12195 -425 12210 -325
rect 12280 -425 12295 -325
rect 12365 -425 12380 -325
rect 12450 -425 12465 -325
rect 12535 -425 12550 -325
rect 12620 -425 12635 -325
rect 12705 -425 12720 -325
rect 12790 -425 12805 -325
rect 12875 -425 12890 -325
rect 12960 -425 12975 -325
rect 13045 -425 13060 -325
rect 13130 -425 13145 -325
rect 13215 -425 13230 -325
rect 13300 -425 13315 -325
rect 13385 -425 13400 -325
rect 13470 -425 13485 -325
rect 13555 -425 13570 -325
rect 13640 -425 13655 -325
rect 13725 -425 13740 -325
rect 13810 -425 13825 -325
rect 13895 -425 13910 -325
rect 13980 -425 13995 -325
rect 14065 -425 14080 -325
rect 14150 -425 14165 -325
rect 14235 -425 14250 -325
rect 14320 -425 14335 -325
rect 14405 -425 14420 -325
rect 14490 -425 14505 -325
rect 14575 -425 14590 -325
rect 14660 -425 14675 -325
rect 14745 -425 14760 -325
rect 14830 -425 14845 -325
rect 14915 -425 14930 -325
rect 15000 -425 15015 -325
rect 15085 -425 15100 -325
rect 15170 -425 15185 -325
rect 15255 -425 15270 -325
rect 15340 -425 15355 -325
rect 15425 -425 15440 -325
rect 15510 -425 15525 -325
rect 15595 -425 15610 -325
rect 15680 -425 15695 -325
rect 15765 -425 15780 -325
rect 15850 -425 15865 -325
rect 15935 -425 15950 -325
rect 16020 -425 16035 -325
rect 16105 -425 16120 -325
rect 16190 -425 16205 -325
rect 16275 -425 16290 -325
rect 16360 -425 16375 -325
rect 16445 -425 16460 -325
rect 16530 -425 16545 -325
rect 16615 -425 16630 -325
rect 16700 -425 16715 -325
rect 16785 -425 16800 -325
rect 16870 -425 16885 -325
rect 16955 -425 16970 -325
rect 17040 -425 17055 -325
rect 17125 -425 17140 -325
rect 17210 -425 17225 -325
rect 17295 -425 17310 -325
rect 17380 -425 17395 -325
rect 17465 -425 17480 -325
rect 17550 -425 17565 -325
rect 17635 -425 17650 -325
rect 17720 -425 17735 -325
rect 17805 -425 17820 -325
rect 17890 -425 17905 -325
rect 17975 -425 17990 -325
rect 18060 -425 18075 -325
rect 18145 -425 18160 -325
rect 18230 -425 18245 -325
rect 18315 -425 18330 -325
rect 18400 -425 18415 -325
rect 18485 -425 18500 -325
rect 18570 -425 18585 -325
rect 18655 -425 18670 -325
rect 18740 -425 18755 -325
rect 18825 -425 18840 -325
rect 18910 -425 18925 -325
rect 18995 -425 19010 -325
rect 19080 -425 19095 -325
rect 19165 -425 19180 -325
rect 19250 -425 19265 -325
rect 19335 -425 19350 -325
rect 19420 -425 19435 -325
rect 19505 -425 19520 -325
rect 19590 -425 19605 -325
rect 19675 -425 19690 -325
rect 19760 -425 19775 -325
rect 19845 -425 19860 -325
rect 19930 -425 19945 -325
rect 20015 -425 20030 -325
rect 20100 -425 20115 -325
rect 20185 -425 20200 -325
rect 20270 -425 20285 -325
rect 20355 -425 20370 -325
rect 20440 -425 20455 -325
rect 20525 -425 20540 -325
rect 20610 -425 20625 -325
rect 20695 -425 20710 -325
rect 20780 -425 20795 -325
rect 20865 -425 20880 -325
rect 20950 -425 20965 -325
rect 21035 -425 21050 -325
rect 21120 -425 21135 -325
rect 21205 -425 21220 -325
rect 21290 -425 21305 -325
rect 21375 -425 21390 -325
rect 21460 -425 21475 -325
rect 21545 -425 21560 -325
rect 21630 -425 21645 -325
rect 21715 -425 21730 -325
rect 21800 -425 21815 -325
rect 21885 -425 21900 -325
rect 21970 -425 21985 -325
rect 22055 -425 22070 -325
rect 22140 -425 22155 -325
rect 22225 -425 22240 -325
rect 22310 -425 22325 -325
rect 22395 -425 22410 -325
rect 22480 -425 22495 -325
rect 22565 -425 22580 -325
rect 22650 -425 22665 -325
rect 22735 -425 22750 -325
rect 22820 -425 22835 -325
rect 22905 -425 22920 -325
rect 22990 -425 23005 -325
rect 23075 -425 23090 -325
rect 23160 -425 23175 -325
rect 23245 -425 23260 -325
rect 23330 -425 23345 -325
rect 23415 -425 23430 -325
rect 23500 -425 23515 -325
rect 23585 -425 23600 -325
rect 23670 -425 23685 -325
rect 23755 -425 23770 -325
rect 23840 -425 23855 -325
rect 23925 -425 23940 -325
rect 24010 -425 24025 -325
rect 24095 -425 24110 -325
rect 24180 -425 24195 -325
rect 24265 -425 24280 -325
rect 24350 -425 24365 -325
rect 24435 -425 24450 -325
rect 24520 -425 24535 -325
rect 24605 -425 24620 -325
rect 24690 -425 24705 -325
rect 24775 -425 24790 -325
rect 24860 -425 24875 -325
rect 24945 -425 24960 -325
rect 25030 -425 25045 -325
rect 25115 -425 25130 -325
rect 25200 -425 25215 -325
rect 25285 -425 25300 -325
rect 25370 -425 25385 -325
rect 25455 -425 25470 -325
rect 25540 -425 25555 -325
rect 25625 -425 25640 -325
rect 25710 -425 25725 -325
rect 25795 -425 25810 -325
rect 25880 -425 25895 -325
rect 25965 -425 25980 -325
rect 26050 -425 26065 -325
rect 26135 -425 26150 -325
rect 26220 -425 26235 -325
rect 26305 -425 26320 -325
rect 26390 -425 26405 -325
rect 26475 -425 26490 -325
rect 26560 -425 26575 -325
rect 26645 -425 26660 -325
rect 26730 -425 26745 -325
rect 26815 -425 26830 -325
rect 26900 -425 26915 -325
rect 26985 -425 27000 -325
rect 27070 -425 27085 -325
rect 27155 -425 27170 -325
rect 27240 -425 27255 -325
rect 27325 -425 27340 -325
rect 27410 -425 27425 -325
rect 27495 -425 27510 -325
rect 27580 -425 27595 -325
rect 27665 -425 27680 -325
rect 27750 -425 27765 -325
rect 27835 -425 27850 -325
rect 27920 -425 27935 -325
rect 28005 -425 28020 -325
rect 28090 -425 28105 -325
rect 28175 -425 28190 -325
rect 28260 -425 28275 -325
rect 28345 -425 28360 -325
rect 28430 -425 28445 -325
rect 28515 -425 28530 -325
rect 28600 -425 28615 -325
rect 28685 -425 28700 -325
rect 28770 -425 28785 -325
rect 28855 -425 28870 -325
rect 28940 -425 28955 -325
rect 29025 -425 29040 -325
rect 29110 -425 29125 -325
rect 29195 -425 29210 -325
rect 29280 -425 29295 -325
rect 29365 -425 29380 -325
rect 29450 -425 29465 -325
rect 29535 -425 29550 -325
rect 29620 -425 29635 -325
rect 29705 -425 29720 -325
rect 29790 -425 29805 -325
rect 29875 -425 29890 -325
rect 29960 -425 29975 -325
rect 30045 -425 30060 -325
rect 30130 -425 30145 -325
rect 30215 -425 30230 -325
rect 30300 -425 30315 -325
rect 30385 -425 30400 -325
rect 30470 -425 30485 -325
rect 30555 -425 30570 -325
rect 30640 -425 30655 -325
rect 30725 -425 30740 -325
rect 30810 -425 30825 -325
rect 30895 -425 30910 -325
rect 30980 -425 30995 -325
rect 31065 -425 31080 -325
rect 31150 -425 31165 -325
rect 31235 -425 31250 -325
rect 31320 -425 31335 -325
rect 31405 -425 31420 -325
rect 31490 -425 31505 -325
rect 31575 -425 31590 -325
rect 31660 -425 31675 -325
rect 31745 -425 31760 -325
rect 31830 -425 31845 -325
rect 31915 -425 31930 -325
rect 32000 -425 32015 -325
rect 32085 -425 32100 -325
rect 32170 -425 32185 -325
rect 32255 -425 32270 -325
rect 32340 -425 32355 -325
rect 32425 -425 32440 -325
rect 32510 -425 32525 -325
rect 32595 -425 32610 -325
rect 32680 -425 32695 -325
rect 32765 -425 32780 -325
rect 32850 -425 32865 -325
rect 32935 -425 32950 -325
rect 33020 -425 33035 -325
rect 33105 -425 33120 -325
rect 33190 -425 33205 -325
rect 33275 -425 33290 -325
rect 33360 -425 33375 -325
rect 33445 -425 33460 -325
rect 33530 -425 33545 -325
rect 33615 -425 33630 -325
rect 33700 -425 33715 -325
rect 33785 -425 33800 -325
rect 33870 -425 33885 -325
rect 33955 -425 33970 -325
rect 34040 -425 34055 -325
rect 34125 -425 34140 -325
rect 34210 -425 34225 -325
rect 34295 -425 34310 -325
rect 34380 -425 34395 -325
rect 34465 -425 34480 -325
rect 34550 -425 34565 -325
rect 34635 -425 34650 -325
rect 34720 -425 34735 -325
rect 34805 -425 34820 -325
rect 34890 -425 34905 -325
rect 34975 -425 34990 -325
rect 35060 -425 35075 -325
rect 35145 -425 35160 -325
rect 35230 -425 35245 -325
rect 35315 -425 35330 -325
rect 35400 -425 35415 -325
rect 35485 -425 35500 -325
rect 35570 -425 35585 -325
rect 35655 -425 35670 -325
rect 35740 -425 35755 -325
rect 35825 -425 35840 -325
rect 35910 -425 35925 -325
rect 35995 -425 36010 -325
rect 36080 -425 36095 -325
rect 36165 -425 36180 -325
rect 36250 -425 36265 -325
rect 36335 -425 36350 -325
rect 36420 -425 36435 -325
rect 36505 -425 36520 -325
rect 36590 -425 36605 -325
rect 36675 -425 36690 -325
rect 36760 -425 36775 -325
rect 36845 -425 36860 -325
rect 36930 -425 36945 -325
rect 37015 -425 37030 -325
rect 37100 -425 37115 -325
rect 37185 -425 37200 -325
rect 37270 -425 37285 -325
rect 37355 -425 37370 -325
rect 37440 -425 37455 -325
rect 37525 -425 37540 -325
rect 37610 -425 37625 -325
rect 37695 -425 37710 -325
rect 37780 -425 37795 -325
rect 37865 -425 37880 -325
rect 37950 -425 37965 -325
rect 38035 -425 38050 -325
rect 38120 -425 38135 -325
rect 38205 -425 38220 -325
rect 38290 -425 38305 -325
rect 38375 -425 38390 -325
rect 38460 -425 38475 -325
rect 38545 -425 38560 -325
rect 38630 -425 38645 -325
rect 38715 -425 38730 -325
rect 38800 -425 38815 -325
rect 38885 -425 38900 -325
rect 38970 -425 38985 -325
rect 39055 -425 39070 -325
rect 39140 -425 39155 -325
rect 39225 -425 39240 -325
rect 39310 -425 39325 -325
rect 39395 -425 39410 -325
rect 39480 -425 39495 -325
rect 39565 -425 39580 -325
rect 39650 -425 39665 -325
rect 39735 -425 39750 -325
rect 39820 -425 39835 -325
rect 39905 -425 39920 -325
rect 39990 -425 40005 -325
rect 40075 -425 40090 -325
rect 40160 -425 40175 -325
rect 40245 -425 40260 -325
rect 40330 -425 40345 -325
rect 40415 -425 40430 -325
rect 40500 -425 40515 -325
rect 40585 -425 40600 -325
rect 40670 -425 40685 -325
rect 40755 -425 40770 -325
rect 40840 -425 40855 -325
rect 40925 -425 40940 -325
rect 41010 -425 41025 -325
rect 41095 -425 41110 -325
rect 41180 -425 41195 -325
rect 41265 -425 41280 -325
rect 41350 -425 41365 -325
rect 41435 -425 41450 -325
rect 41520 -425 41535 -325
rect 41605 -425 41620 -325
rect 41690 -425 41705 -325
rect 41775 -425 41790 -325
rect 41860 -425 41875 -325
rect 41945 -425 41960 -325
rect 42030 -425 42045 -325
rect 42115 -425 42130 -325
rect 42200 -425 42215 -325
rect 42285 -425 42300 -325
rect 42370 -425 42385 -325
rect 42455 -425 42470 -325
rect 42540 -425 42555 -325
rect 42625 -425 42640 -325
rect 42710 -425 42725 -325
rect 42795 -425 42810 -325
rect 42880 -425 42895 -325
rect 42965 -425 42980 -325
rect 43050 -425 43065 -325
rect 43135 -425 43150 -325
rect 43220 -425 43235 -325
rect 43305 -425 43320 -325
rect 43390 -425 43405 -325
rect 43475 -425 43490 -325
rect 43560 -425 43575 -325
<< pmos >>
rect 65 115 80 215
rect 275 115 290 215
rect 360 115 375 215
rect 445 115 460 215
rect 530 115 545 215
rect 810 115 825 215
rect 895 115 910 215
rect 980 115 995 215
rect 1065 115 1080 215
rect 1150 115 1165 215
rect 1235 115 1250 215
rect 1320 115 1335 215
rect 1405 115 1420 215
rect 1490 115 1505 215
rect 1575 115 1590 215
rect 1660 115 1675 215
rect 1745 115 1760 215
rect 1830 115 1845 215
rect 1915 115 1930 215
rect 2000 115 2015 215
rect 2085 115 2100 215
rect 2320 115 2335 215
rect 2405 115 2420 215
rect 2490 115 2505 215
rect 2575 115 2590 215
rect 2660 115 2675 215
rect 2745 115 2760 215
rect 2830 115 2845 215
rect 2915 115 2930 215
rect 3000 115 3015 215
rect 3085 115 3100 215
rect 3170 115 3185 215
rect 3255 115 3270 215
rect 3340 115 3355 215
rect 3425 115 3440 215
rect 3510 115 3525 215
rect 3595 115 3610 215
rect 3680 115 3695 215
rect 3765 115 3780 215
rect 3850 115 3865 215
rect 3935 115 3950 215
rect 4020 115 4035 215
rect 4105 115 4120 215
rect 4190 115 4205 215
rect 4275 115 4290 215
rect 4360 115 4375 215
rect 4445 115 4460 215
rect 4530 115 4545 215
rect 4615 115 4630 215
rect 4700 115 4715 215
rect 4785 115 4800 215
rect 4870 115 4885 215
rect 4955 115 4970 215
rect 5040 115 5055 215
rect 5125 115 5140 215
rect 5210 115 5225 215
rect 5295 115 5310 215
rect 5380 115 5395 215
rect 5465 115 5480 215
rect 5550 115 5565 215
rect 5635 115 5650 215
rect 5720 115 5735 215
rect 5805 115 5820 215
rect 5890 115 5905 215
rect 5975 115 5990 215
rect 6060 115 6075 215
rect 6145 115 6160 215
rect 6230 115 6245 215
rect 6315 115 6330 215
rect 6400 115 6415 215
rect 6485 115 6500 215
rect 6570 115 6585 215
rect 6655 115 6670 215
rect 6740 115 6755 215
rect 6825 115 6840 215
rect 6910 115 6925 215
rect 6995 115 7010 215
rect 7080 115 7095 215
rect 7165 115 7180 215
rect 7250 115 7265 215
rect 7335 115 7350 215
rect 7420 115 7435 215
rect 7505 115 7520 215
rect 7590 115 7605 215
rect 7675 115 7690 215
rect 7910 115 7925 215
rect 7995 115 8010 215
rect 8080 115 8095 215
rect 8165 115 8180 215
rect 8250 115 8265 215
rect 8335 115 8350 215
rect 8420 115 8435 215
rect 8505 115 8520 215
rect 8590 115 8605 215
rect 8675 115 8690 215
rect 8760 115 8775 215
rect 8845 115 8860 215
rect 8930 115 8945 215
rect 9015 115 9030 215
rect 9100 115 9115 215
rect 9185 115 9200 215
rect 9270 115 9285 215
rect 9355 115 9370 215
rect 9440 115 9455 215
rect 9525 115 9540 215
rect 9610 115 9625 215
rect 9695 115 9710 215
rect 9780 115 9795 215
rect 9865 115 9880 215
rect 9950 115 9965 215
rect 10035 115 10050 215
rect 10120 115 10135 215
rect 10205 115 10220 215
rect 10290 115 10305 215
rect 10375 115 10390 215
rect 10460 115 10475 215
rect 10545 115 10560 215
rect 10630 115 10645 215
rect 10715 115 10730 215
rect 10800 115 10815 215
rect 10885 115 10900 215
rect 10970 115 10985 215
rect 11055 115 11070 215
rect 11140 115 11155 215
rect 11225 115 11240 215
rect 11310 115 11325 215
rect 11395 115 11410 215
rect 11480 115 11495 215
rect 11565 115 11580 215
rect 11650 115 11665 215
rect 11735 115 11750 215
rect 11820 115 11835 215
rect 11905 115 11920 215
rect 11990 115 12005 215
rect 12075 115 12090 215
rect 12160 115 12175 215
rect 12245 115 12260 215
rect 12330 115 12345 215
rect 12415 115 12430 215
rect 12500 115 12515 215
rect 12585 115 12600 215
rect 12670 115 12685 215
rect 12755 115 12770 215
rect 12840 115 12855 215
rect 12925 115 12940 215
rect 13010 115 13025 215
rect 13095 115 13110 215
rect 13180 115 13195 215
rect 13265 115 13280 215
rect 13350 115 13365 215
rect 13435 115 13450 215
rect 13520 115 13535 215
rect 13605 115 13620 215
rect 13690 115 13705 215
rect 13775 115 13790 215
rect 13860 115 13875 215
rect 13945 115 13960 215
rect 14030 115 14045 215
rect 14115 115 14130 215
rect 14200 115 14215 215
rect 14285 115 14300 215
rect 14370 115 14385 215
rect 14455 115 14470 215
rect 14540 115 14555 215
rect 14625 115 14640 215
rect 14710 115 14725 215
rect 14795 115 14810 215
rect 14880 115 14895 215
rect 14965 115 14980 215
rect 15050 115 15065 215
rect 15135 115 15150 215
rect 15220 115 15235 215
rect 15305 115 15320 215
rect 15390 115 15405 215
rect 15475 115 15490 215
rect 15560 115 15575 215
rect 15645 115 15660 215
rect 15730 115 15745 215
rect 15815 115 15830 215
rect 15900 115 15915 215
rect 15985 115 16000 215
rect 16070 115 16085 215
rect 16155 115 16170 215
rect 16240 115 16255 215
rect 16325 115 16340 215
rect 16410 115 16425 215
rect 16495 115 16510 215
rect 16580 115 16595 215
rect 16665 115 16680 215
rect 16750 115 16765 215
rect 16835 115 16850 215
rect 16920 115 16935 215
rect 17005 115 17020 215
rect 17090 115 17105 215
rect 17175 115 17190 215
rect 17260 115 17275 215
rect 17345 115 17360 215
rect 17430 115 17445 215
rect 17515 115 17530 215
rect 17600 115 17615 215
rect 17685 115 17700 215
rect 17770 115 17785 215
rect 17855 115 17870 215
rect 17940 115 17955 215
rect 18025 115 18040 215
rect 18110 115 18125 215
rect 18195 115 18210 215
rect 18280 115 18295 215
rect 18365 115 18380 215
rect 18450 115 18465 215
rect 18535 115 18550 215
rect 18620 115 18635 215
rect 18705 115 18720 215
rect 18790 115 18805 215
rect 18875 115 18890 215
rect 18960 115 18975 215
rect 19045 115 19060 215
rect 19130 115 19145 215
rect 19215 115 19230 215
rect 19300 115 19315 215
rect 19385 115 19400 215
rect 19470 115 19485 215
rect 19555 115 19570 215
rect 19640 115 19655 215
rect 19725 115 19740 215
rect 19810 115 19825 215
rect 19895 115 19910 215
rect 19980 115 19995 215
rect 20065 115 20080 215
rect 20150 115 20165 215
rect 20235 115 20250 215
rect 20320 115 20335 215
rect 20405 115 20420 215
rect 20490 115 20505 215
rect 20575 115 20590 215
rect 20660 115 20675 215
rect 20745 115 20760 215
rect 20830 115 20845 215
rect 20915 115 20930 215
rect 21000 115 21015 215
rect 21085 115 21100 215
rect 21170 115 21185 215
rect 21255 115 21270 215
rect 21340 115 21355 215
rect 21425 115 21440 215
rect 21510 115 21525 215
rect 21595 115 21610 215
rect 21680 115 21695 215
rect 21765 115 21780 215
rect 21850 115 21865 215
rect 21935 115 21950 215
rect 22020 115 22035 215
rect 22105 115 22120 215
rect 22190 115 22205 215
rect 22275 115 22290 215
rect 22360 115 22375 215
rect 22445 115 22460 215
rect 22530 115 22545 215
rect 22615 115 22630 215
rect 22700 115 22715 215
rect 22785 115 22800 215
rect 22870 115 22885 215
rect 22955 115 22970 215
rect 23040 115 23055 215
rect 23125 115 23140 215
rect 23210 115 23225 215
rect 23295 115 23310 215
rect 23380 115 23395 215
rect 23465 115 23480 215
rect 23550 115 23565 215
rect 23635 115 23650 215
rect 23720 115 23735 215
rect 23805 115 23820 215
rect 23890 115 23905 215
rect 23975 115 23990 215
rect 24060 115 24075 215
rect 24145 115 24160 215
rect 24230 115 24245 215
rect 24315 115 24330 215
rect 24400 115 24415 215
rect 24485 115 24500 215
rect 24570 115 24585 215
rect 24655 115 24670 215
rect 24740 115 24755 215
rect 24825 115 24840 215
rect 24910 115 24925 215
rect 24995 115 25010 215
rect 25080 115 25095 215
rect 25165 115 25180 215
rect 25250 115 25265 215
rect 25335 115 25350 215
rect 25420 115 25435 215
rect 25505 115 25520 215
rect 25590 115 25605 215
rect 25675 115 25690 215
rect 25760 115 25775 215
rect 25845 115 25860 215
rect 25930 115 25945 215
rect 26015 115 26030 215
rect 26100 115 26115 215
rect 26185 115 26200 215
rect 26270 115 26285 215
rect 26355 115 26370 215
rect 26440 115 26455 215
rect 26525 115 26540 215
rect 26610 115 26625 215
rect 26695 115 26710 215
rect 26780 115 26795 215
rect 26865 115 26880 215
rect 26950 115 26965 215
rect 27035 115 27050 215
rect 27120 115 27135 215
rect 27205 115 27220 215
rect 27290 115 27305 215
rect 27375 115 27390 215
rect 27460 115 27475 215
rect 27545 115 27560 215
rect 27630 115 27645 215
rect 27715 115 27730 215
rect 27800 115 27815 215
rect 27885 115 27900 215
rect 27970 115 27985 215
rect 28055 115 28070 215
rect 28140 115 28155 215
rect 28225 115 28240 215
rect 28310 115 28325 215
rect 28395 115 28410 215
rect 28480 115 28495 215
rect 28565 115 28580 215
rect 28650 115 28665 215
rect 28735 115 28750 215
rect 28820 115 28835 215
rect 28905 115 28920 215
rect 28990 115 29005 215
rect 29075 115 29090 215
rect 29160 115 29175 215
rect 29245 115 29260 215
rect 29330 115 29345 215
rect 29415 115 29430 215
rect 29500 115 29515 215
rect 29585 115 29600 215
rect 125 -690 140 -490
rect 210 -690 225 -490
rect 295 -690 310 -490
rect 380 -690 395 -490
rect 465 -690 480 -490
rect 550 -690 565 -490
rect 635 -690 650 -490
rect 720 -690 735 -490
rect 805 -690 820 -490
rect 890 -690 905 -490
rect 975 -690 990 -490
rect 1060 -690 1075 -490
rect 1145 -690 1160 -490
rect 1230 -690 1245 -490
rect 1315 -690 1330 -490
rect 1400 -690 1415 -490
rect 1485 -690 1500 -490
rect 1570 -690 1585 -490
rect 1655 -690 1670 -490
rect 1740 -690 1755 -490
rect 1825 -690 1840 -490
rect 1910 -690 1925 -490
rect 1995 -690 2010 -490
rect 2080 -690 2095 -490
rect 2165 -690 2180 -490
rect 2250 -690 2265 -490
rect 2335 -690 2350 -490
rect 2420 -690 2435 -490
rect 2505 -690 2520 -490
rect 2590 -690 2605 -490
rect 2675 -690 2690 -490
rect 2760 -690 2775 -490
rect 2845 -690 2860 -490
rect 2930 -690 2945 -490
rect 3015 -690 3030 -490
rect 3100 -690 3115 -490
rect 3185 -690 3200 -490
rect 3270 -690 3285 -490
rect 3355 -690 3370 -490
rect 3440 -690 3455 -490
rect 3525 -690 3540 -490
rect 3610 -690 3625 -490
rect 3695 -690 3710 -490
rect 3780 -690 3795 -490
rect 3865 -690 3880 -490
rect 3950 -690 3965 -490
rect 4035 -690 4050 -490
rect 4120 -690 4135 -490
rect 4205 -690 4220 -490
rect 4290 -690 4305 -490
rect 4375 -690 4390 -490
rect 4460 -690 4475 -490
rect 4545 -690 4560 -490
rect 4630 -690 4645 -490
rect 4715 -690 4730 -490
rect 4800 -690 4815 -490
rect 4885 -690 4900 -490
rect 4970 -690 4985 -490
rect 5055 -690 5070 -490
rect 5140 -690 5155 -490
rect 5225 -690 5240 -490
rect 5310 -690 5325 -490
rect 5395 -690 5410 -490
rect 5480 -690 5495 -490
rect 5565 -690 5580 -490
rect 5650 -690 5665 -490
rect 5735 -690 5750 -490
rect 5820 -690 5835 -490
rect 5905 -690 5920 -490
rect 5990 -690 6005 -490
rect 6075 -690 6090 -490
rect 6160 -690 6175 -490
rect 6245 -690 6260 -490
rect 6330 -690 6345 -490
rect 6415 -690 6430 -490
rect 6500 -690 6515 -490
rect 6585 -690 6600 -490
rect 6670 -690 6685 -490
rect 6755 -690 6770 -490
rect 6840 -690 6855 -490
rect 6925 -690 6940 -490
rect 7010 -690 7025 -490
rect 7095 -690 7110 -490
rect 7180 -690 7195 -490
rect 7265 -690 7280 -490
rect 7350 -690 7365 -490
rect 7435 -690 7450 -490
rect 7520 -690 7535 -490
rect 7605 -690 7620 -490
rect 7690 -690 7705 -490
rect 7775 -690 7790 -490
rect 7860 -690 7875 -490
rect 7945 -690 7960 -490
rect 8030 -690 8045 -490
rect 8115 -690 8130 -490
rect 8200 -690 8215 -490
rect 8285 -690 8300 -490
rect 8370 -690 8385 -490
rect 8455 -690 8470 -490
rect 8540 -690 8555 -490
rect 8625 -690 8640 -490
rect 8710 -690 8725 -490
rect 8795 -690 8810 -490
rect 8880 -690 8895 -490
rect 8965 -690 8980 -490
rect 9050 -690 9065 -490
rect 9135 -690 9150 -490
rect 9220 -690 9235 -490
rect 9305 -690 9320 -490
rect 9390 -690 9405 -490
rect 9475 -690 9490 -490
rect 9560 -690 9575 -490
rect 9645 -690 9660 -490
rect 9730 -690 9745 -490
rect 9815 -690 9830 -490
rect 9900 -690 9915 -490
rect 9985 -690 10000 -490
rect 10070 -690 10085 -490
rect 10155 -690 10170 -490
rect 10240 -690 10255 -490
rect 10325 -690 10340 -490
rect 10410 -690 10425 -490
rect 10495 -690 10510 -490
rect 10580 -690 10595 -490
rect 10665 -690 10680 -490
rect 10750 -690 10765 -490
rect 10835 -690 10850 -490
rect 10920 -690 10935 -490
rect 11005 -690 11020 -490
rect 11090 -690 11105 -490
rect 11175 -690 11190 -490
rect 11260 -690 11275 -490
rect 11345 -690 11360 -490
rect 11430 -690 11445 -490
rect 11515 -690 11530 -490
rect 11600 -690 11615 -490
rect 11685 -690 11700 -490
rect 11770 -690 11785 -490
rect 11855 -690 11870 -490
rect 11940 -690 11955 -490
rect 12025 -690 12040 -490
rect 12110 -690 12125 -490
rect 12195 -690 12210 -490
rect 12280 -690 12295 -490
rect 12365 -690 12380 -490
rect 12450 -690 12465 -490
rect 12535 -690 12550 -490
rect 12620 -690 12635 -490
rect 12705 -690 12720 -490
rect 12790 -690 12805 -490
rect 12875 -690 12890 -490
rect 12960 -690 12975 -490
rect 13045 -690 13060 -490
rect 13130 -690 13145 -490
rect 13215 -690 13230 -490
rect 13300 -690 13315 -490
rect 13385 -690 13400 -490
rect 13470 -690 13485 -490
rect 13555 -690 13570 -490
rect 13640 -690 13655 -490
rect 13725 -690 13740 -490
rect 13810 -690 13825 -490
rect 13895 -690 13910 -490
rect 13980 -690 13995 -490
rect 14065 -690 14080 -490
rect 14150 -690 14165 -490
rect 14235 -690 14250 -490
rect 14320 -690 14335 -490
rect 14405 -690 14420 -490
rect 14490 -690 14505 -490
rect 14575 -690 14590 -490
rect 14660 -690 14675 -490
rect 14745 -690 14760 -490
rect 14830 -690 14845 -490
rect 14915 -690 14930 -490
rect 15000 -690 15015 -490
rect 15085 -690 15100 -490
rect 15170 -690 15185 -490
rect 15255 -690 15270 -490
rect 15340 -690 15355 -490
rect 15425 -690 15440 -490
rect 15510 -690 15525 -490
rect 15595 -690 15610 -490
rect 15680 -690 15695 -490
rect 15765 -690 15780 -490
rect 15850 -690 15865 -490
rect 15935 -690 15950 -490
rect 16020 -690 16035 -490
rect 16105 -690 16120 -490
rect 16190 -690 16205 -490
rect 16275 -690 16290 -490
rect 16360 -690 16375 -490
rect 16445 -690 16460 -490
rect 16530 -690 16545 -490
rect 16615 -690 16630 -490
rect 16700 -690 16715 -490
rect 16785 -690 16800 -490
rect 16870 -690 16885 -490
rect 16955 -690 16970 -490
rect 17040 -690 17055 -490
rect 17125 -690 17140 -490
rect 17210 -690 17225 -490
rect 17295 -690 17310 -490
rect 17380 -690 17395 -490
rect 17465 -690 17480 -490
rect 17550 -690 17565 -490
rect 17635 -690 17650 -490
rect 17720 -690 17735 -490
rect 17805 -690 17820 -490
rect 17890 -690 17905 -490
rect 17975 -690 17990 -490
rect 18060 -690 18075 -490
rect 18145 -690 18160 -490
rect 18230 -690 18245 -490
rect 18315 -690 18330 -490
rect 18400 -690 18415 -490
rect 18485 -690 18500 -490
rect 18570 -690 18585 -490
rect 18655 -690 18670 -490
rect 18740 -690 18755 -490
rect 18825 -690 18840 -490
rect 18910 -690 18925 -490
rect 18995 -690 19010 -490
rect 19080 -690 19095 -490
rect 19165 -690 19180 -490
rect 19250 -690 19265 -490
rect 19335 -690 19350 -490
rect 19420 -690 19435 -490
rect 19505 -690 19520 -490
rect 19590 -690 19605 -490
rect 19675 -690 19690 -490
rect 19760 -690 19775 -490
rect 19845 -690 19860 -490
rect 19930 -690 19945 -490
rect 20015 -690 20030 -490
rect 20100 -690 20115 -490
rect 20185 -690 20200 -490
rect 20270 -690 20285 -490
rect 20355 -690 20370 -490
rect 20440 -690 20455 -490
rect 20525 -690 20540 -490
rect 20610 -690 20625 -490
rect 20695 -690 20710 -490
rect 20780 -690 20795 -490
rect 20865 -690 20880 -490
rect 20950 -690 20965 -490
rect 21035 -690 21050 -490
rect 21120 -690 21135 -490
rect 21205 -690 21220 -490
rect 21290 -690 21305 -490
rect 21375 -690 21390 -490
rect 21460 -690 21475 -490
rect 21545 -690 21560 -490
rect 21630 -690 21645 -490
rect 21715 -690 21730 -490
rect 21800 -690 21815 -490
rect 21885 -690 21900 -490
rect 21970 -690 21985 -490
rect 22055 -690 22070 -490
rect 22140 -690 22155 -490
rect 22225 -690 22240 -490
rect 22310 -690 22325 -490
rect 22395 -690 22410 -490
rect 22480 -690 22495 -490
rect 22565 -690 22580 -490
rect 22650 -690 22665 -490
rect 22735 -690 22750 -490
rect 22820 -690 22835 -490
rect 22905 -690 22920 -490
rect 22990 -690 23005 -490
rect 23075 -690 23090 -490
rect 23160 -690 23175 -490
rect 23245 -690 23260 -490
rect 23330 -690 23345 -490
rect 23415 -690 23430 -490
rect 23500 -690 23515 -490
rect 23585 -690 23600 -490
rect 23670 -690 23685 -490
rect 23755 -690 23770 -490
rect 23840 -690 23855 -490
rect 23925 -690 23940 -490
rect 24010 -690 24025 -490
rect 24095 -690 24110 -490
rect 24180 -690 24195 -490
rect 24265 -690 24280 -490
rect 24350 -690 24365 -490
rect 24435 -690 24450 -490
rect 24520 -690 24535 -490
rect 24605 -690 24620 -490
rect 24690 -690 24705 -490
rect 24775 -690 24790 -490
rect 24860 -690 24875 -490
rect 24945 -690 24960 -490
rect 25030 -690 25045 -490
rect 25115 -690 25130 -490
rect 25200 -690 25215 -490
rect 25285 -690 25300 -490
rect 25370 -690 25385 -490
rect 25455 -690 25470 -490
rect 25540 -690 25555 -490
rect 25625 -690 25640 -490
rect 25710 -690 25725 -490
rect 25795 -690 25810 -490
rect 25880 -690 25895 -490
rect 25965 -690 25980 -490
rect 26050 -690 26065 -490
rect 26135 -690 26150 -490
rect 26220 -690 26235 -490
rect 26305 -690 26320 -490
rect 26390 -690 26405 -490
rect 26475 -690 26490 -490
rect 26560 -690 26575 -490
rect 26645 -690 26660 -490
rect 26730 -690 26745 -490
rect 26815 -690 26830 -490
rect 26900 -690 26915 -490
rect 26985 -690 27000 -490
rect 27070 -690 27085 -490
rect 27155 -690 27170 -490
rect 27240 -690 27255 -490
rect 27325 -690 27340 -490
rect 27410 -690 27425 -490
rect 27495 -690 27510 -490
rect 27580 -690 27595 -490
rect 27665 -690 27680 -490
rect 27750 -690 27765 -490
rect 27835 -690 27850 -490
rect 27920 -690 27935 -490
rect 28005 -690 28020 -490
rect 28090 -690 28105 -490
rect 28175 -690 28190 -490
rect 28260 -690 28275 -490
rect 28345 -690 28360 -490
rect 28430 -690 28445 -490
rect 28515 -690 28530 -490
rect 28600 -690 28615 -490
rect 28685 -690 28700 -490
rect 28770 -690 28785 -490
rect 28855 -690 28870 -490
rect 28940 -690 28955 -490
rect 29025 -690 29040 -490
rect 29110 -690 29125 -490
rect 29195 -690 29210 -490
rect 29280 -690 29295 -490
rect 29365 -690 29380 -490
rect 29450 -690 29465 -490
rect 29535 -690 29550 -490
rect 29620 -690 29635 -490
rect 29705 -690 29720 -490
rect 29790 -690 29805 -490
rect 29875 -690 29890 -490
rect 29960 -690 29975 -490
rect 30045 -690 30060 -490
rect 30130 -690 30145 -490
rect 30215 -690 30230 -490
rect 30300 -690 30315 -490
rect 30385 -690 30400 -490
rect 30470 -690 30485 -490
rect 30555 -690 30570 -490
rect 30640 -690 30655 -490
rect 30725 -690 30740 -490
rect 30810 -690 30825 -490
rect 30895 -690 30910 -490
rect 30980 -690 30995 -490
rect 31065 -690 31080 -490
rect 31150 -690 31165 -490
rect 31235 -690 31250 -490
rect 31320 -690 31335 -490
rect 31405 -690 31420 -490
rect 31490 -690 31505 -490
rect 31575 -690 31590 -490
rect 31660 -690 31675 -490
rect 31745 -690 31760 -490
rect 31830 -690 31845 -490
rect 31915 -690 31930 -490
rect 32000 -690 32015 -490
rect 32085 -690 32100 -490
rect 32170 -690 32185 -490
rect 32255 -690 32270 -490
rect 32340 -690 32355 -490
rect 32425 -690 32440 -490
rect 32510 -690 32525 -490
rect 32595 -690 32610 -490
rect 32680 -690 32695 -490
rect 32765 -690 32780 -490
rect 32850 -690 32865 -490
rect 32935 -690 32950 -490
rect 33020 -690 33035 -490
rect 33105 -690 33120 -490
rect 33190 -690 33205 -490
rect 33275 -690 33290 -490
rect 33360 -690 33375 -490
rect 33445 -690 33460 -490
rect 33530 -690 33545 -490
rect 33615 -690 33630 -490
rect 33700 -690 33715 -490
rect 33785 -690 33800 -490
rect 33870 -690 33885 -490
rect 33955 -690 33970 -490
rect 34040 -690 34055 -490
rect 34125 -690 34140 -490
rect 34210 -690 34225 -490
rect 34295 -690 34310 -490
rect 34380 -690 34395 -490
rect 34465 -690 34480 -490
rect 34550 -690 34565 -490
rect 34635 -690 34650 -490
rect 34720 -690 34735 -490
rect 34805 -690 34820 -490
rect 34890 -690 34905 -490
rect 34975 -690 34990 -490
rect 35060 -690 35075 -490
rect 35145 -690 35160 -490
rect 35230 -690 35245 -490
rect 35315 -690 35330 -490
rect 35400 -690 35415 -490
rect 35485 -690 35500 -490
rect 35570 -690 35585 -490
rect 35655 -690 35670 -490
rect 35740 -690 35755 -490
rect 35825 -690 35840 -490
rect 35910 -690 35925 -490
rect 35995 -690 36010 -490
rect 36080 -690 36095 -490
rect 36165 -690 36180 -490
rect 36250 -690 36265 -490
rect 36335 -690 36350 -490
rect 36420 -690 36435 -490
rect 36505 -690 36520 -490
rect 36590 -690 36605 -490
rect 36675 -690 36690 -490
rect 36760 -690 36775 -490
rect 36845 -690 36860 -490
rect 36930 -690 36945 -490
rect 37015 -690 37030 -490
rect 37100 -690 37115 -490
rect 37185 -690 37200 -490
rect 37270 -690 37285 -490
rect 37355 -690 37370 -490
rect 37440 -690 37455 -490
rect 37525 -690 37540 -490
rect 37610 -690 37625 -490
rect 37695 -690 37710 -490
rect 37780 -690 37795 -490
rect 37865 -690 37880 -490
rect 37950 -690 37965 -490
rect 38035 -690 38050 -490
rect 38120 -690 38135 -490
rect 38205 -690 38220 -490
rect 38290 -690 38305 -490
rect 38375 -690 38390 -490
rect 38460 -690 38475 -490
rect 38545 -690 38560 -490
rect 38630 -690 38645 -490
rect 38715 -690 38730 -490
rect 38800 -690 38815 -490
rect 38885 -690 38900 -490
rect 38970 -690 38985 -490
rect 39055 -690 39070 -490
rect 39140 -690 39155 -490
rect 39225 -690 39240 -490
rect 39310 -690 39325 -490
rect 39395 -690 39410 -490
rect 39480 -690 39495 -490
rect 39565 -690 39580 -490
rect 39650 -690 39665 -490
rect 39735 -690 39750 -490
rect 39820 -690 39835 -490
rect 39905 -690 39920 -490
rect 39990 -690 40005 -490
rect 40075 -690 40090 -490
rect 40160 -690 40175 -490
rect 40245 -690 40260 -490
rect 40330 -690 40345 -490
rect 40415 -690 40430 -490
rect 40500 -690 40515 -490
rect 40585 -690 40600 -490
rect 40670 -690 40685 -490
rect 40755 -690 40770 -490
rect 40840 -690 40855 -490
rect 40925 -690 40940 -490
rect 41010 -690 41025 -490
rect 41095 -690 41110 -490
rect 41180 -690 41195 -490
rect 41265 -690 41280 -490
rect 41350 -690 41365 -490
rect 41435 -690 41450 -490
rect 41520 -690 41535 -490
rect 41605 -690 41620 -490
rect 41690 -690 41705 -490
rect 41775 -690 41790 -490
rect 41860 -690 41875 -490
rect 41945 -690 41960 -490
rect 42030 -690 42045 -490
rect 42115 -690 42130 -490
rect 42200 -690 42215 -490
rect 42285 -690 42300 -490
rect 42370 -690 42385 -490
rect 42455 -690 42470 -490
rect 42540 -690 42555 -490
rect 42625 -690 42640 -490
rect 42710 -690 42725 -490
rect 42795 -690 42810 -490
rect 42880 -690 42895 -490
rect 42965 -690 42980 -490
rect 43050 -690 43065 -490
rect 43135 -690 43150 -490
rect 43220 -690 43235 -490
rect 43305 -690 43320 -490
rect 43390 -690 43405 -490
rect 43475 -690 43490 -490
rect 43560 -690 43575 -490
<< ndiff >>
rect 205 40 275 50
rect 205 10 225 40
rect 255 10 275 40
rect 205 0 275 10
rect 290 40 360 50
rect 290 10 310 40
rect 340 10 360 40
rect 290 0 360 10
rect 375 40 445 50
rect 375 10 395 40
rect 425 10 445 40
rect 375 0 445 10
rect 460 40 530 50
rect 460 10 480 40
rect 510 10 530 40
rect 460 0 530 10
rect 545 40 615 50
rect 545 10 565 40
rect 595 10 615 40
rect 545 0 615 10
rect 740 40 810 50
rect 740 10 760 40
rect 790 10 810 40
rect 740 0 810 10
rect 825 40 895 50
rect 825 10 845 40
rect 875 10 895 40
rect 825 0 895 10
rect 910 40 980 50
rect 910 10 930 40
rect 960 10 980 40
rect 910 0 980 10
rect 995 40 1065 50
rect 995 10 1015 40
rect 1045 10 1065 40
rect 995 0 1065 10
rect 1080 40 1150 50
rect 1080 10 1100 40
rect 1130 10 1150 40
rect 1080 0 1150 10
rect 1165 40 1235 50
rect 1165 10 1185 40
rect 1215 10 1235 40
rect 1165 0 1235 10
rect 1250 40 1320 50
rect 1250 10 1270 40
rect 1300 10 1320 40
rect 1250 0 1320 10
rect 1335 40 1405 50
rect 1335 10 1355 40
rect 1385 10 1405 40
rect 1335 0 1405 10
rect 1420 40 1490 50
rect 1420 10 1440 40
rect 1470 10 1490 40
rect 1420 0 1490 10
rect 1505 40 1575 50
rect 1505 10 1525 40
rect 1555 10 1575 40
rect 1505 0 1575 10
rect 1590 40 1660 50
rect 1590 10 1610 40
rect 1640 10 1660 40
rect 1590 0 1660 10
rect 1675 40 1745 50
rect 1675 10 1695 40
rect 1725 10 1745 40
rect 1675 0 1745 10
rect 1760 40 1830 50
rect 1760 10 1780 40
rect 1810 10 1830 40
rect 1760 0 1830 10
rect 1845 40 1915 50
rect 1845 10 1865 40
rect 1895 10 1915 40
rect 1845 0 1915 10
rect 1930 40 2000 50
rect 1930 10 1950 40
rect 1980 10 2000 40
rect 1930 0 2000 10
rect 2015 40 2085 50
rect 2015 10 2035 40
rect 2065 10 2085 40
rect 2015 0 2085 10
rect 2100 40 2170 50
rect 2100 10 2120 40
rect 2150 10 2170 40
rect 2100 0 2170 10
rect 2250 40 2320 50
rect 2250 10 2270 40
rect 2300 10 2320 40
rect 2250 0 2320 10
rect 2335 40 2405 50
rect 2335 10 2355 40
rect 2385 10 2405 40
rect 2335 0 2405 10
rect 2420 40 2490 50
rect 2420 10 2440 40
rect 2470 10 2490 40
rect 2420 0 2490 10
rect 2505 40 2575 50
rect 2505 10 2525 40
rect 2555 10 2575 40
rect 2505 0 2575 10
rect 2590 40 2660 50
rect 2590 10 2610 40
rect 2640 10 2660 40
rect 2590 0 2660 10
rect 2675 40 2745 50
rect 2675 10 2695 40
rect 2725 10 2745 40
rect 2675 0 2745 10
rect 2760 40 2830 50
rect 2760 10 2780 40
rect 2810 10 2830 40
rect 2760 0 2830 10
rect 2845 40 2915 50
rect 2845 10 2865 40
rect 2895 10 2915 40
rect 2845 0 2915 10
rect 2930 40 3000 50
rect 2930 10 2950 40
rect 2980 10 3000 40
rect 2930 0 3000 10
rect 3015 40 3085 50
rect 3015 10 3035 40
rect 3065 10 3085 40
rect 3015 0 3085 10
rect 3100 40 3170 50
rect 3100 10 3120 40
rect 3150 10 3170 40
rect 3100 0 3170 10
rect 3185 40 3255 50
rect 3185 10 3205 40
rect 3235 10 3255 40
rect 3185 0 3255 10
rect 3270 40 3340 50
rect 3270 10 3290 40
rect 3320 10 3340 40
rect 3270 0 3340 10
rect 3355 40 3425 50
rect 3355 10 3375 40
rect 3405 10 3425 40
rect 3355 0 3425 10
rect 3440 40 3510 50
rect 3440 10 3460 40
rect 3490 10 3510 40
rect 3440 0 3510 10
rect 3525 40 3595 50
rect 3525 10 3545 40
rect 3575 10 3595 40
rect 3525 0 3595 10
rect 3610 40 3680 50
rect 3610 10 3630 40
rect 3660 10 3680 40
rect 3610 0 3680 10
rect 3695 40 3765 50
rect 3695 10 3715 40
rect 3745 10 3765 40
rect 3695 0 3765 10
rect 3780 40 3850 50
rect 3780 10 3800 40
rect 3830 10 3850 40
rect 3780 0 3850 10
rect 3865 40 3935 50
rect 3865 10 3885 40
rect 3915 10 3935 40
rect 3865 0 3935 10
rect 3950 40 4020 50
rect 3950 10 3970 40
rect 4000 10 4020 40
rect 3950 0 4020 10
rect 4035 40 4105 50
rect 4035 10 4055 40
rect 4085 10 4105 40
rect 4035 0 4105 10
rect 4120 40 4190 50
rect 4120 10 4140 40
rect 4170 10 4190 40
rect 4120 0 4190 10
rect 4205 40 4275 50
rect 4205 10 4225 40
rect 4255 10 4275 40
rect 4205 0 4275 10
rect 4290 40 4360 50
rect 4290 10 4310 40
rect 4340 10 4360 40
rect 4290 0 4360 10
rect 4375 40 4445 50
rect 4375 10 4395 40
rect 4425 10 4445 40
rect 4375 0 4445 10
rect 4460 40 4530 50
rect 4460 10 4480 40
rect 4510 10 4530 40
rect 4460 0 4530 10
rect 4545 40 4615 50
rect 4545 10 4565 40
rect 4595 10 4615 40
rect 4545 0 4615 10
rect 4630 40 4700 50
rect 4630 10 4650 40
rect 4680 10 4700 40
rect 4630 0 4700 10
rect 4715 40 4785 50
rect 4715 10 4735 40
rect 4765 10 4785 40
rect 4715 0 4785 10
rect 4800 40 4870 50
rect 4800 10 4820 40
rect 4850 10 4870 40
rect 4800 0 4870 10
rect 4885 40 4955 50
rect 4885 10 4905 40
rect 4935 10 4955 40
rect 4885 0 4955 10
rect 4970 40 5040 50
rect 4970 10 4990 40
rect 5020 10 5040 40
rect 4970 0 5040 10
rect 5055 40 5125 50
rect 5055 10 5075 40
rect 5105 10 5125 40
rect 5055 0 5125 10
rect 5140 40 5210 50
rect 5140 10 5160 40
rect 5190 10 5210 40
rect 5140 0 5210 10
rect 5225 40 5295 50
rect 5225 10 5245 40
rect 5275 10 5295 40
rect 5225 0 5295 10
rect 5310 40 5380 50
rect 5310 10 5330 40
rect 5360 10 5380 40
rect 5310 0 5380 10
rect 5395 40 5465 50
rect 5395 10 5415 40
rect 5445 10 5465 40
rect 5395 0 5465 10
rect 5480 40 5550 50
rect 5480 10 5500 40
rect 5530 10 5550 40
rect 5480 0 5550 10
rect 5565 40 5635 50
rect 5565 10 5585 40
rect 5615 10 5635 40
rect 5565 0 5635 10
rect 5650 40 5720 50
rect 5650 10 5670 40
rect 5700 10 5720 40
rect 5650 0 5720 10
rect 5735 40 5805 50
rect 5735 10 5755 40
rect 5785 10 5805 40
rect 5735 0 5805 10
rect 5820 40 5890 50
rect 5820 10 5840 40
rect 5870 10 5890 40
rect 5820 0 5890 10
rect 5905 40 5975 50
rect 5905 10 5925 40
rect 5955 10 5975 40
rect 5905 0 5975 10
rect 5990 40 6060 50
rect 5990 10 6010 40
rect 6040 10 6060 40
rect 5990 0 6060 10
rect 6075 40 6145 50
rect 6075 10 6095 40
rect 6125 10 6145 40
rect 6075 0 6145 10
rect 6160 40 6230 50
rect 6160 10 6180 40
rect 6210 10 6230 40
rect 6160 0 6230 10
rect 6245 40 6315 50
rect 6245 10 6265 40
rect 6295 10 6315 40
rect 6245 0 6315 10
rect 6330 40 6400 50
rect 6330 10 6350 40
rect 6380 10 6400 40
rect 6330 0 6400 10
rect 6415 40 6485 50
rect 6415 10 6435 40
rect 6465 10 6485 40
rect 6415 0 6485 10
rect 6500 40 6570 50
rect 6500 10 6520 40
rect 6550 10 6570 40
rect 6500 0 6570 10
rect 6585 40 6655 50
rect 6585 10 6605 40
rect 6635 10 6655 40
rect 6585 0 6655 10
rect 6670 40 6740 50
rect 6670 10 6690 40
rect 6720 10 6740 40
rect 6670 0 6740 10
rect 6755 40 6825 50
rect 6755 10 6775 40
rect 6805 10 6825 40
rect 6755 0 6825 10
rect 6840 40 6910 50
rect 6840 10 6860 40
rect 6890 10 6910 40
rect 6840 0 6910 10
rect 6925 40 6995 50
rect 6925 10 6945 40
rect 6975 10 6995 40
rect 6925 0 6995 10
rect 7010 40 7080 50
rect 7010 10 7030 40
rect 7060 10 7080 40
rect 7010 0 7080 10
rect 7095 40 7165 50
rect 7095 10 7115 40
rect 7145 10 7165 40
rect 7095 0 7165 10
rect 7180 40 7250 50
rect 7180 10 7200 40
rect 7230 10 7250 40
rect 7180 0 7250 10
rect 7265 40 7335 50
rect 7265 10 7285 40
rect 7315 10 7335 40
rect 7265 0 7335 10
rect 7350 40 7420 50
rect 7350 10 7370 40
rect 7400 10 7420 40
rect 7350 0 7420 10
rect 7435 40 7505 50
rect 7435 10 7455 40
rect 7485 10 7505 40
rect 7435 0 7505 10
rect 7520 40 7590 50
rect 7520 10 7540 40
rect 7570 10 7590 40
rect 7520 0 7590 10
rect 7605 40 7675 50
rect 7605 10 7625 40
rect 7655 10 7675 40
rect 7605 0 7675 10
rect 7690 40 7760 50
rect 7690 10 7710 40
rect 7740 10 7760 40
rect 7690 0 7760 10
rect 7840 40 7910 50
rect 7840 10 7860 40
rect 7890 10 7910 40
rect 7840 0 7910 10
rect 7925 40 7995 50
rect 7925 10 7945 40
rect 7975 10 7995 40
rect 7925 0 7995 10
rect 8010 40 8080 50
rect 8010 10 8030 40
rect 8060 10 8080 40
rect 8010 0 8080 10
rect 8095 40 8165 50
rect 8095 10 8115 40
rect 8145 10 8165 40
rect 8095 0 8165 10
rect 8180 40 8250 50
rect 8180 10 8200 40
rect 8230 10 8250 40
rect 8180 0 8250 10
rect 8265 40 8335 50
rect 8265 10 8285 40
rect 8315 10 8335 40
rect 8265 0 8335 10
rect 8350 40 8420 50
rect 8350 10 8370 40
rect 8400 10 8420 40
rect 8350 0 8420 10
rect 8435 40 8505 50
rect 8435 10 8455 40
rect 8485 10 8505 40
rect 8435 0 8505 10
rect 8520 40 8590 50
rect 8520 10 8540 40
rect 8570 10 8590 40
rect 8520 0 8590 10
rect 8605 40 8675 50
rect 8605 10 8625 40
rect 8655 10 8675 40
rect 8605 0 8675 10
rect 8690 40 8760 50
rect 8690 10 8710 40
rect 8740 10 8760 40
rect 8690 0 8760 10
rect 8775 40 8845 50
rect 8775 10 8795 40
rect 8825 10 8845 40
rect 8775 0 8845 10
rect 8860 40 8930 50
rect 8860 10 8880 40
rect 8910 10 8930 40
rect 8860 0 8930 10
rect 8945 40 9015 50
rect 8945 10 8965 40
rect 8995 10 9015 40
rect 8945 0 9015 10
rect 9030 40 9100 50
rect 9030 10 9050 40
rect 9080 10 9100 40
rect 9030 0 9100 10
rect 9115 40 9185 50
rect 9115 10 9135 40
rect 9165 10 9185 40
rect 9115 0 9185 10
rect 9200 40 9270 50
rect 9200 10 9220 40
rect 9250 10 9270 40
rect 9200 0 9270 10
rect 9285 40 9355 50
rect 9285 10 9305 40
rect 9335 10 9355 40
rect 9285 0 9355 10
rect 9370 40 9440 50
rect 9370 10 9390 40
rect 9420 10 9440 40
rect 9370 0 9440 10
rect 9455 40 9525 50
rect 9455 10 9475 40
rect 9505 10 9525 40
rect 9455 0 9525 10
rect 9540 40 9610 50
rect 9540 10 9560 40
rect 9590 10 9610 40
rect 9540 0 9610 10
rect 9625 40 9695 50
rect 9625 10 9645 40
rect 9675 10 9695 40
rect 9625 0 9695 10
rect 9710 40 9780 50
rect 9710 10 9730 40
rect 9760 10 9780 40
rect 9710 0 9780 10
rect 9795 40 9865 50
rect 9795 10 9815 40
rect 9845 10 9865 40
rect 9795 0 9865 10
rect 9880 40 9950 50
rect 9880 10 9900 40
rect 9930 10 9950 40
rect 9880 0 9950 10
rect 9965 40 10035 50
rect 9965 10 9985 40
rect 10015 10 10035 40
rect 9965 0 10035 10
rect 10050 40 10120 50
rect 10050 10 10070 40
rect 10100 10 10120 40
rect 10050 0 10120 10
rect 10135 40 10205 50
rect 10135 10 10155 40
rect 10185 10 10205 40
rect 10135 0 10205 10
rect 10220 40 10290 50
rect 10220 10 10240 40
rect 10270 10 10290 40
rect 10220 0 10290 10
rect 10305 40 10375 50
rect 10305 10 10325 40
rect 10355 10 10375 40
rect 10305 0 10375 10
rect 10390 40 10460 50
rect 10390 10 10410 40
rect 10440 10 10460 40
rect 10390 0 10460 10
rect 10475 40 10545 50
rect 10475 10 10495 40
rect 10525 10 10545 40
rect 10475 0 10545 10
rect 10560 40 10630 50
rect 10560 10 10580 40
rect 10610 10 10630 40
rect 10560 0 10630 10
rect 10645 40 10715 50
rect 10645 10 10665 40
rect 10695 10 10715 40
rect 10645 0 10715 10
rect 10730 40 10800 50
rect 10730 10 10750 40
rect 10780 10 10800 40
rect 10730 0 10800 10
rect 10815 40 10885 50
rect 10815 10 10835 40
rect 10865 10 10885 40
rect 10815 0 10885 10
rect 10900 40 10970 50
rect 10900 10 10920 40
rect 10950 10 10970 40
rect 10900 0 10970 10
rect 10985 40 11055 50
rect 10985 10 11005 40
rect 11035 10 11055 40
rect 10985 0 11055 10
rect 11070 40 11140 50
rect 11070 10 11090 40
rect 11120 10 11140 40
rect 11070 0 11140 10
rect 11155 40 11225 50
rect 11155 10 11175 40
rect 11205 10 11225 40
rect 11155 0 11225 10
rect 11240 40 11310 50
rect 11240 10 11260 40
rect 11290 10 11310 40
rect 11240 0 11310 10
rect 11325 40 11395 50
rect 11325 10 11345 40
rect 11375 10 11395 40
rect 11325 0 11395 10
rect 11410 40 11480 50
rect 11410 10 11430 40
rect 11460 10 11480 40
rect 11410 0 11480 10
rect 11495 40 11565 50
rect 11495 10 11515 40
rect 11545 10 11565 40
rect 11495 0 11565 10
rect 11580 40 11650 50
rect 11580 10 11600 40
rect 11630 10 11650 40
rect 11580 0 11650 10
rect 11665 40 11735 50
rect 11665 10 11685 40
rect 11715 10 11735 40
rect 11665 0 11735 10
rect 11750 40 11820 50
rect 11750 10 11770 40
rect 11800 10 11820 40
rect 11750 0 11820 10
rect 11835 40 11905 50
rect 11835 10 11855 40
rect 11885 10 11905 40
rect 11835 0 11905 10
rect 11920 40 11990 50
rect 11920 10 11940 40
rect 11970 10 11990 40
rect 11920 0 11990 10
rect 12005 40 12075 50
rect 12005 10 12025 40
rect 12055 10 12075 40
rect 12005 0 12075 10
rect 12090 40 12160 50
rect 12090 10 12110 40
rect 12140 10 12160 40
rect 12090 0 12160 10
rect 12175 40 12245 50
rect 12175 10 12195 40
rect 12225 10 12245 40
rect 12175 0 12245 10
rect 12260 40 12330 50
rect 12260 10 12280 40
rect 12310 10 12330 40
rect 12260 0 12330 10
rect 12345 40 12415 50
rect 12345 10 12365 40
rect 12395 10 12415 40
rect 12345 0 12415 10
rect 12430 40 12500 50
rect 12430 10 12450 40
rect 12480 10 12500 40
rect 12430 0 12500 10
rect 12515 40 12585 50
rect 12515 10 12535 40
rect 12565 10 12585 40
rect 12515 0 12585 10
rect 12600 40 12670 50
rect 12600 10 12620 40
rect 12650 10 12670 40
rect 12600 0 12670 10
rect 12685 40 12755 50
rect 12685 10 12705 40
rect 12735 10 12755 40
rect 12685 0 12755 10
rect 12770 40 12840 50
rect 12770 10 12790 40
rect 12820 10 12840 40
rect 12770 0 12840 10
rect 12855 40 12925 50
rect 12855 10 12875 40
rect 12905 10 12925 40
rect 12855 0 12925 10
rect 12940 40 13010 50
rect 12940 10 12960 40
rect 12990 10 13010 40
rect 12940 0 13010 10
rect 13025 40 13095 50
rect 13025 10 13045 40
rect 13075 10 13095 40
rect 13025 0 13095 10
rect 13110 40 13180 50
rect 13110 10 13130 40
rect 13160 10 13180 40
rect 13110 0 13180 10
rect 13195 40 13265 50
rect 13195 10 13215 40
rect 13245 10 13265 40
rect 13195 0 13265 10
rect 13280 40 13350 50
rect 13280 10 13300 40
rect 13330 10 13350 40
rect 13280 0 13350 10
rect 13365 40 13435 50
rect 13365 10 13385 40
rect 13415 10 13435 40
rect 13365 0 13435 10
rect 13450 40 13520 50
rect 13450 10 13470 40
rect 13500 10 13520 40
rect 13450 0 13520 10
rect 13535 40 13605 50
rect 13535 10 13555 40
rect 13585 10 13605 40
rect 13535 0 13605 10
rect 13620 40 13690 50
rect 13620 10 13640 40
rect 13670 10 13690 40
rect 13620 0 13690 10
rect 13705 40 13775 50
rect 13705 10 13725 40
rect 13755 10 13775 40
rect 13705 0 13775 10
rect 13790 40 13860 50
rect 13790 10 13810 40
rect 13840 10 13860 40
rect 13790 0 13860 10
rect 13875 40 13945 50
rect 13875 10 13895 40
rect 13925 10 13945 40
rect 13875 0 13945 10
rect 13960 40 14030 50
rect 13960 10 13980 40
rect 14010 10 14030 40
rect 13960 0 14030 10
rect 14045 40 14115 50
rect 14045 10 14065 40
rect 14095 10 14115 40
rect 14045 0 14115 10
rect 14130 40 14200 50
rect 14130 10 14150 40
rect 14180 10 14200 40
rect 14130 0 14200 10
rect 14215 40 14285 50
rect 14215 10 14235 40
rect 14265 10 14285 40
rect 14215 0 14285 10
rect 14300 40 14370 50
rect 14300 10 14320 40
rect 14350 10 14370 40
rect 14300 0 14370 10
rect 14385 40 14455 50
rect 14385 10 14405 40
rect 14435 10 14455 40
rect 14385 0 14455 10
rect 14470 40 14540 50
rect 14470 10 14490 40
rect 14520 10 14540 40
rect 14470 0 14540 10
rect 14555 40 14625 50
rect 14555 10 14575 40
rect 14605 10 14625 40
rect 14555 0 14625 10
rect 14640 40 14710 50
rect 14640 10 14660 40
rect 14690 10 14710 40
rect 14640 0 14710 10
rect 14725 40 14795 50
rect 14725 10 14745 40
rect 14775 10 14795 40
rect 14725 0 14795 10
rect 14810 40 14880 50
rect 14810 10 14830 40
rect 14860 10 14880 40
rect 14810 0 14880 10
rect 14895 40 14965 50
rect 14895 10 14915 40
rect 14945 10 14965 40
rect 14895 0 14965 10
rect 14980 40 15050 50
rect 14980 10 15000 40
rect 15030 10 15050 40
rect 14980 0 15050 10
rect 15065 40 15135 50
rect 15065 10 15085 40
rect 15115 10 15135 40
rect 15065 0 15135 10
rect 15150 40 15220 50
rect 15150 10 15170 40
rect 15200 10 15220 40
rect 15150 0 15220 10
rect 15235 40 15305 50
rect 15235 10 15255 40
rect 15285 10 15305 40
rect 15235 0 15305 10
rect 15320 40 15390 50
rect 15320 10 15340 40
rect 15370 10 15390 40
rect 15320 0 15390 10
rect 15405 40 15475 50
rect 15405 10 15425 40
rect 15455 10 15475 40
rect 15405 0 15475 10
rect 15490 40 15560 50
rect 15490 10 15510 40
rect 15540 10 15560 40
rect 15490 0 15560 10
rect 15575 40 15645 50
rect 15575 10 15595 40
rect 15625 10 15645 40
rect 15575 0 15645 10
rect 15660 40 15730 50
rect 15660 10 15680 40
rect 15710 10 15730 40
rect 15660 0 15730 10
rect 15745 40 15815 50
rect 15745 10 15765 40
rect 15795 10 15815 40
rect 15745 0 15815 10
rect 15830 40 15900 50
rect 15830 10 15850 40
rect 15880 10 15900 40
rect 15830 0 15900 10
rect 15915 40 15985 50
rect 15915 10 15935 40
rect 15965 10 15985 40
rect 15915 0 15985 10
rect 16000 40 16070 50
rect 16000 10 16020 40
rect 16050 10 16070 40
rect 16000 0 16070 10
rect 16085 40 16155 50
rect 16085 10 16105 40
rect 16135 10 16155 40
rect 16085 0 16155 10
rect 16170 40 16240 50
rect 16170 10 16190 40
rect 16220 10 16240 40
rect 16170 0 16240 10
rect 16255 40 16325 50
rect 16255 10 16275 40
rect 16305 10 16325 40
rect 16255 0 16325 10
rect 16340 40 16410 50
rect 16340 10 16360 40
rect 16390 10 16410 40
rect 16340 0 16410 10
rect 16425 40 16495 50
rect 16425 10 16445 40
rect 16475 10 16495 40
rect 16425 0 16495 10
rect 16510 40 16580 50
rect 16510 10 16530 40
rect 16560 10 16580 40
rect 16510 0 16580 10
rect 16595 40 16665 50
rect 16595 10 16615 40
rect 16645 10 16665 40
rect 16595 0 16665 10
rect 16680 40 16750 50
rect 16680 10 16700 40
rect 16730 10 16750 40
rect 16680 0 16750 10
rect 16765 40 16835 50
rect 16765 10 16785 40
rect 16815 10 16835 40
rect 16765 0 16835 10
rect 16850 40 16920 50
rect 16850 10 16870 40
rect 16900 10 16920 40
rect 16850 0 16920 10
rect 16935 40 17005 50
rect 16935 10 16955 40
rect 16985 10 17005 40
rect 16935 0 17005 10
rect 17020 40 17090 50
rect 17020 10 17040 40
rect 17070 10 17090 40
rect 17020 0 17090 10
rect 17105 40 17175 50
rect 17105 10 17125 40
rect 17155 10 17175 40
rect 17105 0 17175 10
rect 17190 40 17260 50
rect 17190 10 17210 40
rect 17240 10 17260 40
rect 17190 0 17260 10
rect 17275 40 17345 50
rect 17275 10 17295 40
rect 17325 10 17345 40
rect 17275 0 17345 10
rect 17360 40 17430 50
rect 17360 10 17380 40
rect 17410 10 17430 40
rect 17360 0 17430 10
rect 17445 40 17515 50
rect 17445 10 17465 40
rect 17495 10 17515 40
rect 17445 0 17515 10
rect 17530 40 17600 50
rect 17530 10 17550 40
rect 17580 10 17600 40
rect 17530 0 17600 10
rect 17615 40 17685 50
rect 17615 10 17635 40
rect 17665 10 17685 40
rect 17615 0 17685 10
rect 17700 40 17770 50
rect 17700 10 17720 40
rect 17750 10 17770 40
rect 17700 0 17770 10
rect 17785 40 17855 50
rect 17785 10 17805 40
rect 17835 10 17855 40
rect 17785 0 17855 10
rect 17870 40 17940 50
rect 17870 10 17890 40
rect 17920 10 17940 40
rect 17870 0 17940 10
rect 17955 40 18025 50
rect 17955 10 17975 40
rect 18005 10 18025 40
rect 17955 0 18025 10
rect 18040 40 18110 50
rect 18040 10 18060 40
rect 18090 10 18110 40
rect 18040 0 18110 10
rect 18125 40 18195 50
rect 18125 10 18145 40
rect 18175 10 18195 40
rect 18125 0 18195 10
rect 18210 40 18280 50
rect 18210 10 18230 40
rect 18260 10 18280 40
rect 18210 0 18280 10
rect 18295 40 18365 50
rect 18295 10 18315 40
rect 18345 10 18365 40
rect 18295 0 18365 10
rect 18380 40 18450 50
rect 18380 10 18400 40
rect 18430 10 18450 40
rect 18380 0 18450 10
rect 18465 40 18535 50
rect 18465 10 18485 40
rect 18515 10 18535 40
rect 18465 0 18535 10
rect 18550 40 18620 50
rect 18550 10 18570 40
rect 18600 10 18620 40
rect 18550 0 18620 10
rect 18635 40 18705 50
rect 18635 10 18655 40
rect 18685 10 18705 40
rect 18635 0 18705 10
rect 18720 40 18790 50
rect 18720 10 18740 40
rect 18770 10 18790 40
rect 18720 0 18790 10
rect 18805 40 18875 50
rect 18805 10 18825 40
rect 18855 10 18875 40
rect 18805 0 18875 10
rect 18890 40 18960 50
rect 18890 10 18910 40
rect 18940 10 18960 40
rect 18890 0 18960 10
rect 18975 40 19045 50
rect 18975 10 18995 40
rect 19025 10 19045 40
rect 18975 0 19045 10
rect 19060 40 19130 50
rect 19060 10 19080 40
rect 19110 10 19130 40
rect 19060 0 19130 10
rect 19145 40 19215 50
rect 19145 10 19165 40
rect 19195 10 19215 40
rect 19145 0 19215 10
rect 19230 40 19300 50
rect 19230 10 19250 40
rect 19280 10 19300 40
rect 19230 0 19300 10
rect 19315 40 19385 50
rect 19315 10 19335 40
rect 19365 10 19385 40
rect 19315 0 19385 10
rect 19400 40 19470 50
rect 19400 10 19420 40
rect 19450 10 19470 40
rect 19400 0 19470 10
rect 19485 40 19555 50
rect 19485 10 19505 40
rect 19535 10 19555 40
rect 19485 0 19555 10
rect 19570 40 19640 50
rect 19570 10 19590 40
rect 19620 10 19640 40
rect 19570 0 19640 10
rect 19655 40 19725 50
rect 19655 10 19675 40
rect 19705 10 19725 40
rect 19655 0 19725 10
rect 19740 40 19810 50
rect 19740 10 19760 40
rect 19790 10 19810 40
rect 19740 0 19810 10
rect 19825 40 19895 50
rect 19825 10 19845 40
rect 19875 10 19895 40
rect 19825 0 19895 10
rect 19910 40 19980 50
rect 19910 10 19930 40
rect 19960 10 19980 40
rect 19910 0 19980 10
rect 19995 40 20065 50
rect 19995 10 20015 40
rect 20045 10 20065 40
rect 19995 0 20065 10
rect 20080 40 20150 50
rect 20080 10 20100 40
rect 20130 10 20150 40
rect 20080 0 20150 10
rect 20165 40 20235 50
rect 20165 10 20185 40
rect 20215 10 20235 40
rect 20165 0 20235 10
rect 20250 40 20320 50
rect 20250 10 20270 40
rect 20300 10 20320 40
rect 20250 0 20320 10
rect 20335 40 20405 50
rect 20335 10 20355 40
rect 20385 10 20405 40
rect 20335 0 20405 10
rect 20420 40 20490 50
rect 20420 10 20440 40
rect 20470 10 20490 40
rect 20420 0 20490 10
rect 20505 40 20575 50
rect 20505 10 20525 40
rect 20555 10 20575 40
rect 20505 0 20575 10
rect 20590 40 20660 50
rect 20590 10 20610 40
rect 20640 10 20660 40
rect 20590 0 20660 10
rect 20675 40 20745 50
rect 20675 10 20695 40
rect 20725 10 20745 40
rect 20675 0 20745 10
rect 20760 40 20830 50
rect 20760 10 20780 40
rect 20810 10 20830 40
rect 20760 0 20830 10
rect 20845 40 20915 50
rect 20845 10 20865 40
rect 20895 10 20915 40
rect 20845 0 20915 10
rect 20930 40 21000 50
rect 20930 10 20950 40
rect 20980 10 21000 40
rect 20930 0 21000 10
rect 21015 40 21085 50
rect 21015 10 21035 40
rect 21065 10 21085 40
rect 21015 0 21085 10
rect 21100 40 21170 50
rect 21100 10 21120 40
rect 21150 10 21170 40
rect 21100 0 21170 10
rect 21185 40 21255 50
rect 21185 10 21205 40
rect 21235 10 21255 40
rect 21185 0 21255 10
rect 21270 40 21340 50
rect 21270 10 21290 40
rect 21320 10 21340 40
rect 21270 0 21340 10
rect 21355 40 21425 50
rect 21355 10 21375 40
rect 21405 10 21425 40
rect 21355 0 21425 10
rect 21440 40 21510 50
rect 21440 10 21460 40
rect 21490 10 21510 40
rect 21440 0 21510 10
rect 21525 40 21595 50
rect 21525 10 21545 40
rect 21575 10 21595 40
rect 21525 0 21595 10
rect 21610 40 21680 50
rect 21610 10 21630 40
rect 21660 10 21680 40
rect 21610 0 21680 10
rect 21695 40 21765 50
rect 21695 10 21715 40
rect 21745 10 21765 40
rect 21695 0 21765 10
rect 21780 40 21850 50
rect 21780 10 21800 40
rect 21830 10 21850 40
rect 21780 0 21850 10
rect 21865 40 21935 50
rect 21865 10 21885 40
rect 21915 10 21935 40
rect 21865 0 21935 10
rect 21950 40 22020 50
rect 21950 10 21970 40
rect 22000 10 22020 40
rect 21950 0 22020 10
rect 22035 40 22105 50
rect 22035 10 22055 40
rect 22085 10 22105 40
rect 22035 0 22105 10
rect 22120 40 22190 50
rect 22120 10 22140 40
rect 22170 10 22190 40
rect 22120 0 22190 10
rect 22205 40 22275 50
rect 22205 10 22225 40
rect 22255 10 22275 40
rect 22205 0 22275 10
rect 22290 40 22360 50
rect 22290 10 22310 40
rect 22340 10 22360 40
rect 22290 0 22360 10
rect 22375 40 22445 50
rect 22375 10 22395 40
rect 22425 10 22445 40
rect 22375 0 22445 10
rect 22460 40 22530 50
rect 22460 10 22480 40
rect 22510 10 22530 40
rect 22460 0 22530 10
rect 22545 40 22615 50
rect 22545 10 22565 40
rect 22595 10 22615 40
rect 22545 0 22615 10
rect 22630 40 22700 50
rect 22630 10 22650 40
rect 22680 10 22700 40
rect 22630 0 22700 10
rect 22715 40 22785 50
rect 22715 10 22735 40
rect 22765 10 22785 40
rect 22715 0 22785 10
rect 22800 40 22870 50
rect 22800 10 22820 40
rect 22850 10 22870 40
rect 22800 0 22870 10
rect 22885 40 22955 50
rect 22885 10 22905 40
rect 22935 10 22955 40
rect 22885 0 22955 10
rect 22970 40 23040 50
rect 22970 10 22990 40
rect 23020 10 23040 40
rect 22970 0 23040 10
rect 23055 40 23125 50
rect 23055 10 23075 40
rect 23105 10 23125 40
rect 23055 0 23125 10
rect 23140 40 23210 50
rect 23140 10 23160 40
rect 23190 10 23210 40
rect 23140 0 23210 10
rect 23225 40 23295 50
rect 23225 10 23245 40
rect 23275 10 23295 40
rect 23225 0 23295 10
rect 23310 40 23380 50
rect 23310 10 23330 40
rect 23360 10 23380 40
rect 23310 0 23380 10
rect 23395 40 23465 50
rect 23395 10 23415 40
rect 23445 10 23465 40
rect 23395 0 23465 10
rect 23480 40 23550 50
rect 23480 10 23500 40
rect 23530 10 23550 40
rect 23480 0 23550 10
rect 23565 40 23635 50
rect 23565 10 23585 40
rect 23615 10 23635 40
rect 23565 0 23635 10
rect 23650 40 23720 50
rect 23650 10 23670 40
rect 23700 10 23720 40
rect 23650 0 23720 10
rect 23735 40 23805 50
rect 23735 10 23755 40
rect 23785 10 23805 40
rect 23735 0 23805 10
rect 23820 40 23890 50
rect 23820 10 23840 40
rect 23870 10 23890 40
rect 23820 0 23890 10
rect 23905 40 23975 50
rect 23905 10 23925 40
rect 23955 10 23975 40
rect 23905 0 23975 10
rect 23990 40 24060 50
rect 23990 10 24010 40
rect 24040 10 24060 40
rect 23990 0 24060 10
rect 24075 40 24145 50
rect 24075 10 24095 40
rect 24125 10 24145 40
rect 24075 0 24145 10
rect 24160 40 24230 50
rect 24160 10 24180 40
rect 24210 10 24230 40
rect 24160 0 24230 10
rect 24245 40 24315 50
rect 24245 10 24265 40
rect 24295 10 24315 40
rect 24245 0 24315 10
rect 24330 40 24400 50
rect 24330 10 24350 40
rect 24380 10 24400 40
rect 24330 0 24400 10
rect 24415 40 24485 50
rect 24415 10 24435 40
rect 24465 10 24485 40
rect 24415 0 24485 10
rect 24500 40 24570 50
rect 24500 10 24520 40
rect 24550 10 24570 40
rect 24500 0 24570 10
rect 24585 40 24655 50
rect 24585 10 24605 40
rect 24635 10 24655 40
rect 24585 0 24655 10
rect 24670 40 24740 50
rect 24670 10 24690 40
rect 24720 10 24740 40
rect 24670 0 24740 10
rect 24755 40 24825 50
rect 24755 10 24775 40
rect 24805 10 24825 40
rect 24755 0 24825 10
rect 24840 40 24910 50
rect 24840 10 24860 40
rect 24890 10 24910 40
rect 24840 0 24910 10
rect 24925 40 24995 50
rect 24925 10 24945 40
rect 24975 10 24995 40
rect 24925 0 24995 10
rect 25010 40 25080 50
rect 25010 10 25030 40
rect 25060 10 25080 40
rect 25010 0 25080 10
rect 25095 40 25165 50
rect 25095 10 25115 40
rect 25145 10 25165 40
rect 25095 0 25165 10
rect 25180 40 25250 50
rect 25180 10 25200 40
rect 25230 10 25250 40
rect 25180 0 25250 10
rect 25265 40 25335 50
rect 25265 10 25285 40
rect 25315 10 25335 40
rect 25265 0 25335 10
rect 25350 40 25420 50
rect 25350 10 25370 40
rect 25400 10 25420 40
rect 25350 0 25420 10
rect 25435 40 25505 50
rect 25435 10 25455 40
rect 25485 10 25505 40
rect 25435 0 25505 10
rect 25520 40 25590 50
rect 25520 10 25540 40
rect 25570 10 25590 40
rect 25520 0 25590 10
rect 25605 40 25675 50
rect 25605 10 25625 40
rect 25655 10 25675 40
rect 25605 0 25675 10
rect 25690 40 25760 50
rect 25690 10 25710 40
rect 25740 10 25760 40
rect 25690 0 25760 10
rect 25775 40 25845 50
rect 25775 10 25795 40
rect 25825 10 25845 40
rect 25775 0 25845 10
rect 25860 40 25930 50
rect 25860 10 25880 40
rect 25910 10 25930 40
rect 25860 0 25930 10
rect 25945 40 26015 50
rect 25945 10 25965 40
rect 25995 10 26015 40
rect 25945 0 26015 10
rect 26030 40 26100 50
rect 26030 10 26050 40
rect 26080 10 26100 40
rect 26030 0 26100 10
rect 26115 40 26185 50
rect 26115 10 26135 40
rect 26165 10 26185 40
rect 26115 0 26185 10
rect 26200 40 26270 50
rect 26200 10 26220 40
rect 26250 10 26270 40
rect 26200 0 26270 10
rect 26285 40 26355 50
rect 26285 10 26305 40
rect 26335 10 26355 40
rect 26285 0 26355 10
rect 26370 40 26440 50
rect 26370 10 26390 40
rect 26420 10 26440 40
rect 26370 0 26440 10
rect 26455 40 26525 50
rect 26455 10 26475 40
rect 26505 10 26525 40
rect 26455 0 26525 10
rect 26540 40 26610 50
rect 26540 10 26560 40
rect 26590 10 26610 40
rect 26540 0 26610 10
rect 26625 40 26695 50
rect 26625 10 26645 40
rect 26675 10 26695 40
rect 26625 0 26695 10
rect 26710 40 26780 50
rect 26710 10 26730 40
rect 26760 10 26780 40
rect 26710 0 26780 10
rect 26795 40 26865 50
rect 26795 10 26815 40
rect 26845 10 26865 40
rect 26795 0 26865 10
rect 26880 40 26950 50
rect 26880 10 26900 40
rect 26930 10 26950 40
rect 26880 0 26950 10
rect 26965 40 27035 50
rect 26965 10 26985 40
rect 27015 10 27035 40
rect 26965 0 27035 10
rect 27050 40 27120 50
rect 27050 10 27070 40
rect 27100 10 27120 40
rect 27050 0 27120 10
rect 27135 40 27205 50
rect 27135 10 27155 40
rect 27185 10 27205 40
rect 27135 0 27205 10
rect 27220 40 27290 50
rect 27220 10 27240 40
rect 27270 10 27290 40
rect 27220 0 27290 10
rect 27305 40 27375 50
rect 27305 10 27325 40
rect 27355 10 27375 40
rect 27305 0 27375 10
rect 27390 40 27460 50
rect 27390 10 27410 40
rect 27440 10 27460 40
rect 27390 0 27460 10
rect 27475 40 27545 50
rect 27475 10 27495 40
rect 27525 10 27545 40
rect 27475 0 27545 10
rect 27560 40 27630 50
rect 27560 10 27580 40
rect 27610 10 27630 40
rect 27560 0 27630 10
rect 27645 40 27715 50
rect 27645 10 27665 40
rect 27695 10 27715 40
rect 27645 0 27715 10
rect 27730 40 27800 50
rect 27730 10 27750 40
rect 27780 10 27800 40
rect 27730 0 27800 10
rect 27815 40 27885 50
rect 27815 10 27835 40
rect 27865 10 27885 40
rect 27815 0 27885 10
rect 27900 40 27970 50
rect 27900 10 27920 40
rect 27950 10 27970 40
rect 27900 0 27970 10
rect 27985 40 28055 50
rect 27985 10 28005 40
rect 28035 10 28055 40
rect 27985 0 28055 10
rect 28070 40 28140 50
rect 28070 10 28090 40
rect 28120 10 28140 40
rect 28070 0 28140 10
rect 28155 40 28225 50
rect 28155 10 28175 40
rect 28205 10 28225 40
rect 28155 0 28225 10
rect 28240 40 28310 50
rect 28240 10 28260 40
rect 28290 10 28310 40
rect 28240 0 28310 10
rect 28325 40 28395 50
rect 28325 10 28345 40
rect 28375 10 28395 40
rect 28325 0 28395 10
rect 28410 40 28480 50
rect 28410 10 28430 40
rect 28460 10 28480 40
rect 28410 0 28480 10
rect 28495 40 28565 50
rect 28495 10 28515 40
rect 28545 10 28565 40
rect 28495 0 28565 10
rect 28580 40 28650 50
rect 28580 10 28600 40
rect 28630 10 28650 40
rect 28580 0 28650 10
rect 28665 40 28735 50
rect 28665 10 28685 40
rect 28715 10 28735 40
rect 28665 0 28735 10
rect 28750 40 28820 50
rect 28750 10 28770 40
rect 28800 10 28820 40
rect 28750 0 28820 10
rect 28835 40 28905 50
rect 28835 10 28855 40
rect 28885 10 28905 40
rect 28835 0 28905 10
rect 28920 40 28990 50
rect 28920 10 28940 40
rect 28970 10 28990 40
rect 28920 0 28990 10
rect 29005 40 29075 50
rect 29005 10 29025 40
rect 29055 10 29075 40
rect 29005 0 29075 10
rect 29090 40 29160 50
rect 29090 10 29110 40
rect 29140 10 29160 40
rect 29090 0 29160 10
rect 29175 40 29245 50
rect 29175 10 29195 40
rect 29225 10 29245 40
rect 29175 0 29245 10
rect 29260 40 29330 50
rect 29260 10 29280 40
rect 29310 10 29330 40
rect 29260 0 29330 10
rect 29345 40 29415 50
rect 29345 10 29365 40
rect 29395 10 29415 40
rect 29345 0 29415 10
rect 29430 40 29500 50
rect 29430 10 29450 40
rect 29480 10 29500 40
rect 29430 0 29500 10
rect 29515 40 29585 50
rect 29515 10 29535 40
rect 29565 10 29585 40
rect 29515 0 29585 10
rect 29600 40 29670 50
rect 29600 10 29620 40
rect 29650 10 29670 40
rect 29600 0 29670 10
rect -5 -30 65 -20
rect -5 -60 15 -30
rect 45 -60 65 -30
rect -5 -70 65 -60
rect 80 -30 150 -20
rect 80 -60 100 -30
rect 130 -60 150 -30
rect 80 -70 150 -60
rect 55 -335 125 -325
rect 55 -365 75 -335
rect 105 -365 125 -335
rect 55 -385 125 -365
rect 55 -415 75 -385
rect 105 -415 125 -385
rect 55 -425 125 -415
rect 140 -335 210 -325
rect 140 -365 160 -335
rect 190 -365 210 -335
rect 140 -385 210 -365
rect 140 -415 160 -385
rect 190 -415 210 -385
rect 140 -425 210 -415
rect 225 -335 295 -325
rect 225 -365 245 -335
rect 275 -365 295 -335
rect 225 -385 295 -365
rect 225 -415 245 -385
rect 275 -415 295 -385
rect 225 -425 295 -415
rect 310 -335 380 -325
rect 310 -365 330 -335
rect 360 -365 380 -335
rect 310 -385 380 -365
rect 310 -415 330 -385
rect 360 -415 380 -385
rect 310 -425 380 -415
rect 395 -335 465 -325
rect 395 -365 415 -335
rect 445 -365 465 -335
rect 395 -385 465 -365
rect 395 -415 415 -385
rect 445 -415 465 -385
rect 395 -425 465 -415
rect 480 -335 550 -325
rect 480 -365 500 -335
rect 530 -365 550 -335
rect 480 -385 550 -365
rect 480 -415 500 -385
rect 530 -415 550 -385
rect 480 -425 550 -415
rect 565 -335 635 -325
rect 565 -365 585 -335
rect 615 -365 635 -335
rect 565 -385 635 -365
rect 565 -415 585 -385
rect 615 -415 635 -385
rect 565 -425 635 -415
rect 650 -335 720 -325
rect 650 -365 670 -335
rect 700 -365 720 -335
rect 650 -385 720 -365
rect 650 -415 670 -385
rect 700 -415 720 -385
rect 650 -425 720 -415
rect 735 -335 805 -325
rect 735 -365 755 -335
rect 785 -365 805 -335
rect 735 -385 805 -365
rect 735 -415 755 -385
rect 785 -415 805 -385
rect 735 -425 805 -415
rect 820 -335 890 -325
rect 820 -365 840 -335
rect 870 -365 890 -335
rect 820 -385 890 -365
rect 820 -415 840 -385
rect 870 -415 890 -385
rect 820 -425 890 -415
rect 905 -335 975 -325
rect 905 -365 925 -335
rect 955 -365 975 -335
rect 905 -385 975 -365
rect 905 -415 925 -385
rect 955 -415 975 -385
rect 905 -425 975 -415
rect 990 -335 1060 -325
rect 990 -365 1010 -335
rect 1040 -365 1060 -335
rect 990 -385 1060 -365
rect 990 -415 1010 -385
rect 1040 -415 1060 -385
rect 990 -425 1060 -415
rect 1075 -335 1145 -325
rect 1075 -365 1095 -335
rect 1125 -365 1145 -335
rect 1075 -385 1145 -365
rect 1075 -415 1095 -385
rect 1125 -415 1145 -385
rect 1075 -425 1145 -415
rect 1160 -335 1230 -325
rect 1160 -365 1180 -335
rect 1210 -365 1230 -335
rect 1160 -385 1230 -365
rect 1160 -415 1180 -385
rect 1210 -415 1230 -385
rect 1160 -425 1230 -415
rect 1245 -335 1315 -325
rect 1245 -365 1265 -335
rect 1295 -365 1315 -335
rect 1245 -385 1315 -365
rect 1245 -415 1265 -385
rect 1295 -415 1315 -385
rect 1245 -425 1315 -415
rect 1330 -335 1400 -325
rect 1330 -365 1350 -335
rect 1380 -365 1400 -335
rect 1330 -385 1400 -365
rect 1330 -415 1350 -385
rect 1380 -415 1400 -385
rect 1330 -425 1400 -415
rect 1415 -335 1485 -325
rect 1415 -365 1435 -335
rect 1465 -365 1485 -335
rect 1415 -385 1485 -365
rect 1415 -415 1435 -385
rect 1465 -415 1485 -385
rect 1415 -425 1485 -415
rect 1500 -335 1570 -325
rect 1500 -365 1520 -335
rect 1550 -365 1570 -335
rect 1500 -385 1570 -365
rect 1500 -415 1520 -385
rect 1550 -415 1570 -385
rect 1500 -425 1570 -415
rect 1585 -335 1655 -325
rect 1585 -365 1605 -335
rect 1635 -365 1655 -335
rect 1585 -385 1655 -365
rect 1585 -415 1605 -385
rect 1635 -415 1655 -385
rect 1585 -425 1655 -415
rect 1670 -335 1740 -325
rect 1670 -365 1690 -335
rect 1720 -365 1740 -335
rect 1670 -385 1740 -365
rect 1670 -415 1690 -385
rect 1720 -415 1740 -385
rect 1670 -425 1740 -415
rect 1755 -335 1825 -325
rect 1755 -365 1775 -335
rect 1805 -365 1825 -335
rect 1755 -385 1825 -365
rect 1755 -415 1775 -385
rect 1805 -415 1825 -385
rect 1755 -425 1825 -415
rect 1840 -335 1910 -325
rect 1840 -365 1860 -335
rect 1890 -365 1910 -335
rect 1840 -385 1910 -365
rect 1840 -415 1860 -385
rect 1890 -415 1910 -385
rect 1840 -425 1910 -415
rect 1925 -335 1995 -325
rect 1925 -365 1945 -335
rect 1975 -365 1995 -335
rect 1925 -385 1995 -365
rect 1925 -415 1945 -385
rect 1975 -415 1995 -385
rect 1925 -425 1995 -415
rect 2010 -335 2080 -325
rect 2010 -365 2030 -335
rect 2060 -365 2080 -335
rect 2010 -385 2080 -365
rect 2010 -415 2030 -385
rect 2060 -415 2080 -385
rect 2010 -425 2080 -415
rect 2095 -335 2165 -325
rect 2095 -365 2115 -335
rect 2145 -365 2165 -335
rect 2095 -385 2165 -365
rect 2095 -415 2115 -385
rect 2145 -415 2165 -385
rect 2095 -425 2165 -415
rect 2180 -335 2250 -325
rect 2180 -365 2200 -335
rect 2230 -365 2250 -335
rect 2180 -385 2250 -365
rect 2180 -415 2200 -385
rect 2230 -415 2250 -385
rect 2180 -425 2250 -415
rect 2265 -335 2335 -325
rect 2265 -365 2285 -335
rect 2315 -365 2335 -335
rect 2265 -385 2335 -365
rect 2265 -415 2285 -385
rect 2315 -415 2335 -385
rect 2265 -425 2335 -415
rect 2350 -335 2420 -325
rect 2350 -365 2370 -335
rect 2400 -365 2420 -335
rect 2350 -385 2420 -365
rect 2350 -415 2370 -385
rect 2400 -415 2420 -385
rect 2350 -425 2420 -415
rect 2435 -335 2505 -325
rect 2435 -365 2455 -335
rect 2485 -365 2505 -335
rect 2435 -385 2505 -365
rect 2435 -415 2455 -385
rect 2485 -415 2505 -385
rect 2435 -425 2505 -415
rect 2520 -335 2590 -325
rect 2520 -365 2540 -335
rect 2570 -365 2590 -335
rect 2520 -385 2590 -365
rect 2520 -415 2540 -385
rect 2570 -415 2590 -385
rect 2520 -425 2590 -415
rect 2605 -335 2675 -325
rect 2605 -365 2625 -335
rect 2655 -365 2675 -335
rect 2605 -385 2675 -365
rect 2605 -415 2625 -385
rect 2655 -415 2675 -385
rect 2605 -425 2675 -415
rect 2690 -335 2760 -325
rect 2690 -365 2710 -335
rect 2740 -365 2760 -335
rect 2690 -385 2760 -365
rect 2690 -415 2710 -385
rect 2740 -415 2760 -385
rect 2690 -425 2760 -415
rect 2775 -335 2845 -325
rect 2775 -365 2795 -335
rect 2825 -365 2845 -335
rect 2775 -385 2845 -365
rect 2775 -415 2795 -385
rect 2825 -415 2845 -385
rect 2775 -425 2845 -415
rect 2860 -335 2930 -325
rect 2860 -365 2880 -335
rect 2910 -365 2930 -335
rect 2860 -385 2930 -365
rect 2860 -415 2880 -385
rect 2910 -415 2930 -385
rect 2860 -425 2930 -415
rect 2945 -335 3015 -325
rect 2945 -365 2965 -335
rect 2995 -365 3015 -335
rect 2945 -385 3015 -365
rect 2945 -415 2965 -385
rect 2995 -415 3015 -385
rect 2945 -425 3015 -415
rect 3030 -335 3100 -325
rect 3030 -365 3050 -335
rect 3080 -365 3100 -335
rect 3030 -385 3100 -365
rect 3030 -415 3050 -385
rect 3080 -415 3100 -385
rect 3030 -425 3100 -415
rect 3115 -335 3185 -325
rect 3115 -365 3135 -335
rect 3165 -365 3185 -335
rect 3115 -385 3185 -365
rect 3115 -415 3135 -385
rect 3165 -415 3185 -385
rect 3115 -425 3185 -415
rect 3200 -335 3270 -325
rect 3200 -365 3220 -335
rect 3250 -365 3270 -335
rect 3200 -385 3270 -365
rect 3200 -415 3220 -385
rect 3250 -415 3270 -385
rect 3200 -425 3270 -415
rect 3285 -335 3355 -325
rect 3285 -365 3305 -335
rect 3335 -365 3355 -335
rect 3285 -385 3355 -365
rect 3285 -415 3305 -385
rect 3335 -415 3355 -385
rect 3285 -425 3355 -415
rect 3370 -335 3440 -325
rect 3370 -365 3390 -335
rect 3420 -365 3440 -335
rect 3370 -385 3440 -365
rect 3370 -415 3390 -385
rect 3420 -415 3440 -385
rect 3370 -425 3440 -415
rect 3455 -335 3525 -325
rect 3455 -365 3475 -335
rect 3505 -365 3525 -335
rect 3455 -385 3525 -365
rect 3455 -415 3475 -385
rect 3505 -415 3525 -385
rect 3455 -425 3525 -415
rect 3540 -335 3610 -325
rect 3540 -365 3560 -335
rect 3590 -365 3610 -335
rect 3540 -385 3610 -365
rect 3540 -415 3560 -385
rect 3590 -415 3610 -385
rect 3540 -425 3610 -415
rect 3625 -335 3695 -325
rect 3625 -365 3645 -335
rect 3675 -365 3695 -335
rect 3625 -385 3695 -365
rect 3625 -415 3645 -385
rect 3675 -415 3695 -385
rect 3625 -425 3695 -415
rect 3710 -335 3780 -325
rect 3710 -365 3730 -335
rect 3760 -365 3780 -335
rect 3710 -385 3780 -365
rect 3710 -415 3730 -385
rect 3760 -415 3780 -385
rect 3710 -425 3780 -415
rect 3795 -335 3865 -325
rect 3795 -365 3815 -335
rect 3845 -365 3865 -335
rect 3795 -385 3865 -365
rect 3795 -415 3815 -385
rect 3845 -415 3865 -385
rect 3795 -425 3865 -415
rect 3880 -335 3950 -325
rect 3880 -365 3900 -335
rect 3930 -365 3950 -335
rect 3880 -385 3950 -365
rect 3880 -415 3900 -385
rect 3930 -415 3950 -385
rect 3880 -425 3950 -415
rect 3965 -335 4035 -325
rect 3965 -365 3985 -335
rect 4015 -365 4035 -335
rect 3965 -385 4035 -365
rect 3965 -415 3985 -385
rect 4015 -415 4035 -385
rect 3965 -425 4035 -415
rect 4050 -335 4120 -325
rect 4050 -365 4070 -335
rect 4100 -365 4120 -335
rect 4050 -385 4120 -365
rect 4050 -415 4070 -385
rect 4100 -415 4120 -385
rect 4050 -425 4120 -415
rect 4135 -335 4205 -325
rect 4135 -365 4155 -335
rect 4185 -365 4205 -335
rect 4135 -385 4205 -365
rect 4135 -415 4155 -385
rect 4185 -415 4205 -385
rect 4135 -425 4205 -415
rect 4220 -335 4290 -325
rect 4220 -365 4240 -335
rect 4270 -365 4290 -335
rect 4220 -385 4290 -365
rect 4220 -415 4240 -385
rect 4270 -415 4290 -385
rect 4220 -425 4290 -415
rect 4305 -335 4375 -325
rect 4305 -365 4325 -335
rect 4355 -365 4375 -335
rect 4305 -385 4375 -365
rect 4305 -415 4325 -385
rect 4355 -415 4375 -385
rect 4305 -425 4375 -415
rect 4390 -335 4460 -325
rect 4390 -365 4410 -335
rect 4440 -365 4460 -335
rect 4390 -385 4460 -365
rect 4390 -415 4410 -385
rect 4440 -415 4460 -385
rect 4390 -425 4460 -415
rect 4475 -335 4545 -325
rect 4475 -365 4495 -335
rect 4525 -365 4545 -335
rect 4475 -385 4545 -365
rect 4475 -415 4495 -385
rect 4525 -415 4545 -385
rect 4475 -425 4545 -415
rect 4560 -335 4630 -325
rect 4560 -365 4580 -335
rect 4610 -365 4630 -335
rect 4560 -385 4630 -365
rect 4560 -415 4580 -385
rect 4610 -415 4630 -385
rect 4560 -425 4630 -415
rect 4645 -335 4715 -325
rect 4645 -365 4665 -335
rect 4695 -365 4715 -335
rect 4645 -385 4715 -365
rect 4645 -415 4665 -385
rect 4695 -415 4715 -385
rect 4645 -425 4715 -415
rect 4730 -335 4800 -325
rect 4730 -365 4750 -335
rect 4780 -365 4800 -335
rect 4730 -385 4800 -365
rect 4730 -415 4750 -385
rect 4780 -415 4800 -385
rect 4730 -425 4800 -415
rect 4815 -335 4885 -325
rect 4815 -365 4835 -335
rect 4865 -365 4885 -335
rect 4815 -385 4885 -365
rect 4815 -415 4835 -385
rect 4865 -415 4885 -385
rect 4815 -425 4885 -415
rect 4900 -335 4970 -325
rect 4900 -365 4920 -335
rect 4950 -365 4970 -335
rect 4900 -385 4970 -365
rect 4900 -415 4920 -385
rect 4950 -415 4970 -385
rect 4900 -425 4970 -415
rect 4985 -335 5055 -325
rect 4985 -365 5005 -335
rect 5035 -365 5055 -335
rect 4985 -385 5055 -365
rect 4985 -415 5005 -385
rect 5035 -415 5055 -385
rect 4985 -425 5055 -415
rect 5070 -335 5140 -325
rect 5070 -365 5090 -335
rect 5120 -365 5140 -335
rect 5070 -385 5140 -365
rect 5070 -415 5090 -385
rect 5120 -415 5140 -385
rect 5070 -425 5140 -415
rect 5155 -335 5225 -325
rect 5155 -365 5175 -335
rect 5205 -365 5225 -335
rect 5155 -385 5225 -365
rect 5155 -415 5175 -385
rect 5205 -415 5225 -385
rect 5155 -425 5225 -415
rect 5240 -335 5310 -325
rect 5240 -365 5260 -335
rect 5290 -365 5310 -335
rect 5240 -385 5310 -365
rect 5240 -415 5260 -385
rect 5290 -415 5310 -385
rect 5240 -425 5310 -415
rect 5325 -335 5395 -325
rect 5325 -365 5345 -335
rect 5375 -365 5395 -335
rect 5325 -385 5395 -365
rect 5325 -415 5345 -385
rect 5375 -415 5395 -385
rect 5325 -425 5395 -415
rect 5410 -335 5480 -325
rect 5410 -365 5430 -335
rect 5460 -365 5480 -335
rect 5410 -385 5480 -365
rect 5410 -415 5430 -385
rect 5460 -415 5480 -385
rect 5410 -425 5480 -415
rect 5495 -335 5565 -325
rect 5495 -365 5515 -335
rect 5545 -365 5565 -335
rect 5495 -385 5565 -365
rect 5495 -415 5515 -385
rect 5545 -415 5565 -385
rect 5495 -425 5565 -415
rect 5580 -335 5650 -325
rect 5580 -365 5600 -335
rect 5630 -365 5650 -335
rect 5580 -385 5650 -365
rect 5580 -415 5600 -385
rect 5630 -415 5650 -385
rect 5580 -425 5650 -415
rect 5665 -335 5735 -325
rect 5665 -365 5685 -335
rect 5715 -365 5735 -335
rect 5665 -385 5735 -365
rect 5665 -415 5685 -385
rect 5715 -415 5735 -385
rect 5665 -425 5735 -415
rect 5750 -335 5820 -325
rect 5750 -365 5770 -335
rect 5800 -365 5820 -335
rect 5750 -385 5820 -365
rect 5750 -415 5770 -385
rect 5800 -415 5820 -385
rect 5750 -425 5820 -415
rect 5835 -335 5905 -325
rect 5835 -365 5855 -335
rect 5885 -365 5905 -335
rect 5835 -385 5905 -365
rect 5835 -415 5855 -385
rect 5885 -415 5905 -385
rect 5835 -425 5905 -415
rect 5920 -335 5990 -325
rect 5920 -365 5940 -335
rect 5970 -365 5990 -335
rect 5920 -385 5990 -365
rect 5920 -415 5940 -385
rect 5970 -415 5990 -385
rect 5920 -425 5990 -415
rect 6005 -335 6075 -325
rect 6005 -365 6025 -335
rect 6055 -365 6075 -335
rect 6005 -385 6075 -365
rect 6005 -415 6025 -385
rect 6055 -415 6075 -385
rect 6005 -425 6075 -415
rect 6090 -335 6160 -325
rect 6090 -365 6110 -335
rect 6140 -365 6160 -335
rect 6090 -385 6160 -365
rect 6090 -415 6110 -385
rect 6140 -415 6160 -385
rect 6090 -425 6160 -415
rect 6175 -335 6245 -325
rect 6175 -365 6195 -335
rect 6225 -365 6245 -335
rect 6175 -385 6245 -365
rect 6175 -415 6195 -385
rect 6225 -415 6245 -385
rect 6175 -425 6245 -415
rect 6260 -335 6330 -325
rect 6260 -365 6280 -335
rect 6310 -365 6330 -335
rect 6260 -385 6330 -365
rect 6260 -415 6280 -385
rect 6310 -415 6330 -385
rect 6260 -425 6330 -415
rect 6345 -335 6415 -325
rect 6345 -365 6365 -335
rect 6395 -365 6415 -335
rect 6345 -385 6415 -365
rect 6345 -415 6365 -385
rect 6395 -415 6415 -385
rect 6345 -425 6415 -415
rect 6430 -335 6500 -325
rect 6430 -365 6450 -335
rect 6480 -365 6500 -335
rect 6430 -385 6500 -365
rect 6430 -415 6450 -385
rect 6480 -415 6500 -385
rect 6430 -425 6500 -415
rect 6515 -335 6585 -325
rect 6515 -365 6535 -335
rect 6565 -365 6585 -335
rect 6515 -385 6585 -365
rect 6515 -415 6535 -385
rect 6565 -415 6585 -385
rect 6515 -425 6585 -415
rect 6600 -335 6670 -325
rect 6600 -365 6620 -335
rect 6650 -365 6670 -335
rect 6600 -385 6670 -365
rect 6600 -415 6620 -385
rect 6650 -415 6670 -385
rect 6600 -425 6670 -415
rect 6685 -335 6755 -325
rect 6685 -365 6705 -335
rect 6735 -365 6755 -335
rect 6685 -385 6755 -365
rect 6685 -415 6705 -385
rect 6735 -415 6755 -385
rect 6685 -425 6755 -415
rect 6770 -335 6840 -325
rect 6770 -365 6790 -335
rect 6820 -365 6840 -335
rect 6770 -385 6840 -365
rect 6770 -415 6790 -385
rect 6820 -415 6840 -385
rect 6770 -425 6840 -415
rect 6855 -335 6925 -325
rect 6855 -365 6875 -335
rect 6905 -365 6925 -335
rect 6855 -385 6925 -365
rect 6855 -415 6875 -385
rect 6905 -415 6925 -385
rect 6855 -425 6925 -415
rect 6940 -335 7010 -325
rect 6940 -365 6960 -335
rect 6990 -365 7010 -335
rect 6940 -385 7010 -365
rect 6940 -415 6960 -385
rect 6990 -415 7010 -385
rect 6940 -425 7010 -415
rect 7025 -335 7095 -325
rect 7025 -365 7045 -335
rect 7075 -365 7095 -335
rect 7025 -385 7095 -365
rect 7025 -415 7045 -385
rect 7075 -415 7095 -385
rect 7025 -425 7095 -415
rect 7110 -335 7180 -325
rect 7110 -365 7130 -335
rect 7160 -365 7180 -335
rect 7110 -385 7180 -365
rect 7110 -415 7130 -385
rect 7160 -415 7180 -385
rect 7110 -425 7180 -415
rect 7195 -335 7265 -325
rect 7195 -365 7215 -335
rect 7245 -365 7265 -335
rect 7195 -385 7265 -365
rect 7195 -415 7215 -385
rect 7245 -415 7265 -385
rect 7195 -425 7265 -415
rect 7280 -335 7350 -325
rect 7280 -365 7300 -335
rect 7330 -365 7350 -335
rect 7280 -385 7350 -365
rect 7280 -415 7300 -385
rect 7330 -415 7350 -385
rect 7280 -425 7350 -415
rect 7365 -335 7435 -325
rect 7365 -365 7385 -335
rect 7415 -365 7435 -335
rect 7365 -385 7435 -365
rect 7365 -415 7385 -385
rect 7415 -415 7435 -385
rect 7365 -425 7435 -415
rect 7450 -335 7520 -325
rect 7450 -365 7470 -335
rect 7500 -365 7520 -335
rect 7450 -385 7520 -365
rect 7450 -415 7470 -385
rect 7500 -415 7520 -385
rect 7450 -425 7520 -415
rect 7535 -335 7605 -325
rect 7535 -365 7555 -335
rect 7585 -365 7605 -335
rect 7535 -385 7605 -365
rect 7535 -415 7555 -385
rect 7585 -415 7605 -385
rect 7535 -425 7605 -415
rect 7620 -335 7690 -325
rect 7620 -365 7640 -335
rect 7670 -365 7690 -335
rect 7620 -385 7690 -365
rect 7620 -415 7640 -385
rect 7670 -415 7690 -385
rect 7620 -425 7690 -415
rect 7705 -335 7775 -325
rect 7705 -365 7725 -335
rect 7755 -365 7775 -335
rect 7705 -385 7775 -365
rect 7705 -415 7725 -385
rect 7755 -415 7775 -385
rect 7705 -425 7775 -415
rect 7790 -335 7860 -325
rect 7790 -365 7810 -335
rect 7840 -365 7860 -335
rect 7790 -385 7860 -365
rect 7790 -415 7810 -385
rect 7840 -415 7860 -385
rect 7790 -425 7860 -415
rect 7875 -335 7945 -325
rect 7875 -365 7895 -335
rect 7925 -365 7945 -335
rect 7875 -385 7945 -365
rect 7875 -415 7895 -385
rect 7925 -415 7945 -385
rect 7875 -425 7945 -415
rect 7960 -335 8030 -325
rect 7960 -365 7980 -335
rect 8010 -365 8030 -335
rect 7960 -385 8030 -365
rect 7960 -415 7980 -385
rect 8010 -415 8030 -385
rect 7960 -425 8030 -415
rect 8045 -335 8115 -325
rect 8045 -365 8065 -335
rect 8095 -365 8115 -335
rect 8045 -385 8115 -365
rect 8045 -415 8065 -385
rect 8095 -415 8115 -385
rect 8045 -425 8115 -415
rect 8130 -335 8200 -325
rect 8130 -365 8150 -335
rect 8180 -365 8200 -335
rect 8130 -385 8200 -365
rect 8130 -415 8150 -385
rect 8180 -415 8200 -385
rect 8130 -425 8200 -415
rect 8215 -335 8285 -325
rect 8215 -365 8235 -335
rect 8265 -365 8285 -335
rect 8215 -385 8285 -365
rect 8215 -415 8235 -385
rect 8265 -415 8285 -385
rect 8215 -425 8285 -415
rect 8300 -335 8370 -325
rect 8300 -365 8320 -335
rect 8350 -365 8370 -335
rect 8300 -385 8370 -365
rect 8300 -415 8320 -385
rect 8350 -415 8370 -385
rect 8300 -425 8370 -415
rect 8385 -335 8455 -325
rect 8385 -365 8405 -335
rect 8435 -365 8455 -335
rect 8385 -385 8455 -365
rect 8385 -415 8405 -385
rect 8435 -415 8455 -385
rect 8385 -425 8455 -415
rect 8470 -335 8540 -325
rect 8470 -365 8490 -335
rect 8520 -365 8540 -335
rect 8470 -385 8540 -365
rect 8470 -415 8490 -385
rect 8520 -415 8540 -385
rect 8470 -425 8540 -415
rect 8555 -335 8625 -325
rect 8555 -365 8575 -335
rect 8605 -365 8625 -335
rect 8555 -385 8625 -365
rect 8555 -415 8575 -385
rect 8605 -415 8625 -385
rect 8555 -425 8625 -415
rect 8640 -335 8710 -325
rect 8640 -365 8660 -335
rect 8690 -365 8710 -335
rect 8640 -385 8710 -365
rect 8640 -415 8660 -385
rect 8690 -415 8710 -385
rect 8640 -425 8710 -415
rect 8725 -335 8795 -325
rect 8725 -365 8745 -335
rect 8775 -365 8795 -335
rect 8725 -385 8795 -365
rect 8725 -415 8745 -385
rect 8775 -415 8795 -385
rect 8725 -425 8795 -415
rect 8810 -335 8880 -325
rect 8810 -365 8830 -335
rect 8860 -365 8880 -335
rect 8810 -385 8880 -365
rect 8810 -415 8830 -385
rect 8860 -415 8880 -385
rect 8810 -425 8880 -415
rect 8895 -335 8965 -325
rect 8895 -365 8915 -335
rect 8945 -365 8965 -335
rect 8895 -385 8965 -365
rect 8895 -415 8915 -385
rect 8945 -415 8965 -385
rect 8895 -425 8965 -415
rect 8980 -335 9050 -325
rect 8980 -365 9000 -335
rect 9030 -365 9050 -335
rect 8980 -385 9050 -365
rect 8980 -415 9000 -385
rect 9030 -415 9050 -385
rect 8980 -425 9050 -415
rect 9065 -335 9135 -325
rect 9065 -365 9085 -335
rect 9115 -365 9135 -335
rect 9065 -385 9135 -365
rect 9065 -415 9085 -385
rect 9115 -415 9135 -385
rect 9065 -425 9135 -415
rect 9150 -335 9220 -325
rect 9150 -365 9170 -335
rect 9200 -365 9220 -335
rect 9150 -385 9220 -365
rect 9150 -415 9170 -385
rect 9200 -415 9220 -385
rect 9150 -425 9220 -415
rect 9235 -335 9305 -325
rect 9235 -365 9255 -335
rect 9285 -365 9305 -335
rect 9235 -385 9305 -365
rect 9235 -415 9255 -385
rect 9285 -415 9305 -385
rect 9235 -425 9305 -415
rect 9320 -335 9390 -325
rect 9320 -365 9340 -335
rect 9370 -365 9390 -335
rect 9320 -385 9390 -365
rect 9320 -415 9340 -385
rect 9370 -415 9390 -385
rect 9320 -425 9390 -415
rect 9405 -335 9475 -325
rect 9405 -365 9425 -335
rect 9455 -365 9475 -335
rect 9405 -385 9475 -365
rect 9405 -415 9425 -385
rect 9455 -415 9475 -385
rect 9405 -425 9475 -415
rect 9490 -335 9560 -325
rect 9490 -365 9510 -335
rect 9540 -365 9560 -335
rect 9490 -385 9560 -365
rect 9490 -415 9510 -385
rect 9540 -415 9560 -385
rect 9490 -425 9560 -415
rect 9575 -335 9645 -325
rect 9575 -365 9595 -335
rect 9625 -365 9645 -335
rect 9575 -385 9645 -365
rect 9575 -415 9595 -385
rect 9625 -415 9645 -385
rect 9575 -425 9645 -415
rect 9660 -335 9730 -325
rect 9660 -365 9680 -335
rect 9710 -365 9730 -335
rect 9660 -385 9730 -365
rect 9660 -415 9680 -385
rect 9710 -415 9730 -385
rect 9660 -425 9730 -415
rect 9745 -335 9815 -325
rect 9745 -365 9765 -335
rect 9795 -365 9815 -335
rect 9745 -385 9815 -365
rect 9745 -415 9765 -385
rect 9795 -415 9815 -385
rect 9745 -425 9815 -415
rect 9830 -335 9900 -325
rect 9830 -365 9850 -335
rect 9880 -365 9900 -335
rect 9830 -385 9900 -365
rect 9830 -415 9850 -385
rect 9880 -415 9900 -385
rect 9830 -425 9900 -415
rect 9915 -335 9985 -325
rect 9915 -365 9935 -335
rect 9965 -365 9985 -335
rect 9915 -385 9985 -365
rect 9915 -415 9935 -385
rect 9965 -415 9985 -385
rect 9915 -425 9985 -415
rect 10000 -335 10070 -325
rect 10000 -365 10020 -335
rect 10050 -365 10070 -335
rect 10000 -385 10070 -365
rect 10000 -415 10020 -385
rect 10050 -415 10070 -385
rect 10000 -425 10070 -415
rect 10085 -335 10155 -325
rect 10085 -365 10105 -335
rect 10135 -365 10155 -335
rect 10085 -385 10155 -365
rect 10085 -415 10105 -385
rect 10135 -415 10155 -385
rect 10085 -425 10155 -415
rect 10170 -335 10240 -325
rect 10170 -365 10190 -335
rect 10220 -365 10240 -335
rect 10170 -385 10240 -365
rect 10170 -415 10190 -385
rect 10220 -415 10240 -385
rect 10170 -425 10240 -415
rect 10255 -335 10325 -325
rect 10255 -365 10275 -335
rect 10305 -365 10325 -335
rect 10255 -385 10325 -365
rect 10255 -415 10275 -385
rect 10305 -415 10325 -385
rect 10255 -425 10325 -415
rect 10340 -335 10410 -325
rect 10340 -365 10360 -335
rect 10390 -365 10410 -335
rect 10340 -385 10410 -365
rect 10340 -415 10360 -385
rect 10390 -415 10410 -385
rect 10340 -425 10410 -415
rect 10425 -335 10495 -325
rect 10425 -365 10445 -335
rect 10475 -365 10495 -335
rect 10425 -385 10495 -365
rect 10425 -415 10445 -385
rect 10475 -415 10495 -385
rect 10425 -425 10495 -415
rect 10510 -335 10580 -325
rect 10510 -365 10530 -335
rect 10560 -365 10580 -335
rect 10510 -385 10580 -365
rect 10510 -415 10530 -385
rect 10560 -415 10580 -385
rect 10510 -425 10580 -415
rect 10595 -335 10665 -325
rect 10595 -365 10615 -335
rect 10645 -365 10665 -335
rect 10595 -385 10665 -365
rect 10595 -415 10615 -385
rect 10645 -415 10665 -385
rect 10595 -425 10665 -415
rect 10680 -335 10750 -325
rect 10680 -365 10700 -335
rect 10730 -365 10750 -335
rect 10680 -385 10750 -365
rect 10680 -415 10700 -385
rect 10730 -415 10750 -385
rect 10680 -425 10750 -415
rect 10765 -335 10835 -325
rect 10765 -365 10785 -335
rect 10815 -365 10835 -335
rect 10765 -385 10835 -365
rect 10765 -415 10785 -385
rect 10815 -415 10835 -385
rect 10765 -425 10835 -415
rect 10850 -335 10920 -325
rect 10850 -365 10870 -335
rect 10900 -365 10920 -335
rect 10850 -385 10920 -365
rect 10850 -415 10870 -385
rect 10900 -415 10920 -385
rect 10850 -425 10920 -415
rect 10935 -335 11005 -325
rect 10935 -365 10955 -335
rect 10985 -365 11005 -335
rect 10935 -385 11005 -365
rect 10935 -415 10955 -385
rect 10985 -415 11005 -385
rect 10935 -425 11005 -415
rect 11020 -335 11090 -325
rect 11020 -365 11040 -335
rect 11070 -365 11090 -335
rect 11020 -385 11090 -365
rect 11020 -415 11040 -385
rect 11070 -415 11090 -385
rect 11020 -425 11090 -415
rect 11105 -335 11175 -325
rect 11105 -365 11125 -335
rect 11155 -365 11175 -335
rect 11105 -385 11175 -365
rect 11105 -415 11125 -385
rect 11155 -415 11175 -385
rect 11105 -425 11175 -415
rect 11190 -335 11260 -325
rect 11190 -365 11210 -335
rect 11240 -365 11260 -335
rect 11190 -385 11260 -365
rect 11190 -415 11210 -385
rect 11240 -415 11260 -385
rect 11190 -425 11260 -415
rect 11275 -335 11345 -325
rect 11275 -365 11295 -335
rect 11325 -365 11345 -335
rect 11275 -385 11345 -365
rect 11275 -415 11295 -385
rect 11325 -415 11345 -385
rect 11275 -425 11345 -415
rect 11360 -335 11430 -325
rect 11360 -365 11380 -335
rect 11410 -365 11430 -335
rect 11360 -385 11430 -365
rect 11360 -415 11380 -385
rect 11410 -415 11430 -385
rect 11360 -425 11430 -415
rect 11445 -335 11515 -325
rect 11445 -365 11465 -335
rect 11495 -365 11515 -335
rect 11445 -385 11515 -365
rect 11445 -415 11465 -385
rect 11495 -415 11515 -385
rect 11445 -425 11515 -415
rect 11530 -335 11600 -325
rect 11530 -365 11550 -335
rect 11580 -365 11600 -335
rect 11530 -385 11600 -365
rect 11530 -415 11550 -385
rect 11580 -415 11600 -385
rect 11530 -425 11600 -415
rect 11615 -335 11685 -325
rect 11615 -365 11635 -335
rect 11665 -365 11685 -335
rect 11615 -385 11685 -365
rect 11615 -415 11635 -385
rect 11665 -415 11685 -385
rect 11615 -425 11685 -415
rect 11700 -335 11770 -325
rect 11700 -365 11720 -335
rect 11750 -365 11770 -335
rect 11700 -385 11770 -365
rect 11700 -415 11720 -385
rect 11750 -415 11770 -385
rect 11700 -425 11770 -415
rect 11785 -335 11855 -325
rect 11785 -365 11805 -335
rect 11835 -365 11855 -335
rect 11785 -385 11855 -365
rect 11785 -415 11805 -385
rect 11835 -415 11855 -385
rect 11785 -425 11855 -415
rect 11870 -335 11940 -325
rect 11870 -365 11890 -335
rect 11920 -365 11940 -335
rect 11870 -385 11940 -365
rect 11870 -415 11890 -385
rect 11920 -415 11940 -385
rect 11870 -425 11940 -415
rect 11955 -335 12025 -325
rect 11955 -365 11975 -335
rect 12005 -365 12025 -335
rect 11955 -385 12025 -365
rect 11955 -415 11975 -385
rect 12005 -415 12025 -385
rect 11955 -425 12025 -415
rect 12040 -335 12110 -325
rect 12040 -365 12060 -335
rect 12090 -365 12110 -335
rect 12040 -385 12110 -365
rect 12040 -415 12060 -385
rect 12090 -415 12110 -385
rect 12040 -425 12110 -415
rect 12125 -335 12195 -325
rect 12125 -365 12145 -335
rect 12175 -365 12195 -335
rect 12125 -385 12195 -365
rect 12125 -415 12145 -385
rect 12175 -415 12195 -385
rect 12125 -425 12195 -415
rect 12210 -335 12280 -325
rect 12210 -365 12230 -335
rect 12260 -365 12280 -335
rect 12210 -385 12280 -365
rect 12210 -415 12230 -385
rect 12260 -415 12280 -385
rect 12210 -425 12280 -415
rect 12295 -335 12365 -325
rect 12295 -365 12315 -335
rect 12345 -365 12365 -335
rect 12295 -385 12365 -365
rect 12295 -415 12315 -385
rect 12345 -415 12365 -385
rect 12295 -425 12365 -415
rect 12380 -335 12450 -325
rect 12380 -365 12400 -335
rect 12430 -365 12450 -335
rect 12380 -385 12450 -365
rect 12380 -415 12400 -385
rect 12430 -415 12450 -385
rect 12380 -425 12450 -415
rect 12465 -335 12535 -325
rect 12465 -365 12485 -335
rect 12515 -365 12535 -335
rect 12465 -385 12535 -365
rect 12465 -415 12485 -385
rect 12515 -415 12535 -385
rect 12465 -425 12535 -415
rect 12550 -335 12620 -325
rect 12550 -365 12570 -335
rect 12600 -365 12620 -335
rect 12550 -385 12620 -365
rect 12550 -415 12570 -385
rect 12600 -415 12620 -385
rect 12550 -425 12620 -415
rect 12635 -335 12705 -325
rect 12635 -365 12655 -335
rect 12685 -365 12705 -335
rect 12635 -385 12705 -365
rect 12635 -415 12655 -385
rect 12685 -415 12705 -385
rect 12635 -425 12705 -415
rect 12720 -335 12790 -325
rect 12720 -365 12740 -335
rect 12770 -365 12790 -335
rect 12720 -385 12790 -365
rect 12720 -415 12740 -385
rect 12770 -415 12790 -385
rect 12720 -425 12790 -415
rect 12805 -335 12875 -325
rect 12805 -365 12825 -335
rect 12855 -365 12875 -335
rect 12805 -385 12875 -365
rect 12805 -415 12825 -385
rect 12855 -415 12875 -385
rect 12805 -425 12875 -415
rect 12890 -335 12960 -325
rect 12890 -365 12910 -335
rect 12940 -365 12960 -335
rect 12890 -385 12960 -365
rect 12890 -415 12910 -385
rect 12940 -415 12960 -385
rect 12890 -425 12960 -415
rect 12975 -335 13045 -325
rect 12975 -365 12995 -335
rect 13025 -365 13045 -335
rect 12975 -385 13045 -365
rect 12975 -415 12995 -385
rect 13025 -415 13045 -385
rect 12975 -425 13045 -415
rect 13060 -335 13130 -325
rect 13060 -365 13080 -335
rect 13110 -365 13130 -335
rect 13060 -385 13130 -365
rect 13060 -415 13080 -385
rect 13110 -415 13130 -385
rect 13060 -425 13130 -415
rect 13145 -335 13215 -325
rect 13145 -365 13165 -335
rect 13195 -365 13215 -335
rect 13145 -385 13215 -365
rect 13145 -415 13165 -385
rect 13195 -415 13215 -385
rect 13145 -425 13215 -415
rect 13230 -335 13300 -325
rect 13230 -365 13250 -335
rect 13280 -365 13300 -335
rect 13230 -385 13300 -365
rect 13230 -415 13250 -385
rect 13280 -415 13300 -385
rect 13230 -425 13300 -415
rect 13315 -335 13385 -325
rect 13315 -365 13335 -335
rect 13365 -365 13385 -335
rect 13315 -385 13385 -365
rect 13315 -415 13335 -385
rect 13365 -415 13385 -385
rect 13315 -425 13385 -415
rect 13400 -335 13470 -325
rect 13400 -365 13420 -335
rect 13450 -365 13470 -335
rect 13400 -385 13470 -365
rect 13400 -415 13420 -385
rect 13450 -415 13470 -385
rect 13400 -425 13470 -415
rect 13485 -335 13555 -325
rect 13485 -365 13505 -335
rect 13535 -365 13555 -335
rect 13485 -385 13555 -365
rect 13485 -415 13505 -385
rect 13535 -415 13555 -385
rect 13485 -425 13555 -415
rect 13570 -335 13640 -325
rect 13570 -365 13590 -335
rect 13620 -365 13640 -335
rect 13570 -385 13640 -365
rect 13570 -415 13590 -385
rect 13620 -415 13640 -385
rect 13570 -425 13640 -415
rect 13655 -335 13725 -325
rect 13655 -365 13675 -335
rect 13705 -365 13725 -335
rect 13655 -385 13725 -365
rect 13655 -415 13675 -385
rect 13705 -415 13725 -385
rect 13655 -425 13725 -415
rect 13740 -335 13810 -325
rect 13740 -365 13760 -335
rect 13790 -365 13810 -335
rect 13740 -385 13810 -365
rect 13740 -415 13760 -385
rect 13790 -415 13810 -385
rect 13740 -425 13810 -415
rect 13825 -335 13895 -325
rect 13825 -365 13845 -335
rect 13875 -365 13895 -335
rect 13825 -385 13895 -365
rect 13825 -415 13845 -385
rect 13875 -415 13895 -385
rect 13825 -425 13895 -415
rect 13910 -335 13980 -325
rect 13910 -365 13930 -335
rect 13960 -365 13980 -335
rect 13910 -385 13980 -365
rect 13910 -415 13930 -385
rect 13960 -415 13980 -385
rect 13910 -425 13980 -415
rect 13995 -335 14065 -325
rect 13995 -365 14015 -335
rect 14045 -365 14065 -335
rect 13995 -385 14065 -365
rect 13995 -415 14015 -385
rect 14045 -415 14065 -385
rect 13995 -425 14065 -415
rect 14080 -335 14150 -325
rect 14080 -365 14100 -335
rect 14130 -365 14150 -335
rect 14080 -385 14150 -365
rect 14080 -415 14100 -385
rect 14130 -415 14150 -385
rect 14080 -425 14150 -415
rect 14165 -335 14235 -325
rect 14165 -365 14185 -335
rect 14215 -365 14235 -335
rect 14165 -385 14235 -365
rect 14165 -415 14185 -385
rect 14215 -415 14235 -385
rect 14165 -425 14235 -415
rect 14250 -335 14320 -325
rect 14250 -365 14270 -335
rect 14300 -365 14320 -335
rect 14250 -385 14320 -365
rect 14250 -415 14270 -385
rect 14300 -415 14320 -385
rect 14250 -425 14320 -415
rect 14335 -335 14405 -325
rect 14335 -365 14355 -335
rect 14385 -365 14405 -335
rect 14335 -385 14405 -365
rect 14335 -415 14355 -385
rect 14385 -415 14405 -385
rect 14335 -425 14405 -415
rect 14420 -335 14490 -325
rect 14420 -365 14440 -335
rect 14470 -365 14490 -335
rect 14420 -385 14490 -365
rect 14420 -415 14440 -385
rect 14470 -415 14490 -385
rect 14420 -425 14490 -415
rect 14505 -335 14575 -325
rect 14505 -365 14525 -335
rect 14555 -365 14575 -335
rect 14505 -385 14575 -365
rect 14505 -415 14525 -385
rect 14555 -415 14575 -385
rect 14505 -425 14575 -415
rect 14590 -335 14660 -325
rect 14590 -365 14610 -335
rect 14640 -365 14660 -335
rect 14590 -385 14660 -365
rect 14590 -415 14610 -385
rect 14640 -415 14660 -385
rect 14590 -425 14660 -415
rect 14675 -335 14745 -325
rect 14675 -365 14695 -335
rect 14725 -365 14745 -335
rect 14675 -385 14745 -365
rect 14675 -415 14695 -385
rect 14725 -415 14745 -385
rect 14675 -425 14745 -415
rect 14760 -335 14830 -325
rect 14760 -365 14780 -335
rect 14810 -365 14830 -335
rect 14760 -385 14830 -365
rect 14760 -415 14780 -385
rect 14810 -415 14830 -385
rect 14760 -425 14830 -415
rect 14845 -335 14915 -325
rect 14845 -365 14865 -335
rect 14895 -365 14915 -335
rect 14845 -385 14915 -365
rect 14845 -415 14865 -385
rect 14895 -415 14915 -385
rect 14845 -425 14915 -415
rect 14930 -335 15000 -325
rect 14930 -365 14950 -335
rect 14980 -365 15000 -335
rect 14930 -385 15000 -365
rect 14930 -415 14950 -385
rect 14980 -415 15000 -385
rect 14930 -425 15000 -415
rect 15015 -335 15085 -325
rect 15015 -365 15035 -335
rect 15065 -365 15085 -335
rect 15015 -385 15085 -365
rect 15015 -415 15035 -385
rect 15065 -415 15085 -385
rect 15015 -425 15085 -415
rect 15100 -335 15170 -325
rect 15100 -365 15120 -335
rect 15150 -365 15170 -335
rect 15100 -385 15170 -365
rect 15100 -415 15120 -385
rect 15150 -415 15170 -385
rect 15100 -425 15170 -415
rect 15185 -335 15255 -325
rect 15185 -365 15205 -335
rect 15235 -365 15255 -335
rect 15185 -385 15255 -365
rect 15185 -415 15205 -385
rect 15235 -415 15255 -385
rect 15185 -425 15255 -415
rect 15270 -335 15340 -325
rect 15270 -365 15290 -335
rect 15320 -365 15340 -335
rect 15270 -385 15340 -365
rect 15270 -415 15290 -385
rect 15320 -415 15340 -385
rect 15270 -425 15340 -415
rect 15355 -335 15425 -325
rect 15355 -365 15375 -335
rect 15405 -365 15425 -335
rect 15355 -385 15425 -365
rect 15355 -415 15375 -385
rect 15405 -415 15425 -385
rect 15355 -425 15425 -415
rect 15440 -335 15510 -325
rect 15440 -365 15460 -335
rect 15490 -365 15510 -335
rect 15440 -385 15510 -365
rect 15440 -415 15460 -385
rect 15490 -415 15510 -385
rect 15440 -425 15510 -415
rect 15525 -335 15595 -325
rect 15525 -365 15545 -335
rect 15575 -365 15595 -335
rect 15525 -385 15595 -365
rect 15525 -415 15545 -385
rect 15575 -415 15595 -385
rect 15525 -425 15595 -415
rect 15610 -335 15680 -325
rect 15610 -365 15630 -335
rect 15660 -365 15680 -335
rect 15610 -385 15680 -365
rect 15610 -415 15630 -385
rect 15660 -415 15680 -385
rect 15610 -425 15680 -415
rect 15695 -335 15765 -325
rect 15695 -365 15715 -335
rect 15745 -365 15765 -335
rect 15695 -385 15765 -365
rect 15695 -415 15715 -385
rect 15745 -415 15765 -385
rect 15695 -425 15765 -415
rect 15780 -335 15850 -325
rect 15780 -365 15800 -335
rect 15830 -365 15850 -335
rect 15780 -385 15850 -365
rect 15780 -415 15800 -385
rect 15830 -415 15850 -385
rect 15780 -425 15850 -415
rect 15865 -335 15935 -325
rect 15865 -365 15885 -335
rect 15915 -365 15935 -335
rect 15865 -385 15935 -365
rect 15865 -415 15885 -385
rect 15915 -415 15935 -385
rect 15865 -425 15935 -415
rect 15950 -335 16020 -325
rect 15950 -365 15970 -335
rect 16000 -365 16020 -335
rect 15950 -385 16020 -365
rect 15950 -415 15970 -385
rect 16000 -415 16020 -385
rect 15950 -425 16020 -415
rect 16035 -335 16105 -325
rect 16035 -365 16055 -335
rect 16085 -365 16105 -335
rect 16035 -385 16105 -365
rect 16035 -415 16055 -385
rect 16085 -415 16105 -385
rect 16035 -425 16105 -415
rect 16120 -335 16190 -325
rect 16120 -365 16140 -335
rect 16170 -365 16190 -335
rect 16120 -385 16190 -365
rect 16120 -415 16140 -385
rect 16170 -415 16190 -385
rect 16120 -425 16190 -415
rect 16205 -335 16275 -325
rect 16205 -365 16225 -335
rect 16255 -365 16275 -335
rect 16205 -385 16275 -365
rect 16205 -415 16225 -385
rect 16255 -415 16275 -385
rect 16205 -425 16275 -415
rect 16290 -335 16360 -325
rect 16290 -365 16310 -335
rect 16340 -365 16360 -335
rect 16290 -385 16360 -365
rect 16290 -415 16310 -385
rect 16340 -415 16360 -385
rect 16290 -425 16360 -415
rect 16375 -335 16445 -325
rect 16375 -365 16395 -335
rect 16425 -365 16445 -335
rect 16375 -385 16445 -365
rect 16375 -415 16395 -385
rect 16425 -415 16445 -385
rect 16375 -425 16445 -415
rect 16460 -335 16530 -325
rect 16460 -365 16480 -335
rect 16510 -365 16530 -335
rect 16460 -385 16530 -365
rect 16460 -415 16480 -385
rect 16510 -415 16530 -385
rect 16460 -425 16530 -415
rect 16545 -335 16615 -325
rect 16545 -365 16565 -335
rect 16595 -365 16615 -335
rect 16545 -385 16615 -365
rect 16545 -415 16565 -385
rect 16595 -415 16615 -385
rect 16545 -425 16615 -415
rect 16630 -335 16700 -325
rect 16630 -365 16650 -335
rect 16680 -365 16700 -335
rect 16630 -385 16700 -365
rect 16630 -415 16650 -385
rect 16680 -415 16700 -385
rect 16630 -425 16700 -415
rect 16715 -335 16785 -325
rect 16715 -365 16735 -335
rect 16765 -365 16785 -335
rect 16715 -385 16785 -365
rect 16715 -415 16735 -385
rect 16765 -415 16785 -385
rect 16715 -425 16785 -415
rect 16800 -335 16870 -325
rect 16800 -365 16820 -335
rect 16850 -365 16870 -335
rect 16800 -385 16870 -365
rect 16800 -415 16820 -385
rect 16850 -415 16870 -385
rect 16800 -425 16870 -415
rect 16885 -335 16955 -325
rect 16885 -365 16905 -335
rect 16935 -365 16955 -335
rect 16885 -385 16955 -365
rect 16885 -415 16905 -385
rect 16935 -415 16955 -385
rect 16885 -425 16955 -415
rect 16970 -335 17040 -325
rect 16970 -365 16990 -335
rect 17020 -365 17040 -335
rect 16970 -385 17040 -365
rect 16970 -415 16990 -385
rect 17020 -415 17040 -385
rect 16970 -425 17040 -415
rect 17055 -335 17125 -325
rect 17055 -365 17075 -335
rect 17105 -365 17125 -335
rect 17055 -385 17125 -365
rect 17055 -415 17075 -385
rect 17105 -415 17125 -385
rect 17055 -425 17125 -415
rect 17140 -335 17210 -325
rect 17140 -365 17160 -335
rect 17190 -365 17210 -335
rect 17140 -385 17210 -365
rect 17140 -415 17160 -385
rect 17190 -415 17210 -385
rect 17140 -425 17210 -415
rect 17225 -335 17295 -325
rect 17225 -365 17245 -335
rect 17275 -365 17295 -335
rect 17225 -385 17295 -365
rect 17225 -415 17245 -385
rect 17275 -415 17295 -385
rect 17225 -425 17295 -415
rect 17310 -335 17380 -325
rect 17310 -365 17330 -335
rect 17360 -365 17380 -335
rect 17310 -385 17380 -365
rect 17310 -415 17330 -385
rect 17360 -415 17380 -385
rect 17310 -425 17380 -415
rect 17395 -335 17465 -325
rect 17395 -365 17415 -335
rect 17445 -365 17465 -335
rect 17395 -385 17465 -365
rect 17395 -415 17415 -385
rect 17445 -415 17465 -385
rect 17395 -425 17465 -415
rect 17480 -335 17550 -325
rect 17480 -365 17500 -335
rect 17530 -365 17550 -335
rect 17480 -385 17550 -365
rect 17480 -415 17500 -385
rect 17530 -415 17550 -385
rect 17480 -425 17550 -415
rect 17565 -335 17635 -325
rect 17565 -365 17585 -335
rect 17615 -365 17635 -335
rect 17565 -385 17635 -365
rect 17565 -415 17585 -385
rect 17615 -415 17635 -385
rect 17565 -425 17635 -415
rect 17650 -335 17720 -325
rect 17650 -365 17670 -335
rect 17700 -365 17720 -335
rect 17650 -385 17720 -365
rect 17650 -415 17670 -385
rect 17700 -415 17720 -385
rect 17650 -425 17720 -415
rect 17735 -335 17805 -325
rect 17735 -365 17755 -335
rect 17785 -365 17805 -335
rect 17735 -385 17805 -365
rect 17735 -415 17755 -385
rect 17785 -415 17805 -385
rect 17735 -425 17805 -415
rect 17820 -335 17890 -325
rect 17820 -365 17840 -335
rect 17870 -365 17890 -335
rect 17820 -385 17890 -365
rect 17820 -415 17840 -385
rect 17870 -415 17890 -385
rect 17820 -425 17890 -415
rect 17905 -335 17975 -325
rect 17905 -365 17925 -335
rect 17955 -365 17975 -335
rect 17905 -385 17975 -365
rect 17905 -415 17925 -385
rect 17955 -415 17975 -385
rect 17905 -425 17975 -415
rect 17990 -335 18060 -325
rect 17990 -365 18010 -335
rect 18040 -365 18060 -335
rect 17990 -385 18060 -365
rect 17990 -415 18010 -385
rect 18040 -415 18060 -385
rect 17990 -425 18060 -415
rect 18075 -335 18145 -325
rect 18075 -365 18095 -335
rect 18125 -365 18145 -335
rect 18075 -385 18145 -365
rect 18075 -415 18095 -385
rect 18125 -415 18145 -385
rect 18075 -425 18145 -415
rect 18160 -335 18230 -325
rect 18160 -365 18180 -335
rect 18210 -365 18230 -335
rect 18160 -385 18230 -365
rect 18160 -415 18180 -385
rect 18210 -415 18230 -385
rect 18160 -425 18230 -415
rect 18245 -335 18315 -325
rect 18245 -365 18265 -335
rect 18295 -365 18315 -335
rect 18245 -385 18315 -365
rect 18245 -415 18265 -385
rect 18295 -415 18315 -385
rect 18245 -425 18315 -415
rect 18330 -335 18400 -325
rect 18330 -365 18350 -335
rect 18380 -365 18400 -335
rect 18330 -385 18400 -365
rect 18330 -415 18350 -385
rect 18380 -415 18400 -385
rect 18330 -425 18400 -415
rect 18415 -335 18485 -325
rect 18415 -365 18435 -335
rect 18465 -365 18485 -335
rect 18415 -385 18485 -365
rect 18415 -415 18435 -385
rect 18465 -415 18485 -385
rect 18415 -425 18485 -415
rect 18500 -335 18570 -325
rect 18500 -365 18520 -335
rect 18550 -365 18570 -335
rect 18500 -385 18570 -365
rect 18500 -415 18520 -385
rect 18550 -415 18570 -385
rect 18500 -425 18570 -415
rect 18585 -335 18655 -325
rect 18585 -365 18605 -335
rect 18635 -365 18655 -335
rect 18585 -385 18655 -365
rect 18585 -415 18605 -385
rect 18635 -415 18655 -385
rect 18585 -425 18655 -415
rect 18670 -335 18740 -325
rect 18670 -365 18690 -335
rect 18720 -365 18740 -335
rect 18670 -385 18740 -365
rect 18670 -415 18690 -385
rect 18720 -415 18740 -385
rect 18670 -425 18740 -415
rect 18755 -335 18825 -325
rect 18755 -365 18775 -335
rect 18805 -365 18825 -335
rect 18755 -385 18825 -365
rect 18755 -415 18775 -385
rect 18805 -415 18825 -385
rect 18755 -425 18825 -415
rect 18840 -335 18910 -325
rect 18840 -365 18860 -335
rect 18890 -365 18910 -335
rect 18840 -385 18910 -365
rect 18840 -415 18860 -385
rect 18890 -415 18910 -385
rect 18840 -425 18910 -415
rect 18925 -335 18995 -325
rect 18925 -365 18945 -335
rect 18975 -365 18995 -335
rect 18925 -385 18995 -365
rect 18925 -415 18945 -385
rect 18975 -415 18995 -385
rect 18925 -425 18995 -415
rect 19010 -335 19080 -325
rect 19010 -365 19030 -335
rect 19060 -365 19080 -335
rect 19010 -385 19080 -365
rect 19010 -415 19030 -385
rect 19060 -415 19080 -385
rect 19010 -425 19080 -415
rect 19095 -335 19165 -325
rect 19095 -365 19115 -335
rect 19145 -365 19165 -335
rect 19095 -385 19165 -365
rect 19095 -415 19115 -385
rect 19145 -415 19165 -385
rect 19095 -425 19165 -415
rect 19180 -335 19250 -325
rect 19180 -365 19200 -335
rect 19230 -365 19250 -335
rect 19180 -385 19250 -365
rect 19180 -415 19200 -385
rect 19230 -415 19250 -385
rect 19180 -425 19250 -415
rect 19265 -335 19335 -325
rect 19265 -365 19285 -335
rect 19315 -365 19335 -335
rect 19265 -385 19335 -365
rect 19265 -415 19285 -385
rect 19315 -415 19335 -385
rect 19265 -425 19335 -415
rect 19350 -335 19420 -325
rect 19350 -365 19370 -335
rect 19400 -365 19420 -335
rect 19350 -385 19420 -365
rect 19350 -415 19370 -385
rect 19400 -415 19420 -385
rect 19350 -425 19420 -415
rect 19435 -335 19505 -325
rect 19435 -365 19455 -335
rect 19485 -365 19505 -335
rect 19435 -385 19505 -365
rect 19435 -415 19455 -385
rect 19485 -415 19505 -385
rect 19435 -425 19505 -415
rect 19520 -335 19590 -325
rect 19520 -365 19540 -335
rect 19570 -365 19590 -335
rect 19520 -385 19590 -365
rect 19520 -415 19540 -385
rect 19570 -415 19590 -385
rect 19520 -425 19590 -415
rect 19605 -335 19675 -325
rect 19605 -365 19625 -335
rect 19655 -365 19675 -335
rect 19605 -385 19675 -365
rect 19605 -415 19625 -385
rect 19655 -415 19675 -385
rect 19605 -425 19675 -415
rect 19690 -335 19760 -325
rect 19690 -365 19710 -335
rect 19740 -365 19760 -335
rect 19690 -385 19760 -365
rect 19690 -415 19710 -385
rect 19740 -415 19760 -385
rect 19690 -425 19760 -415
rect 19775 -335 19845 -325
rect 19775 -365 19795 -335
rect 19825 -365 19845 -335
rect 19775 -385 19845 -365
rect 19775 -415 19795 -385
rect 19825 -415 19845 -385
rect 19775 -425 19845 -415
rect 19860 -335 19930 -325
rect 19860 -365 19880 -335
rect 19910 -365 19930 -335
rect 19860 -385 19930 -365
rect 19860 -415 19880 -385
rect 19910 -415 19930 -385
rect 19860 -425 19930 -415
rect 19945 -335 20015 -325
rect 19945 -365 19965 -335
rect 19995 -365 20015 -335
rect 19945 -385 20015 -365
rect 19945 -415 19965 -385
rect 19995 -415 20015 -385
rect 19945 -425 20015 -415
rect 20030 -335 20100 -325
rect 20030 -365 20050 -335
rect 20080 -365 20100 -335
rect 20030 -385 20100 -365
rect 20030 -415 20050 -385
rect 20080 -415 20100 -385
rect 20030 -425 20100 -415
rect 20115 -335 20185 -325
rect 20115 -365 20135 -335
rect 20165 -365 20185 -335
rect 20115 -385 20185 -365
rect 20115 -415 20135 -385
rect 20165 -415 20185 -385
rect 20115 -425 20185 -415
rect 20200 -335 20270 -325
rect 20200 -365 20220 -335
rect 20250 -365 20270 -335
rect 20200 -385 20270 -365
rect 20200 -415 20220 -385
rect 20250 -415 20270 -385
rect 20200 -425 20270 -415
rect 20285 -335 20355 -325
rect 20285 -365 20305 -335
rect 20335 -365 20355 -335
rect 20285 -385 20355 -365
rect 20285 -415 20305 -385
rect 20335 -415 20355 -385
rect 20285 -425 20355 -415
rect 20370 -335 20440 -325
rect 20370 -365 20390 -335
rect 20420 -365 20440 -335
rect 20370 -385 20440 -365
rect 20370 -415 20390 -385
rect 20420 -415 20440 -385
rect 20370 -425 20440 -415
rect 20455 -335 20525 -325
rect 20455 -365 20475 -335
rect 20505 -365 20525 -335
rect 20455 -385 20525 -365
rect 20455 -415 20475 -385
rect 20505 -415 20525 -385
rect 20455 -425 20525 -415
rect 20540 -335 20610 -325
rect 20540 -365 20560 -335
rect 20590 -365 20610 -335
rect 20540 -385 20610 -365
rect 20540 -415 20560 -385
rect 20590 -415 20610 -385
rect 20540 -425 20610 -415
rect 20625 -335 20695 -325
rect 20625 -365 20645 -335
rect 20675 -365 20695 -335
rect 20625 -385 20695 -365
rect 20625 -415 20645 -385
rect 20675 -415 20695 -385
rect 20625 -425 20695 -415
rect 20710 -335 20780 -325
rect 20710 -365 20730 -335
rect 20760 -365 20780 -335
rect 20710 -385 20780 -365
rect 20710 -415 20730 -385
rect 20760 -415 20780 -385
rect 20710 -425 20780 -415
rect 20795 -335 20865 -325
rect 20795 -365 20815 -335
rect 20845 -365 20865 -335
rect 20795 -385 20865 -365
rect 20795 -415 20815 -385
rect 20845 -415 20865 -385
rect 20795 -425 20865 -415
rect 20880 -335 20950 -325
rect 20880 -365 20900 -335
rect 20930 -365 20950 -335
rect 20880 -385 20950 -365
rect 20880 -415 20900 -385
rect 20930 -415 20950 -385
rect 20880 -425 20950 -415
rect 20965 -335 21035 -325
rect 20965 -365 20985 -335
rect 21015 -365 21035 -335
rect 20965 -385 21035 -365
rect 20965 -415 20985 -385
rect 21015 -415 21035 -385
rect 20965 -425 21035 -415
rect 21050 -335 21120 -325
rect 21050 -365 21070 -335
rect 21100 -365 21120 -335
rect 21050 -385 21120 -365
rect 21050 -415 21070 -385
rect 21100 -415 21120 -385
rect 21050 -425 21120 -415
rect 21135 -335 21205 -325
rect 21135 -365 21155 -335
rect 21185 -365 21205 -335
rect 21135 -385 21205 -365
rect 21135 -415 21155 -385
rect 21185 -415 21205 -385
rect 21135 -425 21205 -415
rect 21220 -335 21290 -325
rect 21220 -365 21240 -335
rect 21270 -365 21290 -335
rect 21220 -385 21290 -365
rect 21220 -415 21240 -385
rect 21270 -415 21290 -385
rect 21220 -425 21290 -415
rect 21305 -335 21375 -325
rect 21305 -365 21325 -335
rect 21355 -365 21375 -335
rect 21305 -385 21375 -365
rect 21305 -415 21325 -385
rect 21355 -415 21375 -385
rect 21305 -425 21375 -415
rect 21390 -335 21460 -325
rect 21390 -365 21410 -335
rect 21440 -365 21460 -335
rect 21390 -385 21460 -365
rect 21390 -415 21410 -385
rect 21440 -415 21460 -385
rect 21390 -425 21460 -415
rect 21475 -335 21545 -325
rect 21475 -365 21495 -335
rect 21525 -365 21545 -335
rect 21475 -385 21545 -365
rect 21475 -415 21495 -385
rect 21525 -415 21545 -385
rect 21475 -425 21545 -415
rect 21560 -335 21630 -325
rect 21560 -365 21580 -335
rect 21610 -365 21630 -335
rect 21560 -385 21630 -365
rect 21560 -415 21580 -385
rect 21610 -415 21630 -385
rect 21560 -425 21630 -415
rect 21645 -335 21715 -325
rect 21645 -365 21665 -335
rect 21695 -365 21715 -335
rect 21645 -385 21715 -365
rect 21645 -415 21665 -385
rect 21695 -415 21715 -385
rect 21645 -425 21715 -415
rect 21730 -335 21800 -325
rect 21730 -365 21750 -335
rect 21780 -365 21800 -335
rect 21730 -385 21800 -365
rect 21730 -415 21750 -385
rect 21780 -415 21800 -385
rect 21730 -425 21800 -415
rect 21815 -335 21885 -325
rect 21815 -365 21835 -335
rect 21865 -365 21885 -335
rect 21815 -385 21885 -365
rect 21815 -415 21835 -385
rect 21865 -415 21885 -385
rect 21815 -425 21885 -415
rect 21900 -335 21970 -325
rect 21900 -365 21920 -335
rect 21950 -365 21970 -335
rect 21900 -385 21970 -365
rect 21900 -415 21920 -385
rect 21950 -415 21970 -385
rect 21900 -425 21970 -415
rect 21985 -335 22055 -325
rect 21985 -365 22005 -335
rect 22035 -365 22055 -335
rect 21985 -385 22055 -365
rect 21985 -415 22005 -385
rect 22035 -415 22055 -385
rect 21985 -425 22055 -415
rect 22070 -335 22140 -325
rect 22070 -365 22090 -335
rect 22120 -365 22140 -335
rect 22070 -385 22140 -365
rect 22070 -415 22090 -385
rect 22120 -415 22140 -385
rect 22070 -425 22140 -415
rect 22155 -335 22225 -325
rect 22155 -365 22175 -335
rect 22205 -365 22225 -335
rect 22155 -385 22225 -365
rect 22155 -415 22175 -385
rect 22205 -415 22225 -385
rect 22155 -425 22225 -415
rect 22240 -335 22310 -325
rect 22240 -365 22260 -335
rect 22290 -365 22310 -335
rect 22240 -385 22310 -365
rect 22240 -415 22260 -385
rect 22290 -415 22310 -385
rect 22240 -425 22310 -415
rect 22325 -335 22395 -325
rect 22325 -365 22345 -335
rect 22375 -365 22395 -335
rect 22325 -385 22395 -365
rect 22325 -415 22345 -385
rect 22375 -415 22395 -385
rect 22325 -425 22395 -415
rect 22410 -335 22480 -325
rect 22410 -365 22430 -335
rect 22460 -365 22480 -335
rect 22410 -385 22480 -365
rect 22410 -415 22430 -385
rect 22460 -415 22480 -385
rect 22410 -425 22480 -415
rect 22495 -335 22565 -325
rect 22495 -365 22515 -335
rect 22545 -365 22565 -335
rect 22495 -385 22565 -365
rect 22495 -415 22515 -385
rect 22545 -415 22565 -385
rect 22495 -425 22565 -415
rect 22580 -335 22650 -325
rect 22580 -365 22600 -335
rect 22630 -365 22650 -335
rect 22580 -385 22650 -365
rect 22580 -415 22600 -385
rect 22630 -415 22650 -385
rect 22580 -425 22650 -415
rect 22665 -335 22735 -325
rect 22665 -365 22685 -335
rect 22715 -365 22735 -335
rect 22665 -385 22735 -365
rect 22665 -415 22685 -385
rect 22715 -415 22735 -385
rect 22665 -425 22735 -415
rect 22750 -335 22820 -325
rect 22750 -365 22770 -335
rect 22800 -365 22820 -335
rect 22750 -385 22820 -365
rect 22750 -415 22770 -385
rect 22800 -415 22820 -385
rect 22750 -425 22820 -415
rect 22835 -335 22905 -325
rect 22835 -365 22855 -335
rect 22885 -365 22905 -335
rect 22835 -385 22905 -365
rect 22835 -415 22855 -385
rect 22885 -415 22905 -385
rect 22835 -425 22905 -415
rect 22920 -335 22990 -325
rect 22920 -365 22940 -335
rect 22970 -365 22990 -335
rect 22920 -385 22990 -365
rect 22920 -415 22940 -385
rect 22970 -415 22990 -385
rect 22920 -425 22990 -415
rect 23005 -335 23075 -325
rect 23005 -365 23025 -335
rect 23055 -365 23075 -335
rect 23005 -385 23075 -365
rect 23005 -415 23025 -385
rect 23055 -415 23075 -385
rect 23005 -425 23075 -415
rect 23090 -335 23160 -325
rect 23090 -365 23110 -335
rect 23140 -365 23160 -335
rect 23090 -385 23160 -365
rect 23090 -415 23110 -385
rect 23140 -415 23160 -385
rect 23090 -425 23160 -415
rect 23175 -335 23245 -325
rect 23175 -365 23195 -335
rect 23225 -365 23245 -335
rect 23175 -385 23245 -365
rect 23175 -415 23195 -385
rect 23225 -415 23245 -385
rect 23175 -425 23245 -415
rect 23260 -335 23330 -325
rect 23260 -365 23280 -335
rect 23310 -365 23330 -335
rect 23260 -385 23330 -365
rect 23260 -415 23280 -385
rect 23310 -415 23330 -385
rect 23260 -425 23330 -415
rect 23345 -335 23415 -325
rect 23345 -365 23365 -335
rect 23395 -365 23415 -335
rect 23345 -385 23415 -365
rect 23345 -415 23365 -385
rect 23395 -415 23415 -385
rect 23345 -425 23415 -415
rect 23430 -335 23500 -325
rect 23430 -365 23450 -335
rect 23480 -365 23500 -335
rect 23430 -385 23500 -365
rect 23430 -415 23450 -385
rect 23480 -415 23500 -385
rect 23430 -425 23500 -415
rect 23515 -335 23585 -325
rect 23515 -365 23535 -335
rect 23565 -365 23585 -335
rect 23515 -385 23585 -365
rect 23515 -415 23535 -385
rect 23565 -415 23585 -385
rect 23515 -425 23585 -415
rect 23600 -335 23670 -325
rect 23600 -365 23620 -335
rect 23650 -365 23670 -335
rect 23600 -385 23670 -365
rect 23600 -415 23620 -385
rect 23650 -415 23670 -385
rect 23600 -425 23670 -415
rect 23685 -335 23755 -325
rect 23685 -365 23705 -335
rect 23735 -365 23755 -335
rect 23685 -385 23755 -365
rect 23685 -415 23705 -385
rect 23735 -415 23755 -385
rect 23685 -425 23755 -415
rect 23770 -335 23840 -325
rect 23770 -365 23790 -335
rect 23820 -365 23840 -335
rect 23770 -385 23840 -365
rect 23770 -415 23790 -385
rect 23820 -415 23840 -385
rect 23770 -425 23840 -415
rect 23855 -335 23925 -325
rect 23855 -365 23875 -335
rect 23905 -365 23925 -335
rect 23855 -385 23925 -365
rect 23855 -415 23875 -385
rect 23905 -415 23925 -385
rect 23855 -425 23925 -415
rect 23940 -335 24010 -325
rect 23940 -365 23960 -335
rect 23990 -365 24010 -335
rect 23940 -385 24010 -365
rect 23940 -415 23960 -385
rect 23990 -415 24010 -385
rect 23940 -425 24010 -415
rect 24025 -335 24095 -325
rect 24025 -365 24045 -335
rect 24075 -365 24095 -335
rect 24025 -385 24095 -365
rect 24025 -415 24045 -385
rect 24075 -415 24095 -385
rect 24025 -425 24095 -415
rect 24110 -335 24180 -325
rect 24110 -365 24130 -335
rect 24160 -365 24180 -335
rect 24110 -385 24180 -365
rect 24110 -415 24130 -385
rect 24160 -415 24180 -385
rect 24110 -425 24180 -415
rect 24195 -335 24265 -325
rect 24195 -365 24215 -335
rect 24245 -365 24265 -335
rect 24195 -385 24265 -365
rect 24195 -415 24215 -385
rect 24245 -415 24265 -385
rect 24195 -425 24265 -415
rect 24280 -335 24350 -325
rect 24280 -365 24300 -335
rect 24330 -365 24350 -335
rect 24280 -385 24350 -365
rect 24280 -415 24300 -385
rect 24330 -415 24350 -385
rect 24280 -425 24350 -415
rect 24365 -335 24435 -325
rect 24365 -365 24385 -335
rect 24415 -365 24435 -335
rect 24365 -385 24435 -365
rect 24365 -415 24385 -385
rect 24415 -415 24435 -385
rect 24365 -425 24435 -415
rect 24450 -335 24520 -325
rect 24450 -365 24470 -335
rect 24500 -365 24520 -335
rect 24450 -385 24520 -365
rect 24450 -415 24470 -385
rect 24500 -415 24520 -385
rect 24450 -425 24520 -415
rect 24535 -335 24605 -325
rect 24535 -365 24555 -335
rect 24585 -365 24605 -335
rect 24535 -385 24605 -365
rect 24535 -415 24555 -385
rect 24585 -415 24605 -385
rect 24535 -425 24605 -415
rect 24620 -335 24690 -325
rect 24620 -365 24640 -335
rect 24670 -365 24690 -335
rect 24620 -385 24690 -365
rect 24620 -415 24640 -385
rect 24670 -415 24690 -385
rect 24620 -425 24690 -415
rect 24705 -335 24775 -325
rect 24705 -365 24725 -335
rect 24755 -365 24775 -335
rect 24705 -385 24775 -365
rect 24705 -415 24725 -385
rect 24755 -415 24775 -385
rect 24705 -425 24775 -415
rect 24790 -335 24860 -325
rect 24790 -365 24810 -335
rect 24840 -365 24860 -335
rect 24790 -385 24860 -365
rect 24790 -415 24810 -385
rect 24840 -415 24860 -385
rect 24790 -425 24860 -415
rect 24875 -335 24945 -325
rect 24875 -365 24895 -335
rect 24925 -365 24945 -335
rect 24875 -385 24945 -365
rect 24875 -415 24895 -385
rect 24925 -415 24945 -385
rect 24875 -425 24945 -415
rect 24960 -335 25030 -325
rect 24960 -365 24980 -335
rect 25010 -365 25030 -335
rect 24960 -385 25030 -365
rect 24960 -415 24980 -385
rect 25010 -415 25030 -385
rect 24960 -425 25030 -415
rect 25045 -335 25115 -325
rect 25045 -365 25065 -335
rect 25095 -365 25115 -335
rect 25045 -385 25115 -365
rect 25045 -415 25065 -385
rect 25095 -415 25115 -385
rect 25045 -425 25115 -415
rect 25130 -335 25200 -325
rect 25130 -365 25150 -335
rect 25180 -365 25200 -335
rect 25130 -385 25200 -365
rect 25130 -415 25150 -385
rect 25180 -415 25200 -385
rect 25130 -425 25200 -415
rect 25215 -335 25285 -325
rect 25215 -365 25235 -335
rect 25265 -365 25285 -335
rect 25215 -385 25285 -365
rect 25215 -415 25235 -385
rect 25265 -415 25285 -385
rect 25215 -425 25285 -415
rect 25300 -335 25370 -325
rect 25300 -365 25320 -335
rect 25350 -365 25370 -335
rect 25300 -385 25370 -365
rect 25300 -415 25320 -385
rect 25350 -415 25370 -385
rect 25300 -425 25370 -415
rect 25385 -335 25455 -325
rect 25385 -365 25405 -335
rect 25435 -365 25455 -335
rect 25385 -385 25455 -365
rect 25385 -415 25405 -385
rect 25435 -415 25455 -385
rect 25385 -425 25455 -415
rect 25470 -335 25540 -325
rect 25470 -365 25490 -335
rect 25520 -365 25540 -335
rect 25470 -385 25540 -365
rect 25470 -415 25490 -385
rect 25520 -415 25540 -385
rect 25470 -425 25540 -415
rect 25555 -335 25625 -325
rect 25555 -365 25575 -335
rect 25605 -365 25625 -335
rect 25555 -385 25625 -365
rect 25555 -415 25575 -385
rect 25605 -415 25625 -385
rect 25555 -425 25625 -415
rect 25640 -335 25710 -325
rect 25640 -365 25660 -335
rect 25690 -365 25710 -335
rect 25640 -385 25710 -365
rect 25640 -415 25660 -385
rect 25690 -415 25710 -385
rect 25640 -425 25710 -415
rect 25725 -335 25795 -325
rect 25725 -365 25745 -335
rect 25775 -365 25795 -335
rect 25725 -385 25795 -365
rect 25725 -415 25745 -385
rect 25775 -415 25795 -385
rect 25725 -425 25795 -415
rect 25810 -335 25880 -325
rect 25810 -365 25830 -335
rect 25860 -365 25880 -335
rect 25810 -385 25880 -365
rect 25810 -415 25830 -385
rect 25860 -415 25880 -385
rect 25810 -425 25880 -415
rect 25895 -335 25965 -325
rect 25895 -365 25915 -335
rect 25945 -365 25965 -335
rect 25895 -385 25965 -365
rect 25895 -415 25915 -385
rect 25945 -415 25965 -385
rect 25895 -425 25965 -415
rect 25980 -335 26050 -325
rect 25980 -365 26000 -335
rect 26030 -365 26050 -335
rect 25980 -385 26050 -365
rect 25980 -415 26000 -385
rect 26030 -415 26050 -385
rect 25980 -425 26050 -415
rect 26065 -335 26135 -325
rect 26065 -365 26085 -335
rect 26115 -365 26135 -335
rect 26065 -385 26135 -365
rect 26065 -415 26085 -385
rect 26115 -415 26135 -385
rect 26065 -425 26135 -415
rect 26150 -335 26220 -325
rect 26150 -365 26170 -335
rect 26200 -365 26220 -335
rect 26150 -385 26220 -365
rect 26150 -415 26170 -385
rect 26200 -415 26220 -385
rect 26150 -425 26220 -415
rect 26235 -335 26305 -325
rect 26235 -365 26255 -335
rect 26285 -365 26305 -335
rect 26235 -385 26305 -365
rect 26235 -415 26255 -385
rect 26285 -415 26305 -385
rect 26235 -425 26305 -415
rect 26320 -335 26390 -325
rect 26320 -365 26340 -335
rect 26370 -365 26390 -335
rect 26320 -385 26390 -365
rect 26320 -415 26340 -385
rect 26370 -415 26390 -385
rect 26320 -425 26390 -415
rect 26405 -335 26475 -325
rect 26405 -365 26425 -335
rect 26455 -365 26475 -335
rect 26405 -385 26475 -365
rect 26405 -415 26425 -385
rect 26455 -415 26475 -385
rect 26405 -425 26475 -415
rect 26490 -335 26560 -325
rect 26490 -365 26510 -335
rect 26540 -365 26560 -335
rect 26490 -385 26560 -365
rect 26490 -415 26510 -385
rect 26540 -415 26560 -385
rect 26490 -425 26560 -415
rect 26575 -335 26645 -325
rect 26575 -365 26595 -335
rect 26625 -365 26645 -335
rect 26575 -385 26645 -365
rect 26575 -415 26595 -385
rect 26625 -415 26645 -385
rect 26575 -425 26645 -415
rect 26660 -335 26730 -325
rect 26660 -365 26680 -335
rect 26710 -365 26730 -335
rect 26660 -385 26730 -365
rect 26660 -415 26680 -385
rect 26710 -415 26730 -385
rect 26660 -425 26730 -415
rect 26745 -335 26815 -325
rect 26745 -365 26765 -335
rect 26795 -365 26815 -335
rect 26745 -385 26815 -365
rect 26745 -415 26765 -385
rect 26795 -415 26815 -385
rect 26745 -425 26815 -415
rect 26830 -335 26900 -325
rect 26830 -365 26850 -335
rect 26880 -365 26900 -335
rect 26830 -385 26900 -365
rect 26830 -415 26850 -385
rect 26880 -415 26900 -385
rect 26830 -425 26900 -415
rect 26915 -335 26985 -325
rect 26915 -365 26935 -335
rect 26965 -365 26985 -335
rect 26915 -385 26985 -365
rect 26915 -415 26935 -385
rect 26965 -415 26985 -385
rect 26915 -425 26985 -415
rect 27000 -335 27070 -325
rect 27000 -365 27020 -335
rect 27050 -365 27070 -335
rect 27000 -385 27070 -365
rect 27000 -415 27020 -385
rect 27050 -415 27070 -385
rect 27000 -425 27070 -415
rect 27085 -335 27155 -325
rect 27085 -365 27105 -335
rect 27135 -365 27155 -335
rect 27085 -385 27155 -365
rect 27085 -415 27105 -385
rect 27135 -415 27155 -385
rect 27085 -425 27155 -415
rect 27170 -335 27240 -325
rect 27170 -365 27190 -335
rect 27220 -365 27240 -335
rect 27170 -385 27240 -365
rect 27170 -415 27190 -385
rect 27220 -415 27240 -385
rect 27170 -425 27240 -415
rect 27255 -335 27325 -325
rect 27255 -365 27275 -335
rect 27305 -365 27325 -335
rect 27255 -385 27325 -365
rect 27255 -415 27275 -385
rect 27305 -415 27325 -385
rect 27255 -425 27325 -415
rect 27340 -335 27410 -325
rect 27340 -365 27360 -335
rect 27390 -365 27410 -335
rect 27340 -385 27410 -365
rect 27340 -415 27360 -385
rect 27390 -415 27410 -385
rect 27340 -425 27410 -415
rect 27425 -335 27495 -325
rect 27425 -365 27445 -335
rect 27475 -365 27495 -335
rect 27425 -385 27495 -365
rect 27425 -415 27445 -385
rect 27475 -415 27495 -385
rect 27425 -425 27495 -415
rect 27510 -335 27580 -325
rect 27510 -365 27530 -335
rect 27560 -365 27580 -335
rect 27510 -385 27580 -365
rect 27510 -415 27530 -385
rect 27560 -415 27580 -385
rect 27510 -425 27580 -415
rect 27595 -335 27665 -325
rect 27595 -365 27615 -335
rect 27645 -365 27665 -335
rect 27595 -385 27665 -365
rect 27595 -415 27615 -385
rect 27645 -415 27665 -385
rect 27595 -425 27665 -415
rect 27680 -335 27750 -325
rect 27680 -365 27700 -335
rect 27730 -365 27750 -335
rect 27680 -385 27750 -365
rect 27680 -415 27700 -385
rect 27730 -415 27750 -385
rect 27680 -425 27750 -415
rect 27765 -335 27835 -325
rect 27765 -365 27785 -335
rect 27815 -365 27835 -335
rect 27765 -385 27835 -365
rect 27765 -415 27785 -385
rect 27815 -415 27835 -385
rect 27765 -425 27835 -415
rect 27850 -335 27920 -325
rect 27850 -365 27870 -335
rect 27900 -365 27920 -335
rect 27850 -385 27920 -365
rect 27850 -415 27870 -385
rect 27900 -415 27920 -385
rect 27850 -425 27920 -415
rect 27935 -335 28005 -325
rect 27935 -365 27955 -335
rect 27985 -365 28005 -335
rect 27935 -385 28005 -365
rect 27935 -415 27955 -385
rect 27985 -415 28005 -385
rect 27935 -425 28005 -415
rect 28020 -335 28090 -325
rect 28020 -365 28040 -335
rect 28070 -365 28090 -335
rect 28020 -385 28090 -365
rect 28020 -415 28040 -385
rect 28070 -415 28090 -385
rect 28020 -425 28090 -415
rect 28105 -335 28175 -325
rect 28105 -365 28125 -335
rect 28155 -365 28175 -335
rect 28105 -385 28175 -365
rect 28105 -415 28125 -385
rect 28155 -415 28175 -385
rect 28105 -425 28175 -415
rect 28190 -335 28260 -325
rect 28190 -365 28210 -335
rect 28240 -365 28260 -335
rect 28190 -385 28260 -365
rect 28190 -415 28210 -385
rect 28240 -415 28260 -385
rect 28190 -425 28260 -415
rect 28275 -335 28345 -325
rect 28275 -365 28295 -335
rect 28325 -365 28345 -335
rect 28275 -385 28345 -365
rect 28275 -415 28295 -385
rect 28325 -415 28345 -385
rect 28275 -425 28345 -415
rect 28360 -335 28430 -325
rect 28360 -365 28380 -335
rect 28410 -365 28430 -335
rect 28360 -385 28430 -365
rect 28360 -415 28380 -385
rect 28410 -415 28430 -385
rect 28360 -425 28430 -415
rect 28445 -335 28515 -325
rect 28445 -365 28465 -335
rect 28495 -365 28515 -335
rect 28445 -385 28515 -365
rect 28445 -415 28465 -385
rect 28495 -415 28515 -385
rect 28445 -425 28515 -415
rect 28530 -335 28600 -325
rect 28530 -365 28550 -335
rect 28580 -365 28600 -335
rect 28530 -385 28600 -365
rect 28530 -415 28550 -385
rect 28580 -415 28600 -385
rect 28530 -425 28600 -415
rect 28615 -335 28685 -325
rect 28615 -365 28635 -335
rect 28665 -365 28685 -335
rect 28615 -385 28685 -365
rect 28615 -415 28635 -385
rect 28665 -415 28685 -385
rect 28615 -425 28685 -415
rect 28700 -335 28770 -325
rect 28700 -365 28720 -335
rect 28750 -365 28770 -335
rect 28700 -385 28770 -365
rect 28700 -415 28720 -385
rect 28750 -415 28770 -385
rect 28700 -425 28770 -415
rect 28785 -335 28855 -325
rect 28785 -365 28805 -335
rect 28835 -365 28855 -335
rect 28785 -385 28855 -365
rect 28785 -415 28805 -385
rect 28835 -415 28855 -385
rect 28785 -425 28855 -415
rect 28870 -335 28940 -325
rect 28870 -365 28890 -335
rect 28920 -365 28940 -335
rect 28870 -385 28940 -365
rect 28870 -415 28890 -385
rect 28920 -415 28940 -385
rect 28870 -425 28940 -415
rect 28955 -335 29025 -325
rect 28955 -365 28975 -335
rect 29005 -365 29025 -335
rect 28955 -385 29025 -365
rect 28955 -415 28975 -385
rect 29005 -415 29025 -385
rect 28955 -425 29025 -415
rect 29040 -335 29110 -325
rect 29040 -365 29060 -335
rect 29090 -365 29110 -335
rect 29040 -385 29110 -365
rect 29040 -415 29060 -385
rect 29090 -415 29110 -385
rect 29040 -425 29110 -415
rect 29125 -335 29195 -325
rect 29125 -365 29145 -335
rect 29175 -365 29195 -335
rect 29125 -385 29195 -365
rect 29125 -415 29145 -385
rect 29175 -415 29195 -385
rect 29125 -425 29195 -415
rect 29210 -335 29280 -325
rect 29210 -365 29230 -335
rect 29260 -365 29280 -335
rect 29210 -385 29280 -365
rect 29210 -415 29230 -385
rect 29260 -415 29280 -385
rect 29210 -425 29280 -415
rect 29295 -335 29365 -325
rect 29295 -365 29315 -335
rect 29345 -365 29365 -335
rect 29295 -385 29365 -365
rect 29295 -415 29315 -385
rect 29345 -415 29365 -385
rect 29295 -425 29365 -415
rect 29380 -335 29450 -325
rect 29380 -365 29400 -335
rect 29430 -365 29450 -335
rect 29380 -385 29450 -365
rect 29380 -415 29400 -385
rect 29430 -415 29450 -385
rect 29380 -425 29450 -415
rect 29465 -335 29535 -325
rect 29465 -365 29485 -335
rect 29515 -365 29535 -335
rect 29465 -385 29535 -365
rect 29465 -415 29485 -385
rect 29515 -415 29535 -385
rect 29465 -425 29535 -415
rect 29550 -335 29620 -325
rect 29550 -365 29570 -335
rect 29600 -365 29620 -335
rect 29550 -385 29620 -365
rect 29550 -415 29570 -385
rect 29600 -415 29620 -385
rect 29550 -425 29620 -415
rect 29635 -335 29705 -325
rect 29635 -365 29655 -335
rect 29685 -365 29705 -335
rect 29635 -385 29705 -365
rect 29635 -415 29655 -385
rect 29685 -415 29705 -385
rect 29635 -425 29705 -415
rect 29720 -335 29790 -325
rect 29720 -365 29740 -335
rect 29770 -365 29790 -335
rect 29720 -385 29790 -365
rect 29720 -415 29740 -385
rect 29770 -415 29790 -385
rect 29720 -425 29790 -415
rect 29805 -335 29875 -325
rect 29805 -365 29825 -335
rect 29855 -365 29875 -335
rect 29805 -385 29875 -365
rect 29805 -415 29825 -385
rect 29855 -415 29875 -385
rect 29805 -425 29875 -415
rect 29890 -335 29960 -325
rect 29890 -365 29910 -335
rect 29940 -365 29960 -335
rect 29890 -385 29960 -365
rect 29890 -415 29910 -385
rect 29940 -415 29960 -385
rect 29890 -425 29960 -415
rect 29975 -335 30045 -325
rect 29975 -365 29995 -335
rect 30025 -365 30045 -335
rect 29975 -385 30045 -365
rect 29975 -415 29995 -385
rect 30025 -415 30045 -385
rect 29975 -425 30045 -415
rect 30060 -335 30130 -325
rect 30060 -365 30080 -335
rect 30110 -365 30130 -335
rect 30060 -385 30130 -365
rect 30060 -415 30080 -385
rect 30110 -415 30130 -385
rect 30060 -425 30130 -415
rect 30145 -335 30215 -325
rect 30145 -365 30165 -335
rect 30195 -365 30215 -335
rect 30145 -385 30215 -365
rect 30145 -415 30165 -385
rect 30195 -415 30215 -385
rect 30145 -425 30215 -415
rect 30230 -335 30300 -325
rect 30230 -365 30250 -335
rect 30280 -365 30300 -335
rect 30230 -385 30300 -365
rect 30230 -415 30250 -385
rect 30280 -415 30300 -385
rect 30230 -425 30300 -415
rect 30315 -335 30385 -325
rect 30315 -365 30335 -335
rect 30365 -365 30385 -335
rect 30315 -385 30385 -365
rect 30315 -415 30335 -385
rect 30365 -415 30385 -385
rect 30315 -425 30385 -415
rect 30400 -335 30470 -325
rect 30400 -365 30420 -335
rect 30450 -365 30470 -335
rect 30400 -385 30470 -365
rect 30400 -415 30420 -385
rect 30450 -415 30470 -385
rect 30400 -425 30470 -415
rect 30485 -335 30555 -325
rect 30485 -365 30505 -335
rect 30535 -365 30555 -335
rect 30485 -385 30555 -365
rect 30485 -415 30505 -385
rect 30535 -415 30555 -385
rect 30485 -425 30555 -415
rect 30570 -335 30640 -325
rect 30570 -365 30590 -335
rect 30620 -365 30640 -335
rect 30570 -385 30640 -365
rect 30570 -415 30590 -385
rect 30620 -415 30640 -385
rect 30570 -425 30640 -415
rect 30655 -335 30725 -325
rect 30655 -365 30675 -335
rect 30705 -365 30725 -335
rect 30655 -385 30725 -365
rect 30655 -415 30675 -385
rect 30705 -415 30725 -385
rect 30655 -425 30725 -415
rect 30740 -335 30810 -325
rect 30740 -365 30760 -335
rect 30790 -365 30810 -335
rect 30740 -385 30810 -365
rect 30740 -415 30760 -385
rect 30790 -415 30810 -385
rect 30740 -425 30810 -415
rect 30825 -335 30895 -325
rect 30825 -365 30845 -335
rect 30875 -365 30895 -335
rect 30825 -385 30895 -365
rect 30825 -415 30845 -385
rect 30875 -415 30895 -385
rect 30825 -425 30895 -415
rect 30910 -335 30980 -325
rect 30910 -365 30930 -335
rect 30960 -365 30980 -335
rect 30910 -385 30980 -365
rect 30910 -415 30930 -385
rect 30960 -415 30980 -385
rect 30910 -425 30980 -415
rect 30995 -335 31065 -325
rect 30995 -365 31015 -335
rect 31045 -365 31065 -335
rect 30995 -385 31065 -365
rect 30995 -415 31015 -385
rect 31045 -415 31065 -385
rect 30995 -425 31065 -415
rect 31080 -335 31150 -325
rect 31080 -365 31100 -335
rect 31130 -365 31150 -335
rect 31080 -385 31150 -365
rect 31080 -415 31100 -385
rect 31130 -415 31150 -385
rect 31080 -425 31150 -415
rect 31165 -335 31235 -325
rect 31165 -365 31185 -335
rect 31215 -365 31235 -335
rect 31165 -385 31235 -365
rect 31165 -415 31185 -385
rect 31215 -415 31235 -385
rect 31165 -425 31235 -415
rect 31250 -335 31320 -325
rect 31250 -365 31270 -335
rect 31300 -365 31320 -335
rect 31250 -385 31320 -365
rect 31250 -415 31270 -385
rect 31300 -415 31320 -385
rect 31250 -425 31320 -415
rect 31335 -335 31405 -325
rect 31335 -365 31355 -335
rect 31385 -365 31405 -335
rect 31335 -385 31405 -365
rect 31335 -415 31355 -385
rect 31385 -415 31405 -385
rect 31335 -425 31405 -415
rect 31420 -335 31490 -325
rect 31420 -365 31440 -335
rect 31470 -365 31490 -335
rect 31420 -385 31490 -365
rect 31420 -415 31440 -385
rect 31470 -415 31490 -385
rect 31420 -425 31490 -415
rect 31505 -335 31575 -325
rect 31505 -365 31525 -335
rect 31555 -365 31575 -335
rect 31505 -385 31575 -365
rect 31505 -415 31525 -385
rect 31555 -415 31575 -385
rect 31505 -425 31575 -415
rect 31590 -335 31660 -325
rect 31590 -365 31610 -335
rect 31640 -365 31660 -335
rect 31590 -385 31660 -365
rect 31590 -415 31610 -385
rect 31640 -415 31660 -385
rect 31590 -425 31660 -415
rect 31675 -335 31745 -325
rect 31675 -365 31695 -335
rect 31725 -365 31745 -335
rect 31675 -385 31745 -365
rect 31675 -415 31695 -385
rect 31725 -415 31745 -385
rect 31675 -425 31745 -415
rect 31760 -335 31830 -325
rect 31760 -365 31780 -335
rect 31810 -365 31830 -335
rect 31760 -385 31830 -365
rect 31760 -415 31780 -385
rect 31810 -415 31830 -385
rect 31760 -425 31830 -415
rect 31845 -335 31915 -325
rect 31845 -365 31865 -335
rect 31895 -365 31915 -335
rect 31845 -385 31915 -365
rect 31845 -415 31865 -385
rect 31895 -415 31915 -385
rect 31845 -425 31915 -415
rect 31930 -335 32000 -325
rect 31930 -365 31950 -335
rect 31980 -365 32000 -335
rect 31930 -385 32000 -365
rect 31930 -415 31950 -385
rect 31980 -415 32000 -385
rect 31930 -425 32000 -415
rect 32015 -335 32085 -325
rect 32015 -365 32035 -335
rect 32065 -365 32085 -335
rect 32015 -385 32085 -365
rect 32015 -415 32035 -385
rect 32065 -415 32085 -385
rect 32015 -425 32085 -415
rect 32100 -335 32170 -325
rect 32100 -365 32120 -335
rect 32150 -365 32170 -335
rect 32100 -385 32170 -365
rect 32100 -415 32120 -385
rect 32150 -415 32170 -385
rect 32100 -425 32170 -415
rect 32185 -335 32255 -325
rect 32185 -365 32205 -335
rect 32235 -365 32255 -335
rect 32185 -385 32255 -365
rect 32185 -415 32205 -385
rect 32235 -415 32255 -385
rect 32185 -425 32255 -415
rect 32270 -335 32340 -325
rect 32270 -365 32290 -335
rect 32320 -365 32340 -335
rect 32270 -385 32340 -365
rect 32270 -415 32290 -385
rect 32320 -415 32340 -385
rect 32270 -425 32340 -415
rect 32355 -335 32425 -325
rect 32355 -365 32375 -335
rect 32405 -365 32425 -335
rect 32355 -385 32425 -365
rect 32355 -415 32375 -385
rect 32405 -415 32425 -385
rect 32355 -425 32425 -415
rect 32440 -335 32510 -325
rect 32440 -365 32460 -335
rect 32490 -365 32510 -335
rect 32440 -385 32510 -365
rect 32440 -415 32460 -385
rect 32490 -415 32510 -385
rect 32440 -425 32510 -415
rect 32525 -335 32595 -325
rect 32525 -365 32545 -335
rect 32575 -365 32595 -335
rect 32525 -385 32595 -365
rect 32525 -415 32545 -385
rect 32575 -415 32595 -385
rect 32525 -425 32595 -415
rect 32610 -335 32680 -325
rect 32610 -365 32630 -335
rect 32660 -365 32680 -335
rect 32610 -385 32680 -365
rect 32610 -415 32630 -385
rect 32660 -415 32680 -385
rect 32610 -425 32680 -415
rect 32695 -335 32765 -325
rect 32695 -365 32715 -335
rect 32745 -365 32765 -335
rect 32695 -385 32765 -365
rect 32695 -415 32715 -385
rect 32745 -415 32765 -385
rect 32695 -425 32765 -415
rect 32780 -335 32850 -325
rect 32780 -365 32800 -335
rect 32830 -365 32850 -335
rect 32780 -385 32850 -365
rect 32780 -415 32800 -385
rect 32830 -415 32850 -385
rect 32780 -425 32850 -415
rect 32865 -335 32935 -325
rect 32865 -365 32885 -335
rect 32915 -365 32935 -335
rect 32865 -385 32935 -365
rect 32865 -415 32885 -385
rect 32915 -415 32935 -385
rect 32865 -425 32935 -415
rect 32950 -335 33020 -325
rect 32950 -365 32970 -335
rect 33000 -365 33020 -335
rect 32950 -385 33020 -365
rect 32950 -415 32970 -385
rect 33000 -415 33020 -385
rect 32950 -425 33020 -415
rect 33035 -335 33105 -325
rect 33035 -365 33055 -335
rect 33085 -365 33105 -335
rect 33035 -385 33105 -365
rect 33035 -415 33055 -385
rect 33085 -415 33105 -385
rect 33035 -425 33105 -415
rect 33120 -335 33190 -325
rect 33120 -365 33140 -335
rect 33170 -365 33190 -335
rect 33120 -385 33190 -365
rect 33120 -415 33140 -385
rect 33170 -415 33190 -385
rect 33120 -425 33190 -415
rect 33205 -335 33275 -325
rect 33205 -365 33225 -335
rect 33255 -365 33275 -335
rect 33205 -385 33275 -365
rect 33205 -415 33225 -385
rect 33255 -415 33275 -385
rect 33205 -425 33275 -415
rect 33290 -335 33360 -325
rect 33290 -365 33310 -335
rect 33340 -365 33360 -335
rect 33290 -385 33360 -365
rect 33290 -415 33310 -385
rect 33340 -415 33360 -385
rect 33290 -425 33360 -415
rect 33375 -335 33445 -325
rect 33375 -365 33395 -335
rect 33425 -365 33445 -335
rect 33375 -385 33445 -365
rect 33375 -415 33395 -385
rect 33425 -415 33445 -385
rect 33375 -425 33445 -415
rect 33460 -335 33530 -325
rect 33460 -365 33480 -335
rect 33510 -365 33530 -335
rect 33460 -385 33530 -365
rect 33460 -415 33480 -385
rect 33510 -415 33530 -385
rect 33460 -425 33530 -415
rect 33545 -335 33615 -325
rect 33545 -365 33565 -335
rect 33595 -365 33615 -335
rect 33545 -385 33615 -365
rect 33545 -415 33565 -385
rect 33595 -415 33615 -385
rect 33545 -425 33615 -415
rect 33630 -335 33700 -325
rect 33630 -365 33650 -335
rect 33680 -365 33700 -335
rect 33630 -385 33700 -365
rect 33630 -415 33650 -385
rect 33680 -415 33700 -385
rect 33630 -425 33700 -415
rect 33715 -335 33785 -325
rect 33715 -365 33735 -335
rect 33765 -365 33785 -335
rect 33715 -385 33785 -365
rect 33715 -415 33735 -385
rect 33765 -415 33785 -385
rect 33715 -425 33785 -415
rect 33800 -335 33870 -325
rect 33800 -365 33820 -335
rect 33850 -365 33870 -335
rect 33800 -385 33870 -365
rect 33800 -415 33820 -385
rect 33850 -415 33870 -385
rect 33800 -425 33870 -415
rect 33885 -335 33955 -325
rect 33885 -365 33905 -335
rect 33935 -365 33955 -335
rect 33885 -385 33955 -365
rect 33885 -415 33905 -385
rect 33935 -415 33955 -385
rect 33885 -425 33955 -415
rect 33970 -335 34040 -325
rect 33970 -365 33990 -335
rect 34020 -365 34040 -335
rect 33970 -385 34040 -365
rect 33970 -415 33990 -385
rect 34020 -415 34040 -385
rect 33970 -425 34040 -415
rect 34055 -335 34125 -325
rect 34055 -365 34075 -335
rect 34105 -365 34125 -335
rect 34055 -385 34125 -365
rect 34055 -415 34075 -385
rect 34105 -415 34125 -385
rect 34055 -425 34125 -415
rect 34140 -335 34210 -325
rect 34140 -365 34160 -335
rect 34190 -365 34210 -335
rect 34140 -385 34210 -365
rect 34140 -415 34160 -385
rect 34190 -415 34210 -385
rect 34140 -425 34210 -415
rect 34225 -335 34295 -325
rect 34225 -365 34245 -335
rect 34275 -365 34295 -335
rect 34225 -385 34295 -365
rect 34225 -415 34245 -385
rect 34275 -415 34295 -385
rect 34225 -425 34295 -415
rect 34310 -335 34380 -325
rect 34310 -365 34330 -335
rect 34360 -365 34380 -335
rect 34310 -385 34380 -365
rect 34310 -415 34330 -385
rect 34360 -415 34380 -385
rect 34310 -425 34380 -415
rect 34395 -335 34465 -325
rect 34395 -365 34415 -335
rect 34445 -365 34465 -335
rect 34395 -385 34465 -365
rect 34395 -415 34415 -385
rect 34445 -415 34465 -385
rect 34395 -425 34465 -415
rect 34480 -335 34550 -325
rect 34480 -365 34500 -335
rect 34530 -365 34550 -335
rect 34480 -385 34550 -365
rect 34480 -415 34500 -385
rect 34530 -415 34550 -385
rect 34480 -425 34550 -415
rect 34565 -335 34635 -325
rect 34565 -365 34585 -335
rect 34615 -365 34635 -335
rect 34565 -385 34635 -365
rect 34565 -415 34585 -385
rect 34615 -415 34635 -385
rect 34565 -425 34635 -415
rect 34650 -335 34720 -325
rect 34650 -365 34670 -335
rect 34700 -365 34720 -335
rect 34650 -385 34720 -365
rect 34650 -415 34670 -385
rect 34700 -415 34720 -385
rect 34650 -425 34720 -415
rect 34735 -335 34805 -325
rect 34735 -365 34755 -335
rect 34785 -365 34805 -335
rect 34735 -385 34805 -365
rect 34735 -415 34755 -385
rect 34785 -415 34805 -385
rect 34735 -425 34805 -415
rect 34820 -335 34890 -325
rect 34820 -365 34840 -335
rect 34870 -365 34890 -335
rect 34820 -385 34890 -365
rect 34820 -415 34840 -385
rect 34870 -415 34890 -385
rect 34820 -425 34890 -415
rect 34905 -335 34975 -325
rect 34905 -365 34925 -335
rect 34955 -365 34975 -335
rect 34905 -385 34975 -365
rect 34905 -415 34925 -385
rect 34955 -415 34975 -385
rect 34905 -425 34975 -415
rect 34990 -335 35060 -325
rect 34990 -365 35010 -335
rect 35040 -365 35060 -335
rect 34990 -385 35060 -365
rect 34990 -415 35010 -385
rect 35040 -415 35060 -385
rect 34990 -425 35060 -415
rect 35075 -335 35145 -325
rect 35075 -365 35095 -335
rect 35125 -365 35145 -335
rect 35075 -385 35145 -365
rect 35075 -415 35095 -385
rect 35125 -415 35145 -385
rect 35075 -425 35145 -415
rect 35160 -335 35230 -325
rect 35160 -365 35180 -335
rect 35210 -365 35230 -335
rect 35160 -385 35230 -365
rect 35160 -415 35180 -385
rect 35210 -415 35230 -385
rect 35160 -425 35230 -415
rect 35245 -335 35315 -325
rect 35245 -365 35265 -335
rect 35295 -365 35315 -335
rect 35245 -385 35315 -365
rect 35245 -415 35265 -385
rect 35295 -415 35315 -385
rect 35245 -425 35315 -415
rect 35330 -335 35400 -325
rect 35330 -365 35350 -335
rect 35380 -365 35400 -335
rect 35330 -385 35400 -365
rect 35330 -415 35350 -385
rect 35380 -415 35400 -385
rect 35330 -425 35400 -415
rect 35415 -335 35485 -325
rect 35415 -365 35435 -335
rect 35465 -365 35485 -335
rect 35415 -385 35485 -365
rect 35415 -415 35435 -385
rect 35465 -415 35485 -385
rect 35415 -425 35485 -415
rect 35500 -335 35570 -325
rect 35500 -365 35520 -335
rect 35550 -365 35570 -335
rect 35500 -385 35570 -365
rect 35500 -415 35520 -385
rect 35550 -415 35570 -385
rect 35500 -425 35570 -415
rect 35585 -335 35655 -325
rect 35585 -365 35605 -335
rect 35635 -365 35655 -335
rect 35585 -385 35655 -365
rect 35585 -415 35605 -385
rect 35635 -415 35655 -385
rect 35585 -425 35655 -415
rect 35670 -335 35740 -325
rect 35670 -365 35690 -335
rect 35720 -365 35740 -335
rect 35670 -385 35740 -365
rect 35670 -415 35690 -385
rect 35720 -415 35740 -385
rect 35670 -425 35740 -415
rect 35755 -335 35825 -325
rect 35755 -365 35775 -335
rect 35805 -365 35825 -335
rect 35755 -385 35825 -365
rect 35755 -415 35775 -385
rect 35805 -415 35825 -385
rect 35755 -425 35825 -415
rect 35840 -335 35910 -325
rect 35840 -365 35860 -335
rect 35890 -365 35910 -335
rect 35840 -385 35910 -365
rect 35840 -415 35860 -385
rect 35890 -415 35910 -385
rect 35840 -425 35910 -415
rect 35925 -335 35995 -325
rect 35925 -365 35945 -335
rect 35975 -365 35995 -335
rect 35925 -385 35995 -365
rect 35925 -415 35945 -385
rect 35975 -415 35995 -385
rect 35925 -425 35995 -415
rect 36010 -335 36080 -325
rect 36010 -365 36030 -335
rect 36060 -365 36080 -335
rect 36010 -385 36080 -365
rect 36010 -415 36030 -385
rect 36060 -415 36080 -385
rect 36010 -425 36080 -415
rect 36095 -335 36165 -325
rect 36095 -365 36115 -335
rect 36145 -365 36165 -335
rect 36095 -385 36165 -365
rect 36095 -415 36115 -385
rect 36145 -415 36165 -385
rect 36095 -425 36165 -415
rect 36180 -335 36250 -325
rect 36180 -365 36200 -335
rect 36230 -365 36250 -335
rect 36180 -385 36250 -365
rect 36180 -415 36200 -385
rect 36230 -415 36250 -385
rect 36180 -425 36250 -415
rect 36265 -335 36335 -325
rect 36265 -365 36285 -335
rect 36315 -365 36335 -335
rect 36265 -385 36335 -365
rect 36265 -415 36285 -385
rect 36315 -415 36335 -385
rect 36265 -425 36335 -415
rect 36350 -335 36420 -325
rect 36350 -365 36370 -335
rect 36400 -365 36420 -335
rect 36350 -385 36420 -365
rect 36350 -415 36370 -385
rect 36400 -415 36420 -385
rect 36350 -425 36420 -415
rect 36435 -335 36505 -325
rect 36435 -365 36455 -335
rect 36485 -365 36505 -335
rect 36435 -385 36505 -365
rect 36435 -415 36455 -385
rect 36485 -415 36505 -385
rect 36435 -425 36505 -415
rect 36520 -335 36590 -325
rect 36520 -365 36540 -335
rect 36570 -365 36590 -335
rect 36520 -385 36590 -365
rect 36520 -415 36540 -385
rect 36570 -415 36590 -385
rect 36520 -425 36590 -415
rect 36605 -335 36675 -325
rect 36605 -365 36625 -335
rect 36655 -365 36675 -335
rect 36605 -385 36675 -365
rect 36605 -415 36625 -385
rect 36655 -415 36675 -385
rect 36605 -425 36675 -415
rect 36690 -335 36760 -325
rect 36690 -365 36710 -335
rect 36740 -365 36760 -335
rect 36690 -385 36760 -365
rect 36690 -415 36710 -385
rect 36740 -415 36760 -385
rect 36690 -425 36760 -415
rect 36775 -335 36845 -325
rect 36775 -365 36795 -335
rect 36825 -365 36845 -335
rect 36775 -385 36845 -365
rect 36775 -415 36795 -385
rect 36825 -415 36845 -385
rect 36775 -425 36845 -415
rect 36860 -335 36930 -325
rect 36860 -365 36880 -335
rect 36910 -365 36930 -335
rect 36860 -385 36930 -365
rect 36860 -415 36880 -385
rect 36910 -415 36930 -385
rect 36860 -425 36930 -415
rect 36945 -335 37015 -325
rect 36945 -365 36965 -335
rect 36995 -365 37015 -335
rect 36945 -385 37015 -365
rect 36945 -415 36965 -385
rect 36995 -415 37015 -385
rect 36945 -425 37015 -415
rect 37030 -335 37100 -325
rect 37030 -365 37050 -335
rect 37080 -365 37100 -335
rect 37030 -385 37100 -365
rect 37030 -415 37050 -385
rect 37080 -415 37100 -385
rect 37030 -425 37100 -415
rect 37115 -335 37185 -325
rect 37115 -365 37135 -335
rect 37165 -365 37185 -335
rect 37115 -385 37185 -365
rect 37115 -415 37135 -385
rect 37165 -415 37185 -385
rect 37115 -425 37185 -415
rect 37200 -335 37270 -325
rect 37200 -365 37220 -335
rect 37250 -365 37270 -335
rect 37200 -385 37270 -365
rect 37200 -415 37220 -385
rect 37250 -415 37270 -385
rect 37200 -425 37270 -415
rect 37285 -335 37355 -325
rect 37285 -365 37305 -335
rect 37335 -365 37355 -335
rect 37285 -385 37355 -365
rect 37285 -415 37305 -385
rect 37335 -415 37355 -385
rect 37285 -425 37355 -415
rect 37370 -335 37440 -325
rect 37370 -365 37390 -335
rect 37420 -365 37440 -335
rect 37370 -385 37440 -365
rect 37370 -415 37390 -385
rect 37420 -415 37440 -385
rect 37370 -425 37440 -415
rect 37455 -335 37525 -325
rect 37455 -365 37475 -335
rect 37505 -365 37525 -335
rect 37455 -385 37525 -365
rect 37455 -415 37475 -385
rect 37505 -415 37525 -385
rect 37455 -425 37525 -415
rect 37540 -335 37610 -325
rect 37540 -365 37560 -335
rect 37590 -365 37610 -335
rect 37540 -385 37610 -365
rect 37540 -415 37560 -385
rect 37590 -415 37610 -385
rect 37540 -425 37610 -415
rect 37625 -335 37695 -325
rect 37625 -365 37645 -335
rect 37675 -365 37695 -335
rect 37625 -385 37695 -365
rect 37625 -415 37645 -385
rect 37675 -415 37695 -385
rect 37625 -425 37695 -415
rect 37710 -335 37780 -325
rect 37710 -365 37730 -335
rect 37760 -365 37780 -335
rect 37710 -385 37780 -365
rect 37710 -415 37730 -385
rect 37760 -415 37780 -385
rect 37710 -425 37780 -415
rect 37795 -335 37865 -325
rect 37795 -365 37815 -335
rect 37845 -365 37865 -335
rect 37795 -385 37865 -365
rect 37795 -415 37815 -385
rect 37845 -415 37865 -385
rect 37795 -425 37865 -415
rect 37880 -335 37950 -325
rect 37880 -365 37900 -335
rect 37930 -365 37950 -335
rect 37880 -385 37950 -365
rect 37880 -415 37900 -385
rect 37930 -415 37950 -385
rect 37880 -425 37950 -415
rect 37965 -335 38035 -325
rect 37965 -365 37985 -335
rect 38015 -365 38035 -335
rect 37965 -385 38035 -365
rect 37965 -415 37985 -385
rect 38015 -415 38035 -385
rect 37965 -425 38035 -415
rect 38050 -335 38120 -325
rect 38050 -365 38070 -335
rect 38100 -365 38120 -335
rect 38050 -385 38120 -365
rect 38050 -415 38070 -385
rect 38100 -415 38120 -385
rect 38050 -425 38120 -415
rect 38135 -335 38205 -325
rect 38135 -365 38155 -335
rect 38185 -365 38205 -335
rect 38135 -385 38205 -365
rect 38135 -415 38155 -385
rect 38185 -415 38205 -385
rect 38135 -425 38205 -415
rect 38220 -335 38290 -325
rect 38220 -365 38240 -335
rect 38270 -365 38290 -335
rect 38220 -385 38290 -365
rect 38220 -415 38240 -385
rect 38270 -415 38290 -385
rect 38220 -425 38290 -415
rect 38305 -335 38375 -325
rect 38305 -365 38325 -335
rect 38355 -365 38375 -335
rect 38305 -385 38375 -365
rect 38305 -415 38325 -385
rect 38355 -415 38375 -385
rect 38305 -425 38375 -415
rect 38390 -335 38460 -325
rect 38390 -365 38410 -335
rect 38440 -365 38460 -335
rect 38390 -385 38460 -365
rect 38390 -415 38410 -385
rect 38440 -415 38460 -385
rect 38390 -425 38460 -415
rect 38475 -335 38545 -325
rect 38475 -365 38495 -335
rect 38525 -365 38545 -335
rect 38475 -385 38545 -365
rect 38475 -415 38495 -385
rect 38525 -415 38545 -385
rect 38475 -425 38545 -415
rect 38560 -335 38630 -325
rect 38560 -365 38580 -335
rect 38610 -365 38630 -335
rect 38560 -385 38630 -365
rect 38560 -415 38580 -385
rect 38610 -415 38630 -385
rect 38560 -425 38630 -415
rect 38645 -335 38715 -325
rect 38645 -365 38665 -335
rect 38695 -365 38715 -335
rect 38645 -385 38715 -365
rect 38645 -415 38665 -385
rect 38695 -415 38715 -385
rect 38645 -425 38715 -415
rect 38730 -335 38800 -325
rect 38730 -365 38750 -335
rect 38780 -365 38800 -335
rect 38730 -385 38800 -365
rect 38730 -415 38750 -385
rect 38780 -415 38800 -385
rect 38730 -425 38800 -415
rect 38815 -335 38885 -325
rect 38815 -365 38835 -335
rect 38865 -365 38885 -335
rect 38815 -385 38885 -365
rect 38815 -415 38835 -385
rect 38865 -415 38885 -385
rect 38815 -425 38885 -415
rect 38900 -335 38970 -325
rect 38900 -365 38920 -335
rect 38950 -365 38970 -335
rect 38900 -385 38970 -365
rect 38900 -415 38920 -385
rect 38950 -415 38970 -385
rect 38900 -425 38970 -415
rect 38985 -335 39055 -325
rect 38985 -365 39005 -335
rect 39035 -365 39055 -335
rect 38985 -385 39055 -365
rect 38985 -415 39005 -385
rect 39035 -415 39055 -385
rect 38985 -425 39055 -415
rect 39070 -335 39140 -325
rect 39070 -365 39090 -335
rect 39120 -365 39140 -335
rect 39070 -385 39140 -365
rect 39070 -415 39090 -385
rect 39120 -415 39140 -385
rect 39070 -425 39140 -415
rect 39155 -335 39225 -325
rect 39155 -365 39175 -335
rect 39205 -365 39225 -335
rect 39155 -385 39225 -365
rect 39155 -415 39175 -385
rect 39205 -415 39225 -385
rect 39155 -425 39225 -415
rect 39240 -335 39310 -325
rect 39240 -365 39260 -335
rect 39290 -365 39310 -335
rect 39240 -385 39310 -365
rect 39240 -415 39260 -385
rect 39290 -415 39310 -385
rect 39240 -425 39310 -415
rect 39325 -335 39395 -325
rect 39325 -365 39345 -335
rect 39375 -365 39395 -335
rect 39325 -385 39395 -365
rect 39325 -415 39345 -385
rect 39375 -415 39395 -385
rect 39325 -425 39395 -415
rect 39410 -335 39480 -325
rect 39410 -365 39430 -335
rect 39460 -365 39480 -335
rect 39410 -385 39480 -365
rect 39410 -415 39430 -385
rect 39460 -415 39480 -385
rect 39410 -425 39480 -415
rect 39495 -335 39565 -325
rect 39495 -365 39515 -335
rect 39545 -365 39565 -335
rect 39495 -385 39565 -365
rect 39495 -415 39515 -385
rect 39545 -415 39565 -385
rect 39495 -425 39565 -415
rect 39580 -335 39650 -325
rect 39580 -365 39600 -335
rect 39630 -365 39650 -335
rect 39580 -385 39650 -365
rect 39580 -415 39600 -385
rect 39630 -415 39650 -385
rect 39580 -425 39650 -415
rect 39665 -335 39735 -325
rect 39665 -365 39685 -335
rect 39715 -365 39735 -335
rect 39665 -385 39735 -365
rect 39665 -415 39685 -385
rect 39715 -415 39735 -385
rect 39665 -425 39735 -415
rect 39750 -335 39820 -325
rect 39750 -365 39770 -335
rect 39800 -365 39820 -335
rect 39750 -385 39820 -365
rect 39750 -415 39770 -385
rect 39800 -415 39820 -385
rect 39750 -425 39820 -415
rect 39835 -335 39905 -325
rect 39835 -365 39855 -335
rect 39885 -365 39905 -335
rect 39835 -385 39905 -365
rect 39835 -415 39855 -385
rect 39885 -415 39905 -385
rect 39835 -425 39905 -415
rect 39920 -335 39990 -325
rect 39920 -365 39940 -335
rect 39970 -365 39990 -335
rect 39920 -385 39990 -365
rect 39920 -415 39940 -385
rect 39970 -415 39990 -385
rect 39920 -425 39990 -415
rect 40005 -335 40075 -325
rect 40005 -365 40025 -335
rect 40055 -365 40075 -335
rect 40005 -385 40075 -365
rect 40005 -415 40025 -385
rect 40055 -415 40075 -385
rect 40005 -425 40075 -415
rect 40090 -335 40160 -325
rect 40090 -365 40110 -335
rect 40140 -365 40160 -335
rect 40090 -385 40160 -365
rect 40090 -415 40110 -385
rect 40140 -415 40160 -385
rect 40090 -425 40160 -415
rect 40175 -335 40245 -325
rect 40175 -365 40195 -335
rect 40225 -365 40245 -335
rect 40175 -385 40245 -365
rect 40175 -415 40195 -385
rect 40225 -415 40245 -385
rect 40175 -425 40245 -415
rect 40260 -335 40330 -325
rect 40260 -365 40280 -335
rect 40310 -365 40330 -335
rect 40260 -385 40330 -365
rect 40260 -415 40280 -385
rect 40310 -415 40330 -385
rect 40260 -425 40330 -415
rect 40345 -335 40415 -325
rect 40345 -365 40365 -335
rect 40395 -365 40415 -335
rect 40345 -385 40415 -365
rect 40345 -415 40365 -385
rect 40395 -415 40415 -385
rect 40345 -425 40415 -415
rect 40430 -335 40500 -325
rect 40430 -365 40450 -335
rect 40480 -365 40500 -335
rect 40430 -385 40500 -365
rect 40430 -415 40450 -385
rect 40480 -415 40500 -385
rect 40430 -425 40500 -415
rect 40515 -335 40585 -325
rect 40515 -365 40535 -335
rect 40565 -365 40585 -335
rect 40515 -385 40585 -365
rect 40515 -415 40535 -385
rect 40565 -415 40585 -385
rect 40515 -425 40585 -415
rect 40600 -335 40670 -325
rect 40600 -365 40620 -335
rect 40650 -365 40670 -335
rect 40600 -385 40670 -365
rect 40600 -415 40620 -385
rect 40650 -415 40670 -385
rect 40600 -425 40670 -415
rect 40685 -335 40755 -325
rect 40685 -365 40705 -335
rect 40735 -365 40755 -335
rect 40685 -385 40755 -365
rect 40685 -415 40705 -385
rect 40735 -415 40755 -385
rect 40685 -425 40755 -415
rect 40770 -335 40840 -325
rect 40770 -365 40790 -335
rect 40820 -365 40840 -335
rect 40770 -385 40840 -365
rect 40770 -415 40790 -385
rect 40820 -415 40840 -385
rect 40770 -425 40840 -415
rect 40855 -335 40925 -325
rect 40855 -365 40875 -335
rect 40905 -365 40925 -335
rect 40855 -385 40925 -365
rect 40855 -415 40875 -385
rect 40905 -415 40925 -385
rect 40855 -425 40925 -415
rect 40940 -335 41010 -325
rect 40940 -365 40960 -335
rect 40990 -365 41010 -335
rect 40940 -385 41010 -365
rect 40940 -415 40960 -385
rect 40990 -415 41010 -385
rect 40940 -425 41010 -415
rect 41025 -335 41095 -325
rect 41025 -365 41045 -335
rect 41075 -365 41095 -335
rect 41025 -385 41095 -365
rect 41025 -415 41045 -385
rect 41075 -415 41095 -385
rect 41025 -425 41095 -415
rect 41110 -335 41180 -325
rect 41110 -365 41130 -335
rect 41160 -365 41180 -335
rect 41110 -385 41180 -365
rect 41110 -415 41130 -385
rect 41160 -415 41180 -385
rect 41110 -425 41180 -415
rect 41195 -335 41265 -325
rect 41195 -365 41215 -335
rect 41245 -365 41265 -335
rect 41195 -385 41265 -365
rect 41195 -415 41215 -385
rect 41245 -415 41265 -385
rect 41195 -425 41265 -415
rect 41280 -335 41350 -325
rect 41280 -365 41300 -335
rect 41330 -365 41350 -335
rect 41280 -385 41350 -365
rect 41280 -415 41300 -385
rect 41330 -415 41350 -385
rect 41280 -425 41350 -415
rect 41365 -335 41435 -325
rect 41365 -365 41385 -335
rect 41415 -365 41435 -335
rect 41365 -385 41435 -365
rect 41365 -415 41385 -385
rect 41415 -415 41435 -385
rect 41365 -425 41435 -415
rect 41450 -335 41520 -325
rect 41450 -365 41470 -335
rect 41500 -365 41520 -335
rect 41450 -385 41520 -365
rect 41450 -415 41470 -385
rect 41500 -415 41520 -385
rect 41450 -425 41520 -415
rect 41535 -335 41605 -325
rect 41535 -365 41555 -335
rect 41585 -365 41605 -335
rect 41535 -385 41605 -365
rect 41535 -415 41555 -385
rect 41585 -415 41605 -385
rect 41535 -425 41605 -415
rect 41620 -335 41690 -325
rect 41620 -365 41640 -335
rect 41670 -365 41690 -335
rect 41620 -385 41690 -365
rect 41620 -415 41640 -385
rect 41670 -415 41690 -385
rect 41620 -425 41690 -415
rect 41705 -335 41775 -325
rect 41705 -365 41725 -335
rect 41755 -365 41775 -335
rect 41705 -385 41775 -365
rect 41705 -415 41725 -385
rect 41755 -415 41775 -385
rect 41705 -425 41775 -415
rect 41790 -335 41860 -325
rect 41790 -365 41810 -335
rect 41840 -365 41860 -335
rect 41790 -385 41860 -365
rect 41790 -415 41810 -385
rect 41840 -415 41860 -385
rect 41790 -425 41860 -415
rect 41875 -335 41945 -325
rect 41875 -365 41895 -335
rect 41925 -365 41945 -335
rect 41875 -385 41945 -365
rect 41875 -415 41895 -385
rect 41925 -415 41945 -385
rect 41875 -425 41945 -415
rect 41960 -335 42030 -325
rect 41960 -365 41980 -335
rect 42010 -365 42030 -335
rect 41960 -385 42030 -365
rect 41960 -415 41980 -385
rect 42010 -415 42030 -385
rect 41960 -425 42030 -415
rect 42045 -335 42115 -325
rect 42045 -365 42065 -335
rect 42095 -365 42115 -335
rect 42045 -385 42115 -365
rect 42045 -415 42065 -385
rect 42095 -415 42115 -385
rect 42045 -425 42115 -415
rect 42130 -335 42200 -325
rect 42130 -365 42150 -335
rect 42180 -365 42200 -335
rect 42130 -385 42200 -365
rect 42130 -415 42150 -385
rect 42180 -415 42200 -385
rect 42130 -425 42200 -415
rect 42215 -335 42285 -325
rect 42215 -365 42235 -335
rect 42265 -365 42285 -335
rect 42215 -385 42285 -365
rect 42215 -415 42235 -385
rect 42265 -415 42285 -385
rect 42215 -425 42285 -415
rect 42300 -335 42370 -325
rect 42300 -365 42320 -335
rect 42350 -365 42370 -335
rect 42300 -385 42370 -365
rect 42300 -415 42320 -385
rect 42350 -415 42370 -385
rect 42300 -425 42370 -415
rect 42385 -335 42455 -325
rect 42385 -365 42405 -335
rect 42435 -365 42455 -335
rect 42385 -385 42455 -365
rect 42385 -415 42405 -385
rect 42435 -415 42455 -385
rect 42385 -425 42455 -415
rect 42470 -335 42540 -325
rect 42470 -365 42490 -335
rect 42520 -365 42540 -335
rect 42470 -385 42540 -365
rect 42470 -415 42490 -385
rect 42520 -415 42540 -385
rect 42470 -425 42540 -415
rect 42555 -335 42625 -325
rect 42555 -365 42575 -335
rect 42605 -365 42625 -335
rect 42555 -385 42625 -365
rect 42555 -415 42575 -385
rect 42605 -415 42625 -385
rect 42555 -425 42625 -415
rect 42640 -335 42710 -325
rect 42640 -365 42660 -335
rect 42690 -365 42710 -335
rect 42640 -385 42710 -365
rect 42640 -415 42660 -385
rect 42690 -415 42710 -385
rect 42640 -425 42710 -415
rect 42725 -335 42795 -325
rect 42725 -365 42745 -335
rect 42775 -365 42795 -335
rect 42725 -385 42795 -365
rect 42725 -415 42745 -385
rect 42775 -415 42795 -385
rect 42725 -425 42795 -415
rect 42810 -335 42880 -325
rect 42810 -365 42830 -335
rect 42860 -365 42880 -335
rect 42810 -385 42880 -365
rect 42810 -415 42830 -385
rect 42860 -415 42880 -385
rect 42810 -425 42880 -415
rect 42895 -335 42965 -325
rect 42895 -365 42915 -335
rect 42945 -365 42965 -335
rect 42895 -385 42965 -365
rect 42895 -415 42915 -385
rect 42945 -415 42965 -385
rect 42895 -425 42965 -415
rect 42980 -335 43050 -325
rect 42980 -365 43000 -335
rect 43030 -365 43050 -335
rect 42980 -385 43050 -365
rect 42980 -415 43000 -385
rect 43030 -415 43050 -385
rect 42980 -425 43050 -415
rect 43065 -335 43135 -325
rect 43065 -365 43085 -335
rect 43115 -365 43135 -335
rect 43065 -385 43135 -365
rect 43065 -415 43085 -385
rect 43115 -415 43135 -385
rect 43065 -425 43135 -415
rect 43150 -335 43220 -325
rect 43150 -365 43170 -335
rect 43200 -365 43220 -335
rect 43150 -385 43220 -365
rect 43150 -415 43170 -385
rect 43200 -415 43220 -385
rect 43150 -425 43220 -415
rect 43235 -335 43305 -325
rect 43235 -365 43255 -335
rect 43285 -365 43305 -335
rect 43235 -385 43305 -365
rect 43235 -415 43255 -385
rect 43285 -415 43305 -385
rect 43235 -425 43305 -415
rect 43320 -335 43390 -325
rect 43320 -365 43340 -335
rect 43370 -365 43390 -335
rect 43320 -385 43390 -365
rect 43320 -415 43340 -385
rect 43370 -415 43390 -385
rect 43320 -425 43390 -415
rect 43405 -335 43475 -325
rect 43405 -365 43425 -335
rect 43455 -365 43475 -335
rect 43405 -385 43475 -365
rect 43405 -415 43425 -385
rect 43455 -415 43475 -385
rect 43405 -425 43475 -415
rect 43490 -335 43560 -325
rect 43490 -365 43510 -335
rect 43540 -365 43560 -335
rect 43490 -385 43560 -365
rect 43490 -415 43510 -385
rect 43540 -415 43560 -385
rect 43490 -425 43560 -415
rect 43575 -335 43645 -325
rect 43575 -365 43595 -335
rect 43625 -365 43645 -335
rect 43575 -385 43645 -365
rect 43575 -415 43595 -385
rect 43625 -415 43645 -385
rect 43575 -425 43645 -415
<< pdiff >>
rect -5 205 65 215
rect -5 175 15 205
rect 45 175 65 205
rect -5 155 65 175
rect -5 125 15 155
rect 45 125 65 155
rect -5 115 65 125
rect 80 205 150 215
rect 80 175 100 205
rect 130 175 150 205
rect 80 155 150 175
rect 80 125 100 155
rect 130 125 150 155
rect 80 115 150 125
rect 205 205 275 215
rect 205 175 225 205
rect 255 175 275 205
rect 205 155 275 175
rect 205 125 225 155
rect 255 125 275 155
rect 205 115 275 125
rect 290 205 360 215
rect 290 175 310 205
rect 340 175 360 205
rect 290 155 360 175
rect 290 125 310 155
rect 340 125 360 155
rect 290 115 360 125
rect 375 205 445 215
rect 375 175 395 205
rect 425 175 445 205
rect 375 155 445 175
rect 375 125 395 155
rect 425 125 445 155
rect 375 115 445 125
rect 460 205 530 215
rect 460 175 480 205
rect 510 175 530 205
rect 460 155 530 175
rect 460 125 480 155
rect 510 125 530 155
rect 460 115 530 125
rect 545 205 615 215
rect 545 175 565 205
rect 595 175 615 205
rect 545 155 615 175
rect 545 125 565 155
rect 595 125 615 155
rect 545 115 615 125
rect 740 205 810 215
rect 740 175 760 205
rect 790 175 810 205
rect 740 155 810 175
rect 740 125 760 155
rect 790 125 810 155
rect 740 115 810 125
rect 825 205 895 215
rect 825 175 845 205
rect 875 175 895 205
rect 825 155 895 175
rect 825 125 845 155
rect 875 125 895 155
rect 825 115 895 125
rect 910 205 980 215
rect 910 175 930 205
rect 960 175 980 205
rect 910 155 980 175
rect 910 125 930 155
rect 960 125 980 155
rect 910 115 980 125
rect 995 205 1065 215
rect 995 175 1015 205
rect 1045 175 1065 205
rect 995 155 1065 175
rect 995 125 1015 155
rect 1045 125 1065 155
rect 995 115 1065 125
rect 1080 205 1150 215
rect 1080 175 1100 205
rect 1130 175 1150 205
rect 1080 155 1150 175
rect 1080 125 1100 155
rect 1130 125 1150 155
rect 1080 115 1150 125
rect 1165 205 1235 215
rect 1165 175 1185 205
rect 1215 175 1235 205
rect 1165 155 1235 175
rect 1165 125 1185 155
rect 1215 125 1235 155
rect 1165 115 1235 125
rect 1250 205 1320 215
rect 1250 175 1270 205
rect 1300 175 1320 205
rect 1250 155 1320 175
rect 1250 125 1270 155
rect 1300 125 1320 155
rect 1250 115 1320 125
rect 1335 205 1405 215
rect 1335 175 1355 205
rect 1385 175 1405 205
rect 1335 155 1405 175
rect 1335 125 1355 155
rect 1385 125 1405 155
rect 1335 115 1405 125
rect 1420 205 1490 215
rect 1420 175 1440 205
rect 1470 175 1490 205
rect 1420 155 1490 175
rect 1420 125 1440 155
rect 1470 125 1490 155
rect 1420 115 1490 125
rect 1505 205 1575 215
rect 1505 175 1525 205
rect 1555 175 1575 205
rect 1505 155 1575 175
rect 1505 125 1525 155
rect 1555 125 1575 155
rect 1505 115 1575 125
rect 1590 205 1660 215
rect 1590 175 1610 205
rect 1640 175 1660 205
rect 1590 155 1660 175
rect 1590 125 1610 155
rect 1640 125 1660 155
rect 1590 115 1660 125
rect 1675 205 1745 215
rect 1675 175 1695 205
rect 1725 175 1745 205
rect 1675 155 1745 175
rect 1675 125 1695 155
rect 1725 125 1745 155
rect 1675 115 1745 125
rect 1760 205 1830 215
rect 1760 175 1780 205
rect 1810 175 1830 205
rect 1760 155 1830 175
rect 1760 125 1780 155
rect 1810 125 1830 155
rect 1760 115 1830 125
rect 1845 205 1915 215
rect 1845 175 1865 205
rect 1895 175 1915 205
rect 1845 155 1915 175
rect 1845 125 1865 155
rect 1895 125 1915 155
rect 1845 115 1915 125
rect 1930 205 2000 215
rect 1930 175 1950 205
rect 1980 175 2000 205
rect 1930 155 2000 175
rect 1930 125 1950 155
rect 1980 125 2000 155
rect 1930 115 2000 125
rect 2015 205 2085 215
rect 2015 175 2035 205
rect 2065 175 2085 205
rect 2015 155 2085 175
rect 2015 125 2035 155
rect 2065 125 2085 155
rect 2015 115 2085 125
rect 2100 205 2170 215
rect 2100 175 2120 205
rect 2150 175 2170 205
rect 2100 155 2170 175
rect 2100 125 2120 155
rect 2150 125 2170 155
rect 2100 115 2170 125
rect 2250 205 2320 215
rect 2250 175 2270 205
rect 2300 175 2320 205
rect 2250 155 2320 175
rect 2250 125 2270 155
rect 2300 125 2320 155
rect 2250 115 2320 125
rect 2335 205 2405 215
rect 2335 175 2355 205
rect 2385 175 2405 205
rect 2335 155 2405 175
rect 2335 125 2355 155
rect 2385 125 2405 155
rect 2335 115 2405 125
rect 2420 205 2490 215
rect 2420 175 2440 205
rect 2470 175 2490 205
rect 2420 155 2490 175
rect 2420 125 2440 155
rect 2470 125 2490 155
rect 2420 115 2490 125
rect 2505 205 2575 215
rect 2505 175 2525 205
rect 2555 175 2575 205
rect 2505 155 2575 175
rect 2505 125 2525 155
rect 2555 125 2575 155
rect 2505 115 2575 125
rect 2590 205 2660 215
rect 2590 175 2610 205
rect 2640 175 2660 205
rect 2590 155 2660 175
rect 2590 125 2610 155
rect 2640 125 2660 155
rect 2590 115 2660 125
rect 2675 205 2745 215
rect 2675 175 2695 205
rect 2725 175 2745 205
rect 2675 155 2745 175
rect 2675 125 2695 155
rect 2725 125 2745 155
rect 2675 115 2745 125
rect 2760 205 2830 215
rect 2760 175 2780 205
rect 2810 175 2830 205
rect 2760 155 2830 175
rect 2760 125 2780 155
rect 2810 125 2830 155
rect 2760 115 2830 125
rect 2845 205 2915 215
rect 2845 175 2865 205
rect 2895 175 2915 205
rect 2845 155 2915 175
rect 2845 125 2865 155
rect 2895 125 2915 155
rect 2845 115 2915 125
rect 2930 205 3000 215
rect 2930 175 2950 205
rect 2980 175 3000 205
rect 2930 155 3000 175
rect 2930 125 2950 155
rect 2980 125 3000 155
rect 2930 115 3000 125
rect 3015 205 3085 215
rect 3015 175 3035 205
rect 3065 175 3085 205
rect 3015 155 3085 175
rect 3015 125 3035 155
rect 3065 125 3085 155
rect 3015 115 3085 125
rect 3100 205 3170 215
rect 3100 175 3120 205
rect 3150 175 3170 205
rect 3100 155 3170 175
rect 3100 125 3120 155
rect 3150 125 3170 155
rect 3100 115 3170 125
rect 3185 205 3255 215
rect 3185 175 3205 205
rect 3235 175 3255 205
rect 3185 155 3255 175
rect 3185 125 3205 155
rect 3235 125 3255 155
rect 3185 115 3255 125
rect 3270 205 3340 215
rect 3270 175 3290 205
rect 3320 175 3340 205
rect 3270 155 3340 175
rect 3270 125 3290 155
rect 3320 125 3340 155
rect 3270 115 3340 125
rect 3355 205 3425 215
rect 3355 175 3375 205
rect 3405 175 3425 205
rect 3355 155 3425 175
rect 3355 125 3375 155
rect 3405 125 3425 155
rect 3355 115 3425 125
rect 3440 205 3510 215
rect 3440 175 3460 205
rect 3490 175 3510 205
rect 3440 155 3510 175
rect 3440 125 3460 155
rect 3490 125 3510 155
rect 3440 115 3510 125
rect 3525 205 3595 215
rect 3525 175 3545 205
rect 3575 175 3595 205
rect 3525 155 3595 175
rect 3525 125 3545 155
rect 3575 125 3595 155
rect 3525 115 3595 125
rect 3610 205 3680 215
rect 3610 175 3630 205
rect 3660 175 3680 205
rect 3610 155 3680 175
rect 3610 125 3630 155
rect 3660 125 3680 155
rect 3610 115 3680 125
rect 3695 205 3765 215
rect 3695 175 3715 205
rect 3745 175 3765 205
rect 3695 155 3765 175
rect 3695 125 3715 155
rect 3745 125 3765 155
rect 3695 115 3765 125
rect 3780 205 3850 215
rect 3780 175 3800 205
rect 3830 175 3850 205
rect 3780 155 3850 175
rect 3780 125 3800 155
rect 3830 125 3850 155
rect 3780 115 3850 125
rect 3865 205 3935 215
rect 3865 175 3885 205
rect 3915 175 3935 205
rect 3865 155 3935 175
rect 3865 125 3885 155
rect 3915 125 3935 155
rect 3865 115 3935 125
rect 3950 205 4020 215
rect 3950 175 3970 205
rect 4000 175 4020 205
rect 3950 155 4020 175
rect 3950 125 3970 155
rect 4000 125 4020 155
rect 3950 115 4020 125
rect 4035 205 4105 215
rect 4035 175 4055 205
rect 4085 175 4105 205
rect 4035 155 4105 175
rect 4035 125 4055 155
rect 4085 125 4105 155
rect 4035 115 4105 125
rect 4120 205 4190 215
rect 4120 175 4140 205
rect 4170 175 4190 205
rect 4120 155 4190 175
rect 4120 125 4140 155
rect 4170 125 4190 155
rect 4120 115 4190 125
rect 4205 205 4275 215
rect 4205 175 4225 205
rect 4255 175 4275 205
rect 4205 155 4275 175
rect 4205 125 4225 155
rect 4255 125 4275 155
rect 4205 115 4275 125
rect 4290 205 4360 215
rect 4290 175 4310 205
rect 4340 175 4360 205
rect 4290 155 4360 175
rect 4290 125 4310 155
rect 4340 125 4360 155
rect 4290 115 4360 125
rect 4375 205 4445 215
rect 4375 175 4395 205
rect 4425 175 4445 205
rect 4375 155 4445 175
rect 4375 125 4395 155
rect 4425 125 4445 155
rect 4375 115 4445 125
rect 4460 205 4530 215
rect 4460 175 4480 205
rect 4510 175 4530 205
rect 4460 155 4530 175
rect 4460 125 4480 155
rect 4510 125 4530 155
rect 4460 115 4530 125
rect 4545 205 4615 215
rect 4545 175 4565 205
rect 4595 175 4615 205
rect 4545 155 4615 175
rect 4545 125 4565 155
rect 4595 125 4615 155
rect 4545 115 4615 125
rect 4630 205 4700 215
rect 4630 175 4650 205
rect 4680 175 4700 205
rect 4630 155 4700 175
rect 4630 125 4650 155
rect 4680 125 4700 155
rect 4630 115 4700 125
rect 4715 205 4785 215
rect 4715 175 4735 205
rect 4765 175 4785 205
rect 4715 155 4785 175
rect 4715 125 4735 155
rect 4765 125 4785 155
rect 4715 115 4785 125
rect 4800 205 4870 215
rect 4800 175 4820 205
rect 4850 175 4870 205
rect 4800 155 4870 175
rect 4800 125 4820 155
rect 4850 125 4870 155
rect 4800 115 4870 125
rect 4885 205 4955 215
rect 4885 175 4905 205
rect 4935 175 4955 205
rect 4885 155 4955 175
rect 4885 125 4905 155
rect 4935 125 4955 155
rect 4885 115 4955 125
rect 4970 205 5040 215
rect 4970 175 4990 205
rect 5020 175 5040 205
rect 4970 155 5040 175
rect 4970 125 4990 155
rect 5020 125 5040 155
rect 4970 115 5040 125
rect 5055 205 5125 215
rect 5055 175 5075 205
rect 5105 175 5125 205
rect 5055 155 5125 175
rect 5055 125 5075 155
rect 5105 125 5125 155
rect 5055 115 5125 125
rect 5140 205 5210 215
rect 5140 175 5160 205
rect 5190 175 5210 205
rect 5140 155 5210 175
rect 5140 125 5160 155
rect 5190 125 5210 155
rect 5140 115 5210 125
rect 5225 205 5295 215
rect 5225 175 5245 205
rect 5275 175 5295 205
rect 5225 155 5295 175
rect 5225 125 5245 155
rect 5275 125 5295 155
rect 5225 115 5295 125
rect 5310 205 5380 215
rect 5310 175 5330 205
rect 5360 175 5380 205
rect 5310 155 5380 175
rect 5310 125 5330 155
rect 5360 125 5380 155
rect 5310 115 5380 125
rect 5395 205 5465 215
rect 5395 175 5415 205
rect 5445 175 5465 205
rect 5395 155 5465 175
rect 5395 125 5415 155
rect 5445 125 5465 155
rect 5395 115 5465 125
rect 5480 205 5550 215
rect 5480 175 5500 205
rect 5530 175 5550 205
rect 5480 155 5550 175
rect 5480 125 5500 155
rect 5530 125 5550 155
rect 5480 115 5550 125
rect 5565 205 5635 215
rect 5565 175 5585 205
rect 5615 175 5635 205
rect 5565 155 5635 175
rect 5565 125 5585 155
rect 5615 125 5635 155
rect 5565 115 5635 125
rect 5650 205 5720 215
rect 5650 175 5670 205
rect 5700 175 5720 205
rect 5650 155 5720 175
rect 5650 125 5670 155
rect 5700 125 5720 155
rect 5650 115 5720 125
rect 5735 205 5805 215
rect 5735 175 5755 205
rect 5785 175 5805 205
rect 5735 155 5805 175
rect 5735 125 5755 155
rect 5785 125 5805 155
rect 5735 115 5805 125
rect 5820 205 5890 215
rect 5820 175 5840 205
rect 5870 175 5890 205
rect 5820 155 5890 175
rect 5820 125 5840 155
rect 5870 125 5890 155
rect 5820 115 5890 125
rect 5905 205 5975 215
rect 5905 175 5925 205
rect 5955 175 5975 205
rect 5905 155 5975 175
rect 5905 125 5925 155
rect 5955 125 5975 155
rect 5905 115 5975 125
rect 5990 205 6060 215
rect 5990 175 6010 205
rect 6040 175 6060 205
rect 5990 155 6060 175
rect 5990 125 6010 155
rect 6040 125 6060 155
rect 5990 115 6060 125
rect 6075 205 6145 215
rect 6075 175 6095 205
rect 6125 175 6145 205
rect 6075 155 6145 175
rect 6075 125 6095 155
rect 6125 125 6145 155
rect 6075 115 6145 125
rect 6160 205 6230 215
rect 6160 175 6180 205
rect 6210 175 6230 205
rect 6160 155 6230 175
rect 6160 125 6180 155
rect 6210 125 6230 155
rect 6160 115 6230 125
rect 6245 205 6315 215
rect 6245 175 6265 205
rect 6295 175 6315 205
rect 6245 155 6315 175
rect 6245 125 6265 155
rect 6295 125 6315 155
rect 6245 115 6315 125
rect 6330 205 6400 215
rect 6330 175 6350 205
rect 6380 175 6400 205
rect 6330 155 6400 175
rect 6330 125 6350 155
rect 6380 125 6400 155
rect 6330 115 6400 125
rect 6415 205 6485 215
rect 6415 175 6435 205
rect 6465 175 6485 205
rect 6415 155 6485 175
rect 6415 125 6435 155
rect 6465 125 6485 155
rect 6415 115 6485 125
rect 6500 205 6570 215
rect 6500 175 6520 205
rect 6550 175 6570 205
rect 6500 155 6570 175
rect 6500 125 6520 155
rect 6550 125 6570 155
rect 6500 115 6570 125
rect 6585 205 6655 215
rect 6585 175 6605 205
rect 6635 175 6655 205
rect 6585 155 6655 175
rect 6585 125 6605 155
rect 6635 125 6655 155
rect 6585 115 6655 125
rect 6670 205 6740 215
rect 6670 175 6690 205
rect 6720 175 6740 205
rect 6670 155 6740 175
rect 6670 125 6690 155
rect 6720 125 6740 155
rect 6670 115 6740 125
rect 6755 205 6825 215
rect 6755 175 6775 205
rect 6805 175 6825 205
rect 6755 155 6825 175
rect 6755 125 6775 155
rect 6805 125 6825 155
rect 6755 115 6825 125
rect 6840 205 6910 215
rect 6840 175 6860 205
rect 6890 175 6910 205
rect 6840 155 6910 175
rect 6840 125 6860 155
rect 6890 125 6910 155
rect 6840 115 6910 125
rect 6925 205 6995 215
rect 6925 175 6945 205
rect 6975 175 6995 205
rect 6925 155 6995 175
rect 6925 125 6945 155
rect 6975 125 6995 155
rect 6925 115 6995 125
rect 7010 205 7080 215
rect 7010 175 7030 205
rect 7060 175 7080 205
rect 7010 155 7080 175
rect 7010 125 7030 155
rect 7060 125 7080 155
rect 7010 115 7080 125
rect 7095 205 7165 215
rect 7095 175 7115 205
rect 7145 175 7165 205
rect 7095 155 7165 175
rect 7095 125 7115 155
rect 7145 125 7165 155
rect 7095 115 7165 125
rect 7180 205 7250 215
rect 7180 175 7200 205
rect 7230 175 7250 205
rect 7180 155 7250 175
rect 7180 125 7200 155
rect 7230 125 7250 155
rect 7180 115 7250 125
rect 7265 205 7335 215
rect 7265 175 7285 205
rect 7315 175 7335 205
rect 7265 155 7335 175
rect 7265 125 7285 155
rect 7315 125 7335 155
rect 7265 115 7335 125
rect 7350 205 7420 215
rect 7350 175 7370 205
rect 7400 175 7420 205
rect 7350 155 7420 175
rect 7350 125 7370 155
rect 7400 125 7420 155
rect 7350 115 7420 125
rect 7435 205 7505 215
rect 7435 175 7455 205
rect 7485 175 7505 205
rect 7435 155 7505 175
rect 7435 125 7455 155
rect 7485 125 7505 155
rect 7435 115 7505 125
rect 7520 205 7590 215
rect 7520 175 7540 205
rect 7570 175 7590 205
rect 7520 155 7590 175
rect 7520 125 7540 155
rect 7570 125 7590 155
rect 7520 115 7590 125
rect 7605 205 7675 215
rect 7605 175 7625 205
rect 7655 175 7675 205
rect 7605 155 7675 175
rect 7605 125 7625 155
rect 7655 125 7675 155
rect 7605 115 7675 125
rect 7690 205 7760 215
rect 7690 175 7710 205
rect 7740 175 7760 205
rect 7690 155 7760 175
rect 7690 125 7710 155
rect 7740 125 7760 155
rect 7690 115 7760 125
rect 7840 205 7910 215
rect 7840 175 7860 205
rect 7890 175 7910 205
rect 7840 155 7910 175
rect 7840 125 7860 155
rect 7890 125 7910 155
rect 7840 115 7910 125
rect 7925 205 7995 215
rect 7925 175 7945 205
rect 7975 175 7995 205
rect 7925 155 7995 175
rect 7925 125 7945 155
rect 7975 125 7995 155
rect 7925 115 7995 125
rect 8010 205 8080 215
rect 8010 175 8030 205
rect 8060 175 8080 205
rect 8010 155 8080 175
rect 8010 125 8030 155
rect 8060 125 8080 155
rect 8010 115 8080 125
rect 8095 205 8165 215
rect 8095 175 8115 205
rect 8145 175 8165 205
rect 8095 155 8165 175
rect 8095 125 8115 155
rect 8145 125 8165 155
rect 8095 115 8165 125
rect 8180 205 8250 215
rect 8180 175 8200 205
rect 8230 175 8250 205
rect 8180 155 8250 175
rect 8180 125 8200 155
rect 8230 125 8250 155
rect 8180 115 8250 125
rect 8265 205 8335 215
rect 8265 175 8285 205
rect 8315 175 8335 205
rect 8265 155 8335 175
rect 8265 125 8285 155
rect 8315 125 8335 155
rect 8265 115 8335 125
rect 8350 205 8420 215
rect 8350 175 8370 205
rect 8400 175 8420 205
rect 8350 155 8420 175
rect 8350 125 8370 155
rect 8400 125 8420 155
rect 8350 115 8420 125
rect 8435 205 8505 215
rect 8435 175 8455 205
rect 8485 175 8505 205
rect 8435 155 8505 175
rect 8435 125 8455 155
rect 8485 125 8505 155
rect 8435 115 8505 125
rect 8520 205 8590 215
rect 8520 175 8540 205
rect 8570 175 8590 205
rect 8520 155 8590 175
rect 8520 125 8540 155
rect 8570 125 8590 155
rect 8520 115 8590 125
rect 8605 205 8675 215
rect 8605 175 8625 205
rect 8655 175 8675 205
rect 8605 155 8675 175
rect 8605 125 8625 155
rect 8655 125 8675 155
rect 8605 115 8675 125
rect 8690 205 8760 215
rect 8690 175 8710 205
rect 8740 175 8760 205
rect 8690 155 8760 175
rect 8690 125 8710 155
rect 8740 125 8760 155
rect 8690 115 8760 125
rect 8775 205 8845 215
rect 8775 175 8795 205
rect 8825 175 8845 205
rect 8775 155 8845 175
rect 8775 125 8795 155
rect 8825 125 8845 155
rect 8775 115 8845 125
rect 8860 205 8930 215
rect 8860 175 8880 205
rect 8910 175 8930 205
rect 8860 155 8930 175
rect 8860 125 8880 155
rect 8910 125 8930 155
rect 8860 115 8930 125
rect 8945 205 9015 215
rect 8945 175 8965 205
rect 8995 175 9015 205
rect 8945 155 9015 175
rect 8945 125 8965 155
rect 8995 125 9015 155
rect 8945 115 9015 125
rect 9030 205 9100 215
rect 9030 175 9050 205
rect 9080 175 9100 205
rect 9030 155 9100 175
rect 9030 125 9050 155
rect 9080 125 9100 155
rect 9030 115 9100 125
rect 9115 205 9185 215
rect 9115 175 9135 205
rect 9165 175 9185 205
rect 9115 155 9185 175
rect 9115 125 9135 155
rect 9165 125 9185 155
rect 9115 115 9185 125
rect 9200 205 9270 215
rect 9200 175 9220 205
rect 9250 175 9270 205
rect 9200 155 9270 175
rect 9200 125 9220 155
rect 9250 125 9270 155
rect 9200 115 9270 125
rect 9285 205 9355 215
rect 9285 175 9305 205
rect 9335 175 9355 205
rect 9285 155 9355 175
rect 9285 125 9305 155
rect 9335 125 9355 155
rect 9285 115 9355 125
rect 9370 205 9440 215
rect 9370 175 9390 205
rect 9420 175 9440 205
rect 9370 155 9440 175
rect 9370 125 9390 155
rect 9420 125 9440 155
rect 9370 115 9440 125
rect 9455 205 9525 215
rect 9455 175 9475 205
rect 9505 175 9525 205
rect 9455 155 9525 175
rect 9455 125 9475 155
rect 9505 125 9525 155
rect 9455 115 9525 125
rect 9540 205 9610 215
rect 9540 175 9560 205
rect 9590 175 9610 205
rect 9540 155 9610 175
rect 9540 125 9560 155
rect 9590 125 9610 155
rect 9540 115 9610 125
rect 9625 205 9695 215
rect 9625 175 9645 205
rect 9675 175 9695 205
rect 9625 155 9695 175
rect 9625 125 9645 155
rect 9675 125 9695 155
rect 9625 115 9695 125
rect 9710 205 9780 215
rect 9710 175 9730 205
rect 9760 175 9780 205
rect 9710 155 9780 175
rect 9710 125 9730 155
rect 9760 125 9780 155
rect 9710 115 9780 125
rect 9795 205 9865 215
rect 9795 175 9815 205
rect 9845 175 9865 205
rect 9795 155 9865 175
rect 9795 125 9815 155
rect 9845 125 9865 155
rect 9795 115 9865 125
rect 9880 205 9950 215
rect 9880 175 9900 205
rect 9930 175 9950 205
rect 9880 155 9950 175
rect 9880 125 9900 155
rect 9930 125 9950 155
rect 9880 115 9950 125
rect 9965 205 10035 215
rect 9965 175 9985 205
rect 10015 175 10035 205
rect 9965 155 10035 175
rect 9965 125 9985 155
rect 10015 125 10035 155
rect 9965 115 10035 125
rect 10050 205 10120 215
rect 10050 175 10070 205
rect 10100 175 10120 205
rect 10050 155 10120 175
rect 10050 125 10070 155
rect 10100 125 10120 155
rect 10050 115 10120 125
rect 10135 205 10205 215
rect 10135 175 10155 205
rect 10185 175 10205 205
rect 10135 155 10205 175
rect 10135 125 10155 155
rect 10185 125 10205 155
rect 10135 115 10205 125
rect 10220 205 10290 215
rect 10220 175 10240 205
rect 10270 175 10290 205
rect 10220 155 10290 175
rect 10220 125 10240 155
rect 10270 125 10290 155
rect 10220 115 10290 125
rect 10305 205 10375 215
rect 10305 175 10325 205
rect 10355 175 10375 205
rect 10305 155 10375 175
rect 10305 125 10325 155
rect 10355 125 10375 155
rect 10305 115 10375 125
rect 10390 205 10460 215
rect 10390 175 10410 205
rect 10440 175 10460 205
rect 10390 155 10460 175
rect 10390 125 10410 155
rect 10440 125 10460 155
rect 10390 115 10460 125
rect 10475 205 10545 215
rect 10475 175 10495 205
rect 10525 175 10545 205
rect 10475 155 10545 175
rect 10475 125 10495 155
rect 10525 125 10545 155
rect 10475 115 10545 125
rect 10560 205 10630 215
rect 10560 175 10580 205
rect 10610 175 10630 205
rect 10560 155 10630 175
rect 10560 125 10580 155
rect 10610 125 10630 155
rect 10560 115 10630 125
rect 10645 205 10715 215
rect 10645 175 10665 205
rect 10695 175 10715 205
rect 10645 155 10715 175
rect 10645 125 10665 155
rect 10695 125 10715 155
rect 10645 115 10715 125
rect 10730 205 10800 215
rect 10730 175 10750 205
rect 10780 175 10800 205
rect 10730 155 10800 175
rect 10730 125 10750 155
rect 10780 125 10800 155
rect 10730 115 10800 125
rect 10815 205 10885 215
rect 10815 175 10835 205
rect 10865 175 10885 205
rect 10815 155 10885 175
rect 10815 125 10835 155
rect 10865 125 10885 155
rect 10815 115 10885 125
rect 10900 205 10970 215
rect 10900 175 10920 205
rect 10950 175 10970 205
rect 10900 155 10970 175
rect 10900 125 10920 155
rect 10950 125 10970 155
rect 10900 115 10970 125
rect 10985 205 11055 215
rect 10985 175 11005 205
rect 11035 175 11055 205
rect 10985 155 11055 175
rect 10985 125 11005 155
rect 11035 125 11055 155
rect 10985 115 11055 125
rect 11070 205 11140 215
rect 11070 175 11090 205
rect 11120 175 11140 205
rect 11070 155 11140 175
rect 11070 125 11090 155
rect 11120 125 11140 155
rect 11070 115 11140 125
rect 11155 205 11225 215
rect 11155 175 11175 205
rect 11205 175 11225 205
rect 11155 155 11225 175
rect 11155 125 11175 155
rect 11205 125 11225 155
rect 11155 115 11225 125
rect 11240 205 11310 215
rect 11240 175 11260 205
rect 11290 175 11310 205
rect 11240 155 11310 175
rect 11240 125 11260 155
rect 11290 125 11310 155
rect 11240 115 11310 125
rect 11325 205 11395 215
rect 11325 175 11345 205
rect 11375 175 11395 205
rect 11325 155 11395 175
rect 11325 125 11345 155
rect 11375 125 11395 155
rect 11325 115 11395 125
rect 11410 205 11480 215
rect 11410 175 11430 205
rect 11460 175 11480 205
rect 11410 155 11480 175
rect 11410 125 11430 155
rect 11460 125 11480 155
rect 11410 115 11480 125
rect 11495 205 11565 215
rect 11495 175 11515 205
rect 11545 175 11565 205
rect 11495 155 11565 175
rect 11495 125 11515 155
rect 11545 125 11565 155
rect 11495 115 11565 125
rect 11580 205 11650 215
rect 11580 175 11600 205
rect 11630 175 11650 205
rect 11580 155 11650 175
rect 11580 125 11600 155
rect 11630 125 11650 155
rect 11580 115 11650 125
rect 11665 205 11735 215
rect 11665 175 11685 205
rect 11715 175 11735 205
rect 11665 155 11735 175
rect 11665 125 11685 155
rect 11715 125 11735 155
rect 11665 115 11735 125
rect 11750 205 11820 215
rect 11750 175 11770 205
rect 11800 175 11820 205
rect 11750 155 11820 175
rect 11750 125 11770 155
rect 11800 125 11820 155
rect 11750 115 11820 125
rect 11835 205 11905 215
rect 11835 175 11855 205
rect 11885 175 11905 205
rect 11835 155 11905 175
rect 11835 125 11855 155
rect 11885 125 11905 155
rect 11835 115 11905 125
rect 11920 205 11990 215
rect 11920 175 11940 205
rect 11970 175 11990 205
rect 11920 155 11990 175
rect 11920 125 11940 155
rect 11970 125 11990 155
rect 11920 115 11990 125
rect 12005 205 12075 215
rect 12005 175 12025 205
rect 12055 175 12075 205
rect 12005 155 12075 175
rect 12005 125 12025 155
rect 12055 125 12075 155
rect 12005 115 12075 125
rect 12090 205 12160 215
rect 12090 175 12110 205
rect 12140 175 12160 205
rect 12090 155 12160 175
rect 12090 125 12110 155
rect 12140 125 12160 155
rect 12090 115 12160 125
rect 12175 205 12245 215
rect 12175 175 12195 205
rect 12225 175 12245 205
rect 12175 155 12245 175
rect 12175 125 12195 155
rect 12225 125 12245 155
rect 12175 115 12245 125
rect 12260 205 12330 215
rect 12260 175 12280 205
rect 12310 175 12330 205
rect 12260 155 12330 175
rect 12260 125 12280 155
rect 12310 125 12330 155
rect 12260 115 12330 125
rect 12345 205 12415 215
rect 12345 175 12365 205
rect 12395 175 12415 205
rect 12345 155 12415 175
rect 12345 125 12365 155
rect 12395 125 12415 155
rect 12345 115 12415 125
rect 12430 205 12500 215
rect 12430 175 12450 205
rect 12480 175 12500 205
rect 12430 155 12500 175
rect 12430 125 12450 155
rect 12480 125 12500 155
rect 12430 115 12500 125
rect 12515 205 12585 215
rect 12515 175 12535 205
rect 12565 175 12585 205
rect 12515 155 12585 175
rect 12515 125 12535 155
rect 12565 125 12585 155
rect 12515 115 12585 125
rect 12600 205 12670 215
rect 12600 175 12620 205
rect 12650 175 12670 205
rect 12600 155 12670 175
rect 12600 125 12620 155
rect 12650 125 12670 155
rect 12600 115 12670 125
rect 12685 205 12755 215
rect 12685 175 12705 205
rect 12735 175 12755 205
rect 12685 155 12755 175
rect 12685 125 12705 155
rect 12735 125 12755 155
rect 12685 115 12755 125
rect 12770 205 12840 215
rect 12770 175 12790 205
rect 12820 175 12840 205
rect 12770 155 12840 175
rect 12770 125 12790 155
rect 12820 125 12840 155
rect 12770 115 12840 125
rect 12855 205 12925 215
rect 12855 175 12875 205
rect 12905 175 12925 205
rect 12855 155 12925 175
rect 12855 125 12875 155
rect 12905 125 12925 155
rect 12855 115 12925 125
rect 12940 205 13010 215
rect 12940 175 12960 205
rect 12990 175 13010 205
rect 12940 155 13010 175
rect 12940 125 12960 155
rect 12990 125 13010 155
rect 12940 115 13010 125
rect 13025 205 13095 215
rect 13025 175 13045 205
rect 13075 175 13095 205
rect 13025 155 13095 175
rect 13025 125 13045 155
rect 13075 125 13095 155
rect 13025 115 13095 125
rect 13110 205 13180 215
rect 13110 175 13130 205
rect 13160 175 13180 205
rect 13110 155 13180 175
rect 13110 125 13130 155
rect 13160 125 13180 155
rect 13110 115 13180 125
rect 13195 205 13265 215
rect 13195 175 13215 205
rect 13245 175 13265 205
rect 13195 155 13265 175
rect 13195 125 13215 155
rect 13245 125 13265 155
rect 13195 115 13265 125
rect 13280 205 13350 215
rect 13280 175 13300 205
rect 13330 175 13350 205
rect 13280 155 13350 175
rect 13280 125 13300 155
rect 13330 125 13350 155
rect 13280 115 13350 125
rect 13365 205 13435 215
rect 13365 175 13385 205
rect 13415 175 13435 205
rect 13365 155 13435 175
rect 13365 125 13385 155
rect 13415 125 13435 155
rect 13365 115 13435 125
rect 13450 205 13520 215
rect 13450 175 13470 205
rect 13500 175 13520 205
rect 13450 155 13520 175
rect 13450 125 13470 155
rect 13500 125 13520 155
rect 13450 115 13520 125
rect 13535 205 13605 215
rect 13535 175 13555 205
rect 13585 175 13605 205
rect 13535 155 13605 175
rect 13535 125 13555 155
rect 13585 125 13605 155
rect 13535 115 13605 125
rect 13620 205 13690 215
rect 13620 175 13640 205
rect 13670 175 13690 205
rect 13620 155 13690 175
rect 13620 125 13640 155
rect 13670 125 13690 155
rect 13620 115 13690 125
rect 13705 205 13775 215
rect 13705 175 13725 205
rect 13755 175 13775 205
rect 13705 155 13775 175
rect 13705 125 13725 155
rect 13755 125 13775 155
rect 13705 115 13775 125
rect 13790 205 13860 215
rect 13790 175 13810 205
rect 13840 175 13860 205
rect 13790 155 13860 175
rect 13790 125 13810 155
rect 13840 125 13860 155
rect 13790 115 13860 125
rect 13875 205 13945 215
rect 13875 175 13895 205
rect 13925 175 13945 205
rect 13875 155 13945 175
rect 13875 125 13895 155
rect 13925 125 13945 155
rect 13875 115 13945 125
rect 13960 205 14030 215
rect 13960 175 13980 205
rect 14010 175 14030 205
rect 13960 155 14030 175
rect 13960 125 13980 155
rect 14010 125 14030 155
rect 13960 115 14030 125
rect 14045 205 14115 215
rect 14045 175 14065 205
rect 14095 175 14115 205
rect 14045 155 14115 175
rect 14045 125 14065 155
rect 14095 125 14115 155
rect 14045 115 14115 125
rect 14130 205 14200 215
rect 14130 175 14150 205
rect 14180 175 14200 205
rect 14130 155 14200 175
rect 14130 125 14150 155
rect 14180 125 14200 155
rect 14130 115 14200 125
rect 14215 205 14285 215
rect 14215 175 14235 205
rect 14265 175 14285 205
rect 14215 155 14285 175
rect 14215 125 14235 155
rect 14265 125 14285 155
rect 14215 115 14285 125
rect 14300 205 14370 215
rect 14300 175 14320 205
rect 14350 175 14370 205
rect 14300 155 14370 175
rect 14300 125 14320 155
rect 14350 125 14370 155
rect 14300 115 14370 125
rect 14385 205 14455 215
rect 14385 175 14405 205
rect 14435 175 14455 205
rect 14385 155 14455 175
rect 14385 125 14405 155
rect 14435 125 14455 155
rect 14385 115 14455 125
rect 14470 205 14540 215
rect 14470 175 14490 205
rect 14520 175 14540 205
rect 14470 155 14540 175
rect 14470 125 14490 155
rect 14520 125 14540 155
rect 14470 115 14540 125
rect 14555 205 14625 215
rect 14555 175 14575 205
rect 14605 175 14625 205
rect 14555 155 14625 175
rect 14555 125 14575 155
rect 14605 125 14625 155
rect 14555 115 14625 125
rect 14640 205 14710 215
rect 14640 175 14660 205
rect 14690 175 14710 205
rect 14640 155 14710 175
rect 14640 125 14660 155
rect 14690 125 14710 155
rect 14640 115 14710 125
rect 14725 205 14795 215
rect 14725 175 14745 205
rect 14775 175 14795 205
rect 14725 155 14795 175
rect 14725 125 14745 155
rect 14775 125 14795 155
rect 14725 115 14795 125
rect 14810 205 14880 215
rect 14810 175 14830 205
rect 14860 175 14880 205
rect 14810 155 14880 175
rect 14810 125 14830 155
rect 14860 125 14880 155
rect 14810 115 14880 125
rect 14895 205 14965 215
rect 14895 175 14915 205
rect 14945 175 14965 205
rect 14895 155 14965 175
rect 14895 125 14915 155
rect 14945 125 14965 155
rect 14895 115 14965 125
rect 14980 205 15050 215
rect 14980 175 15000 205
rect 15030 175 15050 205
rect 14980 155 15050 175
rect 14980 125 15000 155
rect 15030 125 15050 155
rect 14980 115 15050 125
rect 15065 205 15135 215
rect 15065 175 15085 205
rect 15115 175 15135 205
rect 15065 155 15135 175
rect 15065 125 15085 155
rect 15115 125 15135 155
rect 15065 115 15135 125
rect 15150 205 15220 215
rect 15150 175 15170 205
rect 15200 175 15220 205
rect 15150 155 15220 175
rect 15150 125 15170 155
rect 15200 125 15220 155
rect 15150 115 15220 125
rect 15235 205 15305 215
rect 15235 175 15255 205
rect 15285 175 15305 205
rect 15235 155 15305 175
rect 15235 125 15255 155
rect 15285 125 15305 155
rect 15235 115 15305 125
rect 15320 205 15390 215
rect 15320 175 15340 205
rect 15370 175 15390 205
rect 15320 155 15390 175
rect 15320 125 15340 155
rect 15370 125 15390 155
rect 15320 115 15390 125
rect 15405 205 15475 215
rect 15405 175 15425 205
rect 15455 175 15475 205
rect 15405 155 15475 175
rect 15405 125 15425 155
rect 15455 125 15475 155
rect 15405 115 15475 125
rect 15490 205 15560 215
rect 15490 175 15510 205
rect 15540 175 15560 205
rect 15490 155 15560 175
rect 15490 125 15510 155
rect 15540 125 15560 155
rect 15490 115 15560 125
rect 15575 205 15645 215
rect 15575 175 15595 205
rect 15625 175 15645 205
rect 15575 155 15645 175
rect 15575 125 15595 155
rect 15625 125 15645 155
rect 15575 115 15645 125
rect 15660 205 15730 215
rect 15660 175 15680 205
rect 15710 175 15730 205
rect 15660 155 15730 175
rect 15660 125 15680 155
rect 15710 125 15730 155
rect 15660 115 15730 125
rect 15745 205 15815 215
rect 15745 175 15765 205
rect 15795 175 15815 205
rect 15745 155 15815 175
rect 15745 125 15765 155
rect 15795 125 15815 155
rect 15745 115 15815 125
rect 15830 205 15900 215
rect 15830 175 15850 205
rect 15880 175 15900 205
rect 15830 155 15900 175
rect 15830 125 15850 155
rect 15880 125 15900 155
rect 15830 115 15900 125
rect 15915 205 15985 215
rect 15915 175 15935 205
rect 15965 175 15985 205
rect 15915 155 15985 175
rect 15915 125 15935 155
rect 15965 125 15985 155
rect 15915 115 15985 125
rect 16000 205 16070 215
rect 16000 175 16020 205
rect 16050 175 16070 205
rect 16000 155 16070 175
rect 16000 125 16020 155
rect 16050 125 16070 155
rect 16000 115 16070 125
rect 16085 205 16155 215
rect 16085 175 16105 205
rect 16135 175 16155 205
rect 16085 155 16155 175
rect 16085 125 16105 155
rect 16135 125 16155 155
rect 16085 115 16155 125
rect 16170 205 16240 215
rect 16170 175 16190 205
rect 16220 175 16240 205
rect 16170 155 16240 175
rect 16170 125 16190 155
rect 16220 125 16240 155
rect 16170 115 16240 125
rect 16255 205 16325 215
rect 16255 175 16275 205
rect 16305 175 16325 205
rect 16255 155 16325 175
rect 16255 125 16275 155
rect 16305 125 16325 155
rect 16255 115 16325 125
rect 16340 205 16410 215
rect 16340 175 16360 205
rect 16390 175 16410 205
rect 16340 155 16410 175
rect 16340 125 16360 155
rect 16390 125 16410 155
rect 16340 115 16410 125
rect 16425 205 16495 215
rect 16425 175 16445 205
rect 16475 175 16495 205
rect 16425 155 16495 175
rect 16425 125 16445 155
rect 16475 125 16495 155
rect 16425 115 16495 125
rect 16510 205 16580 215
rect 16510 175 16530 205
rect 16560 175 16580 205
rect 16510 155 16580 175
rect 16510 125 16530 155
rect 16560 125 16580 155
rect 16510 115 16580 125
rect 16595 205 16665 215
rect 16595 175 16615 205
rect 16645 175 16665 205
rect 16595 155 16665 175
rect 16595 125 16615 155
rect 16645 125 16665 155
rect 16595 115 16665 125
rect 16680 205 16750 215
rect 16680 175 16700 205
rect 16730 175 16750 205
rect 16680 155 16750 175
rect 16680 125 16700 155
rect 16730 125 16750 155
rect 16680 115 16750 125
rect 16765 205 16835 215
rect 16765 175 16785 205
rect 16815 175 16835 205
rect 16765 155 16835 175
rect 16765 125 16785 155
rect 16815 125 16835 155
rect 16765 115 16835 125
rect 16850 205 16920 215
rect 16850 175 16870 205
rect 16900 175 16920 205
rect 16850 155 16920 175
rect 16850 125 16870 155
rect 16900 125 16920 155
rect 16850 115 16920 125
rect 16935 205 17005 215
rect 16935 175 16955 205
rect 16985 175 17005 205
rect 16935 155 17005 175
rect 16935 125 16955 155
rect 16985 125 17005 155
rect 16935 115 17005 125
rect 17020 205 17090 215
rect 17020 175 17040 205
rect 17070 175 17090 205
rect 17020 155 17090 175
rect 17020 125 17040 155
rect 17070 125 17090 155
rect 17020 115 17090 125
rect 17105 205 17175 215
rect 17105 175 17125 205
rect 17155 175 17175 205
rect 17105 155 17175 175
rect 17105 125 17125 155
rect 17155 125 17175 155
rect 17105 115 17175 125
rect 17190 205 17260 215
rect 17190 175 17210 205
rect 17240 175 17260 205
rect 17190 155 17260 175
rect 17190 125 17210 155
rect 17240 125 17260 155
rect 17190 115 17260 125
rect 17275 205 17345 215
rect 17275 175 17295 205
rect 17325 175 17345 205
rect 17275 155 17345 175
rect 17275 125 17295 155
rect 17325 125 17345 155
rect 17275 115 17345 125
rect 17360 205 17430 215
rect 17360 175 17380 205
rect 17410 175 17430 205
rect 17360 155 17430 175
rect 17360 125 17380 155
rect 17410 125 17430 155
rect 17360 115 17430 125
rect 17445 205 17515 215
rect 17445 175 17465 205
rect 17495 175 17515 205
rect 17445 155 17515 175
rect 17445 125 17465 155
rect 17495 125 17515 155
rect 17445 115 17515 125
rect 17530 205 17600 215
rect 17530 175 17550 205
rect 17580 175 17600 205
rect 17530 155 17600 175
rect 17530 125 17550 155
rect 17580 125 17600 155
rect 17530 115 17600 125
rect 17615 205 17685 215
rect 17615 175 17635 205
rect 17665 175 17685 205
rect 17615 155 17685 175
rect 17615 125 17635 155
rect 17665 125 17685 155
rect 17615 115 17685 125
rect 17700 205 17770 215
rect 17700 175 17720 205
rect 17750 175 17770 205
rect 17700 155 17770 175
rect 17700 125 17720 155
rect 17750 125 17770 155
rect 17700 115 17770 125
rect 17785 205 17855 215
rect 17785 175 17805 205
rect 17835 175 17855 205
rect 17785 155 17855 175
rect 17785 125 17805 155
rect 17835 125 17855 155
rect 17785 115 17855 125
rect 17870 205 17940 215
rect 17870 175 17890 205
rect 17920 175 17940 205
rect 17870 155 17940 175
rect 17870 125 17890 155
rect 17920 125 17940 155
rect 17870 115 17940 125
rect 17955 205 18025 215
rect 17955 175 17975 205
rect 18005 175 18025 205
rect 17955 155 18025 175
rect 17955 125 17975 155
rect 18005 125 18025 155
rect 17955 115 18025 125
rect 18040 205 18110 215
rect 18040 175 18060 205
rect 18090 175 18110 205
rect 18040 155 18110 175
rect 18040 125 18060 155
rect 18090 125 18110 155
rect 18040 115 18110 125
rect 18125 205 18195 215
rect 18125 175 18145 205
rect 18175 175 18195 205
rect 18125 155 18195 175
rect 18125 125 18145 155
rect 18175 125 18195 155
rect 18125 115 18195 125
rect 18210 205 18280 215
rect 18210 175 18230 205
rect 18260 175 18280 205
rect 18210 155 18280 175
rect 18210 125 18230 155
rect 18260 125 18280 155
rect 18210 115 18280 125
rect 18295 205 18365 215
rect 18295 175 18315 205
rect 18345 175 18365 205
rect 18295 155 18365 175
rect 18295 125 18315 155
rect 18345 125 18365 155
rect 18295 115 18365 125
rect 18380 205 18450 215
rect 18380 175 18400 205
rect 18430 175 18450 205
rect 18380 155 18450 175
rect 18380 125 18400 155
rect 18430 125 18450 155
rect 18380 115 18450 125
rect 18465 205 18535 215
rect 18465 175 18485 205
rect 18515 175 18535 205
rect 18465 155 18535 175
rect 18465 125 18485 155
rect 18515 125 18535 155
rect 18465 115 18535 125
rect 18550 205 18620 215
rect 18550 175 18570 205
rect 18600 175 18620 205
rect 18550 155 18620 175
rect 18550 125 18570 155
rect 18600 125 18620 155
rect 18550 115 18620 125
rect 18635 205 18705 215
rect 18635 175 18655 205
rect 18685 175 18705 205
rect 18635 155 18705 175
rect 18635 125 18655 155
rect 18685 125 18705 155
rect 18635 115 18705 125
rect 18720 205 18790 215
rect 18720 175 18740 205
rect 18770 175 18790 205
rect 18720 155 18790 175
rect 18720 125 18740 155
rect 18770 125 18790 155
rect 18720 115 18790 125
rect 18805 205 18875 215
rect 18805 175 18825 205
rect 18855 175 18875 205
rect 18805 155 18875 175
rect 18805 125 18825 155
rect 18855 125 18875 155
rect 18805 115 18875 125
rect 18890 205 18960 215
rect 18890 175 18910 205
rect 18940 175 18960 205
rect 18890 155 18960 175
rect 18890 125 18910 155
rect 18940 125 18960 155
rect 18890 115 18960 125
rect 18975 205 19045 215
rect 18975 175 18995 205
rect 19025 175 19045 205
rect 18975 155 19045 175
rect 18975 125 18995 155
rect 19025 125 19045 155
rect 18975 115 19045 125
rect 19060 205 19130 215
rect 19060 175 19080 205
rect 19110 175 19130 205
rect 19060 155 19130 175
rect 19060 125 19080 155
rect 19110 125 19130 155
rect 19060 115 19130 125
rect 19145 205 19215 215
rect 19145 175 19165 205
rect 19195 175 19215 205
rect 19145 155 19215 175
rect 19145 125 19165 155
rect 19195 125 19215 155
rect 19145 115 19215 125
rect 19230 205 19300 215
rect 19230 175 19250 205
rect 19280 175 19300 205
rect 19230 155 19300 175
rect 19230 125 19250 155
rect 19280 125 19300 155
rect 19230 115 19300 125
rect 19315 205 19385 215
rect 19315 175 19335 205
rect 19365 175 19385 205
rect 19315 155 19385 175
rect 19315 125 19335 155
rect 19365 125 19385 155
rect 19315 115 19385 125
rect 19400 205 19470 215
rect 19400 175 19420 205
rect 19450 175 19470 205
rect 19400 155 19470 175
rect 19400 125 19420 155
rect 19450 125 19470 155
rect 19400 115 19470 125
rect 19485 205 19555 215
rect 19485 175 19505 205
rect 19535 175 19555 205
rect 19485 155 19555 175
rect 19485 125 19505 155
rect 19535 125 19555 155
rect 19485 115 19555 125
rect 19570 205 19640 215
rect 19570 175 19590 205
rect 19620 175 19640 205
rect 19570 155 19640 175
rect 19570 125 19590 155
rect 19620 125 19640 155
rect 19570 115 19640 125
rect 19655 205 19725 215
rect 19655 175 19675 205
rect 19705 175 19725 205
rect 19655 155 19725 175
rect 19655 125 19675 155
rect 19705 125 19725 155
rect 19655 115 19725 125
rect 19740 205 19810 215
rect 19740 175 19760 205
rect 19790 175 19810 205
rect 19740 155 19810 175
rect 19740 125 19760 155
rect 19790 125 19810 155
rect 19740 115 19810 125
rect 19825 205 19895 215
rect 19825 175 19845 205
rect 19875 175 19895 205
rect 19825 155 19895 175
rect 19825 125 19845 155
rect 19875 125 19895 155
rect 19825 115 19895 125
rect 19910 205 19980 215
rect 19910 175 19930 205
rect 19960 175 19980 205
rect 19910 155 19980 175
rect 19910 125 19930 155
rect 19960 125 19980 155
rect 19910 115 19980 125
rect 19995 205 20065 215
rect 19995 175 20015 205
rect 20045 175 20065 205
rect 19995 155 20065 175
rect 19995 125 20015 155
rect 20045 125 20065 155
rect 19995 115 20065 125
rect 20080 205 20150 215
rect 20080 175 20100 205
rect 20130 175 20150 205
rect 20080 155 20150 175
rect 20080 125 20100 155
rect 20130 125 20150 155
rect 20080 115 20150 125
rect 20165 205 20235 215
rect 20165 175 20185 205
rect 20215 175 20235 205
rect 20165 155 20235 175
rect 20165 125 20185 155
rect 20215 125 20235 155
rect 20165 115 20235 125
rect 20250 205 20320 215
rect 20250 175 20270 205
rect 20300 175 20320 205
rect 20250 155 20320 175
rect 20250 125 20270 155
rect 20300 125 20320 155
rect 20250 115 20320 125
rect 20335 205 20405 215
rect 20335 175 20355 205
rect 20385 175 20405 205
rect 20335 155 20405 175
rect 20335 125 20355 155
rect 20385 125 20405 155
rect 20335 115 20405 125
rect 20420 205 20490 215
rect 20420 175 20440 205
rect 20470 175 20490 205
rect 20420 155 20490 175
rect 20420 125 20440 155
rect 20470 125 20490 155
rect 20420 115 20490 125
rect 20505 205 20575 215
rect 20505 175 20525 205
rect 20555 175 20575 205
rect 20505 155 20575 175
rect 20505 125 20525 155
rect 20555 125 20575 155
rect 20505 115 20575 125
rect 20590 205 20660 215
rect 20590 175 20610 205
rect 20640 175 20660 205
rect 20590 155 20660 175
rect 20590 125 20610 155
rect 20640 125 20660 155
rect 20590 115 20660 125
rect 20675 205 20745 215
rect 20675 175 20695 205
rect 20725 175 20745 205
rect 20675 155 20745 175
rect 20675 125 20695 155
rect 20725 125 20745 155
rect 20675 115 20745 125
rect 20760 205 20830 215
rect 20760 175 20780 205
rect 20810 175 20830 205
rect 20760 155 20830 175
rect 20760 125 20780 155
rect 20810 125 20830 155
rect 20760 115 20830 125
rect 20845 205 20915 215
rect 20845 175 20865 205
rect 20895 175 20915 205
rect 20845 155 20915 175
rect 20845 125 20865 155
rect 20895 125 20915 155
rect 20845 115 20915 125
rect 20930 205 21000 215
rect 20930 175 20950 205
rect 20980 175 21000 205
rect 20930 155 21000 175
rect 20930 125 20950 155
rect 20980 125 21000 155
rect 20930 115 21000 125
rect 21015 205 21085 215
rect 21015 175 21035 205
rect 21065 175 21085 205
rect 21015 155 21085 175
rect 21015 125 21035 155
rect 21065 125 21085 155
rect 21015 115 21085 125
rect 21100 205 21170 215
rect 21100 175 21120 205
rect 21150 175 21170 205
rect 21100 155 21170 175
rect 21100 125 21120 155
rect 21150 125 21170 155
rect 21100 115 21170 125
rect 21185 205 21255 215
rect 21185 175 21205 205
rect 21235 175 21255 205
rect 21185 155 21255 175
rect 21185 125 21205 155
rect 21235 125 21255 155
rect 21185 115 21255 125
rect 21270 205 21340 215
rect 21270 175 21290 205
rect 21320 175 21340 205
rect 21270 155 21340 175
rect 21270 125 21290 155
rect 21320 125 21340 155
rect 21270 115 21340 125
rect 21355 205 21425 215
rect 21355 175 21375 205
rect 21405 175 21425 205
rect 21355 155 21425 175
rect 21355 125 21375 155
rect 21405 125 21425 155
rect 21355 115 21425 125
rect 21440 205 21510 215
rect 21440 175 21460 205
rect 21490 175 21510 205
rect 21440 155 21510 175
rect 21440 125 21460 155
rect 21490 125 21510 155
rect 21440 115 21510 125
rect 21525 205 21595 215
rect 21525 175 21545 205
rect 21575 175 21595 205
rect 21525 155 21595 175
rect 21525 125 21545 155
rect 21575 125 21595 155
rect 21525 115 21595 125
rect 21610 205 21680 215
rect 21610 175 21630 205
rect 21660 175 21680 205
rect 21610 155 21680 175
rect 21610 125 21630 155
rect 21660 125 21680 155
rect 21610 115 21680 125
rect 21695 205 21765 215
rect 21695 175 21715 205
rect 21745 175 21765 205
rect 21695 155 21765 175
rect 21695 125 21715 155
rect 21745 125 21765 155
rect 21695 115 21765 125
rect 21780 205 21850 215
rect 21780 175 21800 205
rect 21830 175 21850 205
rect 21780 155 21850 175
rect 21780 125 21800 155
rect 21830 125 21850 155
rect 21780 115 21850 125
rect 21865 205 21935 215
rect 21865 175 21885 205
rect 21915 175 21935 205
rect 21865 155 21935 175
rect 21865 125 21885 155
rect 21915 125 21935 155
rect 21865 115 21935 125
rect 21950 205 22020 215
rect 21950 175 21970 205
rect 22000 175 22020 205
rect 21950 155 22020 175
rect 21950 125 21970 155
rect 22000 125 22020 155
rect 21950 115 22020 125
rect 22035 205 22105 215
rect 22035 175 22055 205
rect 22085 175 22105 205
rect 22035 155 22105 175
rect 22035 125 22055 155
rect 22085 125 22105 155
rect 22035 115 22105 125
rect 22120 205 22190 215
rect 22120 175 22140 205
rect 22170 175 22190 205
rect 22120 155 22190 175
rect 22120 125 22140 155
rect 22170 125 22190 155
rect 22120 115 22190 125
rect 22205 205 22275 215
rect 22205 175 22225 205
rect 22255 175 22275 205
rect 22205 155 22275 175
rect 22205 125 22225 155
rect 22255 125 22275 155
rect 22205 115 22275 125
rect 22290 205 22360 215
rect 22290 175 22310 205
rect 22340 175 22360 205
rect 22290 155 22360 175
rect 22290 125 22310 155
rect 22340 125 22360 155
rect 22290 115 22360 125
rect 22375 205 22445 215
rect 22375 175 22395 205
rect 22425 175 22445 205
rect 22375 155 22445 175
rect 22375 125 22395 155
rect 22425 125 22445 155
rect 22375 115 22445 125
rect 22460 205 22530 215
rect 22460 175 22480 205
rect 22510 175 22530 205
rect 22460 155 22530 175
rect 22460 125 22480 155
rect 22510 125 22530 155
rect 22460 115 22530 125
rect 22545 205 22615 215
rect 22545 175 22565 205
rect 22595 175 22615 205
rect 22545 155 22615 175
rect 22545 125 22565 155
rect 22595 125 22615 155
rect 22545 115 22615 125
rect 22630 205 22700 215
rect 22630 175 22650 205
rect 22680 175 22700 205
rect 22630 155 22700 175
rect 22630 125 22650 155
rect 22680 125 22700 155
rect 22630 115 22700 125
rect 22715 205 22785 215
rect 22715 175 22735 205
rect 22765 175 22785 205
rect 22715 155 22785 175
rect 22715 125 22735 155
rect 22765 125 22785 155
rect 22715 115 22785 125
rect 22800 205 22870 215
rect 22800 175 22820 205
rect 22850 175 22870 205
rect 22800 155 22870 175
rect 22800 125 22820 155
rect 22850 125 22870 155
rect 22800 115 22870 125
rect 22885 205 22955 215
rect 22885 175 22905 205
rect 22935 175 22955 205
rect 22885 155 22955 175
rect 22885 125 22905 155
rect 22935 125 22955 155
rect 22885 115 22955 125
rect 22970 205 23040 215
rect 22970 175 22990 205
rect 23020 175 23040 205
rect 22970 155 23040 175
rect 22970 125 22990 155
rect 23020 125 23040 155
rect 22970 115 23040 125
rect 23055 205 23125 215
rect 23055 175 23075 205
rect 23105 175 23125 205
rect 23055 155 23125 175
rect 23055 125 23075 155
rect 23105 125 23125 155
rect 23055 115 23125 125
rect 23140 205 23210 215
rect 23140 175 23160 205
rect 23190 175 23210 205
rect 23140 155 23210 175
rect 23140 125 23160 155
rect 23190 125 23210 155
rect 23140 115 23210 125
rect 23225 205 23295 215
rect 23225 175 23245 205
rect 23275 175 23295 205
rect 23225 155 23295 175
rect 23225 125 23245 155
rect 23275 125 23295 155
rect 23225 115 23295 125
rect 23310 205 23380 215
rect 23310 175 23330 205
rect 23360 175 23380 205
rect 23310 155 23380 175
rect 23310 125 23330 155
rect 23360 125 23380 155
rect 23310 115 23380 125
rect 23395 205 23465 215
rect 23395 175 23415 205
rect 23445 175 23465 205
rect 23395 155 23465 175
rect 23395 125 23415 155
rect 23445 125 23465 155
rect 23395 115 23465 125
rect 23480 205 23550 215
rect 23480 175 23500 205
rect 23530 175 23550 205
rect 23480 155 23550 175
rect 23480 125 23500 155
rect 23530 125 23550 155
rect 23480 115 23550 125
rect 23565 205 23635 215
rect 23565 175 23585 205
rect 23615 175 23635 205
rect 23565 155 23635 175
rect 23565 125 23585 155
rect 23615 125 23635 155
rect 23565 115 23635 125
rect 23650 205 23720 215
rect 23650 175 23670 205
rect 23700 175 23720 205
rect 23650 155 23720 175
rect 23650 125 23670 155
rect 23700 125 23720 155
rect 23650 115 23720 125
rect 23735 205 23805 215
rect 23735 175 23755 205
rect 23785 175 23805 205
rect 23735 155 23805 175
rect 23735 125 23755 155
rect 23785 125 23805 155
rect 23735 115 23805 125
rect 23820 205 23890 215
rect 23820 175 23840 205
rect 23870 175 23890 205
rect 23820 155 23890 175
rect 23820 125 23840 155
rect 23870 125 23890 155
rect 23820 115 23890 125
rect 23905 205 23975 215
rect 23905 175 23925 205
rect 23955 175 23975 205
rect 23905 155 23975 175
rect 23905 125 23925 155
rect 23955 125 23975 155
rect 23905 115 23975 125
rect 23990 205 24060 215
rect 23990 175 24010 205
rect 24040 175 24060 205
rect 23990 155 24060 175
rect 23990 125 24010 155
rect 24040 125 24060 155
rect 23990 115 24060 125
rect 24075 205 24145 215
rect 24075 175 24095 205
rect 24125 175 24145 205
rect 24075 155 24145 175
rect 24075 125 24095 155
rect 24125 125 24145 155
rect 24075 115 24145 125
rect 24160 205 24230 215
rect 24160 175 24180 205
rect 24210 175 24230 205
rect 24160 155 24230 175
rect 24160 125 24180 155
rect 24210 125 24230 155
rect 24160 115 24230 125
rect 24245 205 24315 215
rect 24245 175 24265 205
rect 24295 175 24315 205
rect 24245 155 24315 175
rect 24245 125 24265 155
rect 24295 125 24315 155
rect 24245 115 24315 125
rect 24330 205 24400 215
rect 24330 175 24350 205
rect 24380 175 24400 205
rect 24330 155 24400 175
rect 24330 125 24350 155
rect 24380 125 24400 155
rect 24330 115 24400 125
rect 24415 205 24485 215
rect 24415 175 24435 205
rect 24465 175 24485 205
rect 24415 155 24485 175
rect 24415 125 24435 155
rect 24465 125 24485 155
rect 24415 115 24485 125
rect 24500 205 24570 215
rect 24500 175 24520 205
rect 24550 175 24570 205
rect 24500 155 24570 175
rect 24500 125 24520 155
rect 24550 125 24570 155
rect 24500 115 24570 125
rect 24585 205 24655 215
rect 24585 175 24605 205
rect 24635 175 24655 205
rect 24585 155 24655 175
rect 24585 125 24605 155
rect 24635 125 24655 155
rect 24585 115 24655 125
rect 24670 205 24740 215
rect 24670 175 24690 205
rect 24720 175 24740 205
rect 24670 155 24740 175
rect 24670 125 24690 155
rect 24720 125 24740 155
rect 24670 115 24740 125
rect 24755 205 24825 215
rect 24755 175 24775 205
rect 24805 175 24825 205
rect 24755 155 24825 175
rect 24755 125 24775 155
rect 24805 125 24825 155
rect 24755 115 24825 125
rect 24840 205 24910 215
rect 24840 175 24860 205
rect 24890 175 24910 205
rect 24840 155 24910 175
rect 24840 125 24860 155
rect 24890 125 24910 155
rect 24840 115 24910 125
rect 24925 205 24995 215
rect 24925 175 24945 205
rect 24975 175 24995 205
rect 24925 155 24995 175
rect 24925 125 24945 155
rect 24975 125 24995 155
rect 24925 115 24995 125
rect 25010 205 25080 215
rect 25010 175 25030 205
rect 25060 175 25080 205
rect 25010 155 25080 175
rect 25010 125 25030 155
rect 25060 125 25080 155
rect 25010 115 25080 125
rect 25095 205 25165 215
rect 25095 175 25115 205
rect 25145 175 25165 205
rect 25095 155 25165 175
rect 25095 125 25115 155
rect 25145 125 25165 155
rect 25095 115 25165 125
rect 25180 205 25250 215
rect 25180 175 25200 205
rect 25230 175 25250 205
rect 25180 155 25250 175
rect 25180 125 25200 155
rect 25230 125 25250 155
rect 25180 115 25250 125
rect 25265 205 25335 215
rect 25265 175 25285 205
rect 25315 175 25335 205
rect 25265 155 25335 175
rect 25265 125 25285 155
rect 25315 125 25335 155
rect 25265 115 25335 125
rect 25350 205 25420 215
rect 25350 175 25370 205
rect 25400 175 25420 205
rect 25350 155 25420 175
rect 25350 125 25370 155
rect 25400 125 25420 155
rect 25350 115 25420 125
rect 25435 205 25505 215
rect 25435 175 25455 205
rect 25485 175 25505 205
rect 25435 155 25505 175
rect 25435 125 25455 155
rect 25485 125 25505 155
rect 25435 115 25505 125
rect 25520 205 25590 215
rect 25520 175 25540 205
rect 25570 175 25590 205
rect 25520 155 25590 175
rect 25520 125 25540 155
rect 25570 125 25590 155
rect 25520 115 25590 125
rect 25605 205 25675 215
rect 25605 175 25625 205
rect 25655 175 25675 205
rect 25605 155 25675 175
rect 25605 125 25625 155
rect 25655 125 25675 155
rect 25605 115 25675 125
rect 25690 205 25760 215
rect 25690 175 25710 205
rect 25740 175 25760 205
rect 25690 155 25760 175
rect 25690 125 25710 155
rect 25740 125 25760 155
rect 25690 115 25760 125
rect 25775 205 25845 215
rect 25775 175 25795 205
rect 25825 175 25845 205
rect 25775 155 25845 175
rect 25775 125 25795 155
rect 25825 125 25845 155
rect 25775 115 25845 125
rect 25860 205 25930 215
rect 25860 175 25880 205
rect 25910 175 25930 205
rect 25860 155 25930 175
rect 25860 125 25880 155
rect 25910 125 25930 155
rect 25860 115 25930 125
rect 25945 205 26015 215
rect 25945 175 25965 205
rect 25995 175 26015 205
rect 25945 155 26015 175
rect 25945 125 25965 155
rect 25995 125 26015 155
rect 25945 115 26015 125
rect 26030 205 26100 215
rect 26030 175 26050 205
rect 26080 175 26100 205
rect 26030 155 26100 175
rect 26030 125 26050 155
rect 26080 125 26100 155
rect 26030 115 26100 125
rect 26115 205 26185 215
rect 26115 175 26135 205
rect 26165 175 26185 205
rect 26115 155 26185 175
rect 26115 125 26135 155
rect 26165 125 26185 155
rect 26115 115 26185 125
rect 26200 205 26270 215
rect 26200 175 26220 205
rect 26250 175 26270 205
rect 26200 155 26270 175
rect 26200 125 26220 155
rect 26250 125 26270 155
rect 26200 115 26270 125
rect 26285 205 26355 215
rect 26285 175 26305 205
rect 26335 175 26355 205
rect 26285 155 26355 175
rect 26285 125 26305 155
rect 26335 125 26355 155
rect 26285 115 26355 125
rect 26370 205 26440 215
rect 26370 175 26390 205
rect 26420 175 26440 205
rect 26370 155 26440 175
rect 26370 125 26390 155
rect 26420 125 26440 155
rect 26370 115 26440 125
rect 26455 205 26525 215
rect 26455 175 26475 205
rect 26505 175 26525 205
rect 26455 155 26525 175
rect 26455 125 26475 155
rect 26505 125 26525 155
rect 26455 115 26525 125
rect 26540 205 26610 215
rect 26540 175 26560 205
rect 26590 175 26610 205
rect 26540 155 26610 175
rect 26540 125 26560 155
rect 26590 125 26610 155
rect 26540 115 26610 125
rect 26625 205 26695 215
rect 26625 175 26645 205
rect 26675 175 26695 205
rect 26625 155 26695 175
rect 26625 125 26645 155
rect 26675 125 26695 155
rect 26625 115 26695 125
rect 26710 205 26780 215
rect 26710 175 26730 205
rect 26760 175 26780 205
rect 26710 155 26780 175
rect 26710 125 26730 155
rect 26760 125 26780 155
rect 26710 115 26780 125
rect 26795 205 26865 215
rect 26795 175 26815 205
rect 26845 175 26865 205
rect 26795 155 26865 175
rect 26795 125 26815 155
rect 26845 125 26865 155
rect 26795 115 26865 125
rect 26880 205 26950 215
rect 26880 175 26900 205
rect 26930 175 26950 205
rect 26880 155 26950 175
rect 26880 125 26900 155
rect 26930 125 26950 155
rect 26880 115 26950 125
rect 26965 205 27035 215
rect 26965 175 26985 205
rect 27015 175 27035 205
rect 26965 155 27035 175
rect 26965 125 26985 155
rect 27015 125 27035 155
rect 26965 115 27035 125
rect 27050 205 27120 215
rect 27050 175 27070 205
rect 27100 175 27120 205
rect 27050 155 27120 175
rect 27050 125 27070 155
rect 27100 125 27120 155
rect 27050 115 27120 125
rect 27135 205 27205 215
rect 27135 175 27155 205
rect 27185 175 27205 205
rect 27135 155 27205 175
rect 27135 125 27155 155
rect 27185 125 27205 155
rect 27135 115 27205 125
rect 27220 205 27290 215
rect 27220 175 27240 205
rect 27270 175 27290 205
rect 27220 155 27290 175
rect 27220 125 27240 155
rect 27270 125 27290 155
rect 27220 115 27290 125
rect 27305 205 27375 215
rect 27305 175 27325 205
rect 27355 175 27375 205
rect 27305 155 27375 175
rect 27305 125 27325 155
rect 27355 125 27375 155
rect 27305 115 27375 125
rect 27390 205 27460 215
rect 27390 175 27410 205
rect 27440 175 27460 205
rect 27390 155 27460 175
rect 27390 125 27410 155
rect 27440 125 27460 155
rect 27390 115 27460 125
rect 27475 205 27545 215
rect 27475 175 27495 205
rect 27525 175 27545 205
rect 27475 155 27545 175
rect 27475 125 27495 155
rect 27525 125 27545 155
rect 27475 115 27545 125
rect 27560 205 27630 215
rect 27560 175 27580 205
rect 27610 175 27630 205
rect 27560 155 27630 175
rect 27560 125 27580 155
rect 27610 125 27630 155
rect 27560 115 27630 125
rect 27645 205 27715 215
rect 27645 175 27665 205
rect 27695 175 27715 205
rect 27645 155 27715 175
rect 27645 125 27665 155
rect 27695 125 27715 155
rect 27645 115 27715 125
rect 27730 205 27800 215
rect 27730 175 27750 205
rect 27780 175 27800 205
rect 27730 155 27800 175
rect 27730 125 27750 155
rect 27780 125 27800 155
rect 27730 115 27800 125
rect 27815 205 27885 215
rect 27815 175 27835 205
rect 27865 175 27885 205
rect 27815 155 27885 175
rect 27815 125 27835 155
rect 27865 125 27885 155
rect 27815 115 27885 125
rect 27900 205 27970 215
rect 27900 175 27920 205
rect 27950 175 27970 205
rect 27900 155 27970 175
rect 27900 125 27920 155
rect 27950 125 27970 155
rect 27900 115 27970 125
rect 27985 205 28055 215
rect 27985 175 28005 205
rect 28035 175 28055 205
rect 27985 155 28055 175
rect 27985 125 28005 155
rect 28035 125 28055 155
rect 27985 115 28055 125
rect 28070 205 28140 215
rect 28070 175 28090 205
rect 28120 175 28140 205
rect 28070 155 28140 175
rect 28070 125 28090 155
rect 28120 125 28140 155
rect 28070 115 28140 125
rect 28155 205 28225 215
rect 28155 175 28175 205
rect 28205 175 28225 205
rect 28155 155 28225 175
rect 28155 125 28175 155
rect 28205 125 28225 155
rect 28155 115 28225 125
rect 28240 205 28310 215
rect 28240 175 28260 205
rect 28290 175 28310 205
rect 28240 155 28310 175
rect 28240 125 28260 155
rect 28290 125 28310 155
rect 28240 115 28310 125
rect 28325 205 28395 215
rect 28325 175 28345 205
rect 28375 175 28395 205
rect 28325 155 28395 175
rect 28325 125 28345 155
rect 28375 125 28395 155
rect 28325 115 28395 125
rect 28410 205 28480 215
rect 28410 175 28430 205
rect 28460 175 28480 205
rect 28410 155 28480 175
rect 28410 125 28430 155
rect 28460 125 28480 155
rect 28410 115 28480 125
rect 28495 205 28565 215
rect 28495 175 28515 205
rect 28545 175 28565 205
rect 28495 155 28565 175
rect 28495 125 28515 155
rect 28545 125 28565 155
rect 28495 115 28565 125
rect 28580 205 28650 215
rect 28580 175 28600 205
rect 28630 175 28650 205
rect 28580 155 28650 175
rect 28580 125 28600 155
rect 28630 125 28650 155
rect 28580 115 28650 125
rect 28665 205 28735 215
rect 28665 175 28685 205
rect 28715 175 28735 205
rect 28665 155 28735 175
rect 28665 125 28685 155
rect 28715 125 28735 155
rect 28665 115 28735 125
rect 28750 205 28820 215
rect 28750 175 28770 205
rect 28800 175 28820 205
rect 28750 155 28820 175
rect 28750 125 28770 155
rect 28800 125 28820 155
rect 28750 115 28820 125
rect 28835 205 28905 215
rect 28835 175 28855 205
rect 28885 175 28905 205
rect 28835 155 28905 175
rect 28835 125 28855 155
rect 28885 125 28905 155
rect 28835 115 28905 125
rect 28920 205 28990 215
rect 28920 175 28940 205
rect 28970 175 28990 205
rect 28920 155 28990 175
rect 28920 125 28940 155
rect 28970 125 28990 155
rect 28920 115 28990 125
rect 29005 205 29075 215
rect 29005 175 29025 205
rect 29055 175 29075 205
rect 29005 155 29075 175
rect 29005 125 29025 155
rect 29055 125 29075 155
rect 29005 115 29075 125
rect 29090 205 29160 215
rect 29090 175 29110 205
rect 29140 175 29160 205
rect 29090 155 29160 175
rect 29090 125 29110 155
rect 29140 125 29160 155
rect 29090 115 29160 125
rect 29175 205 29245 215
rect 29175 175 29195 205
rect 29225 175 29245 205
rect 29175 155 29245 175
rect 29175 125 29195 155
rect 29225 125 29245 155
rect 29175 115 29245 125
rect 29260 205 29330 215
rect 29260 175 29280 205
rect 29310 175 29330 205
rect 29260 155 29330 175
rect 29260 125 29280 155
rect 29310 125 29330 155
rect 29260 115 29330 125
rect 29345 205 29415 215
rect 29345 175 29365 205
rect 29395 175 29415 205
rect 29345 155 29415 175
rect 29345 125 29365 155
rect 29395 125 29415 155
rect 29345 115 29415 125
rect 29430 205 29500 215
rect 29430 175 29450 205
rect 29480 175 29500 205
rect 29430 155 29500 175
rect 29430 125 29450 155
rect 29480 125 29500 155
rect 29430 115 29500 125
rect 29515 205 29585 215
rect 29515 175 29535 205
rect 29565 175 29585 205
rect 29515 155 29585 175
rect 29515 125 29535 155
rect 29565 125 29585 155
rect 29515 115 29585 125
rect 29600 205 29670 215
rect 29600 175 29620 205
rect 29650 175 29670 205
rect 29600 155 29670 175
rect 29600 125 29620 155
rect 29650 125 29670 155
rect 29600 115 29670 125
rect 55 -500 125 -490
rect 55 -530 75 -500
rect 105 -530 125 -500
rect 55 -550 125 -530
rect 55 -580 75 -550
rect 105 -580 125 -550
rect 55 -600 125 -580
rect 55 -630 75 -600
rect 105 -630 125 -600
rect 55 -650 125 -630
rect 55 -680 75 -650
rect 105 -680 125 -650
rect 55 -690 125 -680
rect 140 -500 210 -490
rect 140 -530 160 -500
rect 190 -530 210 -500
rect 140 -550 210 -530
rect 140 -580 160 -550
rect 190 -580 210 -550
rect 140 -600 210 -580
rect 140 -630 160 -600
rect 190 -630 210 -600
rect 140 -650 210 -630
rect 140 -680 160 -650
rect 190 -680 210 -650
rect 140 -690 210 -680
rect 225 -500 295 -490
rect 225 -530 245 -500
rect 275 -530 295 -500
rect 225 -550 295 -530
rect 225 -580 245 -550
rect 275 -580 295 -550
rect 225 -600 295 -580
rect 225 -630 245 -600
rect 275 -630 295 -600
rect 225 -650 295 -630
rect 225 -680 245 -650
rect 275 -680 295 -650
rect 225 -690 295 -680
rect 310 -500 380 -490
rect 310 -530 330 -500
rect 360 -530 380 -500
rect 310 -550 380 -530
rect 310 -580 330 -550
rect 360 -580 380 -550
rect 310 -600 380 -580
rect 310 -630 330 -600
rect 360 -630 380 -600
rect 310 -650 380 -630
rect 310 -680 330 -650
rect 360 -680 380 -650
rect 310 -690 380 -680
rect 395 -500 465 -490
rect 395 -530 415 -500
rect 445 -530 465 -500
rect 395 -550 465 -530
rect 395 -580 415 -550
rect 445 -580 465 -550
rect 395 -600 465 -580
rect 395 -630 415 -600
rect 445 -630 465 -600
rect 395 -650 465 -630
rect 395 -680 415 -650
rect 445 -680 465 -650
rect 395 -690 465 -680
rect 480 -500 550 -490
rect 480 -530 500 -500
rect 530 -530 550 -500
rect 480 -550 550 -530
rect 480 -580 500 -550
rect 530 -580 550 -550
rect 480 -600 550 -580
rect 480 -630 500 -600
rect 530 -630 550 -600
rect 480 -650 550 -630
rect 480 -680 500 -650
rect 530 -680 550 -650
rect 480 -690 550 -680
rect 565 -500 635 -490
rect 565 -530 585 -500
rect 615 -530 635 -500
rect 565 -550 635 -530
rect 565 -580 585 -550
rect 615 -580 635 -550
rect 565 -600 635 -580
rect 565 -630 585 -600
rect 615 -630 635 -600
rect 565 -650 635 -630
rect 565 -680 585 -650
rect 615 -680 635 -650
rect 565 -690 635 -680
rect 650 -500 720 -490
rect 650 -530 670 -500
rect 700 -530 720 -500
rect 650 -550 720 -530
rect 650 -580 670 -550
rect 700 -580 720 -550
rect 650 -600 720 -580
rect 650 -630 670 -600
rect 700 -630 720 -600
rect 650 -650 720 -630
rect 650 -680 670 -650
rect 700 -680 720 -650
rect 650 -690 720 -680
rect 735 -500 805 -490
rect 735 -530 755 -500
rect 785 -530 805 -500
rect 735 -550 805 -530
rect 735 -580 755 -550
rect 785 -580 805 -550
rect 735 -600 805 -580
rect 735 -630 755 -600
rect 785 -630 805 -600
rect 735 -650 805 -630
rect 735 -680 755 -650
rect 785 -680 805 -650
rect 735 -690 805 -680
rect 820 -500 890 -490
rect 820 -530 840 -500
rect 870 -530 890 -500
rect 820 -550 890 -530
rect 820 -580 840 -550
rect 870 -580 890 -550
rect 820 -600 890 -580
rect 820 -630 840 -600
rect 870 -630 890 -600
rect 820 -650 890 -630
rect 820 -680 840 -650
rect 870 -680 890 -650
rect 820 -690 890 -680
rect 905 -500 975 -490
rect 905 -530 925 -500
rect 955 -530 975 -500
rect 905 -550 975 -530
rect 905 -580 925 -550
rect 955 -580 975 -550
rect 905 -600 975 -580
rect 905 -630 925 -600
rect 955 -630 975 -600
rect 905 -650 975 -630
rect 905 -680 925 -650
rect 955 -680 975 -650
rect 905 -690 975 -680
rect 990 -500 1060 -490
rect 990 -530 1010 -500
rect 1040 -530 1060 -500
rect 990 -550 1060 -530
rect 990 -580 1010 -550
rect 1040 -580 1060 -550
rect 990 -600 1060 -580
rect 990 -630 1010 -600
rect 1040 -630 1060 -600
rect 990 -650 1060 -630
rect 990 -680 1010 -650
rect 1040 -680 1060 -650
rect 990 -690 1060 -680
rect 1075 -500 1145 -490
rect 1075 -530 1095 -500
rect 1125 -530 1145 -500
rect 1075 -550 1145 -530
rect 1075 -580 1095 -550
rect 1125 -580 1145 -550
rect 1075 -600 1145 -580
rect 1075 -630 1095 -600
rect 1125 -630 1145 -600
rect 1075 -650 1145 -630
rect 1075 -680 1095 -650
rect 1125 -680 1145 -650
rect 1075 -690 1145 -680
rect 1160 -500 1230 -490
rect 1160 -530 1180 -500
rect 1210 -530 1230 -500
rect 1160 -550 1230 -530
rect 1160 -580 1180 -550
rect 1210 -580 1230 -550
rect 1160 -600 1230 -580
rect 1160 -630 1180 -600
rect 1210 -630 1230 -600
rect 1160 -650 1230 -630
rect 1160 -680 1180 -650
rect 1210 -680 1230 -650
rect 1160 -690 1230 -680
rect 1245 -500 1315 -490
rect 1245 -530 1265 -500
rect 1295 -530 1315 -500
rect 1245 -550 1315 -530
rect 1245 -580 1265 -550
rect 1295 -580 1315 -550
rect 1245 -600 1315 -580
rect 1245 -630 1265 -600
rect 1295 -630 1315 -600
rect 1245 -650 1315 -630
rect 1245 -680 1265 -650
rect 1295 -680 1315 -650
rect 1245 -690 1315 -680
rect 1330 -500 1400 -490
rect 1330 -530 1350 -500
rect 1380 -530 1400 -500
rect 1330 -550 1400 -530
rect 1330 -580 1350 -550
rect 1380 -580 1400 -550
rect 1330 -600 1400 -580
rect 1330 -630 1350 -600
rect 1380 -630 1400 -600
rect 1330 -650 1400 -630
rect 1330 -680 1350 -650
rect 1380 -680 1400 -650
rect 1330 -690 1400 -680
rect 1415 -500 1485 -490
rect 1415 -530 1435 -500
rect 1465 -530 1485 -500
rect 1415 -550 1485 -530
rect 1415 -580 1435 -550
rect 1465 -580 1485 -550
rect 1415 -600 1485 -580
rect 1415 -630 1435 -600
rect 1465 -630 1485 -600
rect 1415 -650 1485 -630
rect 1415 -680 1435 -650
rect 1465 -680 1485 -650
rect 1415 -690 1485 -680
rect 1500 -500 1570 -490
rect 1500 -530 1520 -500
rect 1550 -530 1570 -500
rect 1500 -550 1570 -530
rect 1500 -580 1520 -550
rect 1550 -580 1570 -550
rect 1500 -600 1570 -580
rect 1500 -630 1520 -600
rect 1550 -630 1570 -600
rect 1500 -650 1570 -630
rect 1500 -680 1520 -650
rect 1550 -680 1570 -650
rect 1500 -690 1570 -680
rect 1585 -500 1655 -490
rect 1585 -530 1605 -500
rect 1635 -530 1655 -500
rect 1585 -550 1655 -530
rect 1585 -580 1605 -550
rect 1635 -580 1655 -550
rect 1585 -600 1655 -580
rect 1585 -630 1605 -600
rect 1635 -630 1655 -600
rect 1585 -650 1655 -630
rect 1585 -680 1605 -650
rect 1635 -680 1655 -650
rect 1585 -690 1655 -680
rect 1670 -500 1740 -490
rect 1670 -530 1690 -500
rect 1720 -530 1740 -500
rect 1670 -550 1740 -530
rect 1670 -580 1690 -550
rect 1720 -580 1740 -550
rect 1670 -600 1740 -580
rect 1670 -630 1690 -600
rect 1720 -630 1740 -600
rect 1670 -650 1740 -630
rect 1670 -680 1690 -650
rect 1720 -680 1740 -650
rect 1670 -690 1740 -680
rect 1755 -500 1825 -490
rect 1755 -530 1775 -500
rect 1805 -530 1825 -500
rect 1755 -550 1825 -530
rect 1755 -580 1775 -550
rect 1805 -580 1825 -550
rect 1755 -600 1825 -580
rect 1755 -630 1775 -600
rect 1805 -630 1825 -600
rect 1755 -650 1825 -630
rect 1755 -680 1775 -650
rect 1805 -680 1825 -650
rect 1755 -690 1825 -680
rect 1840 -500 1910 -490
rect 1840 -530 1860 -500
rect 1890 -530 1910 -500
rect 1840 -550 1910 -530
rect 1840 -580 1860 -550
rect 1890 -580 1910 -550
rect 1840 -600 1910 -580
rect 1840 -630 1860 -600
rect 1890 -630 1910 -600
rect 1840 -650 1910 -630
rect 1840 -680 1860 -650
rect 1890 -680 1910 -650
rect 1840 -690 1910 -680
rect 1925 -500 1995 -490
rect 1925 -530 1945 -500
rect 1975 -530 1995 -500
rect 1925 -550 1995 -530
rect 1925 -580 1945 -550
rect 1975 -580 1995 -550
rect 1925 -600 1995 -580
rect 1925 -630 1945 -600
rect 1975 -630 1995 -600
rect 1925 -650 1995 -630
rect 1925 -680 1945 -650
rect 1975 -680 1995 -650
rect 1925 -690 1995 -680
rect 2010 -500 2080 -490
rect 2010 -530 2030 -500
rect 2060 -530 2080 -500
rect 2010 -550 2080 -530
rect 2010 -580 2030 -550
rect 2060 -580 2080 -550
rect 2010 -600 2080 -580
rect 2010 -630 2030 -600
rect 2060 -630 2080 -600
rect 2010 -650 2080 -630
rect 2010 -680 2030 -650
rect 2060 -680 2080 -650
rect 2010 -690 2080 -680
rect 2095 -500 2165 -490
rect 2095 -530 2115 -500
rect 2145 -530 2165 -500
rect 2095 -550 2165 -530
rect 2095 -580 2115 -550
rect 2145 -580 2165 -550
rect 2095 -600 2165 -580
rect 2095 -630 2115 -600
rect 2145 -630 2165 -600
rect 2095 -650 2165 -630
rect 2095 -680 2115 -650
rect 2145 -680 2165 -650
rect 2095 -690 2165 -680
rect 2180 -500 2250 -490
rect 2180 -530 2200 -500
rect 2230 -530 2250 -500
rect 2180 -550 2250 -530
rect 2180 -580 2200 -550
rect 2230 -580 2250 -550
rect 2180 -600 2250 -580
rect 2180 -630 2200 -600
rect 2230 -630 2250 -600
rect 2180 -650 2250 -630
rect 2180 -680 2200 -650
rect 2230 -680 2250 -650
rect 2180 -690 2250 -680
rect 2265 -500 2335 -490
rect 2265 -530 2285 -500
rect 2315 -530 2335 -500
rect 2265 -550 2335 -530
rect 2265 -580 2285 -550
rect 2315 -580 2335 -550
rect 2265 -600 2335 -580
rect 2265 -630 2285 -600
rect 2315 -630 2335 -600
rect 2265 -650 2335 -630
rect 2265 -680 2285 -650
rect 2315 -680 2335 -650
rect 2265 -690 2335 -680
rect 2350 -500 2420 -490
rect 2350 -530 2370 -500
rect 2400 -530 2420 -500
rect 2350 -550 2420 -530
rect 2350 -580 2370 -550
rect 2400 -580 2420 -550
rect 2350 -600 2420 -580
rect 2350 -630 2370 -600
rect 2400 -630 2420 -600
rect 2350 -650 2420 -630
rect 2350 -680 2370 -650
rect 2400 -680 2420 -650
rect 2350 -690 2420 -680
rect 2435 -500 2505 -490
rect 2435 -530 2455 -500
rect 2485 -530 2505 -500
rect 2435 -550 2505 -530
rect 2435 -580 2455 -550
rect 2485 -580 2505 -550
rect 2435 -600 2505 -580
rect 2435 -630 2455 -600
rect 2485 -630 2505 -600
rect 2435 -650 2505 -630
rect 2435 -680 2455 -650
rect 2485 -680 2505 -650
rect 2435 -690 2505 -680
rect 2520 -500 2590 -490
rect 2520 -530 2540 -500
rect 2570 -530 2590 -500
rect 2520 -550 2590 -530
rect 2520 -580 2540 -550
rect 2570 -580 2590 -550
rect 2520 -600 2590 -580
rect 2520 -630 2540 -600
rect 2570 -630 2590 -600
rect 2520 -650 2590 -630
rect 2520 -680 2540 -650
rect 2570 -680 2590 -650
rect 2520 -690 2590 -680
rect 2605 -500 2675 -490
rect 2605 -530 2625 -500
rect 2655 -530 2675 -500
rect 2605 -550 2675 -530
rect 2605 -580 2625 -550
rect 2655 -580 2675 -550
rect 2605 -600 2675 -580
rect 2605 -630 2625 -600
rect 2655 -630 2675 -600
rect 2605 -650 2675 -630
rect 2605 -680 2625 -650
rect 2655 -680 2675 -650
rect 2605 -690 2675 -680
rect 2690 -500 2760 -490
rect 2690 -530 2710 -500
rect 2740 -530 2760 -500
rect 2690 -550 2760 -530
rect 2690 -580 2710 -550
rect 2740 -580 2760 -550
rect 2690 -600 2760 -580
rect 2690 -630 2710 -600
rect 2740 -630 2760 -600
rect 2690 -650 2760 -630
rect 2690 -680 2710 -650
rect 2740 -680 2760 -650
rect 2690 -690 2760 -680
rect 2775 -500 2845 -490
rect 2775 -530 2795 -500
rect 2825 -530 2845 -500
rect 2775 -550 2845 -530
rect 2775 -580 2795 -550
rect 2825 -580 2845 -550
rect 2775 -600 2845 -580
rect 2775 -630 2795 -600
rect 2825 -630 2845 -600
rect 2775 -650 2845 -630
rect 2775 -680 2795 -650
rect 2825 -680 2845 -650
rect 2775 -690 2845 -680
rect 2860 -500 2930 -490
rect 2860 -530 2880 -500
rect 2910 -530 2930 -500
rect 2860 -550 2930 -530
rect 2860 -580 2880 -550
rect 2910 -580 2930 -550
rect 2860 -600 2930 -580
rect 2860 -630 2880 -600
rect 2910 -630 2930 -600
rect 2860 -650 2930 -630
rect 2860 -680 2880 -650
rect 2910 -680 2930 -650
rect 2860 -690 2930 -680
rect 2945 -500 3015 -490
rect 2945 -530 2965 -500
rect 2995 -530 3015 -500
rect 2945 -550 3015 -530
rect 2945 -580 2965 -550
rect 2995 -580 3015 -550
rect 2945 -600 3015 -580
rect 2945 -630 2965 -600
rect 2995 -630 3015 -600
rect 2945 -650 3015 -630
rect 2945 -680 2965 -650
rect 2995 -680 3015 -650
rect 2945 -690 3015 -680
rect 3030 -500 3100 -490
rect 3030 -530 3050 -500
rect 3080 -530 3100 -500
rect 3030 -550 3100 -530
rect 3030 -580 3050 -550
rect 3080 -580 3100 -550
rect 3030 -600 3100 -580
rect 3030 -630 3050 -600
rect 3080 -630 3100 -600
rect 3030 -650 3100 -630
rect 3030 -680 3050 -650
rect 3080 -680 3100 -650
rect 3030 -690 3100 -680
rect 3115 -500 3185 -490
rect 3115 -530 3135 -500
rect 3165 -530 3185 -500
rect 3115 -550 3185 -530
rect 3115 -580 3135 -550
rect 3165 -580 3185 -550
rect 3115 -600 3185 -580
rect 3115 -630 3135 -600
rect 3165 -630 3185 -600
rect 3115 -650 3185 -630
rect 3115 -680 3135 -650
rect 3165 -680 3185 -650
rect 3115 -690 3185 -680
rect 3200 -500 3270 -490
rect 3200 -530 3220 -500
rect 3250 -530 3270 -500
rect 3200 -550 3270 -530
rect 3200 -580 3220 -550
rect 3250 -580 3270 -550
rect 3200 -600 3270 -580
rect 3200 -630 3220 -600
rect 3250 -630 3270 -600
rect 3200 -650 3270 -630
rect 3200 -680 3220 -650
rect 3250 -680 3270 -650
rect 3200 -690 3270 -680
rect 3285 -500 3355 -490
rect 3285 -530 3305 -500
rect 3335 -530 3355 -500
rect 3285 -550 3355 -530
rect 3285 -580 3305 -550
rect 3335 -580 3355 -550
rect 3285 -600 3355 -580
rect 3285 -630 3305 -600
rect 3335 -630 3355 -600
rect 3285 -650 3355 -630
rect 3285 -680 3305 -650
rect 3335 -680 3355 -650
rect 3285 -690 3355 -680
rect 3370 -500 3440 -490
rect 3370 -530 3390 -500
rect 3420 -530 3440 -500
rect 3370 -550 3440 -530
rect 3370 -580 3390 -550
rect 3420 -580 3440 -550
rect 3370 -600 3440 -580
rect 3370 -630 3390 -600
rect 3420 -630 3440 -600
rect 3370 -650 3440 -630
rect 3370 -680 3390 -650
rect 3420 -680 3440 -650
rect 3370 -690 3440 -680
rect 3455 -500 3525 -490
rect 3455 -530 3475 -500
rect 3505 -530 3525 -500
rect 3455 -550 3525 -530
rect 3455 -580 3475 -550
rect 3505 -580 3525 -550
rect 3455 -600 3525 -580
rect 3455 -630 3475 -600
rect 3505 -630 3525 -600
rect 3455 -650 3525 -630
rect 3455 -680 3475 -650
rect 3505 -680 3525 -650
rect 3455 -690 3525 -680
rect 3540 -500 3610 -490
rect 3540 -530 3560 -500
rect 3590 -530 3610 -500
rect 3540 -550 3610 -530
rect 3540 -580 3560 -550
rect 3590 -580 3610 -550
rect 3540 -600 3610 -580
rect 3540 -630 3560 -600
rect 3590 -630 3610 -600
rect 3540 -650 3610 -630
rect 3540 -680 3560 -650
rect 3590 -680 3610 -650
rect 3540 -690 3610 -680
rect 3625 -500 3695 -490
rect 3625 -530 3645 -500
rect 3675 -530 3695 -500
rect 3625 -550 3695 -530
rect 3625 -580 3645 -550
rect 3675 -580 3695 -550
rect 3625 -600 3695 -580
rect 3625 -630 3645 -600
rect 3675 -630 3695 -600
rect 3625 -650 3695 -630
rect 3625 -680 3645 -650
rect 3675 -680 3695 -650
rect 3625 -690 3695 -680
rect 3710 -500 3780 -490
rect 3710 -530 3730 -500
rect 3760 -530 3780 -500
rect 3710 -550 3780 -530
rect 3710 -580 3730 -550
rect 3760 -580 3780 -550
rect 3710 -600 3780 -580
rect 3710 -630 3730 -600
rect 3760 -630 3780 -600
rect 3710 -650 3780 -630
rect 3710 -680 3730 -650
rect 3760 -680 3780 -650
rect 3710 -690 3780 -680
rect 3795 -500 3865 -490
rect 3795 -530 3815 -500
rect 3845 -530 3865 -500
rect 3795 -550 3865 -530
rect 3795 -580 3815 -550
rect 3845 -580 3865 -550
rect 3795 -600 3865 -580
rect 3795 -630 3815 -600
rect 3845 -630 3865 -600
rect 3795 -650 3865 -630
rect 3795 -680 3815 -650
rect 3845 -680 3865 -650
rect 3795 -690 3865 -680
rect 3880 -500 3950 -490
rect 3880 -530 3900 -500
rect 3930 -530 3950 -500
rect 3880 -550 3950 -530
rect 3880 -580 3900 -550
rect 3930 -580 3950 -550
rect 3880 -600 3950 -580
rect 3880 -630 3900 -600
rect 3930 -630 3950 -600
rect 3880 -650 3950 -630
rect 3880 -680 3900 -650
rect 3930 -680 3950 -650
rect 3880 -690 3950 -680
rect 3965 -500 4035 -490
rect 3965 -530 3985 -500
rect 4015 -530 4035 -500
rect 3965 -550 4035 -530
rect 3965 -580 3985 -550
rect 4015 -580 4035 -550
rect 3965 -600 4035 -580
rect 3965 -630 3985 -600
rect 4015 -630 4035 -600
rect 3965 -650 4035 -630
rect 3965 -680 3985 -650
rect 4015 -680 4035 -650
rect 3965 -690 4035 -680
rect 4050 -500 4120 -490
rect 4050 -530 4070 -500
rect 4100 -530 4120 -500
rect 4050 -550 4120 -530
rect 4050 -580 4070 -550
rect 4100 -580 4120 -550
rect 4050 -600 4120 -580
rect 4050 -630 4070 -600
rect 4100 -630 4120 -600
rect 4050 -650 4120 -630
rect 4050 -680 4070 -650
rect 4100 -680 4120 -650
rect 4050 -690 4120 -680
rect 4135 -500 4205 -490
rect 4135 -530 4155 -500
rect 4185 -530 4205 -500
rect 4135 -550 4205 -530
rect 4135 -580 4155 -550
rect 4185 -580 4205 -550
rect 4135 -600 4205 -580
rect 4135 -630 4155 -600
rect 4185 -630 4205 -600
rect 4135 -650 4205 -630
rect 4135 -680 4155 -650
rect 4185 -680 4205 -650
rect 4135 -690 4205 -680
rect 4220 -500 4290 -490
rect 4220 -530 4240 -500
rect 4270 -530 4290 -500
rect 4220 -550 4290 -530
rect 4220 -580 4240 -550
rect 4270 -580 4290 -550
rect 4220 -600 4290 -580
rect 4220 -630 4240 -600
rect 4270 -630 4290 -600
rect 4220 -650 4290 -630
rect 4220 -680 4240 -650
rect 4270 -680 4290 -650
rect 4220 -690 4290 -680
rect 4305 -500 4375 -490
rect 4305 -530 4325 -500
rect 4355 -530 4375 -500
rect 4305 -550 4375 -530
rect 4305 -580 4325 -550
rect 4355 -580 4375 -550
rect 4305 -600 4375 -580
rect 4305 -630 4325 -600
rect 4355 -630 4375 -600
rect 4305 -650 4375 -630
rect 4305 -680 4325 -650
rect 4355 -680 4375 -650
rect 4305 -690 4375 -680
rect 4390 -500 4460 -490
rect 4390 -530 4410 -500
rect 4440 -530 4460 -500
rect 4390 -550 4460 -530
rect 4390 -580 4410 -550
rect 4440 -580 4460 -550
rect 4390 -600 4460 -580
rect 4390 -630 4410 -600
rect 4440 -630 4460 -600
rect 4390 -650 4460 -630
rect 4390 -680 4410 -650
rect 4440 -680 4460 -650
rect 4390 -690 4460 -680
rect 4475 -500 4545 -490
rect 4475 -530 4495 -500
rect 4525 -530 4545 -500
rect 4475 -550 4545 -530
rect 4475 -580 4495 -550
rect 4525 -580 4545 -550
rect 4475 -600 4545 -580
rect 4475 -630 4495 -600
rect 4525 -630 4545 -600
rect 4475 -650 4545 -630
rect 4475 -680 4495 -650
rect 4525 -680 4545 -650
rect 4475 -690 4545 -680
rect 4560 -500 4630 -490
rect 4560 -530 4580 -500
rect 4610 -530 4630 -500
rect 4560 -550 4630 -530
rect 4560 -580 4580 -550
rect 4610 -580 4630 -550
rect 4560 -600 4630 -580
rect 4560 -630 4580 -600
rect 4610 -630 4630 -600
rect 4560 -650 4630 -630
rect 4560 -680 4580 -650
rect 4610 -680 4630 -650
rect 4560 -690 4630 -680
rect 4645 -500 4715 -490
rect 4645 -530 4665 -500
rect 4695 -530 4715 -500
rect 4645 -550 4715 -530
rect 4645 -580 4665 -550
rect 4695 -580 4715 -550
rect 4645 -600 4715 -580
rect 4645 -630 4665 -600
rect 4695 -630 4715 -600
rect 4645 -650 4715 -630
rect 4645 -680 4665 -650
rect 4695 -680 4715 -650
rect 4645 -690 4715 -680
rect 4730 -500 4800 -490
rect 4730 -530 4750 -500
rect 4780 -530 4800 -500
rect 4730 -550 4800 -530
rect 4730 -580 4750 -550
rect 4780 -580 4800 -550
rect 4730 -600 4800 -580
rect 4730 -630 4750 -600
rect 4780 -630 4800 -600
rect 4730 -650 4800 -630
rect 4730 -680 4750 -650
rect 4780 -680 4800 -650
rect 4730 -690 4800 -680
rect 4815 -500 4885 -490
rect 4815 -530 4835 -500
rect 4865 -530 4885 -500
rect 4815 -550 4885 -530
rect 4815 -580 4835 -550
rect 4865 -580 4885 -550
rect 4815 -600 4885 -580
rect 4815 -630 4835 -600
rect 4865 -630 4885 -600
rect 4815 -650 4885 -630
rect 4815 -680 4835 -650
rect 4865 -680 4885 -650
rect 4815 -690 4885 -680
rect 4900 -500 4970 -490
rect 4900 -530 4920 -500
rect 4950 -530 4970 -500
rect 4900 -550 4970 -530
rect 4900 -580 4920 -550
rect 4950 -580 4970 -550
rect 4900 -600 4970 -580
rect 4900 -630 4920 -600
rect 4950 -630 4970 -600
rect 4900 -650 4970 -630
rect 4900 -680 4920 -650
rect 4950 -680 4970 -650
rect 4900 -690 4970 -680
rect 4985 -500 5055 -490
rect 4985 -530 5005 -500
rect 5035 -530 5055 -500
rect 4985 -550 5055 -530
rect 4985 -580 5005 -550
rect 5035 -580 5055 -550
rect 4985 -600 5055 -580
rect 4985 -630 5005 -600
rect 5035 -630 5055 -600
rect 4985 -650 5055 -630
rect 4985 -680 5005 -650
rect 5035 -680 5055 -650
rect 4985 -690 5055 -680
rect 5070 -500 5140 -490
rect 5070 -530 5090 -500
rect 5120 -530 5140 -500
rect 5070 -550 5140 -530
rect 5070 -580 5090 -550
rect 5120 -580 5140 -550
rect 5070 -600 5140 -580
rect 5070 -630 5090 -600
rect 5120 -630 5140 -600
rect 5070 -650 5140 -630
rect 5070 -680 5090 -650
rect 5120 -680 5140 -650
rect 5070 -690 5140 -680
rect 5155 -500 5225 -490
rect 5155 -530 5175 -500
rect 5205 -530 5225 -500
rect 5155 -550 5225 -530
rect 5155 -580 5175 -550
rect 5205 -580 5225 -550
rect 5155 -600 5225 -580
rect 5155 -630 5175 -600
rect 5205 -630 5225 -600
rect 5155 -650 5225 -630
rect 5155 -680 5175 -650
rect 5205 -680 5225 -650
rect 5155 -690 5225 -680
rect 5240 -500 5310 -490
rect 5240 -530 5260 -500
rect 5290 -530 5310 -500
rect 5240 -550 5310 -530
rect 5240 -580 5260 -550
rect 5290 -580 5310 -550
rect 5240 -600 5310 -580
rect 5240 -630 5260 -600
rect 5290 -630 5310 -600
rect 5240 -650 5310 -630
rect 5240 -680 5260 -650
rect 5290 -680 5310 -650
rect 5240 -690 5310 -680
rect 5325 -500 5395 -490
rect 5325 -530 5345 -500
rect 5375 -530 5395 -500
rect 5325 -550 5395 -530
rect 5325 -580 5345 -550
rect 5375 -580 5395 -550
rect 5325 -600 5395 -580
rect 5325 -630 5345 -600
rect 5375 -630 5395 -600
rect 5325 -650 5395 -630
rect 5325 -680 5345 -650
rect 5375 -680 5395 -650
rect 5325 -690 5395 -680
rect 5410 -500 5480 -490
rect 5410 -530 5430 -500
rect 5460 -530 5480 -500
rect 5410 -550 5480 -530
rect 5410 -580 5430 -550
rect 5460 -580 5480 -550
rect 5410 -600 5480 -580
rect 5410 -630 5430 -600
rect 5460 -630 5480 -600
rect 5410 -650 5480 -630
rect 5410 -680 5430 -650
rect 5460 -680 5480 -650
rect 5410 -690 5480 -680
rect 5495 -500 5565 -490
rect 5495 -530 5515 -500
rect 5545 -530 5565 -500
rect 5495 -550 5565 -530
rect 5495 -580 5515 -550
rect 5545 -580 5565 -550
rect 5495 -600 5565 -580
rect 5495 -630 5515 -600
rect 5545 -630 5565 -600
rect 5495 -650 5565 -630
rect 5495 -680 5515 -650
rect 5545 -680 5565 -650
rect 5495 -690 5565 -680
rect 5580 -500 5650 -490
rect 5580 -530 5600 -500
rect 5630 -530 5650 -500
rect 5580 -550 5650 -530
rect 5580 -580 5600 -550
rect 5630 -580 5650 -550
rect 5580 -600 5650 -580
rect 5580 -630 5600 -600
rect 5630 -630 5650 -600
rect 5580 -650 5650 -630
rect 5580 -680 5600 -650
rect 5630 -680 5650 -650
rect 5580 -690 5650 -680
rect 5665 -500 5735 -490
rect 5665 -530 5685 -500
rect 5715 -530 5735 -500
rect 5665 -550 5735 -530
rect 5665 -580 5685 -550
rect 5715 -580 5735 -550
rect 5665 -600 5735 -580
rect 5665 -630 5685 -600
rect 5715 -630 5735 -600
rect 5665 -650 5735 -630
rect 5665 -680 5685 -650
rect 5715 -680 5735 -650
rect 5665 -690 5735 -680
rect 5750 -500 5820 -490
rect 5750 -530 5770 -500
rect 5800 -530 5820 -500
rect 5750 -550 5820 -530
rect 5750 -580 5770 -550
rect 5800 -580 5820 -550
rect 5750 -600 5820 -580
rect 5750 -630 5770 -600
rect 5800 -630 5820 -600
rect 5750 -650 5820 -630
rect 5750 -680 5770 -650
rect 5800 -680 5820 -650
rect 5750 -690 5820 -680
rect 5835 -500 5905 -490
rect 5835 -530 5855 -500
rect 5885 -530 5905 -500
rect 5835 -550 5905 -530
rect 5835 -580 5855 -550
rect 5885 -580 5905 -550
rect 5835 -600 5905 -580
rect 5835 -630 5855 -600
rect 5885 -630 5905 -600
rect 5835 -650 5905 -630
rect 5835 -680 5855 -650
rect 5885 -680 5905 -650
rect 5835 -690 5905 -680
rect 5920 -500 5990 -490
rect 5920 -530 5940 -500
rect 5970 -530 5990 -500
rect 5920 -550 5990 -530
rect 5920 -580 5940 -550
rect 5970 -580 5990 -550
rect 5920 -600 5990 -580
rect 5920 -630 5940 -600
rect 5970 -630 5990 -600
rect 5920 -650 5990 -630
rect 5920 -680 5940 -650
rect 5970 -680 5990 -650
rect 5920 -690 5990 -680
rect 6005 -500 6075 -490
rect 6005 -530 6025 -500
rect 6055 -530 6075 -500
rect 6005 -550 6075 -530
rect 6005 -580 6025 -550
rect 6055 -580 6075 -550
rect 6005 -600 6075 -580
rect 6005 -630 6025 -600
rect 6055 -630 6075 -600
rect 6005 -650 6075 -630
rect 6005 -680 6025 -650
rect 6055 -680 6075 -650
rect 6005 -690 6075 -680
rect 6090 -500 6160 -490
rect 6090 -530 6110 -500
rect 6140 -530 6160 -500
rect 6090 -550 6160 -530
rect 6090 -580 6110 -550
rect 6140 -580 6160 -550
rect 6090 -600 6160 -580
rect 6090 -630 6110 -600
rect 6140 -630 6160 -600
rect 6090 -650 6160 -630
rect 6090 -680 6110 -650
rect 6140 -680 6160 -650
rect 6090 -690 6160 -680
rect 6175 -500 6245 -490
rect 6175 -530 6195 -500
rect 6225 -530 6245 -500
rect 6175 -550 6245 -530
rect 6175 -580 6195 -550
rect 6225 -580 6245 -550
rect 6175 -600 6245 -580
rect 6175 -630 6195 -600
rect 6225 -630 6245 -600
rect 6175 -650 6245 -630
rect 6175 -680 6195 -650
rect 6225 -680 6245 -650
rect 6175 -690 6245 -680
rect 6260 -500 6330 -490
rect 6260 -530 6280 -500
rect 6310 -530 6330 -500
rect 6260 -550 6330 -530
rect 6260 -580 6280 -550
rect 6310 -580 6330 -550
rect 6260 -600 6330 -580
rect 6260 -630 6280 -600
rect 6310 -630 6330 -600
rect 6260 -650 6330 -630
rect 6260 -680 6280 -650
rect 6310 -680 6330 -650
rect 6260 -690 6330 -680
rect 6345 -500 6415 -490
rect 6345 -530 6365 -500
rect 6395 -530 6415 -500
rect 6345 -550 6415 -530
rect 6345 -580 6365 -550
rect 6395 -580 6415 -550
rect 6345 -600 6415 -580
rect 6345 -630 6365 -600
rect 6395 -630 6415 -600
rect 6345 -650 6415 -630
rect 6345 -680 6365 -650
rect 6395 -680 6415 -650
rect 6345 -690 6415 -680
rect 6430 -500 6500 -490
rect 6430 -530 6450 -500
rect 6480 -530 6500 -500
rect 6430 -550 6500 -530
rect 6430 -580 6450 -550
rect 6480 -580 6500 -550
rect 6430 -600 6500 -580
rect 6430 -630 6450 -600
rect 6480 -630 6500 -600
rect 6430 -650 6500 -630
rect 6430 -680 6450 -650
rect 6480 -680 6500 -650
rect 6430 -690 6500 -680
rect 6515 -500 6585 -490
rect 6515 -530 6535 -500
rect 6565 -530 6585 -500
rect 6515 -550 6585 -530
rect 6515 -580 6535 -550
rect 6565 -580 6585 -550
rect 6515 -600 6585 -580
rect 6515 -630 6535 -600
rect 6565 -630 6585 -600
rect 6515 -650 6585 -630
rect 6515 -680 6535 -650
rect 6565 -680 6585 -650
rect 6515 -690 6585 -680
rect 6600 -500 6670 -490
rect 6600 -530 6620 -500
rect 6650 -530 6670 -500
rect 6600 -550 6670 -530
rect 6600 -580 6620 -550
rect 6650 -580 6670 -550
rect 6600 -600 6670 -580
rect 6600 -630 6620 -600
rect 6650 -630 6670 -600
rect 6600 -650 6670 -630
rect 6600 -680 6620 -650
rect 6650 -680 6670 -650
rect 6600 -690 6670 -680
rect 6685 -500 6755 -490
rect 6685 -530 6705 -500
rect 6735 -530 6755 -500
rect 6685 -550 6755 -530
rect 6685 -580 6705 -550
rect 6735 -580 6755 -550
rect 6685 -600 6755 -580
rect 6685 -630 6705 -600
rect 6735 -630 6755 -600
rect 6685 -650 6755 -630
rect 6685 -680 6705 -650
rect 6735 -680 6755 -650
rect 6685 -690 6755 -680
rect 6770 -500 6840 -490
rect 6770 -530 6790 -500
rect 6820 -530 6840 -500
rect 6770 -550 6840 -530
rect 6770 -580 6790 -550
rect 6820 -580 6840 -550
rect 6770 -600 6840 -580
rect 6770 -630 6790 -600
rect 6820 -630 6840 -600
rect 6770 -650 6840 -630
rect 6770 -680 6790 -650
rect 6820 -680 6840 -650
rect 6770 -690 6840 -680
rect 6855 -500 6925 -490
rect 6855 -530 6875 -500
rect 6905 -530 6925 -500
rect 6855 -550 6925 -530
rect 6855 -580 6875 -550
rect 6905 -580 6925 -550
rect 6855 -600 6925 -580
rect 6855 -630 6875 -600
rect 6905 -630 6925 -600
rect 6855 -650 6925 -630
rect 6855 -680 6875 -650
rect 6905 -680 6925 -650
rect 6855 -690 6925 -680
rect 6940 -500 7010 -490
rect 6940 -530 6960 -500
rect 6990 -530 7010 -500
rect 6940 -550 7010 -530
rect 6940 -580 6960 -550
rect 6990 -580 7010 -550
rect 6940 -600 7010 -580
rect 6940 -630 6960 -600
rect 6990 -630 7010 -600
rect 6940 -650 7010 -630
rect 6940 -680 6960 -650
rect 6990 -680 7010 -650
rect 6940 -690 7010 -680
rect 7025 -500 7095 -490
rect 7025 -530 7045 -500
rect 7075 -530 7095 -500
rect 7025 -550 7095 -530
rect 7025 -580 7045 -550
rect 7075 -580 7095 -550
rect 7025 -600 7095 -580
rect 7025 -630 7045 -600
rect 7075 -630 7095 -600
rect 7025 -650 7095 -630
rect 7025 -680 7045 -650
rect 7075 -680 7095 -650
rect 7025 -690 7095 -680
rect 7110 -500 7180 -490
rect 7110 -530 7130 -500
rect 7160 -530 7180 -500
rect 7110 -550 7180 -530
rect 7110 -580 7130 -550
rect 7160 -580 7180 -550
rect 7110 -600 7180 -580
rect 7110 -630 7130 -600
rect 7160 -630 7180 -600
rect 7110 -650 7180 -630
rect 7110 -680 7130 -650
rect 7160 -680 7180 -650
rect 7110 -690 7180 -680
rect 7195 -500 7265 -490
rect 7195 -530 7215 -500
rect 7245 -530 7265 -500
rect 7195 -550 7265 -530
rect 7195 -580 7215 -550
rect 7245 -580 7265 -550
rect 7195 -600 7265 -580
rect 7195 -630 7215 -600
rect 7245 -630 7265 -600
rect 7195 -650 7265 -630
rect 7195 -680 7215 -650
rect 7245 -680 7265 -650
rect 7195 -690 7265 -680
rect 7280 -500 7350 -490
rect 7280 -530 7300 -500
rect 7330 -530 7350 -500
rect 7280 -550 7350 -530
rect 7280 -580 7300 -550
rect 7330 -580 7350 -550
rect 7280 -600 7350 -580
rect 7280 -630 7300 -600
rect 7330 -630 7350 -600
rect 7280 -650 7350 -630
rect 7280 -680 7300 -650
rect 7330 -680 7350 -650
rect 7280 -690 7350 -680
rect 7365 -500 7435 -490
rect 7365 -530 7385 -500
rect 7415 -530 7435 -500
rect 7365 -550 7435 -530
rect 7365 -580 7385 -550
rect 7415 -580 7435 -550
rect 7365 -600 7435 -580
rect 7365 -630 7385 -600
rect 7415 -630 7435 -600
rect 7365 -650 7435 -630
rect 7365 -680 7385 -650
rect 7415 -680 7435 -650
rect 7365 -690 7435 -680
rect 7450 -500 7520 -490
rect 7450 -530 7470 -500
rect 7500 -530 7520 -500
rect 7450 -550 7520 -530
rect 7450 -580 7470 -550
rect 7500 -580 7520 -550
rect 7450 -600 7520 -580
rect 7450 -630 7470 -600
rect 7500 -630 7520 -600
rect 7450 -650 7520 -630
rect 7450 -680 7470 -650
rect 7500 -680 7520 -650
rect 7450 -690 7520 -680
rect 7535 -500 7605 -490
rect 7535 -530 7555 -500
rect 7585 -530 7605 -500
rect 7535 -550 7605 -530
rect 7535 -580 7555 -550
rect 7585 -580 7605 -550
rect 7535 -600 7605 -580
rect 7535 -630 7555 -600
rect 7585 -630 7605 -600
rect 7535 -650 7605 -630
rect 7535 -680 7555 -650
rect 7585 -680 7605 -650
rect 7535 -690 7605 -680
rect 7620 -500 7690 -490
rect 7620 -530 7640 -500
rect 7670 -530 7690 -500
rect 7620 -550 7690 -530
rect 7620 -580 7640 -550
rect 7670 -580 7690 -550
rect 7620 -600 7690 -580
rect 7620 -630 7640 -600
rect 7670 -630 7690 -600
rect 7620 -650 7690 -630
rect 7620 -680 7640 -650
rect 7670 -680 7690 -650
rect 7620 -690 7690 -680
rect 7705 -500 7775 -490
rect 7705 -530 7725 -500
rect 7755 -530 7775 -500
rect 7705 -550 7775 -530
rect 7705 -580 7725 -550
rect 7755 -580 7775 -550
rect 7705 -600 7775 -580
rect 7705 -630 7725 -600
rect 7755 -630 7775 -600
rect 7705 -650 7775 -630
rect 7705 -680 7725 -650
rect 7755 -680 7775 -650
rect 7705 -690 7775 -680
rect 7790 -500 7860 -490
rect 7790 -530 7810 -500
rect 7840 -530 7860 -500
rect 7790 -550 7860 -530
rect 7790 -580 7810 -550
rect 7840 -580 7860 -550
rect 7790 -600 7860 -580
rect 7790 -630 7810 -600
rect 7840 -630 7860 -600
rect 7790 -650 7860 -630
rect 7790 -680 7810 -650
rect 7840 -680 7860 -650
rect 7790 -690 7860 -680
rect 7875 -500 7945 -490
rect 7875 -530 7895 -500
rect 7925 -530 7945 -500
rect 7875 -550 7945 -530
rect 7875 -580 7895 -550
rect 7925 -580 7945 -550
rect 7875 -600 7945 -580
rect 7875 -630 7895 -600
rect 7925 -630 7945 -600
rect 7875 -650 7945 -630
rect 7875 -680 7895 -650
rect 7925 -680 7945 -650
rect 7875 -690 7945 -680
rect 7960 -500 8030 -490
rect 7960 -530 7980 -500
rect 8010 -530 8030 -500
rect 7960 -550 8030 -530
rect 7960 -580 7980 -550
rect 8010 -580 8030 -550
rect 7960 -600 8030 -580
rect 7960 -630 7980 -600
rect 8010 -630 8030 -600
rect 7960 -650 8030 -630
rect 7960 -680 7980 -650
rect 8010 -680 8030 -650
rect 7960 -690 8030 -680
rect 8045 -500 8115 -490
rect 8045 -530 8065 -500
rect 8095 -530 8115 -500
rect 8045 -550 8115 -530
rect 8045 -580 8065 -550
rect 8095 -580 8115 -550
rect 8045 -600 8115 -580
rect 8045 -630 8065 -600
rect 8095 -630 8115 -600
rect 8045 -650 8115 -630
rect 8045 -680 8065 -650
rect 8095 -680 8115 -650
rect 8045 -690 8115 -680
rect 8130 -500 8200 -490
rect 8130 -530 8150 -500
rect 8180 -530 8200 -500
rect 8130 -550 8200 -530
rect 8130 -580 8150 -550
rect 8180 -580 8200 -550
rect 8130 -600 8200 -580
rect 8130 -630 8150 -600
rect 8180 -630 8200 -600
rect 8130 -650 8200 -630
rect 8130 -680 8150 -650
rect 8180 -680 8200 -650
rect 8130 -690 8200 -680
rect 8215 -500 8285 -490
rect 8215 -530 8235 -500
rect 8265 -530 8285 -500
rect 8215 -550 8285 -530
rect 8215 -580 8235 -550
rect 8265 -580 8285 -550
rect 8215 -600 8285 -580
rect 8215 -630 8235 -600
rect 8265 -630 8285 -600
rect 8215 -650 8285 -630
rect 8215 -680 8235 -650
rect 8265 -680 8285 -650
rect 8215 -690 8285 -680
rect 8300 -500 8370 -490
rect 8300 -530 8320 -500
rect 8350 -530 8370 -500
rect 8300 -550 8370 -530
rect 8300 -580 8320 -550
rect 8350 -580 8370 -550
rect 8300 -600 8370 -580
rect 8300 -630 8320 -600
rect 8350 -630 8370 -600
rect 8300 -650 8370 -630
rect 8300 -680 8320 -650
rect 8350 -680 8370 -650
rect 8300 -690 8370 -680
rect 8385 -500 8455 -490
rect 8385 -530 8405 -500
rect 8435 -530 8455 -500
rect 8385 -550 8455 -530
rect 8385 -580 8405 -550
rect 8435 -580 8455 -550
rect 8385 -600 8455 -580
rect 8385 -630 8405 -600
rect 8435 -630 8455 -600
rect 8385 -650 8455 -630
rect 8385 -680 8405 -650
rect 8435 -680 8455 -650
rect 8385 -690 8455 -680
rect 8470 -500 8540 -490
rect 8470 -530 8490 -500
rect 8520 -530 8540 -500
rect 8470 -550 8540 -530
rect 8470 -580 8490 -550
rect 8520 -580 8540 -550
rect 8470 -600 8540 -580
rect 8470 -630 8490 -600
rect 8520 -630 8540 -600
rect 8470 -650 8540 -630
rect 8470 -680 8490 -650
rect 8520 -680 8540 -650
rect 8470 -690 8540 -680
rect 8555 -500 8625 -490
rect 8555 -530 8575 -500
rect 8605 -530 8625 -500
rect 8555 -550 8625 -530
rect 8555 -580 8575 -550
rect 8605 -580 8625 -550
rect 8555 -600 8625 -580
rect 8555 -630 8575 -600
rect 8605 -630 8625 -600
rect 8555 -650 8625 -630
rect 8555 -680 8575 -650
rect 8605 -680 8625 -650
rect 8555 -690 8625 -680
rect 8640 -500 8710 -490
rect 8640 -530 8660 -500
rect 8690 -530 8710 -500
rect 8640 -550 8710 -530
rect 8640 -580 8660 -550
rect 8690 -580 8710 -550
rect 8640 -600 8710 -580
rect 8640 -630 8660 -600
rect 8690 -630 8710 -600
rect 8640 -650 8710 -630
rect 8640 -680 8660 -650
rect 8690 -680 8710 -650
rect 8640 -690 8710 -680
rect 8725 -500 8795 -490
rect 8725 -530 8745 -500
rect 8775 -530 8795 -500
rect 8725 -550 8795 -530
rect 8725 -580 8745 -550
rect 8775 -580 8795 -550
rect 8725 -600 8795 -580
rect 8725 -630 8745 -600
rect 8775 -630 8795 -600
rect 8725 -650 8795 -630
rect 8725 -680 8745 -650
rect 8775 -680 8795 -650
rect 8725 -690 8795 -680
rect 8810 -500 8880 -490
rect 8810 -530 8830 -500
rect 8860 -530 8880 -500
rect 8810 -550 8880 -530
rect 8810 -580 8830 -550
rect 8860 -580 8880 -550
rect 8810 -600 8880 -580
rect 8810 -630 8830 -600
rect 8860 -630 8880 -600
rect 8810 -650 8880 -630
rect 8810 -680 8830 -650
rect 8860 -680 8880 -650
rect 8810 -690 8880 -680
rect 8895 -500 8965 -490
rect 8895 -530 8915 -500
rect 8945 -530 8965 -500
rect 8895 -550 8965 -530
rect 8895 -580 8915 -550
rect 8945 -580 8965 -550
rect 8895 -600 8965 -580
rect 8895 -630 8915 -600
rect 8945 -630 8965 -600
rect 8895 -650 8965 -630
rect 8895 -680 8915 -650
rect 8945 -680 8965 -650
rect 8895 -690 8965 -680
rect 8980 -500 9050 -490
rect 8980 -530 9000 -500
rect 9030 -530 9050 -500
rect 8980 -550 9050 -530
rect 8980 -580 9000 -550
rect 9030 -580 9050 -550
rect 8980 -600 9050 -580
rect 8980 -630 9000 -600
rect 9030 -630 9050 -600
rect 8980 -650 9050 -630
rect 8980 -680 9000 -650
rect 9030 -680 9050 -650
rect 8980 -690 9050 -680
rect 9065 -500 9135 -490
rect 9065 -530 9085 -500
rect 9115 -530 9135 -500
rect 9065 -550 9135 -530
rect 9065 -580 9085 -550
rect 9115 -580 9135 -550
rect 9065 -600 9135 -580
rect 9065 -630 9085 -600
rect 9115 -630 9135 -600
rect 9065 -650 9135 -630
rect 9065 -680 9085 -650
rect 9115 -680 9135 -650
rect 9065 -690 9135 -680
rect 9150 -500 9220 -490
rect 9150 -530 9170 -500
rect 9200 -530 9220 -500
rect 9150 -550 9220 -530
rect 9150 -580 9170 -550
rect 9200 -580 9220 -550
rect 9150 -600 9220 -580
rect 9150 -630 9170 -600
rect 9200 -630 9220 -600
rect 9150 -650 9220 -630
rect 9150 -680 9170 -650
rect 9200 -680 9220 -650
rect 9150 -690 9220 -680
rect 9235 -500 9305 -490
rect 9235 -530 9255 -500
rect 9285 -530 9305 -500
rect 9235 -550 9305 -530
rect 9235 -580 9255 -550
rect 9285 -580 9305 -550
rect 9235 -600 9305 -580
rect 9235 -630 9255 -600
rect 9285 -630 9305 -600
rect 9235 -650 9305 -630
rect 9235 -680 9255 -650
rect 9285 -680 9305 -650
rect 9235 -690 9305 -680
rect 9320 -500 9390 -490
rect 9320 -530 9340 -500
rect 9370 -530 9390 -500
rect 9320 -550 9390 -530
rect 9320 -580 9340 -550
rect 9370 -580 9390 -550
rect 9320 -600 9390 -580
rect 9320 -630 9340 -600
rect 9370 -630 9390 -600
rect 9320 -650 9390 -630
rect 9320 -680 9340 -650
rect 9370 -680 9390 -650
rect 9320 -690 9390 -680
rect 9405 -500 9475 -490
rect 9405 -530 9425 -500
rect 9455 -530 9475 -500
rect 9405 -550 9475 -530
rect 9405 -580 9425 -550
rect 9455 -580 9475 -550
rect 9405 -600 9475 -580
rect 9405 -630 9425 -600
rect 9455 -630 9475 -600
rect 9405 -650 9475 -630
rect 9405 -680 9425 -650
rect 9455 -680 9475 -650
rect 9405 -690 9475 -680
rect 9490 -500 9560 -490
rect 9490 -530 9510 -500
rect 9540 -530 9560 -500
rect 9490 -550 9560 -530
rect 9490 -580 9510 -550
rect 9540 -580 9560 -550
rect 9490 -600 9560 -580
rect 9490 -630 9510 -600
rect 9540 -630 9560 -600
rect 9490 -650 9560 -630
rect 9490 -680 9510 -650
rect 9540 -680 9560 -650
rect 9490 -690 9560 -680
rect 9575 -500 9645 -490
rect 9575 -530 9595 -500
rect 9625 -530 9645 -500
rect 9575 -550 9645 -530
rect 9575 -580 9595 -550
rect 9625 -580 9645 -550
rect 9575 -600 9645 -580
rect 9575 -630 9595 -600
rect 9625 -630 9645 -600
rect 9575 -650 9645 -630
rect 9575 -680 9595 -650
rect 9625 -680 9645 -650
rect 9575 -690 9645 -680
rect 9660 -500 9730 -490
rect 9660 -530 9680 -500
rect 9710 -530 9730 -500
rect 9660 -550 9730 -530
rect 9660 -580 9680 -550
rect 9710 -580 9730 -550
rect 9660 -600 9730 -580
rect 9660 -630 9680 -600
rect 9710 -630 9730 -600
rect 9660 -650 9730 -630
rect 9660 -680 9680 -650
rect 9710 -680 9730 -650
rect 9660 -690 9730 -680
rect 9745 -500 9815 -490
rect 9745 -530 9765 -500
rect 9795 -530 9815 -500
rect 9745 -550 9815 -530
rect 9745 -580 9765 -550
rect 9795 -580 9815 -550
rect 9745 -600 9815 -580
rect 9745 -630 9765 -600
rect 9795 -630 9815 -600
rect 9745 -650 9815 -630
rect 9745 -680 9765 -650
rect 9795 -680 9815 -650
rect 9745 -690 9815 -680
rect 9830 -500 9900 -490
rect 9830 -530 9850 -500
rect 9880 -530 9900 -500
rect 9830 -550 9900 -530
rect 9830 -580 9850 -550
rect 9880 -580 9900 -550
rect 9830 -600 9900 -580
rect 9830 -630 9850 -600
rect 9880 -630 9900 -600
rect 9830 -650 9900 -630
rect 9830 -680 9850 -650
rect 9880 -680 9900 -650
rect 9830 -690 9900 -680
rect 9915 -500 9985 -490
rect 9915 -530 9935 -500
rect 9965 -530 9985 -500
rect 9915 -550 9985 -530
rect 9915 -580 9935 -550
rect 9965 -580 9985 -550
rect 9915 -600 9985 -580
rect 9915 -630 9935 -600
rect 9965 -630 9985 -600
rect 9915 -650 9985 -630
rect 9915 -680 9935 -650
rect 9965 -680 9985 -650
rect 9915 -690 9985 -680
rect 10000 -500 10070 -490
rect 10000 -530 10020 -500
rect 10050 -530 10070 -500
rect 10000 -550 10070 -530
rect 10000 -580 10020 -550
rect 10050 -580 10070 -550
rect 10000 -600 10070 -580
rect 10000 -630 10020 -600
rect 10050 -630 10070 -600
rect 10000 -650 10070 -630
rect 10000 -680 10020 -650
rect 10050 -680 10070 -650
rect 10000 -690 10070 -680
rect 10085 -500 10155 -490
rect 10085 -530 10105 -500
rect 10135 -530 10155 -500
rect 10085 -550 10155 -530
rect 10085 -580 10105 -550
rect 10135 -580 10155 -550
rect 10085 -600 10155 -580
rect 10085 -630 10105 -600
rect 10135 -630 10155 -600
rect 10085 -650 10155 -630
rect 10085 -680 10105 -650
rect 10135 -680 10155 -650
rect 10085 -690 10155 -680
rect 10170 -500 10240 -490
rect 10170 -530 10190 -500
rect 10220 -530 10240 -500
rect 10170 -550 10240 -530
rect 10170 -580 10190 -550
rect 10220 -580 10240 -550
rect 10170 -600 10240 -580
rect 10170 -630 10190 -600
rect 10220 -630 10240 -600
rect 10170 -650 10240 -630
rect 10170 -680 10190 -650
rect 10220 -680 10240 -650
rect 10170 -690 10240 -680
rect 10255 -500 10325 -490
rect 10255 -530 10275 -500
rect 10305 -530 10325 -500
rect 10255 -550 10325 -530
rect 10255 -580 10275 -550
rect 10305 -580 10325 -550
rect 10255 -600 10325 -580
rect 10255 -630 10275 -600
rect 10305 -630 10325 -600
rect 10255 -650 10325 -630
rect 10255 -680 10275 -650
rect 10305 -680 10325 -650
rect 10255 -690 10325 -680
rect 10340 -500 10410 -490
rect 10340 -530 10360 -500
rect 10390 -530 10410 -500
rect 10340 -550 10410 -530
rect 10340 -580 10360 -550
rect 10390 -580 10410 -550
rect 10340 -600 10410 -580
rect 10340 -630 10360 -600
rect 10390 -630 10410 -600
rect 10340 -650 10410 -630
rect 10340 -680 10360 -650
rect 10390 -680 10410 -650
rect 10340 -690 10410 -680
rect 10425 -500 10495 -490
rect 10425 -530 10445 -500
rect 10475 -530 10495 -500
rect 10425 -550 10495 -530
rect 10425 -580 10445 -550
rect 10475 -580 10495 -550
rect 10425 -600 10495 -580
rect 10425 -630 10445 -600
rect 10475 -630 10495 -600
rect 10425 -650 10495 -630
rect 10425 -680 10445 -650
rect 10475 -680 10495 -650
rect 10425 -690 10495 -680
rect 10510 -500 10580 -490
rect 10510 -530 10530 -500
rect 10560 -530 10580 -500
rect 10510 -550 10580 -530
rect 10510 -580 10530 -550
rect 10560 -580 10580 -550
rect 10510 -600 10580 -580
rect 10510 -630 10530 -600
rect 10560 -630 10580 -600
rect 10510 -650 10580 -630
rect 10510 -680 10530 -650
rect 10560 -680 10580 -650
rect 10510 -690 10580 -680
rect 10595 -500 10665 -490
rect 10595 -530 10615 -500
rect 10645 -530 10665 -500
rect 10595 -550 10665 -530
rect 10595 -580 10615 -550
rect 10645 -580 10665 -550
rect 10595 -600 10665 -580
rect 10595 -630 10615 -600
rect 10645 -630 10665 -600
rect 10595 -650 10665 -630
rect 10595 -680 10615 -650
rect 10645 -680 10665 -650
rect 10595 -690 10665 -680
rect 10680 -500 10750 -490
rect 10680 -530 10700 -500
rect 10730 -530 10750 -500
rect 10680 -550 10750 -530
rect 10680 -580 10700 -550
rect 10730 -580 10750 -550
rect 10680 -600 10750 -580
rect 10680 -630 10700 -600
rect 10730 -630 10750 -600
rect 10680 -650 10750 -630
rect 10680 -680 10700 -650
rect 10730 -680 10750 -650
rect 10680 -690 10750 -680
rect 10765 -500 10835 -490
rect 10765 -530 10785 -500
rect 10815 -530 10835 -500
rect 10765 -550 10835 -530
rect 10765 -580 10785 -550
rect 10815 -580 10835 -550
rect 10765 -600 10835 -580
rect 10765 -630 10785 -600
rect 10815 -630 10835 -600
rect 10765 -650 10835 -630
rect 10765 -680 10785 -650
rect 10815 -680 10835 -650
rect 10765 -690 10835 -680
rect 10850 -500 10920 -490
rect 10850 -530 10870 -500
rect 10900 -530 10920 -500
rect 10850 -550 10920 -530
rect 10850 -580 10870 -550
rect 10900 -580 10920 -550
rect 10850 -600 10920 -580
rect 10850 -630 10870 -600
rect 10900 -630 10920 -600
rect 10850 -650 10920 -630
rect 10850 -680 10870 -650
rect 10900 -680 10920 -650
rect 10850 -690 10920 -680
rect 10935 -500 11005 -490
rect 10935 -530 10955 -500
rect 10985 -530 11005 -500
rect 10935 -550 11005 -530
rect 10935 -580 10955 -550
rect 10985 -580 11005 -550
rect 10935 -600 11005 -580
rect 10935 -630 10955 -600
rect 10985 -630 11005 -600
rect 10935 -650 11005 -630
rect 10935 -680 10955 -650
rect 10985 -680 11005 -650
rect 10935 -690 11005 -680
rect 11020 -500 11090 -490
rect 11020 -530 11040 -500
rect 11070 -530 11090 -500
rect 11020 -550 11090 -530
rect 11020 -580 11040 -550
rect 11070 -580 11090 -550
rect 11020 -600 11090 -580
rect 11020 -630 11040 -600
rect 11070 -630 11090 -600
rect 11020 -650 11090 -630
rect 11020 -680 11040 -650
rect 11070 -680 11090 -650
rect 11020 -690 11090 -680
rect 11105 -500 11175 -490
rect 11105 -530 11125 -500
rect 11155 -530 11175 -500
rect 11105 -550 11175 -530
rect 11105 -580 11125 -550
rect 11155 -580 11175 -550
rect 11105 -600 11175 -580
rect 11105 -630 11125 -600
rect 11155 -630 11175 -600
rect 11105 -650 11175 -630
rect 11105 -680 11125 -650
rect 11155 -680 11175 -650
rect 11105 -690 11175 -680
rect 11190 -500 11260 -490
rect 11190 -530 11210 -500
rect 11240 -530 11260 -500
rect 11190 -550 11260 -530
rect 11190 -580 11210 -550
rect 11240 -580 11260 -550
rect 11190 -600 11260 -580
rect 11190 -630 11210 -600
rect 11240 -630 11260 -600
rect 11190 -650 11260 -630
rect 11190 -680 11210 -650
rect 11240 -680 11260 -650
rect 11190 -690 11260 -680
rect 11275 -500 11345 -490
rect 11275 -530 11295 -500
rect 11325 -530 11345 -500
rect 11275 -550 11345 -530
rect 11275 -580 11295 -550
rect 11325 -580 11345 -550
rect 11275 -600 11345 -580
rect 11275 -630 11295 -600
rect 11325 -630 11345 -600
rect 11275 -650 11345 -630
rect 11275 -680 11295 -650
rect 11325 -680 11345 -650
rect 11275 -690 11345 -680
rect 11360 -500 11430 -490
rect 11360 -530 11380 -500
rect 11410 -530 11430 -500
rect 11360 -550 11430 -530
rect 11360 -580 11380 -550
rect 11410 -580 11430 -550
rect 11360 -600 11430 -580
rect 11360 -630 11380 -600
rect 11410 -630 11430 -600
rect 11360 -650 11430 -630
rect 11360 -680 11380 -650
rect 11410 -680 11430 -650
rect 11360 -690 11430 -680
rect 11445 -500 11515 -490
rect 11445 -530 11465 -500
rect 11495 -530 11515 -500
rect 11445 -550 11515 -530
rect 11445 -580 11465 -550
rect 11495 -580 11515 -550
rect 11445 -600 11515 -580
rect 11445 -630 11465 -600
rect 11495 -630 11515 -600
rect 11445 -650 11515 -630
rect 11445 -680 11465 -650
rect 11495 -680 11515 -650
rect 11445 -690 11515 -680
rect 11530 -500 11600 -490
rect 11530 -530 11550 -500
rect 11580 -530 11600 -500
rect 11530 -550 11600 -530
rect 11530 -580 11550 -550
rect 11580 -580 11600 -550
rect 11530 -600 11600 -580
rect 11530 -630 11550 -600
rect 11580 -630 11600 -600
rect 11530 -650 11600 -630
rect 11530 -680 11550 -650
rect 11580 -680 11600 -650
rect 11530 -690 11600 -680
rect 11615 -500 11685 -490
rect 11615 -530 11635 -500
rect 11665 -530 11685 -500
rect 11615 -550 11685 -530
rect 11615 -580 11635 -550
rect 11665 -580 11685 -550
rect 11615 -600 11685 -580
rect 11615 -630 11635 -600
rect 11665 -630 11685 -600
rect 11615 -650 11685 -630
rect 11615 -680 11635 -650
rect 11665 -680 11685 -650
rect 11615 -690 11685 -680
rect 11700 -500 11770 -490
rect 11700 -530 11720 -500
rect 11750 -530 11770 -500
rect 11700 -550 11770 -530
rect 11700 -580 11720 -550
rect 11750 -580 11770 -550
rect 11700 -600 11770 -580
rect 11700 -630 11720 -600
rect 11750 -630 11770 -600
rect 11700 -650 11770 -630
rect 11700 -680 11720 -650
rect 11750 -680 11770 -650
rect 11700 -690 11770 -680
rect 11785 -500 11855 -490
rect 11785 -530 11805 -500
rect 11835 -530 11855 -500
rect 11785 -550 11855 -530
rect 11785 -580 11805 -550
rect 11835 -580 11855 -550
rect 11785 -600 11855 -580
rect 11785 -630 11805 -600
rect 11835 -630 11855 -600
rect 11785 -650 11855 -630
rect 11785 -680 11805 -650
rect 11835 -680 11855 -650
rect 11785 -690 11855 -680
rect 11870 -500 11940 -490
rect 11870 -530 11890 -500
rect 11920 -530 11940 -500
rect 11870 -550 11940 -530
rect 11870 -580 11890 -550
rect 11920 -580 11940 -550
rect 11870 -600 11940 -580
rect 11870 -630 11890 -600
rect 11920 -630 11940 -600
rect 11870 -650 11940 -630
rect 11870 -680 11890 -650
rect 11920 -680 11940 -650
rect 11870 -690 11940 -680
rect 11955 -500 12025 -490
rect 11955 -530 11975 -500
rect 12005 -530 12025 -500
rect 11955 -550 12025 -530
rect 11955 -580 11975 -550
rect 12005 -580 12025 -550
rect 11955 -600 12025 -580
rect 11955 -630 11975 -600
rect 12005 -630 12025 -600
rect 11955 -650 12025 -630
rect 11955 -680 11975 -650
rect 12005 -680 12025 -650
rect 11955 -690 12025 -680
rect 12040 -500 12110 -490
rect 12040 -530 12060 -500
rect 12090 -530 12110 -500
rect 12040 -550 12110 -530
rect 12040 -580 12060 -550
rect 12090 -580 12110 -550
rect 12040 -600 12110 -580
rect 12040 -630 12060 -600
rect 12090 -630 12110 -600
rect 12040 -650 12110 -630
rect 12040 -680 12060 -650
rect 12090 -680 12110 -650
rect 12040 -690 12110 -680
rect 12125 -500 12195 -490
rect 12125 -530 12145 -500
rect 12175 -530 12195 -500
rect 12125 -550 12195 -530
rect 12125 -580 12145 -550
rect 12175 -580 12195 -550
rect 12125 -600 12195 -580
rect 12125 -630 12145 -600
rect 12175 -630 12195 -600
rect 12125 -650 12195 -630
rect 12125 -680 12145 -650
rect 12175 -680 12195 -650
rect 12125 -690 12195 -680
rect 12210 -500 12280 -490
rect 12210 -530 12230 -500
rect 12260 -530 12280 -500
rect 12210 -550 12280 -530
rect 12210 -580 12230 -550
rect 12260 -580 12280 -550
rect 12210 -600 12280 -580
rect 12210 -630 12230 -600
rect 12260 -630 12280 -600
rect 12210 -650 12280 -630
rect 12210 -680 12230 -650
rect 12260 -680 12280 -650
rect 12210 -690 12280 -680
rect 12295 -500 12365 -490
rect 12295 -530 12315 -500
rect 12345 -530 12365 -500
rect 12295 -550 12365 -530
rect 12295 -580 12315 -550
rect 12345 -580 12365 -550
rect 12295 -600 12365 -580
rect 12295 -630 12315 -600
rect 12345 -630 12365 -600
rect 12295 -650 12365 -630
rect 12295 -680 12315 -650
rect 12345 -680 12365 -650
rect 12295 -690 12365 -680
rect 12380 -500 12450 -490
rect 12380 -530 12400 -500
rect 12430 -530 12450 -500
rect 12380 -550 12450 -530
rect 12380 -580 12400 -550
rect 12430 -580 12450 -550
rect 12380 -600 12450 -580
rect 12380 -630 12400 -600
rect 12430 -630 12450 -600
rect 12380 -650 12450 -630
rect 12380 -680 12400 -650
rect 12430 -680 12450 -650
rect 12380 -690 12450 -680
rect 12465 -500 12535 -490
rect 12465 -530 12485 -500
rect 12515 -530 12535 -500
rect 12465 -550 12535 -530
rect 12465 -580 12485 -550
rect 12515 -580 12535 -550
rect 12465 -600 12535 -580
rect 12465 -630 12485 -600
rect 12515 -630 12535 -600
rect 12465 -650 12535 -630
rect 12465 -680 12485 -650
rect 12515 -680 12535 -650
rect 12465 -690 12535 -680
rect 12550 -500 12620 -490
rect 12550 -530 12570 -500
rect 12600 -530 12620 -500
rect 12550 -550 12620 -530
rect 12550 -580 12570 -550
rect 12600 -580 12620 -550
rect 12550 -600 12620 -580
rect 12550 -630 12570 -600
rect 12600 -630 12620 -600
rect 12550 -650 12620 -630
rect 12550 -680 12570 -650
rect 12600 -680 12620 -650
rect 12550 -690 12620 -680
rect 12635 -500 12705 -490
rect 12635 -530 12655 -500
rect 12685 -530 12705 -500
rect 12635 -550 12705 -530
rect 12635 -580 12655 -550
rect 12685 -580 12705 -550
rect 12635 -600 12705 -580
rect 12635 -630 12655 -600
rect 12685 -630 12705 -600
rect 12635 -650 12705 -630
rect 12635 -680 12655 -650
rect 12685 -680 12705 -650
rect 12635 -690 12705 -680
rect 12720 -500 12790 -490
rect 12720 -530 12740 -500
rect 12770 -530 12790 -500
rect 12720 -550 12790 -530
rect 12720 -580 12740 -550
rect 12770 -580 12790 -550
rect 12720 -600 12790 -580
rect 12720 -630 12740 -600
rect 12770 -630 12790 -600
rect 12720 -650 12790 -630
rect 12720 -680 12740 -650
rect 12770 -680 12790 -650
rect 12720 -690 12790 -680
rect 12805 -500 12875 -490
rect 12805 -530 12825 -500
rect 12855 -530 12875 -500
rect 12805 -550 12875 -530
rect 12805 -580 12825 -550
rect 12855 -580 12875 -550
rect 12805 -600 12875 -580
rect 12805 -630 12825 -600
rect 12855 -630 12875 -600
rect 12805 -650 12875 -630
rect 12805 -680 12825 -650
rect 12855 -680 12875 -650
rect 12805 -690 12875 -680
rect 12890 -500 12960 -490
rect 12890 -530 12910 -500
rect 12940 -530 12960 -500
rect 12890 -550 12960 -530
rect 12890 -580 12910 -550
rect 12940 -580 12960 -550
rect 12890 -600 12960 -580
rect 12890 -630 12910 -600
rect 12940 -630 12960 -600
rect 12890 -650 12960 -630
rect 12890 -680 12910 -650
rect 12940 -680 12960 -650
rect 12890 -690 12960 -680
rect 12975 -500 13045 -490
rect 12975 -530 12995 -500
rect 13025 -530 13045 -500
rect 12975 -550 13045 -530
rect 12975 -580 12995 -550
rect 13025 -580 13045 -550
rect 12975 -600 13045 -580
rect 12975 -630 12995 -600
rect 13025 -630 13045 -600
rect 12975 -650 13045 -630
rect 12975 -680 12995 -650
rect 13025 -680 13045 -650
rect 12975 -690 13045 -680
rect 13060 -500 13130 -490
rect 13060 -530 13080 -500
rect 13110 -530 13130 -500
rect 13060 -550 13130 -530
rect 13060 -580 13080 -550
rect 13110 -580 13130 -550
rect 13060 -600 13130 -580
rect 13060 -630 13080 -600
rect 13110 -630 13130 -600
rect 13060 -650 13130 -630
rect 13060 -680 13080 -650
rect 13110 -680 13130 -650
rect 13060 -690 13130 -680
rect 13145 -500 13215 -490
rect 13145 -530 13165 -500
rect 13195 -530 13215 -500
rect 13145 -550 13215 -530
rect 13145 -580 13165 -550
rect 13195 -580 13215 -550
rect 13145 -600 13215 -580
rect 13145 -630 13165 -600
rect 13195 -630 13215 -600
rect 13145 -650 13215 -630
rect 13145 -680 13165 -650
rect 13195 -680 13215 -650
rect 13145 -690 13215 -680
rect 13230 -500 13300 -490
rect 13230 -530 13250 -500
rect 13280 -530 13300 -500
rect 13230 -550 13300 -530
rect 13230 -580 13250 -550
rect 13280 -580 13300 -550
rect 13230 -600 13300 -580
rect 13230 -630 13250 -600
rect 13280 -630 13300 -600
rect 13230 -650 13300 -630
rect 13230 -680 13250 -650
rect 13280 -680 13300 -650
rect 13230 -690 13300 -680
rect 13315 -500 13385 -490
rect 13315 -530 13335 -500
rect 13365 -530 13385 -500
rect 13315 -550 13385 -530
rect 13315 -580 13335 -550
rect 13365 -580 13385 -550
rect 13315 -600 13385 -580
rect 13315 -630 13335 -600
rect 13365 -630 13385 -600
rect 13315 -650 13385 -630
rect 13315 -680 13335 -650
rect 13365 -680 13385 -650
rect 13315 -690 13385 -680
rect 13400 -500 13470 -490
rect 13400 -530 13420 -500
rect 13450 -530 13470 -500
rect 13400 -550 13470 -530
rect 13400 -580 13420 -550
rect 13450 -580 13470 -550
rect 13400 -600 13470 -580
rect 13400 -630 13420 -600
rect 13450 -630 13470 -600
rect 13400 -650 13470 -630
rect 13400 -680 13420 -650
rect 13450 -680 13470 -650
rect 13400 -690 13470 -680
rect 13485 -500 13555 -490
rect 13485 -530 13505 -500
rect 13535 -530 13555 -500
rect 13485 -550 13555 -530
rect 13485 -580 13505 -550
rect 13535 -580 13555 -550
rect 13485 -600 13555 -580
rect 13485 -630 13505 -600
rect 13535 -630 13555 -600
rect 13485 -650 13555 -630
rect 13485 -680 13505 -650
rect 13535 -680 13555 -650
rect 13485 -690 13555 -680
rect 13570 -500 13640 -490
rect 13570 -530 13590 -500
rect 13620 -530 13640 -500
rect 13570 -550 13640 -530
rect 13570 -580 13590 -550
rect 13620 -580 13640 -550
rect 13570 -600 13640 -580
rect 13570 -630 13590 -600
rect 13620 -630 13640 -600
rect 13570 -650 13640 -630
rect 13570 -680 13590 -650
rect 13620 -680 13640 -650
rect 13570 -690 13640 -680
rect 13655 -500 13725 -490
rect 13655 -530 13675 -500
rect 13705 -530 13725 -500
rect 13655 -550 13725 -530
rect 13655 -580 13675 -550
rect 13705 -580 13725 -550
rect 13655 -600 13725 -580
rect 13655 -630 13675 -600
rect 13705 -630 13725 -600
rect 13655 -650 13725 -630
rect 13655 -680 13675 -650
rect 13705 -680 13725 -650
rect 13655 -690 13725 -680
rect 13740 -500 13810 -490
rect 13740 -530 13760 -500
rect 13790 -530 13810 -500
rect 13740 -550 13810 -530
rect 13740 -580 13760 -550
rect 13790 -580 13810 -550
rect 13740 -600 13810 -580
rect 13740 -630 13760 -600
rect 13790 -630 13810 -600
rect 13740 -650 13810 -630
rect 13740 -680 13760 -650
rect 13790 -680 13810 -650
rect 13740 -690 13810 -680
rect 13825 -500 13895 -490
rect 13825 -530 13845 -500
rect 13875 -530 13895 -500
rect 13825 -550 13895 -530
rect 13825 -580 13845 -550
rect 13875 -580 13895 -550
rect 13825 -600 13895 -580
rect 13825 -630 13845 -600
rect 13875 -630 13895 -600
rect 13825 -650 13895 -630
rect 13825 -680 13845 -650
rect 13875 -680 13895 -650
rect 13825 -690 13895 -680
rect 13910 -500 13980 -490
rect 13910 -530 13930 -500
rect 13960 -530 13980 -500
rect 13910 -550 13980 -530
rect 13910 -580 13930 -550
rect 13960 -580 13980 -550
rect 13910 -600 13980 -580
rect 13910 -630 13930 -600
rect 13960 -630 13980 -600
rect 13910 -650 13980 -630
rect 13910 -680 13930 -650
rect 13960 -680 13980 -650
rect 13910 -690 13980 -680
rect 13995 -500 14065 -490
rect 13995 -530 14015 -500
rect 14045 -530 14065 -500
rect 13995 -550 14065 -530
rect 13995 -580 14015 -550
rect 14045 -580 14065 -550
rect 13995 -600 14065 -580
rect 13995 -630 14015 -600
rect 14045 -630 14065 -600
rect 13995 -650 14065 -630
rect 13995 -680 14015 -650
rect 14045 -680 14065 -650
rect 13995 -690 14065 -680
rect 14080 -500 14150 -490
rect 14080 -530 14100 -500
rect 14130 -530 14150 -500
rect 14080 -550 14150 -530
rect 14080 -580 14100 -550
rect 14130 -580 14150 -550
rect 14080 -600 14150 -580
rect 14080 -630 14100 -600
rect 14130 -630 14150 -600
rect 14080 -650 14150 -630
rect 14080 -680 14100 -650
rect 14130 -680 14150 -650
rect 14080 -690 14150 -680
rect 14165 -500 14235 -490
rect 14165 -530 14185 -500
rect 14215 -530 14235 -500
rect 14165 -550 14235 -530
rect 14165 -580 14185 -550
rect 14215 -580 14235 -550
rect 14165 -600 14235 -580
rect 14165 -630 14185 -600
rect 14215 -630 14235 -600
rect 14165 -650 14235 -630
rect 14165 -680 14185 -650
rect 14215 -680 14235 -650
rect 14165 -690 14235 -680
rect 14250 -500 14320 -490
rect 14250 -530 14270 -500
rect 14300 -530 14320 -500
rect 14250 -550 14320 -530
rect 14250 -580 14270 -550
rect 14300 -580 14320 -550
rect 14250 -600 14320 -580
rect 14250 -630 14270 -600
rect 14300 -630 14320 -600
rect 14250 -650 14320 -630
rect 14250 -680 14270 -650
rect 14300 -680 14320 -650
rect 14250 -690 14320 -680
rect 14335 -500 14405 -490
rect 14335 -530 14355 -500
rect 14385 -530 14405 -500
rect 14335 -550 14405 -530
rect 14335 -580 14355 -550
rect 14385 -580 14405 -550
rect 14335 -600 14405 -580
rect 14335 -630 14355 -600
rect 14385 -630 14405 -600
rect 14335 -650 14405 -630
rect 14335 -680 14355 -650
rect 14385 -680 14405 -650
rect 14335 -690 14405 -680
rect 14420 -500 14490 -490
rect 14420 -530 14440 -500
rect 14470 -530 14490 -500
rect 14420 -550 14490 -530
rect 14420 -580 14440 -550
rect 14470 -580 14490 -550
rect 14420 -600 14490 -580
rect 14420 -630 14440 -600
rect 14470 -630 14490 -600
rect 14420 -650 14490 -630
rect 14420 -680 14440 -650
rect 14470 -680 14490 -650
rect 14420 -690 14490 -680
rect 14505 -500 14575 -490
rect 14505 -530 14525 -500
rect 14555 -530 14575 -500
rect 14505 -550 14575 -530
rect 14505 -580 14525 -550
rect 14555 -580 14575 -550
rect 14505 -600 14575 -580
rect 14505 -630 14525 -600
rect 14555 -630 14575 -600
rect 14505 -650 14575 -630
rect 14505 -680 14525 -650
rect 14555 -680 14575 -650
rect 14505 -690 14575 -680
rect 14590 -500 14660 -490
rect 14590 -530 14610 -500
rect 14640 -530 14660 -500
rect 14590 -550 14660 -530
rect 14590 -580 14610 -550
rect 14640 -580 14660 -550
rect 14590 -600 14660 -580
rect 14590 -630 14610 -600
rect 14640 -630 14660 -600
rect 14590 -650 14660 -630
rect 14590 -680 14610 -650
rect 14640 -680 14660 -650
rect 14590 -690 14660 -680
rect 14675 -500 14745 -490
rect 14675 -530 14695 -500
rect 14725 -530 14745 -500
rect 14675 -550 14745 -530
rect 14675 -580 14695 -550
rect 14725 -580 14745 -550
rect 14675 -600 14745 -580
rect 14675 -630 14695 -600
rect 14725 -630 14745 -600
rect 14675 -650 14745 -630
rect 14675 -680 14695 -650
rect 14725 -680 14745 -650
rect 14675 -690 14745 -680
rect 14760 -500 14830 -490
rect 14760 -530 14780 -500
rect 14810 -530 14830 -500
rect 14760 -550 14830 -530
rect 14760 -580 14780 -550
rect 14810 -580 14830 -550
rect 14760 -600 14830 -580
rect 14760 -630 14780 -600
rect 14810 -630 14830 -600
rect 14760 -650 14830 -630
rect 14760 -680 14780 -650
rect 14810 -680 14830 -650
rect 14760 -690 14830 -680
rect 14845 -500 14915 -490
rect 14845 -530 14865 -500
rect 14895 -530 14915 -500
rect 14845 -550 14915 -530
rect 14845 -580 14865 -550
rect 14895 -580 14915 -550
rect 14845 -600 14915 -580
rect 14845 -630 14865 -600
rect 14895 -630 14915 -600
rect 14845 -650 14915 -630
rect 14845 -680 14865 -650
rect 14895 -680 14915 -650
rect 14845 -690 14915 -680
rect 14930 -500 15000 -490
rect 14930 -530 14950 -500
rect 14980 -530 15000 -500
rect 14930 -550 15000 -530
rect 14930 -580 14950 -550
rect 14980 -580 15000 -550
rect 14930 -600 15000 -580
rect 14930 -630 14950 -600
rect 14980 -630 15000 -600
rect 14930 -650 15000 -630
rect 14930 -680 14950 -650
rect 14980 -680 15000 -650
rect 14930 -690 15000 -680
rect 15015 -500 15085 -490
rect 15015 -530 15035 -500
rect 15065 -530 15085 -500
rect 15015 -550 15085 -530
rect 15015 -580 15035 -550
rect 15065 -580 15085 -550
rect 15015 -600 15085 -580
rect 15015 -630 15035 -600
rect 15065 -630 15085 -600
rect 15015 -650 15085 -630
rect 15015 -680 15035 -650
rect 15065 -680 15085 -650
rect 15015 -690 15085 -680
rect 15100 -500 15170 -490
rect 15100 -530 15120 -500
rect 15150 -530 15170 -500
rect 15100 -550 15170 -530
rect 15100 -580 15120 -550
rect 15150 -580 15170 -550
rect 15100 -600 15170 -580
rect 15100 -630 15120 -600
rect 15150 -630 15170 -600
rect 15100 -650 15170 -630
rect 15100 -680 15120 -650
rect 15150 -680 15170 -650
rect 15100 -690 15170 -680
rect 15185 -500 15255 -490
rect 15185 -530 15205 -500
rect 15235 -530 15255 -500
rect 15185 -550 15255 -530
rect 15185 -580 15205 -550
rect 15235 -580 15255 -550
rect 15185 -600 15255 -580
rect 15185 -630 15205 -600
rect 15235 -630 15255 -600
rect 15185 -650 15255 -630
rect 15185 -680 15205 -650
rect 15235 -680 15255 -650
rect 15185 -690 15255 -680
rect 15270 -500 15340 -490
rect 15270 -530 15290 -500
rect 15320 -530 15340 -500
rect 15270 -550 15340 -530
rect 15270 -580 15290 -550
rect 15320 -580 15340 -550
rect 15270 -600 15340 -580
rect 15270 -630 15290 -600
rect 15320 -630 15340 -600
rect 15270 -650 15340 -630
rect 15270 -680 15290 -650
rect 15320 -680 15340 -650
rect 15270 -690 15340 -680
rect 15355 -500 15425 -490
rect 15355 -530 15375 -500
rect 15405 -530 15425 -500
rect 15355 -550 15425 -530
rect 15355 -580 15375 -550
rect 15405 -580 15425 -550
rect 15355 -600 15425 -580
rect 15355 -630 15375 -600
rect 15405 -630 15425 -600
rect 15355 -650 15425 -630
rect 15355 -680 15375 -650
rect 15405 -680 15425 -650
rect 15355 -690 15425 -680
rect 15440 -500 15510 -490
rect 15440 -530 15460 -500
rect 15490 -530 15510 -500
rect 15440 -550 15510 -530
rect 15440 -580 15460 -550
rect 15490 -580 15510 -550
rect 15440 -600 15510 -580
rect 15440 -630 15460 -600
rect 15490 -630 15510 -600
rect 15440 -650 15510 -630
rect 15440 -680 15460 -650
rect 15490 -680 15510 -650
rect 15440 -690 15510 -680
rect 15525 -500 15595 -490
rect 15525 -530 15545 -500
rect 15575 -530 15595 -500
rect 15525 -550 15595 -530
rect 15525 -580 15545 -550
rect 15575 -580 15595 -550
rect 15525 -600 15595 -580
rect 15525 -630 15545 -600
rect 15575 -630 15595 -600
rect 15525 -650 15595 -630
rect 15525 -680 15545 -650
rect 15575 -680 15595 -650
rect 15525 -690 15595 -680
rect 15610 -500 15680 -490
rect 15610 -530 15630 -500
rect 15660 -530 15680 -500
rect 15610 -550 15680 -530
rect 15610 -580 15630 -550
rect 15660 -580 15680 -550
rect 15610 -600 15680 -580
rect 15610 -630 15630 -600
rect 15660 -630 15680 -600
rect 15610 -650 15680 -630
rect 15610 -680 15630 -650
rect 15660 -680 15680 -650
rect 15610 -690 15680 -680
rect 15695 -500 15765 -490
rect 15695 -530 15715 -500
rect 15745 -530 15765 -500
rect 15695 -550 15765 -530
rect 15695 -580 15715 -550
rect 15745 -580 15765 -550
rect 15695 -600 15765 -580
rect 15695 -630 15715 -600
rect 15745 -630 15765 -600
rect 15695 -650 15765 -630
rect 15695 -680 15715 -650
rect 15745 -680 15765 -650
rect 15695 -690 15765 -680
rect 15780 -500 15850 -490
rect 15780 -530 15800 -500
rect 15830 -530 15850 -500
rect 15780 -550 15850 -530
rect 15780 -580 15800 -550
rect 15830 -580 15850 -550
rect 15780 -600 15850 -580
rect 15780 -630 15800 -600
rect 15830 -630 15850 -600
rect 15780 -650 15850 -630
rect 15780 -680 15800 -650
rect 15830 -680 15850 -650
rect 15780 -690 15850 -680
rect 15865 -500 15935 -490
rect 15865 -530 15885 -500
rect 15915 -530 15935 -500
rect 15865 -550 15935 -530
rect 15865 -580 15885 -550
rect 15915 -580 15935 -550
rect 15865 -600 15935 -580
rect 15865 -630 15885 -600
rect 15915 -630 15935 -600
rect 15865 -650 15935 -630
rect 15865 -680 15885 -650
rect 15915 -680 15935 -650
rect 15865 -690 15935 -680
rect 15950 -500 16020 -490
rect 15950 -530 15970 -500
rect 16000 -530 16020 -500
rect 15950 -550 16020 -530
rect 15950 -580 15970 -550
rect 16000 -580 16020 -550
rect 15950 -600 16020 -580
rect 15950 -630 15970 -600
rect 16000 -630 16020 -600
rect 15950 -650 16020 -630
rect 15950 -680 15970 -650
rect 16000 -680 16020 -650
rect 15950 -690 16020 -680
rect 16035 -500 16105 -490
rect 16035 -530 16055 -500
rect 16085 -530 16105 -500
rect 16035 -550 16105 -530
rect 16035 -580 16055 -550
rect 16085 -580 16105 -550
rect 16035 -600 16105 -580
rect 16035 -630 16055 -600
rect 16085 -630 16105 -600
rect 16035 -650 16105 -630
rect 16035 -680 16055 -650
rect 16085 -680 16105 -650
rect 16035 -690 16105 -680
rect 16120 -500 16190 -490
rect 16120 -530 16140 -500
rect 16170 -530 16190 -500
rect 16120 -550 16190 -530
rect 16120 -580 16140 -550
rect 16170 -580 16190 -550
rect 16120 -600 16190 -580
rect 16120 -630 16140 -600
rect 16170 -630 16190 -600
rect 16120 -650 16190 -630
rect 16120 -680 16140 -650
rect 16170 -680 16190 -650
rect 16120 -690 16190 -680
rect 16205 -500 16275 -490
rect 16205 -530 16225 -500
rect 16255 -530 16275 -500
rect 16205 -550 16275 -530
rect 16205 -580 16225 -550
rect 16255 -580 16275 -550
rect 16205 -600 16275 -580
rect 16205 -630 16225 -600
rect 16255 -630 16275 -600
rect 16205 -650 16275 -630
rect 16205 -680 16225 -650
rect 16255 -680 16275 -650
rect 16205 -690 16275 -680
rect 16290 -500 16360 -490
rect 16290 -530 16310 -500
rect 16340 -530 16360 -500
rect 16290 -550 16360 -530
rect 16290 -580 16310 -550
rect 16340 -580 16360 -550
rect 16290 -600 16360 -580
rect 16290 -630 16310 -600
rect 16340 -630 16360 -600
rect 16290 -650 16360 -630
rect 16290 -680 16310 -650
rect 16340 -680 16360 -650
rect 16290 -690 16360 -680
rect 16375 -500 16445 -490
rect 16375 -530 16395 -500
rect 16425 -530 16445 -500
rect 16375 -550 16445 -530
rect 16375 -580 16395 -550
rect 16425 -580 16445 -550
rect 16375 -600 16445 -580
rect 16375 -630 16395 -600
rect 16425 -630 16445 -600
rect 16375 -650 16445 -630
rect 16375 -680 16395 -650
rect 16425 -680 16445 -650
rect 16375 -690 16445 -680
rect 16460 -500 16530 -490
rect 16460 -530 16480 -500
rect 16510 -530 16530 -500
rect 16460 -550 16530 -530
rect 16460 -580 16480 -550
rect 16510 -580 16530 -550
rect 16460 -600 16530 -580
rect 16460 -630 16480 -600
rect 16510 -630 16530 -600
rect 16460 -650 16530 -630
rect 16460 -680 16480 -650
rect 16510 -680 16530 -650
rect 16460 -690 16530 -680
rect 16545 -500 16615 -490
rect 16545 -530 16565 -500
rect 16595 -530 16615 -500
rect 16545 -550 16615 -530
rect 16545 -580 16565 -550
rect 16595 -580 16615 -550
rect 16545 -600 16615 -580
rect 16545 -630 16565 -600
rect 16595 -630 16615 -600
rect 16545 -650 16615 -630
rect 16545 -680 16565 -650
rect 16595 -680 16615 -650
rect 16545 -690 16615 -680
rect 16630 -500 16700 -490
rect 16630 -530 16650 -500
rect 16680 -530 16700 -500
rect 16630 -550 16700 -530
rect 16630 -580 16650 -550
rect 16680 -580 16700 -550
rect 16630 -600 16700 -580
rect 16630 -630 16650 -600
rect 16680 -630 16700 -600
rect 16630 -650 16700 -630
rect 16630 -680 16650 -650
rect 16680 -680 16700 -650
rect 16630 -690 16700 -680
rect 16715 -500 16785 -490
rect 16715 -530 16735 -500
rect 16765 -530 16785 -500
rect 16715 -550 16785 -530
rect 16715 -580 16735 -550
rect 16765 -580 16785 -550
rect 16715 -600 16785 -580
rect 16715 -630 16735 -600
rect 16765 -630 16785 -600
rect 16715 -650 16785 -630
rect 16715 -680 16735 -650
rect 16765 -680 16785 -650
rect 16715 -690 16785 -680
rect 16800 -500 16870 -490
rect 16800 -530 16820 -500
rect 16850 -530 16870 -500
rect 16800 -550 16870 -530
rect 16800 -580 16820 -550
rect 16850 -580 16870 -550
rect 16800 -600 16870 -580
rect 16800 -630 16820 -600
rect 16850 -630 16870 -600
rect 16800 -650 16870 -630
rect 16800 -680 16820 -650
rect 16850 -680 16870 -650
rect 16800 -690 16870 -680
rect 16885 -500 16955 -490
rect 16885 -530 16905 -500
rect 16935 -530 16955 -500
rect 16885 -550 16955 -530
rect 16885 -580 16905 -550
rect 16935 -580 16955 -550
rect 16885 -600 16955 -580
rect 16885 -630 16905 -600
rect 16935 -630 16955 -600
rect 16885 -650 16955 -630
rect 16885 -680 16905 -650
rect 16935 -680 16955 -650
rect 16885 -690 16955 -680
rect 16970 -500 17040 -490
rect 16970 -530 16990 -500
rect 17020 -530 17040 -500
rect 16970 -550 17040 -530
rect 16970 -580 16990 -550
rect 17020 -580 17040 -550
rect 16970 -600 17040 -580
rect 16970 -630 16990 -600
rect 17020 -630 17040 -600
rect 16970 -650 17040 -630
rect 16970 -680 16990 -650
rect 17020 -680 17040 -650
rect 16970 -690 17040 -680
rect 17055 -500 17125 -490
rect 17055 -530 17075 -500
rect 17105 -530 17125 -500
rect 17055 -550 17125 -530
rect 17055 -580 17075 -550
rect 17105 -580 17125 -550
rect 17055 -600 17125 -580
rect 17055 -630 17075 -600
rect 17105 -630 17125 -600
rect 17055 -650 17125 -630
rect 17055 -680 17075 -650
rect 17105 -680 17125 -650
rect 17055 -690 17125 -680
rect 17140 -500 17210 -490
rect 17140 -530 17160 -500
rect 17190 -530 17210 -500
rect 17140 -550 17210 -530
rect 17140 -580 17160 -550
rect 17190 -580 17210 -550
rect 17140 -600 17210 -580
rect 17140 -630 17160 -600
rect 17190 -630 17210 -600
rect 17140 -650 17210 -630
rect 17140 -680 17160 -650
rect 17190 -680 17210 -650
rect 17140 -690 17210 -680
rect 17225 -500 17295 -490
rect 17225 -530 17245 -500
rect 17275 -530 17295 -500
rect 17225 -550 17295 -530
rect 17225 -580 17245 -550
rect 17275 -580 17295 -550
rect 17225 -600 17295 -580
rect 17225 -630 17245 -600
rect 17275 -630 17295 -600
rect 17225 -650 17295 -630
rect 17225 -680 17245 -650
rect 17275 -680 17295 -650
rect 17225 -690 17295 -680
rect 17310 -500 17380 -490
rect 17310 -530 17330 -500
rect 17360 -530 17380 -500
rect 17310 -550 17380 -530
rect 17310 -580 17330 -550
rect 17360 -580 17380 -550
rect 17310 -600 17380 -580
rect 17310 -630 17330 -600
rect 17360 -630 17380 -600
rect 17310 -650 17380 -630
rect 17310 -680 17330 -650
rect 17360 -680 17380 -650
rect 17310 -690 17380 -680
rect 17395 -500 17465 -490
rect 17395 -530 17415 -500
rect 17445 -530 17465 -500
rect 17395 -550 17465 -530
rect 17395 -580 17415 -550
rect 17445 -580 17465 -550
rect 17395 -600 17465 -580
rect 17395 -630 17415 -600
rect 17445 -630 17465 -600
rect 17395 -650 17465 -630
rect 17395 -680 17415 -650
rect 17445 -680 17465 -650
rect 17395 -690 17465 -680
rect 17480 -500 17550 -490
rect 17480 -530 17500 -500
rect 17530 -530 17550 -500
rect 17480 -550 17550 -530
rect 17480 -580 17500 -550
rect 17530 -580 17550 -550
rect 17480 -600 17550 -580
rect 17480 -630 17500 -600
rect 17530 -630 17550 -600
rect 17480 -650 17550 -630
rect 17480 -680 17500 -650
rect 17530 -680 17550 -650
rect 17480 -690 17550 -680
rect 17565 -500 17635 -490
rect 17565 -530 17585 -500
rect 17615 -530 17635 -500
rect 17565 -550 17635 -530
rect 17565 -580 17585 -550
rect 17615 -580 17635 -550
rect 17565 -600 17635 -580
rect 17565 -630 17585 -600
rect 17615 -630 17635 -600
rect 17565 -650 17635 -630
rect 17565 -680 17585 -650
rect 17615 -680 17635 -650
rect 17565 -690 17635 -680
rect 17650 -500 17720 -490
rect 17650 -530 17670 -500
rect 17700 -530 17720 -500
rect 17650 -550 17720 -530
rect 17650 -580 17670 -550
rect 17700 -580 17720 -550
rect 17650 -600 17720 -580
rect 17650 -630 17670 -600
rect 17700 -630 17720 -600
rect 17650 -650 17720 -630
rect 17650 -680 17670 -650
rect 17700 -680 17720 -650
rect 17650 -690 17720 -680
rect 17735 -500 17805 -490
rect 17735 -530 17755 -500
rect 17785 -530 17805 -500
rect 17735 -550 17805 -530
rect 17735 -580 17755 -550
rect 17785 -580 17805 -550
rect 17735 -600 17805 -580
rect 17735 -630 17755 -600
rect 17785 -630 17805 -600
rect 17735 -650 17805 -630
rect 17735 -680 17755 -650
rect 17785 -680 17805 -650
rect 17735 -690 17805 -680
rect 17820 -500 17890 -490
rect 17820 -530 17840 -500
rect 17870 -530 17890 -500
rect 17820 -550 17890 -530
rect 17820 -580 17840 -550
rect 17870 -580 17890 -550
rect 17820 -600 17890 -580
rect 17820 -630 17840 -600
rect 17870 -630 17890 -600
rect 17820 -650 17890 -630
rect 17820 -680 17840 -650
rect 17870 -680 17890 -650
rect 17820 -690 17890 -680
rect 17905 -500 17975 -490
rect 17905 -530 17925 -500
rect 17955 -530 17975 -500
rect 17905 -550 17975 -530
rect 17905 -580 17925 -550
rect 17955 -580 17975 -550
rect 17905 -600 17975 -580
rect 17905 -630 17925 -600
rect 17955 -630 17975 -600
rect 17905 -650 17975 -630
rect 17905 -680 17925 -650
rect 17955 -680 17975 -650
rect 17905 -690 17975 -680
rect 17990 -500 18060 -490
rect 17990 -530 18010 -500
rect 18040 -530 18060 -500
rect 17990 -550 18060 -530
rect 17990 -580 18010 -550
rect 18040 -580 18060 -550
rect 17990 -600 18060 -580
rect 17990 -630 18010 -600
rect 18040 -630 18060 -600
rect 17990 -650 18060 -630
rect 17990 -680 18010 -650
rect 18040 -680 18060 -650
rect 17990 -690 18060 -680
rect 18075 -500 18145 -490
rect 18075 -530 18095 -500
rect 18125 -530 18145 -500
rect 18075 -550 18145 -530
rect 18075 -580 18095 -550
rect 18125 -580 18145 -550
rect 18075 -600 18145 -580
rect 18075 -630 18095 -600
rect 18125 -630 18145 -600
rect 18075 -650 18145 -630
rect 18075 -680 18095 -650
rect 18125 -680 18145 -650
rect 18075 -690 18145 -680
rect 18160 -500 18230 -490
rect 18160 -530 18180 -500
rect 18210 -530 18230 -500
rect 18160 -550 18230 -530
rect 18160 -580 18180 -550
rect 18210 -580 18230 -550
rect 18160 -600 18230 -580
rect 18160 -630 18180 -600
rect 18210 -630 18230 -600
rect 18160 -650 18230 -630
rect 18160 -680 18180 -650
rect 18210 -680 18230 -650
rect 18160 -690 18230 -680
rect 18245 -500 18315 -490
rect 18245 -530 18265 -500
rect 18295 -530 18315 -500
rect 18245 -550 18315 -530
rect 18245 -580 18265 -550
rect 18295 -580 18315 -550
rect 18245 -600 18315 -580
rect 18245 -630 18265 -600
rect 18295 -630 18315 -600
rect 18245 -650 18315 -630
rect 18245 -680 18265 -650
rect 18295 -680 18315 -650
rect 18245 -690 18315 -680
rect 18330 -500 18400 -490
rect 18330 -530 18350 -500
rect 18380 -530 18400 -500
rect 18330 -550 18400 -530
rect 18330 -580 18350 -550
rect 18380 -580 18400 -550
rect 18330 -600 18400 -580
rect 18330 -630 18350 -600
rect 18380 -630 18400 -600
rect 18330 -650 18400 -630
rect 18330 -680 18350 -650
rect 18380 -680 18400 -650
rect 18330 -690 18400 -680
rect 18415 -500 18485 -490
rect 18415 -530 18435 -500
rect 18465 -530 18485 -500
rect 18415 -550 18485 -530
rect 18415 -580 18435 -550
rect 18465 -580 18485 -550
rect 18415 -600 18485 -580
rect 18415 -630 18435 -600
rect 18465 -630 18485 -600
rect 18415 -650 18485 -630
rect 18415 -680 18435 -650
rect 18465 -680 18485 -650
rect 18415 -690 18485 -680
rect 18500 -500 18570 -490
rect 18500 -530 18520 -500
rect 18550 -530 18570 -500
rect 18500 -550 18570 -530
rect 18500 -580 18520 -550
rect 18550 -580 18570 -550
rect 18500 -600 18570 -580
rect 18500 -630 18520 -600
rect 18550 -630 18570 -600
rect 18500 -650 18570 -630
rect 18500 -680 18520 -650
rect 18550 -680 18570 -650
rect 18500 -690 18570 -680
rect 18585 -500 18655 -490
rect 18585 -530 18605 -500
rect 18635 -530 18655 -500
rect 18585 -550 18655 -530
rect 18585 -580 18605 -550
rect 18635 -580 18655 -550
rect 18585 -600 18655 -580
rect 18585 -630 18605 -600
rect 18635 -630 18655 -600
rect 18585 -650 18655 -630
rect 18585 -680 18605 -650
rect 18635 -680 18655 -650
rect 18585 -690 18655 -680
rect 18670 -500 18740 -490
rect 18670 -530 18690 -500
rect 18720 -530 18740 -500
rect 18670 -550 18740 -530
rect 18670 -580 18690 -550
rect 18720 -580 18740 -550
rect 18670 -600 18740 -580
rect 18670 -630 18690 -600
rect 18720 -630 18740 -600
rect 18670 -650 18740 -630
rect 18670 -680 18690 -650
rect 18720 -680 18740 -650
rect 18670 -690 18740 -680
rect 18755 -500 18825 -490
rect 18755 -530 18775 -500
rect 18805 -530 18825 -500
rect 18755 -550 18825 -530
rect 18755 -580 18775 -550
rect 18805 -580 18825 -550
rect 18755 -600 18825 -580
rect 18755 -630 18775 -600
rect 18805 -630 18825 -600
rect 18755 -650 18825 -630
rect 18755 -680 18775 -650
rect 18805 -680 18825 -650
rect 18755 -690 18825 -680
rect 18840 -500 18910 -490
rect 18840 -530 18860 -500
rect 18890 -530 18910 -500
rect 18840 -550 18910 -530
rect 18840 -580 18860 -550
rect 18890 -580 18910 -550
rect 18840 -600 18910 -580
rect 18840 -630 18860 -600
rect 18890 -630 18910 -600
rect 18840 -650 18910 -630
rect 18840 -680 18860 -650
rect 18890 -680 18910 -650
rect 18840 -690 18910 -680
rect 18925 -500 18995 -490
rect 18925 -530 18945 -500
rect 18975 -530 18995 -500
rect 18925 -550 18995 -530
rect 18925 -580 18945 -550
rect 18975 -580 18995 -550
rect 18925 -600 18995 -580
rect 18925 -630 18945 -600
rect 18975 -630 18995 -600
rect 18925 -650 18995 -630
rect 18925 -680 18945 -650
rect 18975 -680 18995 -650
rect 18925 -690 18995 -680
rect 19010 -500 19080 -490
rect 19010 -530 19030 -500
rect 19060 -530 19080 -500
rect 19010 -550 19080 -530
rect 19010 -580 19030 -550
rect 19060 -580 19080 -550
rect 19010 -600 19080 -580
rect 19010 -630 19030 -600
rect 19060 -630 19080 -600
rect 19010 -650 19080 -630
rect 19010 -680 19030 -650
rect 19060 -680 19080 -650
rect 19010 -690 19080 -680
rect 19095 -500 19165 -490
rect 19095 -530 19115 -500
rect 19145 -530 19165 -500
rect 19095 -550 19165 -530
rect 19095 -580 19115 -550
rect 19145 -580 19165 -550
rect 19095 -600 19165 -580
rect 19095 -630 19115 -600
rect 19145 -630 19165 -600
rect 19095 -650 19165 -630
rect 19095 -680 19115 -650
rect 19145 -680 19165 -650
rect 19095 -690 19165 -680
rect 19180 -500 19250 -490
rect 19180 -530 19200 -500
rect 19230 -530 19250 -500
rect 19180 -550 19250 -530
rect 19180 -580 19200 -550
rect 19230 -580 19250 -550
rect 19180 -600 19250 -580
rect 19180 -630 19200 -600
rect 19230 -630 19250 -600
rect 19180 -650 19250 -630
rect 19180 -680 19200 -650
rect 19230 -680 19250 -650
rect 19180 -690 19250 -680
rect 19265 -500 19335 -490
rect 19265 -530 19285 -500
rect 19315 -530 19335 -500
rect 19265 -550 19335 -530
rect 19265 -580 19285 -550
rect 19315 -580 19335 -550
rect 19265 -600 19335 -580
rect 19265 -630 19285 -600
rect 19315 -630 19335 -600
rect 19265 -650 19335 -630
rect 19265 -680 19285 -650
rect 19315 -680 19335 -650
rect 19265 -690 19335 -680
rect 19350 -500 19420 -490
rect 19350 -530 19370 -500
rect 19400 -530 19420 -500
rect 19350 -550 19420 -530
rect 19350 -580 19370 -550
rect 19400 -580 19420 -550
rect 19350 -600 19420 -580
rect 19350 -630 19370 -600
rect 19400 -630 19420 -600
rect 19350 -650 19420 -630
rect 19350 -680 19370 -650
rect 19400 -680 19420 -650
rect 19350 -690 19420 -680
rect 19435 -500 19505 -490
rect 19435 -530 19455 -500
rect 19485 -530 19505 -500
rect 19435 -550 19505 -530
rect 19435 -580 19455 -550
rect 19485 -580 19505 -550
rect 19435 -600 19505 -580
rect 19435 -630 19455 -600
rect 19485 -630 19505 -600
rect 19435 -650 19505 -630
rect 19435 -680 19455 -650
rect 19485 -680 19505 -650
rect 19435 -690 19505 -680
rect 19520 -500 19590 -490
rect 19520 -530 19540 -500
rect 19570 -530 19590 -500
rect 19520 -550 19590 -530
rect 19520 -580 19540 -550
rect 19570 -580 19590 -550
rect 19520 -600 19590 -580
rect 19520 -630 19540 -600
rect 19570 -630 19590 -600
rect 19520 -650 19590 -630
rect 19520 -680 19540 -650
rect 19570 -680 19590 -650
rect 19520 -690 19590 -680
rect 19605 -500 19675 -490
rect 19605 -530 19625 -500
rect 19655 -530 19675 -500
rect 19605 -550 19675 -530
rect 19605 -580 19625 -550
rect 19655 -580 19675 -550
rect 19605 -600 19675 -580
rect 19605 -630 19625 -600
rect 19655 -630 19675 -600
rect 19605 -650 19675 -630
rect 19605 -680 19625 -650
rect 19655 -680 19675 -650
rect 19605 -690 19675 -680
rect 19690 -500 19760 -490
rect 19690 -530 19710 -500
rect 19740 -530 19760 -500
rect 19690 -550 19760 -530
rect 19690 -580 19710 -550
rect 19740 -580 19760 -550
rect 19690 -600 19760 -580
rect 19690 -630 19710 -600
rect 19740 -630 19760 -600
rect 19690 -650 19760 -630
rect 19690 -680 19710 -650
rect 19740 -680 19760 -650
rect 19690 -690 19760 -680
rect 19775 -500 19845 -490
rect 19775 -530 19795 -500
rect 19825 -530 19845 -500
rect 19775 -550 19845 -530
rect 19775 -580 19795 -550
rect 19825 -580 19845 -550
rect 19775 -600 19845 -580
rect 19775 -630 19795 -600
rect 19825 -630 19845 -600
rect 19775 -650 19845 -630
rect 19775 -680 19795 -650
rect 19825 -680 19845 -650
rect 19775 -690 19845 -680
rect 19860 -500 19930 -490
rect 19860 -530 19880 -500
rect 19910 -530 19930 -500
rect 19860 -550 19930 -530
rect 19860 -580 19880 -550
rect 19910 -580 19930 -550
rect 19860 -600 19930 -580
rect 19860 -630 19880 -600
rect 19910 -630 19930 -600
rect 19860 -650 19930 -630
rect 19860 -680 19880 -650
rect 19910 -680 19930 -650
rect 19860 -690 19930 -680
rect 19945 -500 20015 -490
rect 19945 -530 19965 -500
rect 19995 -530 20015 -500
rect 19945 -550 20015 -530
rect 19945 -580 19965 -550
rect 19995 -580 20015 -550
rect 19945 -600 20015 -580
rect 19945 -630 19965 -600
rect 19995 -630 20015 -600
rect 19945 -650 20015 -630
rect 19945 -680 19965 -650
rect 19995 -680 20015 -650
rect 19945 -690 20015 -680
rect 20030 -500 20100 -490
rect 20030 -530 20050 -500
rect 20080 -530 20100 -500
rect 20030 -550 20100 -530
rect 20030 -580 20050 -550
rect 20080 -580 20100 -550
rect 20030 -600 20100 -580
rect 20030 -630 20050 -600
rect 20080 -630 20100 -600
rect 20030 -650 20100 -630
rect 20030 -680 20050 -650
rect 20080 -680 20100 -650
rect 20030 -690 20100 -680
rect 20115 -500 20185 -490
rect 20115 -530 20135 -500
rect 20165 -530 20185 -500
rect 20115 -550 20185 -530
rect 20115 -580 20135 -550
rect 20165 -580 20185 -550
rect 20115 -600 20185 -580
rect 20115 -630 20135 -600
rect 20165 -630 20185 -600
rect 20115 -650 20185 -630
rect 20115 -680 20135 -650
rect 20165 -680 20185 -650
rect 20115 -690 20185 -680
rect 20200 -500 20270 -490
rect 20200 -530 20220 -500
rect 20250 -530 20270 -500
rect 20200 -550 20270 -530
rect 20200 -580 20220 -550
rect 20250 -580 20270 -550
rect 20200 -600 20270 -580
rect 20200 -630 20220 -600
rect 20250 -630 20270 -600
rect 20200 -650 20270 -630
rect 20200 -680 20220 -650
rect 20250 -680 20270 -650
rect 20200 -690 20270 -680
rect 20285 -500 20355 -490
rect 20285 -530 20305 -500
rect 20335 -530 20355 -500
rect 20285 -550 20355 -530
rect 20285 -580 20305 -550
rect 20335 -580 20355 -550
rect 20285 -600 20355 -580
rect 20285 -630 20305 -600
rect 20335 -630 20355 -600
rect 20285 -650 20355 -630
rect 20285 -680 20305 -650
rect 20335 -680 20355 -650
rect 20285 -690 20355 -680
rect 20370 -500 20440 -490
rect 20370 -530 20390 -500
rect 20420 -530 20440 -500
rect 20370 -550 20440 -530
rect 20370 -580 20390 -550
rect 20420 -580 20440 -550
rect 20370 -600 20440 -580
rect 20370 -630 20390 -600
rect 20420 -630 20440 -600
rect 20370 -650 20440 -630
rect 20370 -680 20390 -650
rect 20420 -680 20440 -650
rect 20370 -690 20440 -680
rect 20455 -500 20525 -490
rect 20455 -530 20475 -500
rect 20505 -530 20525 -500
rect 20455 -550 20525 -530
rect 20455 -580 20475 -550
rect 20505 -580 20525 -550
rect 20455 -600 20525 -580
rect 20455 -630 20475 -600
rect 20505 -630 20525 -600
rect 20455 -650 20525 -630
rect 20455 -680 20475 -650
rect 20505 -680 20525 -650
rect 20455 -690 20525 -680
rect 20540 -500 20610 -490
rect 20540 -530 20560 -500
rect 20590 -530 20610 -500
rect 20540 -550 20610 -530
rect 20540 -580 20560 -550
rect 20590 -580 20610 -550
rect 20540 -600 20610 -580
rect 20540 -630 20560 -600
rect 20590 -630 20610 -600
rect 20540 -650 20610 -630
rect 20540 -680 20560 -650
rect 20590 -680 20610 -650
rect 20540 -690 20610 -680
rect 20625 -500 20695 -490
rect 20625 -530 20645 -500
rect 20675 -530 20695 -500
rect 20625 -550 20695 -530
rect 20625 -580 20645 -550
rect 20675 -580 20695 -550
rect 20625 -600 20695 -580
rect 20625 -630 20645 -600
rect 20675 -630 20695 -600
rect 20625 -650 20695 -630
rect 20625 -680 20645 -650
rect 20675 -680 20695 -650
rect 20625 -690 20695 -680
rect 20710 -500 20780 -490
rect 20710 -530 20730 -500
rect 20760 -530 20780 -500
rect 20710 -550 20780 -530
rect 20710 -580 20730 -550
rect 20760 -580 20780 -550
rect 20710 -600 20780 -580
rect 20710 -630 20730 -600
rect 20760 -630 20780 -600
rect 20710 -650 20780 -630
rect 20710 -680 20730 -650
rect 20760 -680 20780 -650
rect 20710 -690 20780 -680
rect 20795 -500 20865 -490
rect 20795 -530 20815 -500
rect 20845 -530 20865 -500
rect 20795 -550 20865 -530
rect 20795 -580 20815 -550
rect 20845 -580 20865 -550
rect 20795 -600 20865 -580
rect 20795 -630 20815 -600
rect 20845 -630 20865 -600
rect 20795 -650 20865 -630
rect 20795 -680 20815 -650
rect 20845 -680 20865 -650
rect 20795 -690 20865 -680
rect 20880 -500 20950 -490
rect 20880 -530 20900 -500
rect 20930 -530 20950 -500
rect 20880 -550 20950 -530
rect 20880 -580 20900 -550
rect 20930 -580 20950 -550
rect 20880 -600 20950 -580
rect 20880 -630 20900 -600
rect 20930 -630 20950 -600
rect 20880 -650 20950 -630
rect 20880 -680 20900 -650
rect 20930 -680 20950 -650
rect 20880 -690 20950 -680
rect 20965 -500 21035 -490
rect 20965 -530 20985 -500
rect 21015 -530 21035 -500
rect 20965 -550 21035 -530
rect 20965 -580 20985 -550
rect 21015 -580 21035 -550
rect 20965 -600 21035 -580
rect 20965 -630 20985 -600
rect 21015 -630 21035 -600
rect 20965 -650 21035 -630
rect 20965 -680 20985 -650
rect 21015 -680 21035 -650
rect 20965 -690 21035 -680
rect 21050 -500 21120 -490
rect 21050 -530 21070 -500
rect 21100 -530 21120 -500
rect 21050 -550 21120 -530
rect 21050 -580 21070 -550
rect 21100 -580 21120 -550
rect 21050 -600 21120 -580
rect 21050 -630 21070 -600
rect 21100 -630 21120 -600
rect 21050 -650 21120 -630
rect 21050 -680 21070 -650
rect 21100 -680 21120 -650
rect 21050 -690 21120 -680
rect 21135 -500 21205 -490
rect 21135 -530 21155 -500
rect 21185 -530 21205 -500
rect 21135 -550 21205 -530
rect 21135 -580 21155 -550
rect 21185 -580 21205 -550
rect 21135 -600 21205 -580
rect 21135 -630 21155 -600
rect 21185 -630 21205 -600
rect 21135 -650 21205 -630
rect 21135 -680 21155 -650
rect 21185 -680 21205 -650
rect 21135 -690 21205 -680
rect 21220 -500 21290 -490
rect 21220 -530 21240 -500
rect 21270 -530 21290 -500
rect 21220 -550 21290 -530
rect 21220 -580 21240 -550
rect 21270 -580 21290 -550
rect 21220 -600 21290 -580
rect 21220 -630 21240 -600
rect 21270 -630 21290 -600
rect 21220 -650 21290 -630
rect 21220 -680 21240 -650
rect 21270 -680 21290 -650
rect 21220 -690 21290 -680
rect 21305 -500 21375 -490
rect 21305 -530 21325 -500
rect 21355 -530 21375 -500
rect 21305 -550 21375 -530
rect 21305 -580 21325 -550
rect 21355 -580 21375 -550
rect 21305 -600 21375 -580
rect 21305 -630 21325 -600
rect 21355 -630 21375 -600
rect 21305 -650 21375 -630
rect 21305 -680 21325 -650
rect 21355 -680 21375 -650
rect 21305 -690 21375 -680
rect 21390 -500 21460 -490
rect 21390 -530 21410 -500
rect 21440 -530 21460 -500
rect 21390 -550 21460 -530
rect 21390 -580 21410 -550
rect 21440 -580 21460 -550
rect 21390 -600 21460 -580
rect 21390 -630 21410 -600
rect 21440 -630 21460 -600
rect 21390 -650 21460 -630
rect 21390 -680 21410 -650
rect 21440 -680 21460 -650
rect 21390 -690 21460 -680
rect 21475 -500 21545 -490
rect 21475 -530 21495 -500
rect 21525 -530 21545 -500
rect 21475 -550 21545 -530
rect 21475 -580 21495 -550
rect 21525 -580 21545 -550
rect 21475 -600 21545 -580
rect 21475 -630 21495 -600
rect 21525 -630 21545 -600
rect 21475 -650 21545 -630
rect 21475 -680 21495 -650
rect 21525 -680 21545 -650
rect 21475 -690 21545 -680
rect 21560 -500 21630 -490
rect 21560 -530 21580 -500
rect 21610 -530 21630 -500
rect 21560 -550 21630 -530
rect 21560 -580 21580 -550
rect 21610 -580 21630 -550
rect 21560 -600 21630 -580
rect 21560 -630 21580 -600
rect 21610 -630 21630 -600
rect 21560 -650 21630 -630
rect 21560 -680 21580 -650
rect 21610 -680 21630 -650
rect 21560 -690 21630 -680
rect 21645 -500 21715 -490
rect 21645 -530 21665 -500
rect 21695 -530 21715 -500
rect 21645 -550 21715 -530
rect 21645 -580 21665 -550
rect 21695 -580 21715 -550
rect 21645 -600 21715 -580
rect 21645 -630 21665 -600
rect 21695 -630 21715 -600
rect 21645 -650 21715 -630
rect 21645 -680 21665 -650
rect 21695 -680 21715 -650
rect 21645 -690 21715 -680
rect 21730 -500 21800 -490
rect 21730 -530 21750 -500
rect 21780 -530 21800 -500
rect 21730 -550 21800 -530
rect 21730 -580 21750 -550
rect 21780 -580 21800 -550
rect 21730 -600 21800 -580
rect 21730 -630 21750 -600
rect 21780 -630 21800 -600
rect 21730 -650 21800 -630
rect 21730 -680 21750 -650
rect 21780 -680 21800 -650
rect 21730 -690 21800 -680
rect 21815 -500 21885 -490
rect 21815 -530 21835 -500
rect 21865 -530 21885 -500
rect 21815 -550 21885 -530
rect 21815 -580 21835 -550
rect 21865 -580 21885 -550
rect 21815 -600 21885 -580
rect 21815 -630 21835 -600
rect 21865 -630 21885 -600
rect 21815 -650 21885 -630
rect 21815 -680 21835 -650
rect 21865 -680 21885 -650
rect 21815 -690 21885 -680
rect 21900 -500 21970 -490
rect 21900 -530 21920 -500
rect 21950 -530 21970 -500
rect 21900 -550 21970 -530
rect 21900 -580 21920 -550
rect 21950 -580 21970 -550
rect 21900 -600 21970 -580
rect 21900 -630 21920 -600
rect 21950 -630 21970 -600
rect 21900 -650 21970 -630
rect 21900 -680 21920 -650
rect 21950 -680 21970 -650
rect 21900 -690 21970 -680
rect 21985 -500 22055 -490
rect 21985 -530 22005 -500
rect 22035 -530 22055 -500
rect 21985 -550 22055 -530
rect 21985 -580 22005 -550
rect 22035 -580 22055 -550
rect 21985 -600 22055 -580
rect 21985 -630 22005 -600
rect 22035 -630 22055 -600
rect 21985 -650 22055 -630
rect 21985 -680 22005 -650
rect 22035 -680 22055 -650
rect 21985 -690 22055 -680
rect 22070 -500 22140 -490
rect 22070 -530 22090 -500
rect 22120 -530 22140 -500
rect 22070 -550 22140 -530
rect 22070 -580 22090 -550
rect 22120 -580 22140 -550
rect 22070 -600 22140 -580
rect 22070 -630 22090 -600
rect 22120 -630 22140 -600
rect 22070 -650 22140 -630
rect 22070 -680 22090 -650
rect 22120 -680 22140 -650
rect 22070 -690 22140 -680
rect 22155 -500 22225 -490
rect 22155 -530 22175 -500
rect 22205 -530 22225 -500
rect 22155 -550 22225 -530
rect 22155 -580 22175 -550
rect 22205 -580 22225 -550
rect 22155 -600 22225 -580
rect 22155 -630 22175 -600
rect 22205 -630 22225 -600
rect 22155 -650 22225 -630
rect 22155 -680 22175 -650
rect 22205 -680 22225 -650
rect 22155 -690 22225 -680
rect 22240 -500 22310 -490
rect 22240 -530 22260 -500
rect 22290 -530 22310 -500
rect 22240 -550 22310 -530
rect 22240 -580 22260 -550
rect 22290 -580 22310 -550
rect 22240 -600 22310 -580
rect 22240 -630 22260 -600
rect 22290 -630 22310 -600
rect 22240 -650 22310 -630
rect 22240 -680 22260 -650
rect 22290 -680 22310 -650
rect 22240 -690 22310 -680
rect 22325 -500 22395 -490
rect 22325 -530 22345 -500
rect 22375 -530 22395 -500
rect 22325 -550 22395 -530
rect 22325 -580 22345 -550
rect 22375 -580 22395 -550
rect 22325 -600 22395 -580
rect 22325 -630 22345 -600
rect 22375 -630 22395 -600
rect 22325 -650 22395 -630
rect 22325 -680 22345 -650
rect 22375 -680 22395 -650
rect 22325 -690 22395 -680
rect 22410 -500 22480 -490
rect 22410 -530 22430 -500
rect 22460 -530 22480 -500
rect 22410 -550 22480 -530
rect 22410 -580 22430 -550
rect 22460 -580 22480 -550
rect 22410 -600 22480 -580
rect 22410 -630 22430 -600
rect 22460 -630 22480 -600
rect 22410 -650 22480 -630
rect 22410 -680 22430 -650
rect 22460 -680 22480 -650
rect 22410 -690 22480 -680
rect 22495 -500 22565 -490
rect 22495 -530 22515 -500
rect 22545 -530 22565 -500
rect 22495 -550 22565 -530
rect 22495 -580 22515 -550
rect 22545 -580 22565 -550
rect 22495 -600 22565 -580
rect 22495 -630 22515 -600
rect 22545 -630 22565 -600
rect 22495 -650 22565 -630
rect 22495 -680 22515 -650
rect 22545 -680 22565 -650
rect 22495 -690 22565 -680
rect 22580 -500 22650 -490
rect 22580 -530 22600 -500
rect 22630 -530 22650 -500
rect 22580 -550 22650 -530
rect 22580 -580 22600 -550
rect 22630 -580 22650 -550
rect 22580 -600 22650 -580
rect 22580 -630 22600 -600
rect 22630 -630 22650 -600
rect 22580 -650 22650 -630
rect 22580 -680 22600 -650
rect 22630 -680 22650 -650
rect 22580 -690 22650 -680
rect 22665 -500 22735 -490
rect 22665 -530 22685 -500
rect 22715 -530 22735 -500
rect 22665 -550 22735 -530
rect 22665 -580 22685 -550
rect 22715 -580 22735 -550
rect 22665 -600 22735 -580
rect 22665 -630 22685 -600
rect 22715 -630 22735 -600
rect 22665 -650 22735 -630
rect 22665 -680 22685 -650
rect 22715 -680 22735 -650
rect 22665 -690 22735 -680
rect 22750 -500 22820 -490
rect 22750 -530 22770 -500
rect 22800 -530 22820 -500
rect 22750 -550 22820 -530
rect 22750 -580 22770 -550
rect 22800 -580 22820 -550
rect 22750 -600 22820 -580
rect 22750 -630 22770 -600
rect 22800 -630 22820 -600
rect 22750 -650 22820 -630
rect 22750 -680 22770 -650
rect 22800 -680 22820 -650
rect 22750 -690 22820 -680
rect 22835 -500 22905 -490
rect 22835 -530 22855 -500
rect 22885 -530 22905 -500
rect 22835 -550 22905 -530
rect 22835 -580 22855 -550
rect 22885 -580 22905 -550
rect 22835 -600 22905 -580
rect 22835 -630 22855 -600
rect 22885 -630 22905 -600
rect 22835 -650 22905 -630
rect 22835 -680 22855 -650
rect 22885 -680 22905 -650
rect 22835 -690 22905 -680
rect 22920 -500 22990 -490
rect 22920 -530 22940 -500
rect 22970 -530 22990 -500
rect 22920 -550 22990 -530
rect 22920 -580 22940 -550
rect 22970 -580 22990 -550
rect 22920 -600 22990 -580
rect 22920 -630 22940 -600
rect 22970 -630 22990 -600
rect 22920 -650 22990 -630
rect 22920 -680 22940 -650
rect 22970 -680 22990 -650
rect 22920 -690 22990 -680
rect 23005 -500 23075 -490
rect 23005 -530 23025 -500
rect 23055 -530 23075 -500
rect 23005 -550 23075 -530
rect 23005 -580 23025 -550
rect 23055 -580 23075 -550
rect 23005 -600 23075 -580
rect 23005 -630 23025 -600
rect 23055 -630 23075 -600
rect 23005 -650 23075 -630
rect 23005 -680 23025 -650
rect 23055 -680 23075 -650
rect 23005 -690 23075 -680
rect 23090 -500 23160 -490
rect 23090 -530 23110 -500
rect 23140 -530 23160 -500
rect 23090 -550 23160 -530
rect 23090 -580 23110 -550
rect 23140 -580 23160 -550
rect 23090 -600 23160 -580
rect 23090 -630 23110 -600
rect 23140 -630 23160 -600
rect 23090 -650 23160 -630
rect 23090 -680 23110 -650
rect 23140 -680 23160 -650
rect 23090 -690 23160 -680
rect 23175 -500 23245 -490
rect 23175 -530 23195 -500
rect 23225 -530 23245 -500
rect 23175 -550 23245 -530
rect 23175 -580 23195 -550
rect 23225 -580 23245 -550
rect 23175 -600 23245 -580
rect 23175 -630 23195 -600
rect 23225 -630 23245 -600
rect 23175 -650 23245 -630
rect 23175 -680 23195 -650
rect 23225 -680 23245 -650
rect 23175 -690 23245 -680
rect 23260 -500 23330 -490
rect 23260 -530 23280 -500
rect 23310 -530 23330 -500
rect 23260 -550 23330 -530
rect 23260 -580 23280 -550
rect 23310 -580 23330 -550
rect 23260 -600 23330 -580
rect 23260 -630 23280 -600
rect 23310 -630 23330 -600
rect 23260 -650 23330 -630
rect 23260 -680 23280 -650
rect 23310 -680 23330 -650
rect 23260 -690 23330 -680
rect 23345 -500 23415 -490
rect 23345 -530 23365 -500
rect 23395 -530 23415 -500
rect 23345 -550 23415 -530
rect 23345 -580 23365 -550
rect 23395 -580 23415 -550
rect 23345 -600 23415 -580
rect 23345 -630 23365 -600
rect 23395 -630 23415 -600
rect 23345 -650 23415 -630
rect 23345 -680 23365 -650
rect 23395 -680 23415 -650
rect 23345 -690 23415 -680
rect 23430 -500 23500 -490
rect 23430 -530 23450 -500
rect 23480 -530 23500 -500
rect 23430 -550 23500 -530
rect 23430 -580 23450 -550
rect 23480 -580 23500 -550
rect 23430 -600 23500 -580
rect 23430 -630 23450 -600
rect 23480 -630 23500 -600
rect 23430 -650 23500 -630
rect 23430 -680 23450 -650
rect 23480 -680 23500 -650
rect 23430 -690 23500 -680
rect 23515 -500 23585 -490
rect 23515 -530 23535 -500
rect 23565 -530 23585 -500
rect 23515 -550 23585 -530
rect 23515 -580 23535 -550
rect 23565 -580 23585 -550
rect 23515 -600 23585 -580
rect 23515 -630 23535 -600
rect 23565 -630 23585 -600
rect 23515 -650 23585 -630
rect 23515 -680 23535 -650
rect 23565 -680 23585 -650
rect 23515 -690 23585 -680
rect 23600 -500 23670 -490
rect 23600 -530 23620 -500
rect 23650 -530 23670 -500
rect 23600 -550 23670 -530
rect 23600 -580 23620 -550
rect 23650 -580 23670 -550
rect 23600 -600 23670 -580
rect 23600 -630 23620 -600
rect 23650 -630 23670 -600
rect 23600 -650 23670 -630
rect 23600 -680 23620 -650
rect 23650 -680 23670 -650
rect 23600 -690 23670 -680
rect 23685 -500 23755 -490
rect 23685 -530 23705 -500
rect 23735 -530 23755 -500
rect 23685 -550 23755 -530
rect 23685 -580 23705 -550
rect 23735 -580 23755 -550
rect 23685 -600 23755 -580
rect 23685 -630 23705 -600
rect 23735 -630 23755 -600
rect 23685 -650 23755 -630
rect 23685 -680 23705 -650
rect 23735 -680 23755 -650
rect 23685 -690 23755 -680
rect 23770 -500 23840 -490
rect 23770 -530 23790 -500
rect 23820 -530 23840 -500
rect 23770 -550 23840 -530
rect 23770 -580 23790 -550
rect 23820 -580 23840 -550
rect 23770 -600 23840 -580
rect 23770 -630 23790 -600
rect 23820 -630 23840 -600
rect 23770 -650 23840 -630
rect 23770 -680 23790 -650
rect 23820 -680 23840 -650
rect 23770 -690 23840 -680
rect 23855 -500 23925 -490
rect 23855 -530 23875 -500
rect 23905 -530 23925 -500
rect 23855 -550 23925 -530
rect 23855 -580 23875 -550
rect 23905 -580 23925 -550
rect 23855 -600 23925 -580
rect 23855 -630 23875 -600
rect 23905 -630 23925 -600
rect 23855 -650 23925 -630
rect 23855 -680 23875 -650
rect 23905 -680 23925 -650
rect 23855 -690 23925 -680
rect 23940 -500 24010 -490
rect 23940 -530 23960 -500
rect 23990 -530 24010 -500
rect 23940 -550 24010 -530
rect 23940 -580 23960 -550
rect 23990 -580 24010 -550
rect 23940 -600 24010 -580
rect 23940 -630 23960 -600
rect 23990 -630 24010 -600
rect 23940 -650 24010 -630
rect 23940 -680 23960 -650
rect 23990 -680 24010 -650
rect 23940 -690 24010 -680
rect 24025 -500 24095 -490
rect 24025 -530 24045 -500
rect 24075 -530 24095 -500
rect 24025 -550 24095 -530
rect 24025 -580 24045 -550
rect 24075 -580 24095 -550
rect 24025 -600 24095 -580
rect 24025 -630 24045 -600
rect 24075 -630 24095 -600
rect 24025 -650 24095 -630
rect 24025 -680 24045 -650
rect 24075 -680 24095 -650
rect 24025 -690 24095 -680
rect 24110 -500 24180 -490
rect 24110 -530 24130 -500
rect 24160 -530 24180 -500
rect 24110 -550 24180 -530
rect 24110 -580 24130 -550
rect 24160 -580 24180 -550
rect 24110 -600 24180 -580
rect 24110 -630 24130 -600
rect 24160 -630 24180 -600
rect 24110 -650 24180 -630
rect 24110 -680 24130 -650
rect 24160 -680 24180 -650
rect 24110 -690 24180 -680
rect 24195 -500 24265 -490
rect 24195 -530 24215 -500
rect 24245 -530 24265 -500
rect 24195 -550 24265 -530
rect 24195 -580 24215 -550
rect 24245 -580 24265 -550
rect 24195 -600 24265 -580
rect 24195 -630 24215 -600
rect 24245 -630 24265 -600
rect 24195 -650 24265 -630
rect 24195 -680 24215 -650
rect 24245 -680 24265 -650
rect 24195 -690 24265 -680
rect 24280 -500 24350 -490
rect 24280 -530 24300 -500
rect 24330 -530 24350 -500
rect 24280 -550 24350 -530
rect 24280 -580 24300 -550
rect 24330 -580 24350 -550
rect 24280 -600 24350 -580
rect 24280 -630 24300 -600
rect 24330 -630 24350 -600
rect 24280 -650 24350 -630
rect 24280 -680 24300 -650
rect 24330 -680 24350 -650
rect 24280 -690 24350 -680
rect 24365 -500 24435 -490
rect 24365 -530 24385 -500
rect 24415 -530 24435 -500
rect 24365 -550 24435 -530
rect 24365 -580 24385 -550
rect 24415 -580 24435 -550
rect 24365 -600 24435 -580
rect 24365 -630 24385 -600
rect 24415 -630 24435 -600
rect 24365 -650 24435 -630
rect 24365 -680 24385 -650
rect 24415 -680 24435 -650
rect 24365 -690 24435 -680
rect 24450 -500 24520 -490
rect 24450 -530 24470 -500
rect 24500 -530 24520 -500
rect 24450 -550 24520 -530
rect 24450 -580 24470 -550
rect 24500 -580 24520 -550
rect 24450 -600 24520 -580
rect 24450 -630 24470 -600
rect 24500 -630 24520 -600
rect 24450 -650 24520 -630
rect 24450 -680 24470 -650
rect 24500 -680 24520 -650
rect 24450 -690 24520 -680
rect 24535 -500 24605 -490
rect 24535 -530 24555 -500
rect 24585 -530 24605 -500
rect 24535 -550 24605 -530
rect 24535 -580 24555 -550
rect 24585 -580 24605 -550
rect 24535 -600 24605 -580
rect 24535 -630 24555 -600
rect 24585 -630 24605 -600
rect 24535 -650 24605 -630
rect 24535 -680 24555 -650
rect 24585 -680 24605 -650
rect 24535 -690 24605 -680
rect 24620 -500 24690 -490
rect 24620 -530 24640 -500
rect 24670 -530 24690 -500
rect 24620 -550 24690 -530
rect 24620 -580 24640 -550
rect 24670 -580 24690 -550
rect 24620 -600 24690 -580
rect 24620 -630 24640 -600
rect 24670 -630 24690 -600
rect 24620 -650 24690 -630
rect 24620 -680 24640 -650
rect 24670 -680 24690 -650
rect 24620 -690 24690 -680
rect 24705 -500 24775 -490
rect 24705 -530 24725 -500
rect 24755 -530 24775 -500
rect 24705 -550 24775 -530
rect 24705 -580 24725 -550
rect 24755 -580 24775 -550
rect 24705 -600 24775 -580
rect 24705 -630 24725 -600
rect 24755 -630 24775 -600
rect 24705 -650 24775 -630
rect 24705 -680 24725 -650
rect 24755 -680 24775 -650
rect 24705 -690 24775 -680
rect 24790 -500 24860 -490
rect 24790 -530 24810 -500
rect 24840 -530 24860 -500
rect 24790 -550 24860 -530
rect 24790 -580 24810 -550
rect 24840 -580 24860 -550
rect 24790 -600 24860 -580
rect 24790 -630 24810 -600
rect 24840 -630 24860 -600
rect 24790 -650 24860 -630
rect 24790 -680 24810 -650
rect 24840 -680 24860 -650
rect 24790 -690 24860 -680
rect 24875 -500 24945 -490
rect 24875 -530 24895 -500
rect 24925 -530 24945 -500
rect 24875 -550 24945 -530
rect 24875 -580 24895 -550
rect 24925 -580 24945 -550
rect 24875 -600 24945 -580
rect 24875 -630 24895 -600
rect 24925 -630 24945 -600
rect 24875 -650 24945 -630
rect 24875 -680 24895 -650
rect 24925 -680 24945 -650
rect 24875 -690 24945 -680
rect 24960 -500 25030 -490
rect 24960 -530 24980 -500
rect 25010 -530 25030 -500
rect 24960 -550 25030 -530
rect 24960 -580 24980 -550
rect 25010 -580 25030 -550
rect 24960 -600 25030 -580
rect 24960 -630 24980 -600
rect 25010 -630 25030 -600
rect 24960 -650 25030 -630
rect 24960 -680 24980 -650
rect 25010 -680 25030 -650
rect 24960 -690 25030 -680
rect 25045 -500 25115 -490
rect 25045 -530 25065 -500
rect 25095 -530 25115 -500
rect 25045 -550 25115 -530
rect 25045 -580 25065 -550
rect 25095 -580 25115 -550
rect 25045 -600 25115 -580
rect 25045 -630 25065 -600
rect 25095 -630 25115 -600
rect 25045 -650 25115 -630
rect 25045 -680 25065 -650
rect 25095 -680 25115 -650
rect 25045 -690 25115 -680
rect 25130 -500 25200 -490
rect 25130 -530 25150 -500
rect 25180 -530 25200 -500
rect 25130 -550 25200 -530
rect 25130 -580 25150 -550
rect 25180 -580 25200 -550
rect 25130 -600 25200 -580
rect 25130 -630 25150 -600
rect 25180 -630 25200 -600
rect 25130 -650 25200 -630
rect 25130 -680 25150 -650
rect 25180 -680 25200 -650
rect 25130 -690 25200 -680
rect 25215 -500 25285 -490
rect 25215 -530 25235 -500
rect 25265 -530 25285 -500
rect 25215 -550 25285 -530
rect 25215 -580 25235 -550
rect 25265 -580 25285 -550
rect 25215 -600 25285 -580
rect 25215 -630 25235 -600
rect 25265 -630 25285 -600
rect 25215 -650 25285 -630
rect 25215 -680 25235 -650
rect 25265 -680 25285 -650
rect 25215 -690 25285 -680
rect 25300 -500 25370 -490
rect 25300 -530 25320 -500
rect 25350 -530 25370 -500
rect 25300 -550 25370 -530
rect 25300 -580 25320 -550
rect 25350 -580 25370 -550
rect 25300 -600 25370 -580
rect 25300 -630 25320 -600
rect 25350 -630 25370 -600
rect 25300 -650 25370 -630
rect 25300 -680 25320 -650
rect 25350 -680 25370 -650
rect 25300 -690 25370 -680
rect 25385 -500 25455 -490
rect 25385 -530 25405 -500
rect 25435 -530 25455 -500
rect 25385 -550 25455 -530
rect 25385 -580 25405 -550
rect 25435 -580 25455 -550
rect 25385 -600 25455 -580
rect 25385 -630 25405 -600
rect 25435 -630 25455 -600
rect 25385 -650 25455 -630
rect 25385 -680 25405 -650
rect 25435 -680 25455 -650
rect 25385 -690 25455 -680
rect 25470 -500 25540 -490
rect 25470 -530 25490 -500
rect 25520 -530 25540 -500
rect 25470 -550 25540 -530
rect 25470 -580 25490 -550
rect 25520 -580 25540 -550
rect 25470 -600 25540 -580
rect 25470 -630 25490 -600
rect 25520 -630 25540 -600
rect 25470 -650 25540 -630
rect 25470 -680 25490 -650
rect 25520 -680 25540 -650
rect 25470 -690 25540 -680
rect 25555 -500 25625 -490
rect 25555 -530 25575 -500
rect 25605 -530 25625 -500
rect 25555 -550 25625 -530
rect 25555 -580 25575 -550
rect 25605 -580 25625 -550
rect 25555 -600 25625 -580
rect 25555 -630 25575 -600
rect 25605 -630 25625 -600
rect 25555 -650 25625 -630
rect 25555 -680 25575 -650
rect 25605 -680 25625 -650
rect 25555 -690 25625 -680
rect 25640 -500 25710 -490
rect 25640 -530 25660 -500
rect 25690 -530 25710 -500
rect 25640 -550 25710 -530
rect 25640 -580 25660 -550
rect 25690 -580 25710 -550
rect 25640 -600 25710 -580
rect 25640 -630 25660 -600
rect 25690 -630 25710 -600
rect 25640 -650 25710 -630
rect 25640 -680 25660 -650
rect 25690 -680 25710 -650
rect 25640 -690 25710 -680
rect 25725 -500 25795 -490
rect 25725 -530 25745 -500
rect 25775 -530 25795 -500
rect 25725 -550 25795 -530
rect 25725 -580 25745 -550
rect 25775 -580 25795 -550
rect 25725 -600 25795 -580
rect 25725 -630 25745 -600
rect 25775 -630 25795 -600
rect 25725 -650 25795 -630
rect 25725 -680 25745 -650
rect 25775 -680 25795 -650
rect 25725 -690 25795 -680
rect 25810 -500 25880 -490
rect 25810 -530 25830 -500
rect 25860 -530 25880 -500
rect 25810 -550 25880 -530
rect 25810 -580 25830 -550
rect 25860 -580 25880 -550
rect 25810 -600 25880 -580
rect 25810 -630 25830 -600
rect 25860 -630 25880 -600
rect 25810 -650 25880 -630
rect 25810 -680 25830 -650
rect 25860 -680 25880 -650
rect 25810 -690 25880 -680
rect 25895 -500 25965 -490
rect 25895 -530 25915 -500
rect 25945 -530 25965 -500
rect 25895 -550 25965 -530
rect 25895 -580 25915 -550
rect 25945 -580 25965 -550
rect 25895 -600 25965 -580
rect 25895 -630 25915 -600
rect 25945 -630 25965 -600
rect 25895 -650 25965 -630
rect 25895 -680 25915 -650
rect 25945 -680 25965 -650
rect 25895 -690 25965 -680
rect 25980 -500 26050 -490
rect 25980 -530 26000 -500
rect 26030 -530 26050 -500
rect 25980 -550 26050 -530
rect 25980 -580 26000 -550
rect 26030 -580 26050 -550
rect 25980 -600 26050 -580
rect 25980 -630 26000 -600
rect 26030 -630 26050 -600
rect 25980 -650 26050 -630
rect 25980 -680 26000 -650
rect 26030 -680 26050 -650
rect 25980 -690 26050 -680
rect 26065 -500 26135 -490
rect 26065 -530 26085 -500
rect 26115 -530 26135 -500
rect 26065 -550 26135 -530
rect 26065 -580 26085 -550
rect 26115 -580 26135 -550
rect 26065 -600 26135 -580
rect 26065 -630 26085 -600
rect 26115 -630 26135 -600
rect 26065 -650 26135 -630
rect 26065 -680 26085 -650
rect 26115 -680 26135 -650
rect 26065 -690 26135 -680
rect 26150 -500 26220 -490
rect 26150 -530 26170 -500
rect 26200 -530 26220 -500
rect 26150 -550 26220 -530
rect 26150 -580 26170 -550
rect 26200 -580 26220 -550
rect 26150 -600 26220 -580
rect 26150 -630 26170 -600
rect 26200 -630 26220 -600
rect 26150 -650 26220 -630
rect 26150 -680 26170 -650
rect 26200 -680 26220 -650
rect 26150 -690 26220 -680
rect 26235 -500 26305 -490
rect 26235 -530 26255 -500
rect 26285 -530 26305 -500
rect 26235 -550 26305 -530
rect 26235 -580 26255 -550
rect 26285 -580 26305 -550
rect 26235 -600 26305 -580
rect 26235 -630 26255 -600
rect 26285 -630 26305 -600
rect 26235 -650 26305 -630
rect 26235 -680 26255 -650
rect 26285 -680 26305 -650
rect 26235 -690 26305 -680
rect 26320 -500 26390 -490
rect 26320 -530 26340 -500
rect 26370 -530 26390 -500
rect 26320 -550 26390 -530
rect 26320 -580 26340 -550
rect 26370 -580 26390 -550
rect 26320 -600 26390 -580
rect 26320 -630 26340 -600
rect 26370 -630 26390 -600
rect 26320 -650 26390 -630
rect 26320 -680 26340 -650
rect 26370 -680 26390 -650
rect 26320 -690 26390 -680
rect 26405 -500 26475 -490
rect 26405 -530 26425 -500
rect 26455 -530 26475 -500
rect 26405 -550 26475 -530
rect 26405 -580 26425 -550
rect 26455 -580 26475 -550
rect 26405 -600 26475 -580
rect 26405 -630 26425 -600
rect 26455 -630 26475 -600
rect 26405 -650 26475 -630
rect 26405 -680 26425 -650
rect 26455 -680 26475 -650
rect 26405 -690 26475 -680
rect 26490 -500 26560 -490
rect 26490 -530 26510 -500
rect 26540 -530 26560 -500
rect 26490 -550 26560 -530
rect 26490 -580 26510 -550
rect 26540 -580 26560 -550
rect 26490 -600 26560 -580
rect 26490 -630 26510 -600
rect 26540 -630 26560 -600
rect 26490 -650 26560 -630
rect 26490 -680 26510 -650
rect 26540 -680 26560 -650
rect 26490 -690 26560 -680
rect 26575 -500 26645 -490
rect 26575 -530 26595 -500
rect 26625 -530 26645 -500
rect 26575 -550 26645 -530
rect 26575 -580 26595 -550
rect 26625 -580 26645 -550
rect 26575 -600 26645 -580
rect 26575 -630 26595 -600
rect 26625 -630 26645 -600
rect 26575 -650 26645 -630
rect 26575 -680 26595 -650
rect 26625 -680 26645 -650
rect 26575 -690 26645 -680
rect 26660 -500 26730 -490
rect 26660 -530 26680 -500
rect 26710 -530 26730 -500
rect 26660 -550 26730 -530
rect 26660 -580 26680 -550
rect 26710 -580 26730 -550
rect 26660 -600 26730 -580
rect 26660 -630 26680 -600
rect 26710 -630 26730 -600
rect 26660 -650 26730 -630
rect 26660 -680 26680 -650
rect 26710 -680 26730 -650
rect 26660 -690 26730 -680
rect 26745 -500 26815 -490
rect 26745 -530 26765 -500
rect 26795 -530 26815 -500
rect 26745 -550 26815 -530
rect 26745 -580 26765 -550
rect 26795 -580 26815 -550
rect 26745 -600 26815 -580
rect 26745 -630 26765 -600
rect 26795 -630 26815 -600
rect 26745 -650 26815 -630
rect 26745 -680 26765 -650
rect 26795 -680 26815 -650
rect 26745 -690 26815 -680
rect 26830 -500 26900 -490
rect 26830 -530 26850 -500
rect 26880 -530 26900 -500
rect 26830 -550 26900 -530
rect 26830 -580 26850 -550
rect 26880 -580 26900 -550
rect 26830 -600 26900 -580
rect 26830 -630 26850 -600
rect 26880 -630 26900 -600
rect 26830 -650 26900 -630
rect 26830 -680 26850 -650
rect 26880 -680 26900 -650
rect 26830 -690 26900 -680
rect 26915 -500 26985 -490
rect 26915 -530 26935 -500
rect 26965 -530 26985 -500
rect 26915 -550 26985 -530
rect 26915 -580 26935 -550
rect 26965 -580 26985 -550
rect 26915 -600 26985 -580
rect 26915 -630 26935 -600
rect 26965 -630 26985 -600
rect 26915 -650 26985 -630
rect 26915 -680 26935 -650
rect 26965 -680 26985 -650
rect 26915 -690 26985 -680
rect 27000 -500 27070 -490
rect 27000 -530 27020 -500
rect 27050 -530 27070 -500
rect 27000 -550 27070 -530
rect 27000 -580 27020 -550
rect 27050 -580 27070 -550
rect 27000 -600 27070 -580
rect 27000 -630 27020 -600
rect 27050 -630 27070 -600
rect 27000 -650 27070 -630
rect 27000 -680 27020 -650
rect 27050 -680 27070 -650
rect 27000 -690 27070 -680
rect 27085 -500 27155 -490
rect 27085 -530 27105 -500
rect 27135 -530 27155 -500
rect 27085 -550 27155 -530
rect 27085 -580 27105 -550
rect 27135 -580 27155 -550
rect 27085 -600 27155 -580
rect 27085 -630 27105 -600
rect 27135 -630 27155 -600
rect 27085 -650 27155 -630
rect 27085 -680 27105 -650
rect 27135 -680 27155 -650
rect 27085 -690 27155 -680
rect 27170 -500 27240 -490
rect 27170 -530 27190 -500
rect 27220 -530 27240 -500
rect 27170 -550 27240 -530
rect 27170 -580 27190 -550
rect 27220 -580 27240 -550
rect 27170 -600 27240 -580
rect 27170 -630 27190 -600
rect 27220 -630 27240 -600
rect 27170 -650 27240 -630
rect 27170 -680 27190 -650
rect 27220 -680 27240 -650
rect 27170 -690 27240 -680
rect 27255 -500 27325 -490
rect 27255 -530 27275 -500
rect 27305 -530 27325 -500
rect 27255 -550 27325 -530
rect 27255 -580 27275 -550
rect 27305 -580 27325 -550
rect 27255 -600 27325 -580
rect 27255 -630 27275 -600
rect 27305 -630 27325 -600
rect 27255 -650 27325 -630
rect 27255 -680 27275 -650
rect 27305 -680 27325 -650
rect 27255 -690 27325 -680
rect 27340 -500 27410 -490
rect 27340 -530 27360 -500
rect 27390 -530 27410 -500
rect 27340 -550 27410 -530
rect 27340 -580 27360 -550
rect 27390 -580 27410 -550
rect 27340 -600 27410 -580
rect 27340 -630 27360 -600
rect 27390 -630 27410 -600
rect 27340 -650 27410 -630
rect 27340 -680 27360 -650
rect 27390 -680 27410 -650
rect 27340 -690 27410 -680
rect 27425 -500 27495 -490
rect 27425 -530 27445 -500
rect 27475 -530 27495 -500
rect 27425 -550 27495 -530
rect 27425 -580 27445 -550
rect 27475 -580 27495 -550
rect 27425 -600 27495 -580
rect 27425 -630 27445 -600
rect 27475 -630 27495 -600
rect 27425 -650 27495 -630
rect 27425 -680 27445 -650
rect 27475 -680 27495 -650
rect 27425 -690 27495 -680
rect 27510 -500 27580 -490
rect 27510 -530 27530 -500
rect 27560 -530 27580 -500
rect 27510 -550 27580 -530
rect 27510 -580 27530 -550
rect 27560 -580 27580 -550
rect 27510 -600 27580 -580
rect 27510 -630 27530 -600
rect 27560 -630 27580 -600
rect 27510 -650 27580 -630
rect 27510 -680 27530 -650
rect 27560 -680 27580 -650
rect 27510 -690 27580 -680
rect 27595 -500 27665 -490
rect 27595 -530 27615 -500
rect 27645 -530 27665 -500
rect 27595 -550 27665 -530
rect 27595 -580 27615 -550
rect 27645 -580 27665 -550
rect 27595 -600 27665 -580
rect 27595 -630 27615 -600
rect 27645 -630 27665 -600
rect 27595 -650 27665 -630
rect 27595 -680 27615 -650
rect 27645 -680 27665 -650
rect 27595 -690 27665 -680
rect 27680 -500 27750 -490
rect 27680 -530 27700 -500
rect 27730 -530 27750 -500
rect 27680 -550 27750 -530
rect 27680 -580 27700 -550
rect 27730 -580 27750 -550
rect 27680 -600 27750 -580
rect 27680 -630 27700 -600
rect 27730 -630 27750 -600
rect 27680 -650 27750 -630
rect 27680 -680 27700 -650
rect 27730 -680 27750 -650
rect 27680 -690 27750 -680
rect 27765 -500 27835 -490
rect 27765 -530 27785 -500
rect 27815 -530 27835 -500
rect 27765 -550 27835 -530
rect 27765 -580 27785 -550
rect 27815 -580 27835 -550
rect 27765 -600 27835 -580
rect 27765 -630 27785 -600
rect 27815 -630 27835 -600
rect 27765 -650 27835 -630
rect 27765 -680 27785 -650
rect 27815 -680 27835 -650
rect 27765 -690 27835 -680
rect 27850 -500 27920 -490
rect 27850 -530 27870 -500
rect 27900 -530 27920 -500
rect 27850 -550 27920 -530
rect 27850 -580 27870 -550
rect 27900 -580 27920 -550
rect 27850 -600 27920 -580
rect 27850 -630 27870 -600
rect 27900 -630 27920 -600
rect 27850 -650 27920 -630
rect 27850 -680 27870 -650
rect 27900 -680 27920 -650
rect 27850 -690 27920 -680
rect 27935 -500 28005 -490
rect 27935 -530 27955 -500
rect 27985 -530 28005 -500
rect 27935 -550 28005 -530
rect 27935 -580 27955 -550
rect 27985 -580 28005 -550
rect 27935 -600 28005 -580
rect 27935 -630 27955 -600
rect 27985 -630 28005 -600
rect 27935 -650 28005 -630
rect 27935 -680 27955 -650
rect 27985 -680 28005 -650
rect 27935 -690 28005 -680
rect 28020 -500 28090 -490
rect 28020 -530 28040 -500
rect 28070 -530 28090 -500
rect 28020 -550 28090 -530
rect 28020 -580 28040 -550
rect 28070 -580 28090 -550
rect 28020 -600 28090 -580
rect 28020 -630 28040 -600
rect 28070 -630 28090 -600
rect 28020 -650 28090 -630
rect 28020 -680 28040 -650
rect 28070 -680 28090 -650
rect 28020 -690 28090 -680
rect 28105 -500 28175 -490
rect 28105 -530 28125 -500
rect 28155 -530 28175 -500
rect 28105 -550 28175 -530
rect 28105 -580 28125 -550
rect 28155 -580 28175 -550
rect 28105 -600 28175 -580
rect 28105 -630 28125 -600
rect 28155 -630 28175 -600
rect 28105 -650 28175 -630
rect 28105 -680 28125 -650
rect 28155 -680 28175 -650
rect 28105 -690 28175 -680
rect 28190 -500 28260 -490
rect 28190 -530 28210 -500
rect 28240 -530 28260 -500
rect 28190 -550 28260 -530
rect 28190 -580 28210 -550
rect 28240 -580 28260 -550
rect 28190 -600 28260 -580
rect 28190 -630 28210 -600
rect 28240 -630 28260 -600
rect 28190 -650 28260 -630
rect 28190 -680 28210 -650
rect 28240 -680 28260 -650
rect 28190 -690 28260 -680
rect 28275 -500 28345 -490
rect 28275 -530 28295 -500
rect 28325 -530 28345 -500
rect 28275 -550 28345 -530
rect 28275 -580 28295 -550
rect 28325 -580 28345 -550
rect 28275 -600 28345 -580
rect 28275 -630 28295 -600
rect 28325 -630 28345 -600
rect 28275 -650 28345 -630
rect 28275 -680 28295 -650
rect 28325 -680 28345 -650
rect 28275 -690 28345 -680
rect 28360 -500 28430 -490
rect 28360 -530 28380 -500
rect 28410 -530 28430 -500
rect 28360 -550 28430 -530
rect 28360 -580 28380 -550
rect 28410 -580 28430 -550
rect 28360 -600 28430 -580
rect 28360 -630 28380 -600
rect 28410 -630 28430 -600
rect 28360 -650 28430 -630
rect 28360 -680 28380 -650
rect 28410 -680 28430 -650
rect 28360 -690 28430 -680
rect 28445 -500 28515 -490
rect 28445 -530 28465 -500
rect 28495 -530 28515 -500
rect 28445 -550 28515 -530
rect 28445 -580 28465 -550
rect 28495 -580 28515 -550
rect 28445 -600 28515 -580
rect 28445 -630 28465 -600
rect 28495 -630 28515 -600
rect 28445 -650 28515 -630
rect 28445 -680 28465 -650
rect 28495 -680 28515 -650
rect 28445 -690 28515 -680
rect 28530 -500 28600 -490
rect 28530 -530 28550 -500
rect 28580 -530 28600 -500
rect 28530 -550 28600 -530
rect 28530 -580 28550 -550
rect 28580 -580 28600 -550
rect 28530 -600 28600 -580
rect 28530 -630 28550 -600
rect 28580 -630 28600 -600
rect 28530 -650 28600 -630
rect 28530 -680 28550 -650
rect 28580 -680 28600 -650
rect 28530 -690 28600 -680
rect 28615 -500 28685 -490
rect 28615 -530 28635 -500
rect 28665 -530 28685 -500
rect 28615 -550 28685 -530
rect 28615 -580 28635 -550
rect 28665 -580 28685 -550
rect 28615 -600 28685 -580
rect 28615 -630 28635 -600
rect 28665 -630 28685 -600
rect 28615 -650 28685 -630
rect 28615 -680 28635 -650
rect 28665 -680 28685 -650
rect 28615 -690 28685 -680
rect 28700 -500 28770 -490
rect 28700 -530 28720 -500
rect 28750 -530 28770 -500
rect 28700 -550 28770 -530
rect 28700 -580 28720 -550
rect 28750 -580 28770 -550
rect 28700 -600 28770 -580
rect 28700 -630 28720 -600
rect 28750 -630 28770 -600
rect 28700 -650 28770 -630
rect 28700 -680 28720 -650
rect 28750 -680 28770 -650
rect 28700 -690 28770 -680
rect 28785 -500 28855 -490
rect 28785 -530 28805 -500
rect 28835 -530 28855 -500
rect 28785 -550 28855 -530
rect 28785 -580 28805 -550
rect 28835 -580 28855 -550
rect 28785 -600 28855 -580
rect 28785 -630 28805 -600
rect 28835 -630 28855 -600
rect 28785 -650 28855 -630
rect 28785 -680 28805 -650
rect 28835 -680 28855 -650
rect 28785 -690 28855 -680
rect 28870 -500 28940 -490
rect 28870 -530 28890 -500
rect 28920 -530 28940 -500
rect 28870 -550 28940 -530
rect 28870 -580 28890 -550
rect 28920 -580 28940 -550
rect 28870 -600 28940 -580
rect 28870 -630 28890 -600
rect 28920 -630 28940 -600
rect 28870 -650 28940 -630
rect 28870 -680 28890 -650
rect 28920 -680 28940 -650
rect 28870 -690 28940 -680
rect 28955 -500 29025 -490
rect 28955 -530 28975 -500
rect 29005 -530 29025 -500
rect 28955 -550 29025 -530
rect 28955 -580 28975 -550
rect 29005 -580 29025 -550
rect 28955 -600 29025 -580
rect 28955 -630 28975 -600
rect 29005 -630 29025 -600
rect 28955 -650 29025 -630
rect 28955 -680 28975 -650
rect 29005 -680 29025 -650
rect 28955 -690 29025 -680
rect 29040 -500 29110 -490
rect 29040 -530 29060 -500
rect 29090 -530 29110 -500
rect 29040 -550 29110 -530
rect 29040 -580 29060 -550
rect 29090 -580 29110 -550
rect 29040 -600 29110 -580
rect 29040 -630 29060 -600
rect 29090 -630 29110 -600
rect 29040 -650 29110 -630
rect 29040 -680 29060 -650
rect 29090 -680 29110 -650
rect 29040 -690 29110 -680
rect 29125 -500 29195 -490
rect 29125 -530 29145 -500
rect 29175 -530 29195 -500
rect 29125 -550 29195 -530
rect 29125 -580 29145 -550
rect 29175 -580 29195 -550
rect 29125 -600 29195 -580
rect 29125 -630 29145 -600
rect 29175 -630 29195 -600
rect 29125 -650 29195 -630
rect 29125 -680 29145 -650
rect 29175 -680 29195 -650
rect 29125 -690 29195 -680
rect 29210 -500 29280 -490
rect 29210 -530 29230 -500
rect 29260 -530 29280 -500
rect 29210 -550 29280 -530
rect 29210 -580 29230 -550
rect 29260 -580 29280 -550
rect 29210 -600 29280 -580
rect 29210 -630 29230 -600
rect 29260 -630 29280 -600
rect 29210 -650 29280 -630
rect 29210 -680 29230 -650
rect 29260 -680 29280 -650
rect 29210 -690 29280 -680
rect 29295 -500 29365 -490
rect 29295 -530 29315 -500
rect 29345 -530 29365 -500
rect 29295 -550 29365 -530
rect 29295 -580 29315 -550
rect 29345 -580 29365 -550
rect 29295 -600 29365 -580
rect 29295 -630 29315 -600
rect 29345 -630 29365 -600
rect 29295 -650 29365 -630
rect 29295 -680 29315 -650
rect 29345 -680 29365 -650
rect 29295 -690 29365 -680
rect 29380 -500 29450 -490
rect 29380 -530 29400 -500
rect 29430 -530 29450 -500
rect 29380 -550 29450 -530
rect 29380 -580 29400 -550
rect 29430 -580 29450 -550
rect 29380 -600 29450 -580
rect 29380 -630 29400 -600
rect 29430 -630 29450 -600
rect 29380 -650 29450 -630
rect 29380 -680 29400 -650
rect 29430 -680 29450 -650
rect 29380 -690 29450 -680
rect 29465 -500 29535 -490
rect 29465 -530 29485 -500
rect 29515 -530 29535 -500
rect 29465 -550 29535 -530
rect 29465 -580 29485 -550
rect 29515 -580 29535 -550
rect 29465 -600 29535 -580
rect 29465 -630 29485 -600
rect 29515 -630 29535 -600
rect 29465 -650 29535 -630
rect 29465 -680 29485 -650
rect 29515 -680 29535 -650
rect 29465 -690 29535 -680
rect 29550 -500 29620 -490
rect 29550 -530 29570 -500
rect 29600 -530 29620 -500
rect 29550 -550 29620 -530
rect 29550 -580 29570 -550
rect 29600 -580 29620 -550
rect 29550 -600 29620 -580
rect 29550 -630 29570 -600
rect 29600 -630 29620 -600
rect 29550 -650 29620 -630
rect 29550 -680 29570 -650
rect 29600 -680 29620 -650
rect 29550 -690 29620 -680
rect 29635 -500 29705 -490
rect 29635 -530 29655 -500
rect 29685 -530 29705 -500
rect 29635 -550 29705 -530
rect 29635 -580 29655 -550
rect 29685 -580 29705 -550
rect 29635 -600 29705 -580
rect 29635 -630 29655 -600
rect 29685 -630 29705 -600
rect 29635 -650 29705 -630
rect 29635 -680 29655 -650
rect 29685 -680 29705 -650
rect 29635 -690 29705 -680
rect 29720 -500 29790 -490
rect 29720 -530 29740 -500
rect 29770 -530 29790 -500
rect 29720 -550 29790 -530
rect 29720 -580 29740 -550
rect 29770 -580 29790 -550
rect 29720 -600 29790 -580
rect 29720 -630 29740 -600
rect 29770 -630 29790 -600
rect 29720 -650 29790 -630
rect 29720 -680 29740 -650
rect 29770 -680 29790 -650
rect 29720 -690 29790 -680
rect 29805 -500 29875 -490
rect 29805 -530 29825 -500
rect 29855 -530 29875 -500
rect 29805 -550 29875 -530
rect 29805 -580 29825 -550
rect 29855 -580 29875 -550
rect 29805 -600 29875 -580
rect 29805 -630 29825 -600
rect 29855 -630 29875 -600
rect 29805 -650 29875 -630
rect 29805 -680 29825 -650
rect 29855 -680 29875 -650
rect 29805 -690 29875 -680
rect 29890 -500 29960 -490
rect 29890 -530 29910 -500
rect 29940 -530 29960 -500
rect 29890 -550 29960 -530
rect 29890 -580 29910 -550
rect 29940 -580 29960 -550
rect 29890 -600 29960 -580
rect 29890 -630 29910 -600
rect 29940 -630 29960 -600
rect 29890 -650 29960 -630
rect 29890 -680 29910 -650
rect 29940 -680 29960 -650
rect 29890 -690 29960 -680
rect 29975 -500 30045 -490
rect 29975 -530 29995 -500
rect 30025 -530 30045 -500
rect 29975 -550 30045 -530
rect 29975 -580 29995 -550
rect 30025 -580 30045 -550
rect 29975 -600 30045 -580
rect 29975 -630 29995 -600
rect 30025 -630 30045 -600
rect 29975 -650 30045 -630
rect 29975 -680 29995 -650
rect 30025 -680 30045 -650
rect 29975 -690 30045 -680
rect 30060 -500 30130 -490
rect 30060 -530 30080 -500
rect 30110 -530 30130 -500
rect 30060 -550 30130 -530
rect 30060 -580 30080 -550
rect 30110 -580 30130 -550
rect 30060 -600 30130 -580
rect 30060 -630 30080 -600
rect 30110 -630 30130 -600
rect 30060 -650 30130 -630
rect 30060 -680 30080 -650
rect 30110 -680 30130 -650
rect 30060 -690 30130 -680
rect 30145 -500 30215 -490
rect 30145 -530 30165 -500
rect 30195 -530 30215 -500
rect 30145 -550 30215 -530
rect 30145 -580 30165 -550
rect 30195 -580 30215 -550
rect 30145 -600 30215 -580
rect 30145 -630 30165 -600
rect 30195 -630 30215 -600
rect 30145 -650 30215 -630
rect 30145 -680 30165 -650
rect 30195 -680 30215 -650
rect 30145 -690 30215 -680
rect 30230 -500 30300 -490
rect 30230 -530 30250 -500
rect 30280 -530 30300 -500
rect 30230 -550 30300 -530
rect 30230 -580 30250 -550
rect 30280 -580 30300 -550
rect 30230 -600 30300 -580
rect 30230 -630 30250 -600
rect 30280 -630 30300 -600
rect 30230 -650 30300 -630
rect 30230 -680 30250 -650
rect 30280 -680 30300 -650
rect 30230 -690 30300 -680
rect 30315 -500 30385 -490
rect 30315 -530 30335 -500
rect 30365 -530 30385 -500
rect 30315 -550 30385 -530
rect 30315 -580 30335 -550
rect 30365 -580 30385 -550
rect 30315 -600 30385 -580
rect 30315 -630 30335 -600
rect 30365 -630 30385 -600
rect 30315 -650 30385 -630
rect 30315 -680 30335 -650
rect 30365 -680 30385 -650
rect 30315 -690 30385 -680
rect 30400 -500 30470 -490
rect 30400 -530 30420 -500
rect 30450 -530 30470 -500
rect 30400 -550 30470 -530
rect 30400 -580 30420 -550
rect 30450 -580 30470 -550
rect 30400 -600 30470 -580
rect 30400 -630 30420 -600
rect 30450 -630 30470 -600
rect 30400 -650 30470 -630
rect 30400 -680 30420 -650
rect 30450 -680 30470 -650
rect 30400 -690 30470 -680
rect 30485 -500 30555 -490
rect 30485 -530 30505 -500
rect 30535 -530 30555 -500
rect 30485 -550 30555 -530
rect 30485 -580 30505 -550
rect 30535 -580 30555 -550
rect 30485 -600 30555 -580
rect 30485 -630 30505 -600
rect 30535 -630 30555 -600
rect 30485 -650 30555 -630
rect 30485 -680 30505 -650
rect 30535 -680 30555 -650
rect 30485 -690 30555 -680
rect 30570 -500 30640 -490
rect 30570 -530 30590 -500
rect 30620 -530 30640 -500
rect 30570 -550 30640 -530
rect 30570 -580 30590 -550
rect 30620 -580 30640 -550
rect 30570 -600 30640 -580
rect 30570 -630 30590 -600
rect 30620 -630 30640 -600
rect 30570 -650 30640 -630
rect 30570 -680 30590 -650
rect 30620 -680 30640 -650
rect 30570 -690 30640 -680
rect 30655 -500 30725 -490
rect 30655 -530 30675 -500
rect 30705 -530 30725 -500
rect 30655 -550 30725 -530
rect 30655 -580 30675 -550
rect 30705 -580 30725 -550
rect 30655 -600 30725 -580
rect 30655 -630 30675 -600
rect 30705 -630 30725 -600
rect 30655 -650 30725 -630
rect 30655 -680 30675 -650
rect 30705 -680 30725 -650
rect 30655 -690 30725 -680
rect 30740 -500 30810 -490
rect 30740 -530 30760 -500
rect 30790 -530 30810 -500
rect 30740 -550 30810 -530
rect 30740 -580 30760 -550
rect 30790 -580 30810 -550
rect 30740 -600 30810 -580
rect 30740 -630 30760 -600
rect 30790 -630 30810 -600
rect 30740 -650 30810 -630
rect 30740 -680 30760 -650
rect 30790 -680 30810 -650
rect 30740 -690 30810 -680
rect 30825 -500 30895 -490
rect 30825 -530 30845 -500
rect 30875 -530 30895 -500
rect 30825 -550 30895 -530
rect 30825 -580 30845 -550
rect 30875 -580 30895 -550
rect 30825 -600 30895 -580
rect 30825 -630 30845 -600
rect 30875 -630 30895 -600
rect 30825 -650 30895 -630
rect 30825 -680 30845 -650
rect 30875 -680 30895 -650
rect 30825 -690 30895 -680
rect 30910 -500 30980 -490
rect 30910 -530 30930 -500
rect 30960 -530 30980 -500
rect 30910 -550 30980 -530
rect 30910 -580 30930 -550
rect 30960 -580 30980 -550
rect 30910 -600 30980 -580
rect 30910 -630 30930 -600
rect 30960 -630 30980 -600
rect 30910 -650 30980 -630
rect 30910 -680 30930 -650
rect 30960 -680 30980 -650
rect 30910 -690 30980 -680
rect 30995 -500 31065 -490
rect 30995 -530 31015 -500
rect 31045 -530 31065 -500
rect 30995 -550 31065 -530
rect 30995 -580 31015 -550
rect 31045 -580 31065 -550
rect 30995 -600 31065 -580
rect 30995 -630 31015 -600
rect 31045 -630 31065 -600
rect 30995 -650 31065 -630
rect 30995 -680 31015 -650
rect 31045 -680 31065 -650
rect 30995 -690 31065 -680
rect 31080 -500 31150 -490
rect 31080 -530 31100 -500
rect 31130 -530 31150 -500
rect 31080 -550 31150 -530
rect 31080 -580 31100 -550
rect 31130 -580 31150 -550
rect 31080 -600 31150 -580
rect 31080 -630 31100 -600
rect 31130 -630 31150 -600
rect 31080 -650 31150 -630
rect 31080 -680 31100 -650
rect 31130 -680 31150 -650
rect 31080 -690 31150 -680
rect 31165 -500 31235 -490
rect 31165 -530 31185 -500
rect 31215 -530 31235 -500
rect 31165 -550 31235 -530
rect 31165 -580 31185 -550
rect 31215 -580 31235 -550
rect 31165 -600 31235 -580
rect 31165 -630 31185 -600
rect 31215 -630 31235 -600
rect 31165 -650 31235 -630
rect 31165 -680 31185 -650
rect 31215 -680 31235 -650
rect 31165 -690 31235 -680
rect 31250 -500 31320 -490
rect 31250 -530 31270 -500
rect 31300 -530 31320 -500
rect 31250 -550 31320 -530
rect 31250 -580 31270 -550
rect 31300 -580 31320 -550
rect 31250 -600 31320 -580
rect 31250 -630 31270 -600
rect 31300 -630 31320 -600
rect 31250 -650 31320 -630
rect 31250 -680 31270 -650
rect 31300 -680 31320 -650
rect 31250 -690 31320 -680
rect 31335 -500 31405 -490
rect 31335 -530 31355 -500
rect 31385 -530 31405 -500
rect 31335 -550 31405 -530
rect 31335 -580 31355 -550
rect 31385 -580 31405 -550
rect 31335 -600 31405 -580
rect 31335 -630 31355 -600
rect 31385 -630 31405 -600
rect 31335 -650 31405 -630
rect 31335 -680 31355 -650
rect 31385 -680 31405 -650
rect 31335 -690 31405 -680
rect 31420 -500 31490 -490
rect 31420 -530 31440 -500
rect 31470 -530 31490 -500
rect 31420 -550 31490 -530
rect 31420 -580 31440 -550
rect 31470 -580 31490 -550
rect 31420 -600 31490 -580
rect 31420 -630 31440 -600
rect 31470 -630 31490 -600
rect 31420 -650 31490 -630
rect 31420 -680 31440 -650
rect 31470 -680 31490 -650
rect 31420 -690 31490 -680
rect 31505 -500 31575 -490
rect 31505 -530 31525 -500
rect 31555 -530 31575 -500
rect 31505 -550 31575 -530
rect 31505 -580 31525 -550
rect 31555 -580 31575 -550
rect 31505 -600 31575 -580
rect 31505 -630 31525 -600
rect 31555 -630 31575 -600
rect 31505 -650 31575 -630
rect 31505 -680 31525 -650
rect 31555 -680 31575 -650
rect 31505 -690 31575 -680
rect 31590 -500 31660 -490
rect 31590 -530 31610 -500
rect 31640 -530 31660 -500
rect 31590 -550 31660 -530
rect 31590 -580 31610 -550
rect 31640 -580 31660 -550
rect 31590 -600 31660 -580
rect 31590 -630 31610 -600
rect 31640 -630 31660 -600
rect 31590 -650 31660 -630
rect 31590 -680 31610 -650
rect 31640 -680 31660 -650
rect 31590 -690 31660 -680
rect 31675 -500 31745 -490
rect 31675 -530 31695 -500
rect 31725 -530 31745 -500
rect 31675 -550 31745 -530
rect 31675 -580 31695 -550
rect 31725 -580 31745 -550
rect 31675 -600 31745 -580
rect 31675 -630 31695 -600
rect 31725 -630 31745 -600
rect 31675 -650 31745 -630
rect 31675 -680 31695 -650
rect 31725 -680 31745 -650
rect 31675 -690 31745 -680
rect 31760 -500 31830 -490
rect 31760 -530 31780 -500
rect 31810 -530 31830 -500
rect 31760 -550 31830 -530
rect 31760 -580 31780 -550
rect 31810 -580 31830 -550
rect 31760 -600 31830 -580
rect 31760 -630 31780 -600
rect 31810 -630 31830 -600
rect 31760 -650 31830 -630
rect 31760 -680 31780 -650
rect 31810 -680 31830 -650
rect 31760 -690 31830 -680
rect 31845 -500 31915 -490
rect 31845 -530 31865 -500
rect 31895 -530 31915 -500
rect 31845 -550 31915 -530
rect 31845 -580 31865 -550
rect 31895 -580 31915 -550
rect 31845 -600 31915 -580
rect 31845 -630 31865 -600
rect 31895 -630 31915 -600
rect 31845 -650 31915 -630
rect 31845 -680 31865 -650
rect 31895 -680 31915 -650
rect 31845 -690 31915 -680
rect 31930 -500 32000 -490
rect 31930 -530 31950 -500
rect 31980 -530 32000 -500
rect 31930 -550 32000 -530
rect 31930 -580 31950 -550
rect 31980 -580 32000 -550
rect 31930 -600 32000 -580
rect 31930 -630 31950 -600
rect 31980 -630 32000 -600
rect 31930 -650 32000 -630
rect 31930 -680 31950 -650
rect 31980 -680 32000 -650
rect 31930 -690 32000 -680
rect 32015 -500 32085 -490
rect 32015 -530 32035 -500
rect 32065 -530 32085 -500
rect 32015 -550 32085 -530
rect 32015 -580 32035 -550
rect 32065 -580 32085 -550
rect 32015 -600 32085 -580
rect 32015 -630 32035 -600
rect 32065 -630 32085 -600
rect 32015 -650 32085 -630
rect 32015 -680 32035 -650
rect 32065 -680 32085 -650
rect 32015 -690 32085 -680
rect 32100 -500 32170 -490
rect 32100 -530 32120 -500
rect 32150 -530 32170 -500
rect 32100 -550 32170 -530
rect 32100 -580 32120 -550
rect 32150 -580 32170 -550
rect 32100 -600 32170 -580
rect 32100 -630 32120 -600
rect 32150 -630 32170 -600
rect 32100 -650 32170 -630
rect 32100 -680 32120 -650
rect 32150 -680 32170 -650
rect 32100 -690 32170 -680
rect 32185 -500 32255 -490
rect 32185 -530 32205 -500
rect 32235 -530 32255 -500
rect 32185 -550 32255 -530
rect 32185 -580 32205 -550
rect 32235 -580 32255 -550
rect 32185 -600 32255 -580
rect 32185 -630 32205 -600
rect 32235 -630 32255 -600
rect 32185 -650 32255 -630
rect 32185 -680 32205 -650
rect 32235 -680 32255 -650
rect 32185 -690 32255 -680
rect 32270 -500 32340 -490
rect 32270 -530 32290 -500
rect 32320 -530 32340 -500
rect 32270 -550 32340 -530
rect 32270 -580 32290 -550
rect 32320 -580 32340 -550
rect 32270 -600 32340 -580
rect 32270 -630 32290 -600
rect 32320 -630 32340 -600
rect 32270 -650 32340 -630
rect 32270 -680 32290 -650
rect 32320 -680 32340 -650
rect 32270 -690 32340 -680
rect 32355 -500 32425 -490
rect 32355 -530 32375 -500
rect 32405 -530 32425 -500
rect 32355 -550 32425 -530
rect 32355 -580 32375 -550
rect 32405 -580 32425 -550
rect 32355 -600 32425 -580
rect 32355 -630 32375 -600
rect 32405 -630 32425 -600
rect 32355 -650 32425 -630
rect 32355 -680 32375 -650
rect 32405 -680 32425 -650
rect 32355 -690 32425 -680
rect 32440 -500 32510 -490
rect 32440 -530 32460 -500
rect 32490 -530 32510 -500
rect 32440 -550 32510 -530
rect 32440 -580 32460 -550
rect 32490 -580 32510 -550
rect 32440 -600 32510 -580
rect 32440 -630 32460 -600
rect 32490 -630 32510 -600
rect 32440 -650 32510 -630
rect 32440 -680 32460 -650
rect 32490 -680 32510 -650
rect 32440 -690 32510 -680
rect 32525 -500 32595 -490
rect 32525 -530 32545 -500
rect 32575 -530 32595 -500
rect 32525 -550 32595 -530
rect 32525 -580 32545 -550
rect 32575 -580 32595 -550
rect 32525 -600 32595 -580
rect 32525 -630 32545 -600
rect 32575 -630 32595 -600
rect 32525 -650 32595 -630
rect 32525 -680 32545 -650
rect 32575 -680 32595 -650
rect 32525 -690 32595 -680
rect 32610 -500 32680 -490
rect 32610 -530 32630 -500
rect 32660 -530 32680 -500
rect 32610 -550 32680 -530
rect 32610 -580 32630 -550
rect 32660 -580 32680 -550
rect 32610 -600 32680 -580
rect 32610 -630 32630 -600
rect 32660 -630 32680 -600
rect 32610 -650 32680 -630
rect 32610 -680 32630 -650
rect 32660 -680 32680 -650
rect 32610 -690 32680 -680
rect 32695 -500 32765 -490
rect 32695 -530 32715 -500
rect 32745 -530 32765 -500
rect 32695 -550 32765 -530
rect 32695 -580 32715 -550
rect 32745 -580 32765 -550
rect 32695 -600 32765 -580
rect 32695 -630 32715 -600
rect 32745 -630 32765 -600
rect 32695 -650 32765 -630
rect 32695 -680 32715 -650
rect 32745 -680 32765 -650
rect 32695 -690 32765 -680
rect 32780 -500 32850 -490
rect 32780 -530 32800 -500
rect 32830 -530 32850 -500
rect 32780 -550 32850 -530
rect 32780 -580 32800 -550
rect 32830 -580 32850 -550
rect 32780 -600 32850 -580
rect 32780 -630 32800 -600
rect 32830 -630 32850 -600
rect 32780 -650 32850 -630
rect 32780 -680 32800 -650
rect 32830 -680 32850 -650
rect 32780 -690 32850 -680
rect 32865 -500 32935 -490
rect 32865 -530 32885 -500
rect 32915 -530 32935 -500
rect 32865 -550 32935 -530
rect 32865 -580 32885 -550
rect 32915 -580 32935 -550
rect 32865 -600 32935 -580
rect 32865 -630 32885 -600
rect 32915 -630 32935 -600
rect 32865 -650 32935 -630
rect 32865 -680 32885 -650
rect 32915 -680 32935 -650
rect 32865 -690 32935 -680
rect 32950 -500 33020 -490
rect 32950 -530 32970 -500
rect 33000 -530 33020 -500
rect 32950 -550 33020 -530
rect 32950 -580 32970 -550
rect 33000 -580 33020 -550
rect 32950 -600 33020 -580
rect 32950 -630 32970 -600
rect 33000 -630 33020 -600
rect 32950 -650 33020 -630
rect 32950 -680 32970 -650
rect 33000 -680 33020 -650
rect 32950 -690 33020 -680
rect 33035 -500 33105 -490
rect 33035 -530 33055 -500
rect 33085 -530 33105 -500
rect 33035 -550 33105 -530
rect 33035 -580 33055 -550
rect 33085 -580 33105 -550
rect 33035 -600 33105 -580
rect 33035 -630 33055 -600
rect 33085 -630 33105 -600
rect 33035 -650 33105 -630
rect 33035 -680 33055 -650
rect 33085 -680 33105 -650
rect 33035 -690 33105 -680
rect 33120 -500 33190 -490
rect 33120 -530 33140 -500
rect 33170 -530 33190 -500
rect 33120 -550 33190 -530
rect 33120 -580 33140 -550
rect 33170 -580 33190 -550
rect 33120 -600 33190 -580
rect 33120 -630 33140 -600
rect 33170 -630 33190 -600
rect 33120 -650 33190 -630
rect 33120 -680 33140 -650
rect 33170 -680 33190 -650
rect 33120 -690 33190 -680
rect 33205 -500 33275 -490
rect 33205 -530 33225 -500
rect 33255 -530 33275 -500
rect 33205 -550 33275 -530
rect 33205 -580 33225 -550
rect 33255 -580 33275 -550
rect 33205 -600 33275 -580
rect 33205 -630 33225 -600
rect 33255 -630 33275 -600
rect 33205 -650 33275 -630
rect 33205 -680 33225 -650
rect 33255 -680 33275 -650
rect 33205 -690 33275 -680
rect 33290 -500 33360 -490
rect 33290 -530 33310 -500
rect 33340 -530 33360 -500
rect 33290 -550 33360 -530
rect 33290 -580 33310 -550
rect 33340 -580 33360 -550
rect 33290 -600 33360 -580
rect 33290 -630 33310 -600
rect 33340 -630 33360 -600
rect 33290 -650 33360 -630
rect 33290 -680 33310 -650
rect 33340 -680 33360 -650
rect 33290 -690 33360 -680
rect 33375 -500 33445 -490
rect 33375 -530 33395 -500
rect 33425 -530 33445 -500
rect 33375 -550 33445 -530
rect 33375 -580 33395 -550
rect 33425 -580 33445 -550
rect 33375 -600 33445 -580
rect 33375 -630 33395 -600
rect 33425 -630 33445 -600
rect 33375 -650 33445 -630
rect 33375 -680 33395 -650
rect 33425 -680 33445 -650
rect 33375 -690 33445 -680
rect 33460 -500 33530 -490
rect 33460 -530 33480 -500
rect 33510 -530 33530 -500
rect 33460 -550 33530 -530
rect 33460 -580 33480 -550
rect 33510 -580 33530 -550
rect 33460 -600 33530 -580
rect 33460 -630 33480 -600
rect 33510 -630 33530 -600
rect 33460 -650 33530 -630
rect 33460 -680 33480 -650
rect 33510 -680 33530 -650
rect 33460 -690 33530 -680
rect 33545 -500 33615 -490
rect 33545 -530 33565 -500
rect 33595 -530 33615 -500
rect 33545 -550 33615 -530
rect 33545 -580 33565 -550
rect 33595 -580 33615 -550
rect 33545 -600 33615 -580
rect 33545 -630 33565 -600
rect 33595 -630 33615 -600
rect 33545 -650 33615 -630
rect 33545 -680 33565 -650
rect 33595 -680 33615 -650
rect 33545 -690 33615 -680
rect 33630 -500 33700 -490
rect 33630 -530 33650 -500
rect 33680 -530 33700 -500
rect 33630 -550 33700 -530
rect 33630 -580 33650 -550
rect 33680 -580 33700 -550
rect 33630 -600 33700 -580
rect 33630 -630 33650 -600
rect 33680 -630 33700 -600
rect 33630 -650 33700 -630
rect 33630 -680 33650 -650
rect 33680 -680 33700 -650
rect 33630 -690 33700 -680
rect 33715 -500 33785 -490
rect 33715 -530 33735 -500
rect 33765 -530 33785 -500
rect 33715 -550 33785 -530
rect 33715 -580 33735 -550
rect 33765 -580 33785 -550
rect 33715 -600 33785 -580
rect 33715 -630 33735 -600
rect 33765 -630 33785 -600
rect 33715 -650 33785 -630
rect 33715 -680 33735 -650
rect 33765 -680 33785 -650
rect 33715 -690 33785 -680
rect 33800 -500 33870 -490
rect 33800 -530 33820 -500
rect 33850 -530 33870 -500
rect 33800 -550 33870 -530
rect 33800 -580 33820 -550
rect 33850 -580 33870 -550
rect 33800 -600 33870 -580
rect 33800 -630 33820 -600
rect 33850 -630 33870 -600
rect 33800 -650 33870 -630
rect 33800 -680 33820 -650
rect 33850 -680 33870 -650
rect 33800 -690 33870 -680
rect 33885 -500 33955 -490
rect 33885 -530 33905 -500
rect 33935 -530 33955 -500
rect 33885 -550 33955 -530
rect 33885 -580 33905 -550
rect 33935 -580 33955 -550
rect 33885 -600 33955 -580
rect 33885 -630 33905 -600
rect 33935 -630 33955 -600
rect 33885 -650 33955 -630
rect 33885 -680 33905 -650
rect 33935 -680 33955 -650
rect 33885 -690 33955 -680
rect 33970 -500 34040 -490
rect 33970 -530 33990 -500
rect 34020 -530 34040 -500
rect 33970 -550 34040 -530
rect 33970 -580 33990 -550
rect 34020 -580 34040 -550
rect 33970 -600 34040 -580
rect 33970 -630 33990 -600
rect 34020 -630 34040 -600
rect 33970 -650 34040 -630
rect 33970 -680 33990 -650
rect 34020 -680 34040 -650
rect 33970 -690 34040 -680
rect 34055 -500 34125 -490
rect 34055 -530 34075 -500
rect 34105 -530 34125 -500
rect 34055 -550 34125 -530
rect 34055 -580 34075 -550
rect 34105 -580 34125 -550
rect 34055 -600 34125 -580
rect 34055 -630 34075 -600
rect 34105 -630 34125 -600
rect 34055 -650 34125 -630
rect 34055 -680 34075 -650
rect 34105 -680 34125 -650
rect 34055 -690 34125 -680
rect 34140 -500 34210 -490
rect 34140 -530 34160 -500
rect 34190 -530 34210 -500
rect 34140 -550 34210 -530
rect 34140 -580 34160 -550
rect 34190 -580 34210 -550
rect 34140 -600 34210 -580
rect 34140 -630 34160 -600
rect 34190 -630 34210 -600
rect 34140 -650 34210 -630
rect 34140 -680 34160 -650
rect 34190 -680 34210 -650
rect 34140 -690 34210 -680
rect 34225 -500 34295 -490
rect 34225 -530 34245 -500
rect 34275 -530 34295 -500
rect 34225 -550 34295 -530
rect 34225 -580 34245 -550
rect 34275 -580 34295 -550
rect 34225 -600 34295 -580
rect 34225 -630 34245 -600
rect 34275 -630 34295 -600
rect 34225 -650 34295 -630
rect 34225 -680 34245 -650
rect 34275 -680 34295 -650
rect 34225 -690 34295 -680
rect 34310 -500 34380 -490
rect 34310 -530 34330 -500
rect 34360 -530 34380 -500
rect 34310 -550 34380 -530
rect 34310 -580 34330 -550
rect 34360 -580 34380 -550
rect 34310 -600 34380 -580
rect 34310 -630 34330 -600
rect 34360 -630 34380 -600
rect 34310 -650 34380 -630
rect 34310 -680 34330 -650
rect 34360 -680 34380 -650
rect 34310 -690 34380 -680
rect 34395 -500 34465 -490
rect 34395 -530 34415 -500
rect 34445 -530 34465 -500
rect 34395 -550 34465 -530
rect 34395 -580 34415 -550
rect 34445 -580 34465 -550
rect 34395 -600 34465 -580
rect 34395 -630 34415 -600
rect 34445 -630 34465 -600
rect 34395 -650 34465 -630
rect 34395 -680 34415 -650
rect 34445 -680 34465 -650
rect 34395 -690 34465 -680
rect 34480 -500 34550 -490
rect 34480 -530 34500 -500
rect 34530 -530 34550 -500
rect 34480 -550 34550 -530
rect 34480 -580 34500 -550
rect 34530 -580 34550 -550
rect 34480 -600 34550 -580
rect 34480 -630 34500 -600
rect 34530 -630 34550 -600
rect 34480 -650 34550 -630
rect 34480 -680 34500 -650
rect 34530 -680 34550 -650
rect 34480 -690 34550 -680
rect 34565 -500 34635 -490
rect 34565 -530 34585 -500
rect 34615 -530 34635 -500
rect 34565 -550 34635 -530
rect 34565 -580 34585 -550
rect 34615 -580 34635 -550
rect 34565 -600 34635 -580
rect 34565 -630 34585 -600
rect 34615 -630 34635 -600
rect 34565 -650 34635 -630
rect 34565 -680 34585 -650
rect 34615 -680 34635 -650
rect 34565 -690 34635 -680
rect 34650 -500 34720 -490
rect 34650 -530 34670 -500
rect 34700 -530 34720 -500
rect 34650 -550 34720 -530
rect 34650 -580 34670 -550
rect 34700 -580 34720 -550
rect 34650 -600 34720 -580
rect 34650 -630 34670 -600
rect 34700 -630 34720 -600
rect 34650 -650 34720 -630
rect 34650 -680 34670 -650
rect 34700 -680 34720 -650
rect 34650 -690 34720 -680
rect 34735 -500 34805 -490
rect 34735 -530 34755 -500
rect 34785 -530 34805 -500
rect 34735 -550 34805 -530
rect 34735 -580 34755 -550
rect 34785 -580 34805 -550
rect 34735 -600 34805 -580
rect 34735 -630 34755 -600
rect 34785 -630 34805 -600
rect 34735 -650 34805 -630
rect 34735 -680 34755 -650
rect 34785 -680 34805 -650
rect 34735 -690 34805 -680
rect 34820 -500 34890 -490
rect 34820 -530 34840 -500
rect 34870 -530 34890 -500
rect 34820 -550 34890 -530
rect 34820 -580 34840 -550
rect 34870 -580 34890 -550
rect 34820 -600 34890 -580
rect 34820 -630 34840 -600
rect 34870 -630 34890 -600
rect 34820 -650 34890 -630
rect 34820 -680 34840 -650
rect 34870 -680 34890 -650
rect 34820 -690 34890 -680
rect 34905 -500 34975 -490
rect 34905 -530 34925 -500
rect 34955 -530 34975 -500
rect 34905 -550 34975 -530
rect 34905 -580 34925 -550
rect 34955 -580 34975 -550
rect 34905 -600 34975 -580
rect 34905 -630 34925 -600
rect 34955 -630 34975 -600
rect 34905 -650 34975 -630
rect 34905 -680 34925 -650
rect 34955 -680 34975 -650
rect 34905 -690 34975 -680
rect 34990 -500 35060 -490
rect 34990 -530 35010 -500
rect 35040 -530 35060 -500
rect 34990 -550 35060 -530
rect 34990 -580 35010 -550
rect 35040 -580 35060 -550
rect 34990 -600 35060 -580
rect 34990 -630 35010 -600
rect 35040 -630 35060 -600
rect 34990 -650 35060 -630
rect 34990 -680 35010 -650
rect 35040 -680 35060 -650
rect 34990 -690 35060 -680
rect 35075 -500 35145 -490
rect 35075 -530 35095 -500
rect 35125 -530 35145 -500
rect 35075 -550 35145 -530
rect 35075 -580 35095 -550
rect 35125 -580 35145 -550
rect 35075 -600 35145 -580
rect 35075 -630 35095 -600
rect 35125 -630 35145 -600
rect 35075 -650 35145 -630
rect 35075 -680 35095 -650
rect 35125 -680 35145 -650
rect 35075 -690 35145 -680
rect 35160 -500 35230 -490
rect 35160 -530 35180 -500
rect 35210 -530 35230 -500
rect 35160 -550 35230 -530
rect 35160 -580 35180 -550
rect 35210 -580 35230 -550
rect 35160 -600 35230 -580
rect 35160 -630 35180 -600
rect 35210 -630 35230 -600
rect 35160 -650 35230 -630
rect 35160 -680 35180 -650
rect 35210 -680 35230 -650
rect 35160 -690 35230 -680
rect 35245 -500 35315 -490
rect 35245 -530 35265 -500
rect 35295 -530 35315 -500
rect 35245 -550 35315 -530
rect 35245 -580 35265 -550
rect 35295 -580 35315 -550
rect 35245 -600 35315 -580
rect 35245 -630 35265 -600
rect 35295 -630 35315 -600
rect 35245 -650 35315 -630
rect 35245 -680 35265 -650
rect 35295 -680 35315 -650
rect 35245 -690 35315 -680
rect 35330 -500 35400 -490
rect 35330 -530 35350 -500
rect 35380 -530 35400 -500
rect 35330 -550 35400 -530
rect 35330 -580 35350 -550
rect 35380 -580 35400 -550
rect 35330 -600 35400 -580
rect 35330 -630 35350 -600
rect 35380 -630 35400 -600
rect 35330 -650 35400 -630
rect 35330 -680 35350 -650
rect 35380 -680 35400 -650
rect 35330 -690 35400 -680
rect 35415 -500 35485 -490
rect 35415 -530 35435 -500
rect 35465 -530 35485 -500
rect 35415 -550 35485 -530
rect 35415 -580 35435 -550
rect 35465 -580 35485 -550
rect 35415 -600 35485 -580
rect 35415 -630 35435 -600
rect 35465 -630 35485 -600
rect 35415 -650 35485 -630
rect 35415 -680 35435 -650
rect 35465 -680 35485 -650
rect 35415 -690 35485 -680
rect 35500 -500 35570 -490
rect 35500 -530 35520 -500
rect 35550 -530 35570 -500
rect 35500 -550 35570 -530
rect 35500 -580 35520 -550
rect 35550 -580 35570 -550
rect 35500 -600 35570 -580
rect 35500 -630 35520 -600
rect 35550 -630 35570 -600
rect 35500 -650 35570 -630
rect 35500 -680 35520 -650
rect 35550 -680 35570 -650
rect 35500 -690 35570 -680
rect 35585 -500 35655 -490
rect 35585 -530 35605 -500
rect 35635 -530 35655 -500
rect 35585 -550 35655 -530
rect 35585 -580 35605 -550
rect 35635 -580 35655 -550
rect 35585 -600 35655 -580
rect 35585 -630 35605 -600
rect 35635 -630 35655 -600
rect 35585 -650 35655 -630
rect 35585 -680 35605 -650
rect 35635 -680 35655 -650
rect 35585 -690 35655 -680
rect 35670 -500 35740 -490
rect 35670 -530 35690 -500
rect 35720 -530 35740 -500
rect 35670 -550 35740 -530
rect 35670 -580 35690 -550
rect 35720 -580 35740 -550
rect 35670 -600 35740 -580
rect 35670 -630 35690 -600
rect 35720 -630 35740 -600
rect 35670 -650 35740 -630
rect 35670 -680 35690 -650
rect 35720 -680 35740 -650
rect 35670 -690 35740 -680
rect 35755 -500 35825 -490
rect 35755 -530 35775 -500
rect 35805 -530 35825 -500
rect 35755 -550 35825 -530
rect 35755 -580 35775 -550
rect 35805 -580 35825 -550
rect 35755 -600 35825 -580
rect 35755 -630 35775 -600
rect 35805 -630 35825 -600
rect 35755 -650 35825 -630
rect 35755 -680 35775 -650
rect 35805 -680 35825 -650
rect 35755 -690 35825 -680
rect 35840 -500 35910 -490
rect 35840 -530 35860 -500
rect 35890 -530 35910 -500
rect 35840 -550 35910 -530
rect 35840 -580 35860 -550
rect 35890 -580 35910 -550
rect 35840 -600 35910 -580
rect 35840 -630 35860 -600
rect 35890 -630 35910 -600
rect 35840 -650 35910 -630
rect 35840 -680 35860 -650
rect 35890 -680 35910 -650
rect 35840 -690 35910 -680
rect 35925 -500 35995 -490
rect 35925 -530 35945 -500
rect 35975 -530 35995 -500
rect 35925 -550 35995 -530
rect 35925 -580 35945 -550
rect 35975 -580 35995 -550
rect 35925 -600 35995 -580
rect 35925 -630 35945 -600
rect 35975 -630 35995 -600
rect 35925 -650 35995 -630
rect 35925 -680 35945 -650
rect 35975 -680 35995 -650
rect 35925 -690 35995 -680
rect 36010 -500 36080 -490
rect 36010 -530 36030 -500
rect 36060 -530 36080 -500
rect 36010 -550 36080 -530
rect 36010 -580 36030 -550
rect 36060 -580 36080 -550
rect 36010 -600 36080 -580
rect 36010 -630 36030 -600
rect 36060 -630 36080 -600
rect 36010 -650 36080 -630
rect 36010 -680 36030 -650
rect 36060 -680 36080 -650
rect 36010 -690 36080 -680
rect 36095 -500 36165 -490
rect 36095 -530 36115 -500
rect 36145 -530 36165 -500
rect 36095 -550 36165 -530
rect 36095 -580 36115 -550
rect 36145 -580 36165 -550
rect 36095 -600 36165 -580
rect 36095 -630 36115 -600
rect 36145 -630 36165 -600
rect 36095 -650 36165 -630
rect 36095 -680 36115 -650
rect 36145 -680 36165 -650
rect 36095 -690 36165 -680
rect 36180 -500 36250 -490
rect 36180 -530 36200 -500
rect 36230 -530 36250 -500
rect 36180 -550 36250 -530
rect 36180 -580 36200 -550
rect 36230 -580 36250 -550
rect 36180 -600 36250 -580
rect 36180 -630 36200 -600
rect 36230 -630 36250 -600
rect 36180 -650 36250 -630
rect 36180 -680 36200 -650
rect 36230 -680 36250 -650
rect 36180 -690 36250 -680
rect 36265 -500 36335 -490
rect 36265 -530 36285 -500
rect 36315 -530 36335 -500
rect 36265 -550 36335 -530
rect 36265 -580 36285 -550
rect 36315 -580 36335 -550
rect 36265 -600 36335 -580
rect 36265 -630 36285 -600
rect 36315 -630 36335 -600
rect 36265 -650 36335 -630
rect 36265 -680 36285 -650
rect 36315 -680 36335 -650
rect 36265 -690 36335 -680
rect 36350 -500 36420 -490
rect 36350 -530 36370 -500
rect 36400 -530 36420 -500
rect 36350 -550 36420 -530
rect 36350 -580 36370 -550
rect 36400 -580 36420 -550
rect 36350 -600 36420 -580
rect 36350 -630 36370 -600
rect 36400 -630 36420 -600
rect 36350 -650 36420 -630
rect 36350 -680 36370 -650
rect 36400 -680 36420 -650
rect 36350 -690 36420 -680
rect 36435 -500 36505 -490
rect 36435 -530 36455 -500
rect 36485 -530 36505 -500
rect 36435 -550 36505 -530
rect 36435 -580 36455 -550
rect 36485 -580 36505 -550
rect 36435 -600 36505 -580
rect 36435 -630 36455 -600
rect 36485 -630 36505 -600
rect 36435 -650 36505 -630
rect 36435 -680 36455 -650
rect 36485 -680 36505 -650
rect 36435 -690 36505 -680
rect 36520 -500 36590 -490
rect 36520 -530 36540 -500
rect 36570 -530 36590 -500
rect 36520 -550 36590 -530
rect 36520 -580 36540 -550
rect 36570 -580 36590 -550
rect 36520 -600 36590 -580
rect 36520 -630 36540 -600
rect 36570 -630 36590 -600
rect 36520 -650 36590 -630
rect 36520 -680 36540 -650
rect 36570 -680 36590 -650
rect 36520 -690 36590 -680
rect 36605 -500 36675 -490
rect 36605 -530 36625 -500
rect 36655 -530 36675 -500
rect 36605 -550 36675 -530
rect 36605 -580 36625 -550
rect 36655 -580 36675 -550
rect 36605 -600 36675 -580
rect 36605 -630 36625 -600
rect 36655 -630 36675 -600
rect 36605 -650 36675 -630
rect 36605 -680 36625 -650
rect 36655 -680 36675 -650
rect 36605 -690 36675 -680
rect 36690 -500 36760 -490
rect 36690 -530 36710 -500
rect 36740 -530 36760 -500
rect 36690 -550 36760 -530
rect 36690 -580 36710 -550
rect 36740 -580 36760 -550
rect 36690 -600 36760 -580
rect 36690 -630 36710 -600
rect 36740 -630 36760 -600
rect 36690 -650 36760 -630
rect 36690 -680 36710 -650
rect 36740 -680 36760 -650
rect 36690 -690 36760 -680
rect 36775 -500 36845 -490
rect 36775 -530 36795 -500
rect 36825 -530 36845 -500
rect 36775 -550 36845 -530
rect 36775 -580 36795 -550
rect 36825 -580 36845 -550
rect 36775 -600 36845 -580
rect 36775 -630 36795 -600
rect 36825 -630 36845 -600
rect 36775 -650 36845 -630
rect 36775 -680 36795 -650
rect 36825 -680 36845 -650
rect 36775 -690 36845 -680
rect 36860 -500 36930 -490
rect 36860 -530 36880 -500
rect 36910 -530 36930 -500
rect 36860 -550 36930 -530
rect 36860 -580 36880 -550
rect 36910 -580 36930 -550
rect 36860 -600 36930 -580
rect 36860 -630 36880 -600
rect 36910 -630 36930 -600
rect 36860 -650 36930 -630
rect 36860 -680 36880 -650
rect 36910 -680 36930 -650
rect 36860 -690 36930 -680
rect 36945 -500 37015 -490
rect 36945 -530 36965 -500
rect 36995 -530 37015 -500
rect 36945 -550 37015 -530
rect 36945 -580 36965 -550
rect 36995 -580 37015 -550
rect 36945 -600 37015 -580
rect 36945 -630 36965 -600
rect 36995 -630 37015 -600
rect 36945 -650 37015 -630
rect 36945 -680 36965 -650
rect 36995 -680 37015 -650
rect 36945 -690 37015 -680
rect 37030 -500 37100 -490
rect 37030 -530 37050 -500
rect 37080 -530 37100 -500
rect 37030 -550 37100 -530
rect 37030 -580 37050 -550
rect 37080 -580 37100 -550
rect 37030 -600 37100 -580
rect 37030 -630 37050 -600
rect 37080 -630 37100 -600
rect 37030 -650 37100 -630
rect 37030 -680 37050 -650
rect 37080 -680 37100 -650
rect 37030 -690 37100 -680
rect 37115 -500 37185 -490
rect 37115 -530 37135 -500
rect 37165 -530 37185 -500
rect 37115 -550 37185 -530
rect 37115 -580 37135 -550
rect 37165 -580 37185 -550
rect 37115 -600 37185 -580
rect 37115 -630 37135 -600
rect 37165 -630 37185 -600
rect 37115 -650 37185 -630
rect 37115 -680 37135 -650
rect 37165 -680 37185 -650
rect 37115 -690 37185 -680
rect 37200 -500 37270 -490
rect 37200 -530 37220 -500
rect 37250 -530 37270 -500
rect 37200 -550 37270 -530
rect 37200 -580 37220 -550
rect 37250 -580 37270 -550
rect 37200 -600 37270 -580
rect 37200 -630 37220 -600
rect 37250 -630 37270 -600
rect 37200 -650 37270 -630
rect 37200 -680 37220 -650
rect 37250 -680 37270 -650
rect 37200 -690 37270 -680
rect 37285 -500 37355 -490
rect 37285 -530 37305 -500
rect 37335 -530 37355 -500
rect 37285 -550 37355 -530
rect 37285 -580 37305 -550
rect 37335 -580 37355 -550
rect 37285 -600 37355 -580
rect 37285 -630 37305 -600
rect 37335 -630 37355 -600
rect 37285 -650 37355 -630
rect 37285 -680 37305 -650
rect 37335 -680 37355 -650
rect 37285 -690 37355 -680
rect 37370 -500 37440 -490
rect 37370 -530 37390 -500
rect 37420 -530 37440 -500
rect 37370 -550 37440 -530
rect 37370 -580 37390 -550
rect 37420 -580 37440 -550
rect 37370 -600 37440 -580
rect 37370 -630 37390 -600
rect 37420 -630 37440 -600
rect 37370 -650 37440 -630
rect 37370 -680 37390 -650
rect 37420 -680 37440 -650
rect 37370 -690 37440 -680
rect 37455 -500 37525 -490
rect 37455 -530 37475 -500
rect 37505 -530 37525 -500
rect 37455 -550 37525 -530
rect 37455 -580 37475 -550
rect 37505 -580 37525 -550
rect 37455 -600 37525 -580
rect 37455 -630 37475 -600
rect 37505 -630 37525 -600
rect 37455 -650 37525 -630
rect 37455 -680 37475 -650
rect 37505 -680 37525 -650
rect 37455 -690 37525 -680
rect 37540 -500 37610 -490
rect 37540 -530 37560 -500
rect 37590 -530 37610 -500
rect 37540 -550 37610 -530
rect 37540 -580 37560 -550
rect 37590 -580 37610 -550
rect 37540 -600 37610 -580
rect 37540 -630 37560 -600
rect 37590 -630 37610 -600
rect 37540 -650 37610 -630
rect 37540 -680 37560 -650
rect 37590 -680 37610 -650
rect 37540 -690 37610 -680
rect 37625 -500 37695 -490
rect 37625 -530 37645 -500
rect 37675 -530 37695 -500
rect 37625 -550 37695 -530
rect 37625 -580 37645 -550
rect 37675 -580 37695 -550
rect 37625 -600 37695 -580
rect 37625 -630 37645 -600
rect 37675 -630 37695 -600
rect 37625 -650 37695 -630
rect 37625 -680 37645 -650
rect 37675 -680 37695 -650
rect 37625 -690 37695 -680
rect 37710 -500 37780 -490
rect 37710 -530 37730 -500
rect 37760 -530 37780 -500
rect 37710 -550 37780 -530
rect 37710 -580 37730 -550
rect 37760 -580 37780 -550
rect 37710 -600 37780 -580
rect 37710 -630 37730 -600
rect 37760 -630 37780 -600
rect 37710 -650 37780 -630
rect 37710 -680 37730 -650
rect 37760 -680 37780 -650
rect 37710 -690 37780 -680
rect 37795 -500 37865 -490
rect 37795 -530 37815 -500
rect 37845 -530 37865 -500
rect 37795 -550 37865 -530
rect 37795 -580 37815 -550
rect 37845 -580 37865 -550
rect 37795 -600 37865 -580
rect 37795 -630 37815 -600
rect 37845 -630 37865 -600
rect 37795 -650 37865 -630
rect 37795 -680 37815 -650
rect 37845 -680 37865 -650
rect 37795 -690 37865 -680
rect 37880 -500 37950 -490
rect 37880 -530 37900 -500
rect 37930 -530 37950 -500
rect 37880 -550 37950 -530
rect 37880 -580 37900 -550
rect 37930 -580 37950 -550
rect 37880 -600 37950 -580
rect 37880 -630 37900 -600
rect 37930 -630 37950 -600
rect 37880 -650 37950 -630
rect 37880 -680 37900 -650
rect 37930 -680 37950 -650
rect 37880 -690 37950 -680
rect 37965 -500 38035 -490
rect 37965 -530 37985 -500
rect 38015 -530 38035 -500
rect 37965 -550 38035 -530
rect 37965 -580 37985 -550
rect 38015 -580 38035 -550
rect 37965 -600 38035 -580
rect 37965 -630 37985 -600
rect 38015 -630 38035 -600
rect 37965 -650 38035 -630
rect 37965 -680 37985 -650
rect 38015 -680 38035 -650
rect 37965 -690 38035 -680
rect 38050 -500 38120 -490
rect 38050 -530 38070 -500
rect 38100 -530 38120 -500
rect 38050 -550 38120 -530
rect 38050 -580 38070 -550
rect 38100 -580 38120 -550
rect 38050 -600 38120 -580
rect 38050 -630 38070 -600
rect 38100 -630 38120 -600
rect 38050 -650 38120 -630
rect 38050 -680 38070 -650
rect 38100 -680 38120 -650
rect 38050 -690 38120 -680
rect 38135 -500 38205 -490
rect 38135 -530 38155 -500
rect 38185 -530 38205 -500
rect 38135 -550 38205 -530
rect 38135 -580 38155 -550
rect 38185 -580 38205 -550
rect 38135 -600 38205 -580
rect 38135 -630 38155 -600
rect 38185 -630 38205 -600
rect 38135 -650 38205 -630
rect 38135 -680 38155 -650
rect 38185 -680 38205 -650
rect 38135 -690 38205 -680
rect 38220 -500 38290 -490
rect 38220 -530 38240 -500
rect 38270 -530 38290 -500
rect 38220 -550 38290 -530
rect 38220 -580 38240 -550
rect 38270 -580 38290 -550
rect 38220 -600 38290 -580
rect 38220 -630 38240 -600
rect 38270 -630 38290 -600
rect 38220 -650 38290 -630
rect 38220 -680 38240 -650
rect 38270 -680 38290 -650
rect 38220 -690 38290 -680
rect 38305 -500 38375 -490
rect 38305 -530 38325 -500
rect 38355 -530 38375 -500
rect 38305 -550 38375 -530
rect 38305 -580 38325 -550
rect 38355 -580 38375 -550
rect 38305 -600 38375 -580
rect 38305 -630 38325 -600
rect 38355 -630 38375 -600
rect 38305 -650 38375 -630
rect 38305 -680 38325 -650
rect 38355 -680 38375 -650
rect 38305 -690 38375 -680
rect 38390 -500 38460 -490
rect 38390 -530 38410 -500
rect 38440 -530 38460 -500
rect 38390 -550 38460 -530
rect 38390 -580 38410 -550
rect 38440 -580 38460 -550
rect 38390 -600 38460 -580
rect 38390 -630 38410 -600
rect 38440 -630 38460 -600
rect 38390 -650 38460 -630
rect 38390 -680 38410 -650
rect 38440 -680 38460 -650
rect 38390 -690 38460 -680
rect 38475 -500 38545 -490
rect 38475 -530 38495 -500
rect 38525 -530 38545 -500
rect 38475 -550 38545 -530
rect 38475 -580 38495 -550
rect 38525 -580 38545 -550
rect 38475 -600 38545 -580
rect 38475 -630 38495 -600
rect 38525 -630 38545 -600
rect 38475 -650 38545 -630
rect 38475 -680 38495 -650
rect 38525 -680 38545 -650
rect 38475 -690 38545 -680
rect 38560 -500 38630 -490
rect 38560 -530 38580 -500
rect 38610 -530 38630 -500
rect 38560 -550 38630 -530
rect 38560 -580 38580 -550
rect 38610 -580 38630 -550
rect 38560 -600 38630 -580
rect 38560 -630 38580 -600
rect 38610 -630 38630 -600
rect 38560 -650 38630 -630
rect 38560 -680 38580 -650
rect 38610 -680 38630 -650
rect 38560 -690 38630 -680
rect 38645 -500 38715 -490
rect 38645 -530 38665 -500
rect 38695 -530 38715 -500
rect 38645 -550 38715 -530
rect 38645 -580 38665 -550
rect 38695 -580 38715 -550
rect 38645 -600 38715 -580
rect 38645 -630 38665 -600
rect 38695 -630 38715 -600
rect 38645 -650 38715 -630
rect 38645 -680 38665 -650
rect 38695 -680 38715 -650
rect 38645 -690 38715 -680
rect 38730 -500 38800 -490
rect 38730 -530 38750 -500
rect 38780 -530 38800 -500
rect 38730 -550 38800 -530
rect 38730 -580 38750 -550
rect 38780 -580 38800 -550
rect 38730 -600 38800 -580
rect 38730 -630 38750 -600
rect 38780 -630 38800 -600
rect 38730 -650 38800 -630
rect 38730 -680 38750 -650
rect 38780 -680 38800 -650
rect 38730 -690 38800 -680
rect 38815 -500 38885 -490
rect 38815 -530 38835 -500
rect 38865 -530 38885 -500
rect 38815 -550 38885 -530
rect 38815 -580 38835 -550
rect 38865 -580 38885 -550
rect 38815 -600 38885 -580
rect 38815 -630 38835 -600
rect 38865 -630 38885 -600
rect 38815 -650 38885 -630
rect 38815 -680 38835 -650
rect 38865 -680 38885 -650
rect 38815 -690 38885 -680
rect 38900 -500 38970 -490
rect 38900 -530 38920 -500
rect 38950 -530 38970 -500
rect 38900 -550 38970 -530
rect 38900 -580 38920 -550
rect 38950 -580 38970 -550
rect 38900 -600 38970 -580
rect 38900 -630 38920 -600
rect 38950 -630 38970 -600
rect 38900 -650 38970 -630
rect 38900 -680 38920 -650
rect 38950 -680 38970 -650
rect 38900 -690 38970 -680
rect 38985 -500 39055 -490
rect 38985 -530 39005 -500
rect 39035 -530 39055 -500
rect 38985 -550 39055 -530
rect 38985 -580 39005 -550
rect 39035 -580 39055 -550
rect 38985 -600 39055 -580
rect 38985 -630 39005 -600
rect 39035 -630 39055 -600
rect 38985 -650 39055 -630
rect 38985 -680 39005 -650
rect 39035 -680 39055 -650
rect 38985 -690 39055 -680
rect 39070 -500 39140 -490
rect 39070 -530 39090 -500
rect 39120 -530 39140 -500
rect 39070 -550 39140 -530
rect 39070 -580 39090 -550
rect 39120 -580 39140 -550
rect 39070 -600 39140 -580
rect 39070 -630 39090 -600
rect 39120 -630 39140 -600
rect 39070 -650 39140 -630
rect 39070 -680 39090 -650
rect 39120 -680 39140 -650
rect 39070 -690 39140 -680
rect 39155 -500 39225 -490
rect 39155 -530 39175 -500
rect 39205 -530 39225 -500
rect 39155 -550 39225 -530
rect 39155 -580 39175 -550
rect 39205 -580 39225 -550
rect 39155 -600 39225 -580
rect 39155 -630 39175 -600
rect 39205 -630 39225 -600
rect 39155 -650 39225 -630
rect 39155 -680 39175 -650
rect 39205 -680 39225 -650
rect 39155 -690 39225 -680
rect 39240 -500 39310 -490
rect 39240 -530 39260 -500
rect 39290 -530 39310 -500
rect 39240 -550 39310 -530
rect 39240 -580 39260 -550
rect 39290 -580 39310 -550
rect 39240 -600 39310 -580
rect 39240 -630 39260 -600
rect 39290 -630 39310 -600
rect 39240 -650 39310 -630
rect 39240 -680 39260 -650
rect 39290 -680 39310 -650
rect 39240 -690 39310 -680
rect 39325 -500 39395 -490
rect 39325 -530 39345 -500
rect 39375 -530 39395 -500
rect 39325 -550 39395 -530
rect 39325 -580 39345 -550
rect 39375 -580 39395 -550
rect 39325 -600 39395 -580
rect 39325 -630 39345 -600
rect 39375 -630 39395 -600
rect 39325 -650 39395 -630
rect 39325 -680 39345 -650
rect 39375 -680 39395 -650
rect 39325 -690 39395 -680
rect 39410 -500 39480 -490
rect 39410 -530 39430 -500
rect 39460 -530 39480 -500
rect 39410 -550 39480 -530
rect 39410 -580 39430 -550
rect 39460 -580 39480 -550
rect 39410 -600 39480 -580
rect 39410 -630 39430 -600
rect 39460 -630 39480 -600
rect 39410 -650 39480 -630
rect 39410 -680 39430 -650
rect 39460 -680 39480 -650
rect 39410 -690 39480 -680
rect 39495 -500 39565 -490
rect 39495 -530 39515 -500
rect 39545 -530 39565 -500
rect 39495 -550 39565 -530
rect 39495 -580 39515 -550
rect 39545 -580 39565 -550
rect 39495 -600 39565 -580
rect 39495 -630 39515 -600
rect 39545 -630 39565 -600
rect 39495 -650 39565 -630
rect 39495 -680 39515 -650
rect 39545 -680 39565 -650
rect 39495 -690 39565 -680
rect 39580 -500 39650 -490
rect 39580 -530 39600 -500
rect 39630 -530 39650 -500
rect 39580 -550 39650 -530
rect 39580 -580 39600 -550
rect 39630 -580 39650 -550
rect 39580 -600 39650 -580
rect 39580 -630 39600 -600
rect 39630 -630 39650 -600
rect 39580 -650 39650 -630
rect 39580 -680 39600 -650
rect 39630 -680 39650 -650
rect 39580 -690 39650 -680
rect 39665 -500 39735 -490
rect 39665 -530 39685 -500
rect 39715 -530 39735 -500
rect 39665 -550 39735 -530
rect 39665 -580 39685 -550
rect 39715 -580 39735 -550
rect 39665 -600 39735 -580
rect 39665 -630 39685 -600
rect 39715 -630 39735 -600
rect 39665 -650 39735 -630
rect 39665 -680 39685 -650
rect 39715 -680 39735 -650
rect 39665 -690 39735 -680
rect 39750 -500 39820 -490
rect 39750 -530 39770 -500
rect 39800 -530 39820 -500
rect 39750 -550 39820 -530
rect 39750 -580 39770 -550
rect 39800 -580 39820 -550
rect 39750 -600 39820 -580
rect 39750 -630 39770 -600
rect 39800 -630 39820 -600
rect 39750 -650 39820 -630
rect 39750 -680 39770 -650
rect 39800 -680 39820 -650
rect 39750 -690 39820 -680
rect 39835 -500 39905 -490
rect 39835 -530 39855 -500
rect 39885 -530 39905 -500
rect 39835 -550 39905 -530
rect 39835 -580 39855 -550
rect 39885 -580 39905 -550
rect 39835 -600 39905 -580
rect 39835 -630 39855 -600
rect 39885 -630 39905 -600
rect 39835 -650 39905 -630
rect 39835 -680 39855 -650
rect 39885 -680 39905 -650
rect 39835 -690 39905 -680
rect 39920 -500 39990 -490
rect 39920 -530 39940 -500
rect 39970 -530 39990 -500
rect 39920 -550 39990 -530
rect 39920 -580 39940 -550
rect 39970 -580 39990 -550
rect 39920 -600 39990 -580
rect 39920 -630 39940 -600
rect 39970 -630 39990 -600
rect 39920 -650 39990 -630
rect 39920 -680 39940 -650
rect 39970 -680 39990 -650
rect 39920 -690 39990 -680
rect 40005 -500 40075 -490
rect 40005 -530 40025 -500
rect 40055 -530 40075 -500
rect 40005 -550 40075 -530
rect 40005 -580 40025 -550
rect 40055 -580 40075 -550
rect 40005 -600 40075 -580
rect 40005 -630 40025 -600
rect 40055 -630 40075 -600
rect 40005 -650 40075 -630
rect 40005 -680 40025 -650
rect 40055 -680 40075 -650
rect 40005 -690 40075 -680
rect 40090 -500 40160 -490
rect 40090 -530 40110 -500
rect 40140 -530 40160 -500
rect 40090 -550 40160 -530
rect 40090 -580 40110 -550
rect 40140 -580 40160 -550
rect 40090 -600 40160 -580
rect 40090 -630 40110 -600
rect 40140 -630 40160 -600
rect 40090 -650 40160 -630
rect 40090 -680 40110 -650
rect 40140 -680 40160 -650
rect 40090 -690 40160 -680
rect 40175 -500 40245 -490
rect 40175 -530 40195 -500
rect 40225 -530 40245 -500
rect 40175 -550 40245 -530
rect 40175 -580 40195 -550
rect 40225 -580 40245 -550
rect 40175 -600 40245 -580
rect 40175 -630 40195 -600
rect 40225 -630 40245 -600
rect 40175 -650 40245 -630
rect 40175 -680 40195 -650
rect 40225 -680 40245 -650
rect 40175 -690 40245 -680
rect 40260 -500 40330 -490
rect 40260 -530 40280 -500
rect 40310 -530 40330 -500
rect 40260 -550 40330 -530
rect 40260 -580 40280 -550
rect 40310 -580 40330 -550
rect 40260 -600 40330 -580
rect 40260 -630 40280 -600
rect 40310 -630 40330 -600
rect 40260 -650 40330 -630
rect 40260 -680 40280 -650
rect 40310 -680 40330 -650
rect 40260 -690 40330 -680
rect 40345 -500 40415 -490
rect 40345 -530 40365 -500
rect 40395 -530 40415 -500
rect 40345 -550 40415 -530
rect 40345 -580 40365 -550
rect 40395 -580 40415 -550
rect 40345 -600 40415 -580
rect 40345 -630 40365 -600
rect 40395 -630 40415 -600
rect 40345 -650 40415 -630
rect 40345 -680 40365 -650
rect 40395 -680 40415 -650
rect 40345 -690 40415 -680
rect 40430 -500 40500 -490
rect 40430 -530 40450 -500
rect 40480 -530 40500 -500
rect 40430 -550 40500 -530
rect 40430 -580 40450 -550
rect 40480 -580 40500 -550
rect 40430 -600 40500 -580
rect 40430 -630 40450 -600
rect 40480 -630 40500 -600
rect 40430 -650 40500 -630
rect 40430 -680 40450 -650
rect 40480 -680 40500 -650
rect 40430 -690 40500 -680
rect 40515 -500 40585 -490
rect 40515 -530 40535 -500
rect 40565 -530 40585 -500
rect 40515 -550 40585 -530
rect 40515 -580 40535 -550
rect 40565 -580 40585 -550
rect 40515 -600 40585 -580
rect 40515 -630 40535 -600
rect 40565 -630 40585 -600
rect 40515 -650 40585 -630
rect 40515 -680 40535 -650
rect 40565 -680 40585 -650
rect 40515 -690 40585 -680
rect 40600 -500 40670 -490
rect 40600 -530 40620 -500
rect 40650 -530 40670 -500
rect 40600 -550 40670 -530
rect 40600 -580 40620 -550
rect 40650 -580 40670 -550
rect 40600 -600 40670 -580
rect 40600 -630 40620 -600
rect 40650 -630 40670 -600
rect 40600 -650 40670 -630
rect 40600 -680 40620 -650
rect 40650 -680 40670 -650
rect 40600 -690 40670 -680
rect 40685 -500 40755 -490
rect 40685 -530 40705 -500
rect 40735 -530 40755 -500
rect 40685 -550 40755 -530
rect 40685 -580 40705 -550
rect 40735 -580 40755 -550
rect 40685 -600 40755 -580
rect 40685 -630 40705 -600
rect 40735 -630 40755 -600
rect 40685 -650 40755 -630
rect 40685 -680 40705 -650
rect 40735 -680 40755 -650
rect 40685 -690 40755 -680
rect 40770 -500 40840 -490
rect 40770 -530 40790 -500
rect 40820 -530 40840 -500
rect 40770 -550 40840 -530
rect 40770 -580 40790 -550
rect 40820 -580 40840 -550
rect 40770 -600 40840 -580
rect 40770 -630 40790 -600
rect 40820 -630 40840 -600
rect 40770 -650 40840 -630
rect 40770 -680 40790 -650
rect 40820 -680 40840 -650
rect 40770 -690 40840 -680
rect 40855 -500 40925 -490
rect 40855 -530 40875 -500
rect 40905 -530 40925 -500
rect 40855 -550 40925 -530
rect 40855 -580 40875 -550
rect 40905 -580 40925 -550
rect 40855 -600 40925 -580
rect 40855 -630 40875 -600
rect 40905 -630 40925 -600
rect 40855 -650 40925 -630
rect 40855 -680 40875 -650
rect 40905 -680 40925 -650
rect 40855 -690 40925 -680
rect 40940 -500 41010 -490
rect 40940 -530 40960 -500
rect 40990 -530 41010 -500
rect 40940 -550 41010 -530
rect 40940 -580 40960 -550
rect 40990 -580 41010 -550
rect 40940 -600 41010 -580
rect 40940 -630 40960 -600
rect 40990 -630 41010 -600
rect 40940 -650 41010 -630
rect 40940 -680 40960 -650
rect 40990 -680 41010 -650
rect 40940 -690 41010 -680
rect 41025 -500 41095 -490
rect 41025 -530 41045 -500
rect 41075 -530 41095 -500
rect 41025 -550 41095 -530
rect 41025 -580 41045 -550
rect 41075 -580 41095 -550
rect 41025 -600 41095 -580
rect 41025 -630 41045 -600
rect 41075 -630 41095 -600
rect 41025 -650 41095 -630
rect 41025 -680 41045 -650
rect 41075 -680 41095 -650
rect 41025 -690 41095 -680
rect 41110 -500 41180 -490
rect 41110 -530 41130 -500
rect 41160 -530 41180 -500
rect 41110 -550 41180 -530
rect 41110 -580 41130 -550
rect 41160 -580 41180 -550
rect 41110 -600 41180 -580
rect 41110 -630 41130 -600
rect 41160 -630 41180 -600
rect 41110 -650 41180 -630
rect 41110 -680 41130 -650
rect 41160 -680 41180 -650
rect 41110 -690 41180 -680
rect 41195 -500 41265 -490
rect 41195 -530 41215 -500
rect 41245 -530 41265 -500
rect 41195 -550 41265 -530
rect 41195 -580 41215 -550
rect 41245 -580 41265 -550
rect 41195 -600 41265 -580
rect 41195 -630 41215 -600
rect 41245 -630 41265 -600
rect 41195 -650 41265 -630
rect 41195 -680 41215 -650
rect 41245 -680 41265 -650
rect 41195 -690 41265 -680
rect 41280 -500 41350 -490
rect 41280 -530 41300 -500
rect 41330 -530 41350 -500
rect 41280 -550 41350 -530
rect 41280 -580 41300 -550
rect 41330 -580 41350 -550
rect 41280 -600 41350 -580
rect 41280 -630 41300 -600
rect 41330 -630 41350 -600
rect 41280 -650 41350 -630
rect 41280 -680 41300 -650
rect 41330 -680 41350 -650
rect 41280 -690 41350 -680
rect 41365 -500 41435 -490
rect 41365 -530 41385 -500
rect 41415 -530 41435 -500
rect 41365 -550 41435 -530
rect 41365 -580 41385 -550
rect 41415 -580 41435 -550
rect 41365 -600 41435 -580
rect 41365 -630 41385 -600
rect 41415 -630 41435 -600
rect 41365 -650 41435 -630
rect 41365 -680 41385 -650
rect 41415 -680 41435 -650
rect 41365 -690 41435 -680
rect 41450 -500 41520 -490
rect 41450 -530 41470 -500
rect 41500 -530 41520 -500
rect 41450 -550 41520 -530
rect 41450 -580 41470 -550
rect 41500 -580 41520 -550
rect 41450 -600 41520 -580
rect 41450 -630 41470 -600
rect 41500 -630 41520 -600
rect 41450 -650 41520 -630
rect 41450 -680 41470 -650
rect 41500 -680 41520 -650
rect 41450 -690 41520 -680
rect 41535 -500 41605 -490
rect 41535 -530 41555 -500
rect 41585 -530 41605 -500
rect 41535 -550 41605 -530
rect 41535 -580 41555 -550
rect 41585 -580 41605 -550
rect 41535 -600 41605 -580
rect 41535 -630 41555 -600
rect 41585 -630 41605 -600
rect 41535 -650 41605 -630
rect 41535 -680 41555 -650
rect 41585 -680 41605 -650
rect 41535 -690 41605 -680
rect 41620 -500 41690 -490
rect 41620 -530 41640 -500
rect 41670 -530 41690 -500
rect 41620 -550 41690 -530
rect 41620 -580 41640 -550
rect 41670 -580 41690 -550
rect 41620 -600 41690 -580
rect 41620 -630 41640 -600
rect 41670 -630 41690 -600
rect 41620 -650 41690 -630
rect 41620 -680 41640 -650
rect 41670 -680 41690 -650
rect 41620 -690 41690 -680
rect 41705 -500 41775 -490
rect 41705 -530 41725 -500
rect 41755 -530 41775 -500
rect 41705 -550 41775 -530
rect 41705 -580 41725 -550
rect 41755 -580 41775 -550
rect 41705 -600 41775 -580
rect 41705 -630 41725 -600
rect 41755 -630 41775 -600
rect 41705 -650 41775 -630
rect 41705 -680 41725 -650
rect 41755 -680 41775 -650
rect 41705 -690 41775 -680
rect 41790 -500 41860 -490
rect 41790 -530 41810 -500
rect 41840 -530 41860 -500
rect 41790 -550 41860 -530
rect 41790 -580 41810 -550
rect 41840 -580 41860 -550
rect 41790 -600 41860 -580
rect 41790 -630 41810 -600
rect 41840 -630 41860 -600
rect 41790 -650 41860 -630
rect 41790 -680 41810 -650
rect 41840 -680 41860 -650
rect 41790 -690 41860 -680
rect 41875 -500 41945 -490
rect 41875 -530 41895 -500
rect 41925 -530 41945 -500
rect 41875 -550 41945 -530
rect 41875 -580 41895 -550
rect 41925 -580 41945 -550
rect 41875 -600 41945 -580
rect 41875 -630 41895 -600
rect 41925 -630 41945 -600
rect 41875 -650 41945 -630
rect 41875 -680 41895 -650
rect 41925 -680 41945 -650
rect 41875 -690 41945 -680
rect 41960 -500 42030 -490
rect 41960 -530 41980 -500
rect 42010 -530 42030 -500
rect 41960 -550 42030 -530
rect 41960 -580 41980 -550
rect 42010 -580 42030 -550
rect 41960 -600 42030 -580
rect 41960 -630 41980 -600
rect 42010 -630 42030 -600
rect 41960 -650 42030 -630
rect 41960 -680 41980 -650
rect 42010 -680 42030 -650
rect 41960 -690 42030 -680
rect 42045 -500 42115 -490
rect 42045 -530 42065 -500
rect 42095 -530 42115 -500
rect 42045 -550 42115 -530
rect 42045 -580 42065 -550
rect 42095 -580 42115 -550
rect 42045 -600 42115 -580
rect 42045 -630 42065 -600
rect 42095 -630 42115 -600
rect 42045 -650 42115 -630
rect 42045 -680 42065 -650
rect 42095 -680 42115 -650
rect 42045 -690 42115 -680
rect 42130 -500 42200 -490
rect 42130 -530 42150 -500
rect 42180 -530 42200 -500
rect 42130 -550 42200 -530
rect 42130 -580 42150 -550
rect 42180 -580 42200 -550
rect 42130 -600 42200 -580
rect 42130 -630 42150 -600
rect 42180 -630 42200 -600
rect 42130 -650 42200 -630
rect 42130 -680 42150 -650
rect 42180 -680 42200 -650
rect 42130 -690 42200 -680
rect 42215 -500 42285 -490
rect 42215 -530 42235 -500
rect 42265 -530 42285 -500
rect 42215 -550 42285 -530
rect 42215 -580 42235 -550
rect 42265 -580 42285 -550
rect 42215 -600 42285 -580
rect 42215 -630 42235 -600
rect 42265 -630 42285 -600
rect 42215 -650 42285 -630
rect 42215 -680 42235 -650
rect 42265 -680 42285 -650
rect 42215 -690 42285 -680
rect 42300 -500 42370 -490
rect 42300 -530 42320 -500
rect 42350 -530 42370 -500
rect 42300 -550 42370 -530
rect 42300 -580 42320 -550
rect 42350 -580 42370 -550
rect 42300 -600 42370 -580
rect 42300 -630 42320 -600
rect 42350 -630 42370 -600
rect 42300 -650 42370 -630
rect 42300 -680 42320 -650
rect 42350 -680 42370 -650
rect 42300 -690 42370 -680
rect 42385 -500 42455 -490
rect 42385 -530 42405 -500
rect 42435 -530 42455 -500
rect 42385 -550 42455 -530
rect 42385 -580 42405 -550
rect 42435 -580 42455 -550
rect 42385 -600 42455 -580
rect 42385 -630 42405 -600
rect 42435 -630 42455 -600
rect 42385 -650 42455 -630
rect 42385 -680 42405 -650
rect 42435 -680 42455 -650
rect 42385 -690 42455 -680
rect 42470 -500 42540 -490
rect 42470 -530 42490 -500
rect 42520 -530 42540 -500
rect 42470 -550 42540 -530
rect 42470 -580 42490 -550
rect 42520 -580 42540 -550
rect 42470 -600 42540 -580
rect 42470 -630 42490 -600
rect 42520 -630 42540 -600
rect 42470 -650 42540 -630
rect 42470 -680 42490 -650
rect 42520 -680 42540 -650
rect 42470 -690 42540 -680
rect 42555 -500 42625 -490
rect 42555 -530 42575 -500
rect 42605 -530 42625 -500
rect 42555 -550 42625 -530
rect 42555 -580 42575 -550
rect 42605 -580 42625 -550
rect 42555 -600 42625 -580
rect 42555 -630 42575 -600
rect 42605 -630 42625 -600
rect 42555 -650 42625 -630
rect 42555 -680 42575 -650
rect 42605 -680 42625 -650
rect 42555 -690 42625 -680
rect 42640 -500 42710 -490
rect 42640 -530 42660 -500
rect 42690 -530 42710 -500
rect 42640 -550 42710 -530
rect 42640 -580 42660 -550
rect 42690 -580 42710 -550
rect 42640 -600 42710 -580
rect 42640 -630 42660 -600
rect 42690 -630 42710 -600
rect 42640 -650 42710 -630
rect 42640 -680 42660 -650
rect 42690 -680 42710 -650
rect 42640 -690 42710 -680
rect 42725 -500 42795 -490
rect 42725 -530 42745 -500
rect 42775 -530 42795 -500
rect 42725 -550 42795 -530
rect 42725 -580 42745 -550
rect 42775 -580 42795 -550
rect 42725 -600 42795 -580
rect 42725 -630 42745 -600
rect 42775 -630 42795 -600
rect 42725 -650 42795 -630
rect 42725 -680 42745 -650
rect 42775 -680 42795 -650
rect 42725 -690 42795 -680
rect 42810 -500 42880 -490
rect 42810 -530 42830 -500
rect 42860 -530 42880 -500
rect 42810 -550 42880 -530
rect 42810 -580 42830 -550
rect 42860 -580 42880 -550
rect 42810 -600 42880 -580
rect 42810 -630 42830 -600
rect 42860 -630 42880 -600
rect 42810 -650 42880 -630
rect 42810 -680 42830 -650
rect 42860 -680 42880 -650
rect 42810 -690 42880 -680
rect 42895 -500 42965 -490
rect 42895 -530 42915 -500
rect 42945 -530 42965 -500
rect 42895 -550 42965 -530
rect 42895 -580 42915 -550
rect 42945 -580 42965 -550
rect 42895 -600 42965 -580
rect 42895 -630 42915 -600
rect 42945 -630 42965 -600
rect 42895 -650 42965 -630
rect 42895 -680 42915 -650
rect 42945 -680 42965 -650
rect 42895 -690 42965 -680
rect 42980 -500 43050 -490
rect 42980 -530 43000 -500
rect 43030 -530 43050 -500
rect 42980 -550 43050 -530
rect 42980 -580 43000 -550
rect 43030 -580 43050 -550
rect 42980 -600 43050 -580
rect 42980 -630 43000 -600
rect 43030 -630 43050 -600
rect 42980 -650 43050 -630
rect 42980 -680 43000 -650
rect 43030 -680 43050 -650
rect 42980 -690 43050 -680
rect 43065 -500 43135 -490
rect 43065 -530 43085 -500
rect 43115 -530 43135 -500
rect 43065 -550 43135 -530
rect 43065 -580 43085 -550
rect 43115 -580 43135 -550
rect 43065 -600 43135 -580
rect 43065 -630 43085 -600
rect 43115 -630 43135 -600
rect 43065 -650 43135 -630
rect 43065 -680 43085 -650
rect 43115 -680 43135 -650
rect 43065 -690 43135 -680
rect 43150 -500 43220 -490
rect 43150 -530 43170 -500
rect 43200 -530 43220 -500
rect 43150 -550 43220 -530
rect 43150 -580 43170 -550
rect 43200 -580 43220 -550
rect 43150 -600 43220 -580
rect 43150 -630 43170 -600
rect 43200 -630 43220 -600
rect 43150 -650 43220 -630
rect 43150 -680 43170 -650
rect 43200 -680 43220 -650
rect 43150 -690 43220 -680
rect 43235 -500 43305 -490
rect 43235 -530 43255 -500
rect 43285 -530 43305 -500
rect 43235 -550 43305 -530
rect 43235 -580 43255 -550
rect 43285 -580 43305 -550
rect 43235 -600 43305 -580
rect 43235 -630 43255 -600
rect 43285 -630 43305 -600
rect 43235 -650 43305 -630
rect 43235 -680 43255 -650
rect 43285 -680 43305 -650
rect 43235 -690 43305 -680
rect 43320 -500 43390 -490
rect 43320 -530 43340 -500
rect 43370 -530 43390 -500
rect 43320 -550 43390 -530
rect 43320 -580 43340 -550
rect 43370 -580 43390 -550
rect 43320 -600 43390 -580
rect 43320 -630 43340 -600
rect 43370 -630 43390 -600
rect 43320 -650 43390 -630
rect 43320 -680 43340 -650
rect 43370 -680 43390 -650
rect 43320 -690 43390 -680
rect 43405 -500 43475 -490
rect 43405 -530 43425 -500
rect 43455 -530 43475 -500
rect 43405 -550 43475 -530
rect 43405 -580 43425 -550
rect 43455 -580 43475 -550
rect 43405 -600 43475 -580
rect 43405 -630 43425 -600
rect 43455 -630 43475 -600
rect 43405 -650 43475 -630
rect 43405 -680 43425 -650
rect 43455 -680 43475 -650
rect 43405 -690 43475 -680
rect 43490 -500 43560 -490
rect 43490 -530 43510 -500
rect 43540 -530 43560 -500
rect 43490 -550 43560 -530
rect 43490 -580 43510 -550
rect 43540 -580 43560 -550
rect 43490 -600 43560 -580
rect 43490 -630 43510 -600
rect 43540 -630 43560 -600
rect 43490 -650 43560 -630
rect 43490 -680 43510 -650
rect 43540 -680 43560 -650
rect 43490 -690 43560 -680
rect 43575 -500 43645 -490
rect 43575 -530 43595 -500
rect 43625 -530 43645 -500
rect 43575 -550 43645 -530
rect 43575 -580 43595 -550
rect 43625 -580 43645 -550
rect 43575 -600 43645 -580
rect 43575 -630 43595 -600
rect 43625 -630 43645 -600
rect 43575 -650 43645 -630
rect 43575 -680 43595 -650
rect 43625 -680 43645 -650
rect 43575 -690 43645 -680
<< ndiffc >>
rect 225 10 255 40
rect 310 10 340 40
rect 395 10 425 40
rect 480 10 510 40
rect 565 10 595 40
rect 760 10 790 40
rect 845 10 875 40
rect 930 10 960 40
rect 1015 10 1045 40
rect 1100 10 1130 40
rect 1185 10 1215 40
rect 1270 10 1300 40
rect 1355 10 1385 40
rect 1440 10 1470 40
rect 1525 10 1555 40
rect 1610 10 1640 40
rect 1695 10 1725 40
rect 1780 10 1810 40
rect 1865 10 1895 40
rect 1950 10 1980 40
rect 2035 10 2065 40
rect 2120 10 2150 40
rect 2270 10 2300 40
rect 2355 10 2385 40
rect 2440 10 2470 40
rect 2525 10 2555 40
rect 2610 10 2640 40
rect 2695 10 2725 40
rect 2780 10 2810 40
rect 2865 10 2895 40
rect 2950 10 2980 40
rect 3035 10 3065 40
rect 3120 10 3150 40
rect 3205 10 3235 40
rect 3290 10 3320 40
rect 3375 10 3405 40
rect 3460 10 3490 40
rect 3545 10 3575 40
rect 3630 10 3660 40
rect 3715 10 3745 40
rect 3800 10 3830 40
rect 3885 10 3915 40
rect 3970 10 4000 40
rect 4055 10 4085 40
rect 4140 10 4170 40
rect 4225 10 4255 40
rect 4310 10 4340 40
rect 4395 10 4425 40
rect 4480 10 4510 40
rect 4565 10 4595 40
rect 4650 10 4680 40
rect 4735 10 4765 40
rect 4820 10 4850 40
rect 4905 10 4935 40
rect 4990 10 5020 40
rect 5075 10 5105 40
rect 5160 10 5190 40
rect 5245 10 5275 40
rect 5330 10 5360 40
rect 5415 10 5445 40
rect 5500 10 5530 40
rect 5585 10 5615 40
rect 5670 10 5700 40
rect 5755 10 5785 40
rect 5840 10 5870 40
rect 5925 10 5955 40
rect 6010 10 6040 40
rect 6095 10 6125 40
rect 6180 10 6210 40
rect 6265 10 6295 40
rect 6350 10 6380 40
rect 6435 10 6465 40
rect 6520 10 6550 40
rect 6605 10 6635 40
rect 6690 10 6720 40
rect 6775 10 6805 40
rect 6860 10 6890 40
rect 6945 10 6975 40
rect 7030 10 7060 40
rect 7115 10 7145 40
rect 7200 10 7230 40
rect 7285 10 7315 40
rect 7370 10 7400 40
rect 7455 10 7485 40
rect 7540 10 7570 40
rect 7625 10 7655 40
rect 7710 10 7740 40
rect 7860 10 7890 40
rect 7945 10 7975 40
rect 8030 10 8060 40
rect 8115 10 8145 40
rect 8200 10 8230 40
rect 8285 10 8315 40
rect 8370 10 8400 40
rect 8455 10 8485 40
rect 8540 10 8570 40
rect 8625 10 8655 40
rect 8710 10 8740 40
rect 8795 10 8825 40
rect 8880 10 8910 40
rect 8965 10 8995 40
rect 9050 10 9080 40
rect 9135 10 9165 40
rect 9220 10 9250 40
rect 9305 10 9335 40
rect 9390 10 9420 40
rect 9475 10 9505 40
rect 9560 10 9590 40
rect 9645 10 9675 40
rect 9730 10 9760 40
rect 9815 10 9845 40
rect 9900 10 9930 40
rect 9985 10 10015 40
rect 10070 10 10100 40
rect 10155 10 10185 40
rect 10240 10 10270 40
rect 10325 10 10355 40
rect 10410 10 10440 40
rect 10495 10 10525 40
rect 10580 10 10610 40
rect 10665 10 10695 40
rect 10750 10 10780 40
rect 10835 10 10865 40
rect 10920 10 10950 40
rect 11005 10 11035 40
rect 11090 10 11120 40
rect 11175 10 11205 40
rect 11260 10 11290 40
rect 11345 10 11375 40
rect 11430 10 11460 40
rect 11515 10 11545 40
rect 11600 10 11630 40
rect 11685 10 11715 40
rect 11770 10 11800 40
rect 11855 10 11885 40
rect 11940 10 11970 40
rect 12025 10 12055 40
rect 12110 10 12140 40
rect 12195 10 12225 40
rect 12280 10 12310 40
rect 12365 10 12395 40
rect 12450 10 12480 40
rect 12535 10 12565 40
rect 12620 10 12650 40
rect 12705 10 12735 40
rect 12790 10 12820 40
rect 12875 10 12905 40
rect 12960 10 12990 40
rect 13045 10 13075 40
rect 13130 10 13160 40
rect 13215 10 13245 40
rect 13300 10 13330 40
rect 13385 10 13415 40
rect 13470 10 13500 40
rect 13555 10 13585 40
rect 13640 10 13670 40
rect 13725 10 13755 40
rect 13810 10 13840 40
rect 13895 10 13925 40
rect 13980 10 14010 40
rect 14065 10 14095 40
rect 14150 10 14180 40
rect 14235 10 14265 40
rect 14320 10 14350 40
rect 14405 10 14435 40
rect 14490 10 14520 40
rect 14575 10 14605 40
rect 14660 10 14690 40
rect 14745 10 14775 40
rect 14830 10 14860 40
rect 14915 10 14945 40
rect 15000 10 15030 40
rect 15085 10 15115 40
rect 15170 10 15200 40
rect 15255 10 15285 40
rect 15340 10 15370 40
rect 15425 10 15455 40
rect 15510 10 15540 40
rect 15595 10 15625 40
rect 15680 10 15710 40
rect 15765 10 15795 40
rect 15850 10 15880 40
rect 15935 10 15965 40
rect 16020 10 16050 40
rect 16105 10 16135 40
rect 16190 10 16220 40
rect 16275 10 16305 40
rect 16360 10 16390 40
rect 16445 10 16475 40
rect 16530 10 16560 40
rect 16615 10 16645 40
rect 16700 10 16730 40
rect 16785 10 16815 40
rect 16870 10 16900 40
rect 16955 10 16985 40
rect 17040 10 17070 40
rect 17125 10 17155 40
rect 17210 10 17240 40
rect 17295 10 17325 40
rect 17380 10 17410 40
rect 17465 10 17495 40
rect 17550 10 17580 40
rect 17635 10 17665 40
rect 17720 10 17750 40
rect 17805 10 17835 40
rect 17890 10 17920 40
rect 17975 10 18005 40
rect 18060 10 18090 40
rect 18145 10 18175 40
rect 18230 10 18260 40
rect 18315 10 18345 40
rect 18400 10 18430 40
rect 18485 10 18515 40
rect 18570 10 18600 40
rect 18655 10 18685 40
rect 18740 10 18770 40
rect 18825 10 18855 40
rect 18910 10 18940 40
rect 18995 10 19025 40
rect 19080 10 19110 40
rect 19165 10 19195 40
rect 19250 10 19280 40
rect 19335 10 19365 40
rect 19420 10 19450 40
rect 19505 10 19535 40
rect 19590 10 19620 40
rect 19675 10 19705 40
rect 19760 10 19790 40
rect 19845 10 19875 40
rect 19930 10 19960 40
rect 20015 10 20045 40
rect 20100 10 20130 40
rect 20185 10 20215 40
rect 20270 10 20300 40
rect 20355 10 20385 40
rect 20440 10 20470 40
rect 20525 10 20555 40
rect 20610 10 20640 40
rect 20695 10 20725 40
rect 20780 10 20810 40
rect 20865 10 20895 40
rect 20950 10 20980 40
rect 21035 10 21065 40
rect 21120 10 21150 40
rect 21205 10 21235 40
rect 21290 10 21320 40
rect 21375 10 21405 40
rect 21460 10 21490 40
rect 21545 10 21575 40
rect 21630 10 21660 40
rect 21715 10 21745 40
rect 21800 10 21830 40
rect 21885 10 21915 40
rect 21970 10 22000 40
rect 22055 10 22085 40
rect 22140 10 22170 40
rect 22225 10 22255 40
rect 22310 10 22340 40
rect 22395 10 22425 40
rect 22480 10 22510 40
rect 22565 10 22595 40
rect 22650 10 22680 40
rect 22735 10 22765 40
rect 22820 10 22850 40
rect 22905 10 22935 40
rect 22990 10 23020 40
rect 23075 10 23105 40
rect 23160 10 23190 40
rect 23245 10 23275 40
rect 23330 10 23360 40
rect 23415 10 23445 40
rect 23500 10 23530 40
rect 23585 10 23615 40
rect 23670 10 23700 40
rect 23755 10 23785 40
rect 23840 10 23870 40
rect 23925 10 23955 40
rect 24010 10 24040 40
rect 24095 10 24125 40
rect 24180 10 24210 40
rect 24265 10 24295 40
rect 24350 10 24380 40
rect 24435 10 24465 40
rect 24520 10 24550 40
rect 24605 10 24635 40
rect 24690 10 24720 40
rect 24775 10 24805 40
rect 24860 10 24890 40
rect 24945 10 24975 40
rect 25030 10 25060 40
rect 25115 10 25145 40
rect 25200 10 25230 40
rect 25285 10 25315 40
rect 25370 10 25400 40
rect 25455 10 25485 40
rect 25540 10 25570 40
rect 25625 10 25655 40
rect 25710 10 25740 40
rect 25795 10 25825 40
rect 25880 10 25910 40
rect 25965 10 25995 40
rect 26050 10 26080 40
rect 26135 10 26165 40
rect 26220 10 26250 40
rect 26305 10 26335 40
rect 26390 10 26420 40
rect 26475 10 26505 40
rect 26560 10 26590 40
rect 26645 10 26675 40
rect 26730 10 26760 40
rect 26815 10 26845 40
rect 26900 10 26930 40
rect 26985 10 27015 40
rect 27070 10 27100 40
rect 27155 10 27185 40
rect 27240 10 27270 40
rect 27325 10 27355 40
rect 27410 10 27440 40
rect 27495 10 27525 40
rect 27580 10 27610 40
rect 27665 10 27695 40
rect 27750 10 27780 40
rect 27835 10 27865 40
rect 27920 10 27950 40
rect 28005 10 28035 40
rect 28090 10 28120 40
rect 28175 10 28205 40
rect 28260 10 28290 40
rect 28345 10 28375 40
rect 28430 10 28460 40
rect 28515 10 28545 40
rect 28600 10 28630 40
rect 28685 10 28715 40
rect 28770 10 28800 40
rect 28855 10 28885 40
rect 28940 10 28970 40
rect 29025 10 29055 40
rect 29110 10 29140 40
rect 29195 10 29225 40
rect 29280 10 29310 40
rect 29365 10 29395 40
rect 29450 10 29480 40
rect 29535 10 29565 40
rect 29620 10 29650 40
rect 15 -60 45 -30
rect 100 -60 130 -30
rect 75 -365 105 -335
rect 75 -415 105 -385
rect 160 -365 190 -335
rect 160 -415 190 -385
rect 245 -365 275 -335
rect 245 -415 275 -385
rect 330 -365 360 -335
rect 330 -415 360 -385
rect 415 -365 445 -335
rect 415 -415 445 -385
rect 500 -365 530 -335
rect 500 -415 530 -385
rect 585 -365 615 -335
rect 585 -415 615 -385
rect 670 -365 700 -335
rect 670 -415 700 -385
rect 755 -365 785 -335
rect 755 -415 785 -385
rect 840 -365 870 -335
rect 840 -415 870 -385
rect 925 -365 955 -335
rect 925 -415 955 -385
rect 1010 -365 1040 -335
rect 1010 -415 1040 -385
rect 1095 -365 1125 -335
rect 1095 -415 1125 -385
rect 1180 -365 1210 -335
rect 1180 -415 1210 -385
rect 1265 -365 1295 -335
rect 1265 -415 1295 -385
rect 1350 -365 1380 -335
rect 1350 -415 1380 -385
rect 1435 -365 1465 -335
rect 1435 -415 1465 -385
rect 1520 -365 1550 -335
rect 1520 -415 1550 -385
rect 1605 -365 1635 -335
rect 1605 -415 1635 -385
rect 1690 -365 1720 -335
rect 1690 -415 1720 -385
rect 1775 -365 1805 -335
rect 1775 -415 1805 -385
rect 1860 -365 1890 -335
rect 1860 -415 1890 -385
rect 1945 -365 1975 -335
rect 1945 -415 1975 -385
rect 2030 -365 2060 -335
rect 2030 -415 2060 -385
rect 2115 -365 2145 -335
rect 2115 -415 2145 -385
rect 2200 -365 2230 -335
rect 2200 -415 2230 -385
rect 2285 -365 2315 -335
rect 2285 -415 2315 -385
rect 2370 -365 2400 -335
rect 2370 -415 2400 -385
rect 2455 -365 2485 -335
rect 2455 -415 2485 -385
rect 2540 -365 2570 -335
rect 2540 -415 2570 -385
rect 2625 -365 2655 -335
rect 2625 -415 2655 -385
rect 2710 -365 2740 -335
rect 2710 -415 2740 -385
rect 2795 -365 2825 -335
rect 2795 -415 2825 -385
rect 2880 -365 2910 -335
rect 2880 -415 2910 -385
rect 2965 -365 2995 -335
rect 2965 -415 2995 -385
rect 3050 -365 3080 -335
rect 3050 -415 3080 -385
rect 3135 -365 3165 -335
rect 3135 -415 3165 -385
rect 3220 -365 3250 -335
rect 3220 -415 3250 -385
rect 3305 -365 3335 -335
rect 3305 -415 3335 -385
rect 3390 -365 3420 -335
rect 3390 -415 3420 -385
rect 3475 -365 3505 -335
rect 3475 -415 3505 -385
rect 3560 -365 3590 -335
rect 3560 -415 3590 -385
rect 3645 -365 3675 -335
rect 3645 -415 3675 -385
rect 3730 -365 3760 -335
rect 3730 -415 3760 -385
rect 3815 -365 3845 -335
rect 3815 -415 3845 -385
rect 3900 -365 3930 -335
rect 3900 -415 3930 -385
rect 3985 -365 4015 -335
rect 3985 -415 4015 -385
rect 4070 -365 4100 -335
rect 4070 -415 4100 -385
rect 4155 -365 4185 -335
rect 4155 -415 4185 -385
rect 4240 -365 4270 -335
rect 4240 -415 4270 -385
rect 4325 -365 4355 -335
rect 4325 -415 4355 -385
rect 4410 -365 4440 -335
rect 4410 -415 4440 -385
rect 4495 -365 4525 -335
rect 4495 -415 4525 -385
rect 4580 -365 4610 -335
rect 4580 -415 4610 -385
rect 4665 -365 4695 -335
rect 4665 -415 4695 -385
rect 4750 -365 4780 -335
rect 4750 -415 4780 -385
rect 4835 -365 4865 -335
rect 4835 -415 4865 -385
rect 4920 -365 4950 -335
rect 4920 -415 4950 -385
rect 5005 -365 5035 -335
rect 5005 -415 5035 -385
rect 5090 -365 5120 -335
rect 5090 -415 5120 -385
rect 5175 -365 5205 -335
rect 5175 -415 5205 -385
rect 5260 -365 5290 -335
rect 5260 -415 5290 -385
rect 5345 -365 5375 -335
rect 5345 -415 5375 -385
rect 5430 -365 5460 -335
rect 5430 -415 5460 -385
rect 5515 -365 5545 -335
rect 5515 -415 5545 -385
rect 5600 -365 5630 -335
rect 5600 -415 5630 -385
rect 5685 -365 5715 -335
rect 5685 -415 5715 -385
rect 5770 -365 5800 -335
rect 5770 -415 5800 -385
rect 5855 -365 5885 -335
rect 5855 -415 5885 -385
rect 5940 -365 5970 -335
rect 5940 -415 5970 -385
rect 6025 -365 6055 -335
rect 6025 -415 6055 -385
rect 6110 -365 6140 -335
rect 6110 -415 6140 -385
rect 6195 -365 6225 -335
rect 6195 -415 6225 -385
rect 6280 -365 6310 -335
rect 6280 -415 6310 -385
rect 6365 -365 6395 -335
rect 6365 -415 6395 -385
rect 6450 -365 6480 -335
rect 6450 -415 6480 -385
rect 6535 -365 6565 -335
rect 6535 -415 6565 -385
rect 6620 -365 6650 -335
rect 6620 -415 6650 -385
rect 6705 -365 6735 -335
rect 6705 -415 6735 -385
rect 6790 -365 6820 -335
rect 6790 -415 6820 -385
rect 6875 -365 6905 -335
rect 6875 -415 6905 -385
rect 6960 -365 6990 -335
rect 6960 -415 6990 -385
rect 7045 -365 7075 -335
rect 7045 -415 7075 -385
rect 7130 -365 7160 -335
rect 7130 -415 7160 -385
rect 7215 -365 7245 -335
rect 7215 -415 7245 -385
rect 7300 -365 7330 -335
rect 7300 -415 7330 -385
rect 7385 -365 7415 -335
rect 7385 -415 7415 -385
rect 7470 -365 7500 -335
rect 7470 -415 7500 -385
rect 7555 -365 7585 -335
rect 7555 -415 7585 -385
rect 7640 -365 7670 -335
rect 7640 -415 7670 -385
rect 7725 -365 7755 -335
rect 7725 -415 7755 -385
rect 7810 -365 7840 -335
rect 7810 -415 7840 -385
rect 7895 -365 7925 -335
rect 7895 -415 7925 -385
rect 7980 -365 8010 -335
rect 7980 -415 8010 -385
rect 8065 -365 8095 -335
rect 8065 -415 8095 -385
rect 8150 -365 8180 -335
rect 8150 -415 8180 -385
rect 8235 -365 8265 -335
rect 8235 -415 8265 -385
rect 8320 -365 8350 -335
rect 8320 -415 8350 -385
rect 8405 -365 8435 -335
rect 8405 -415 8435 -385
rect 8490 -365 8520 -335
rect 8490 -415 8520 -385
rect 8575 -365 8605 -335
rect 8575 -415 8605 -385
rect 8660 -365 8690 -335
rect 8660 -415 8690 -385
rect 8745 -365 8775 -335
rect 8745 -415 8775 -385
rect 8830 -365 8860 -335
rect 8830 -415 8860 -385
rect 8915 -365 8945 -335
rect 8915 -415 8945 -385
rect 9000 -365 9030 -335
rect 9000 -415 9030 -385
rect 9085 -365 9115 -335
rect 9085 -415 9115 -385
rect 9170 -365 9200 -335
rect 9170 -415 9200 -385
rect 9255 -365 9285 -335
rect 9255 -415 9285 -385
rect 9340 -365 9370 -335
rect 9340 -415 9370 -385
rect 9425 -365 9455 -335
rect 9425 -415 9455 -385
rect 9510 -365 9540 -335
rect 9510 -415 9540 -385
rect 9595 -365 9625 -335
rect 9595 -415 9625 -385
rect 9680 -365 9710 -335
rect 9680 -415 9710 -385
rect 9765 -365 9795 -335
rect 9765 -415 9795 -385
rect 9850 -365 9880 -335
rect 9850 -415 9880 -385
rect 9935 -365 9965 -335
rect 9935 -415 9965 -385
rect 10020 -365 10050 -335
rect 10020 -415 10050 -385
rect 10105 -365 10135 -335
rect 10105 -415 10135 -385
rect 10190 -365 10220 -335
rect 10190 -415 10220 -385
rect 10275 -365 10305 -335
rect 10275 -415 10305 -385
rect 10360 -365 10390 -335
rect 10360 -415 10390 -385
rect 10445 -365 10475 -335
rect 10445 -415 10475 -385
rect 10530 -365 10560 -335
rect 10530 -415 10560 -385
rect 10615 -365 10645 -335
rect 10615 -415 10645 -385
rect 10700 -365 10730 -335
rect 10700 -415 10730 -385
rect 10785 -365 10815 -335
rect 10785 -415 10815 -385
rect 10870 -365 10900 -335
rect 10870 -415 10900 -385
rect 10955 -365 10985 -335
rect 10955 -415 10985 -385
rect 11040 -365 11070 -335
rect 11040 -415 11070 -385
rect 11125 -365 11155 -335
rect 11125 -415 11155 -385
rect 11210 -365 11240 -335
rect 11210 -415 11240 -385
rect 11295 -365 11325 -335
rect 11295 -415 11325 -385
rect 11380 -365 11410 -335
rect 11380 -415 11410 -385
rect 11465 -365 11495 -335
rect 11465 -415 11495 -385
rect 11550 -365 11580 -335
rect 11550 -415 11580 -385
rect 11635 -365 11665 -335
rect 11635 -415 11665 -385
rect 11720 -365 11750 -335
rect 11720 -415 11750 -385
rect 11805 -365 11835 -335
rect 11805 -415 11835 -385
rect 11890 -365 11920 -335
rect 11890 -415 11920 -385
rect 11975 -365 12005 -335
rect 11975 -415 12005 -385
rect 12060 -365 12090 -335
rect 12060 -415 12090 -385
rect 12145 -365 12175 -335
rect 12145 -415 12175 -385
rect 12230 -365 12260 -335
rect 12230 -415 12260 -385
rect 12315 -365 12345 -335
rect 12315 -415 12345 -385
rect 12400 -365 12430 -335
rect 12400 -415 12430 -385
rect 12485 -365 12515 -335
rect 12485 -415 12515 -385
rect 12570 -365 12600 -335
rect 12570 -415 12600 -385
rect 12655 -365 12685 -335
rect 12655 -415 12685 -385
rect 12740 -365 12770 -335
rect 12740 -415 12770 -385
rect 12825 -365 12855 -335
rect 12825 -415 12855 -385
rect 12910 -365 12940 -335
rect 12910 -415 12940 -385
rect 12995 -365 13025 -335
rect 12995 -415 13025 -385
rect 13080 -365 13110 -335
rect 13080 -415 13110 -385
rect 13165 -365 13195 -335
rect 13165 -415 13195 -385
rect 13250 -365 13280 -335
rect 13250 -415 13280 -385
rect 13335 -365 13365 -335
rect 13335 -415 13365 -385
rect 13420 -365 13450 -335
rect 13420 -415 13450 -385
rect 13505 -365 13535 -335
rect 13505 -415 13535 -385
rect 13590 -365 13620 -335
rect 13590 -415 13620 -385
rect 13675 -365 13705 -335
rect 13675 -415 13705 -385
rect 13760 -365 13790 -335
rect 13760 -415 13790 -385
rect 13845 -365 13875 -335
rect 13845 -415 13875 -385
rect 13930 -365 13960 -335
rect 13930 -415 13960 -385
rect 14015 -365 14045 -335
rect 14015 -415 14045 -385
rect 14100 -365 14130 -335
rect 14100 -415 14130 -385
rect 14185 -365 14215 -335
rect 14185 -415 14215 -385
rect 14270 -365 14300 -335
rect 14270 -415 14300 -385
rect 14355 -365 14385 -335
rect 14355 -415 14385 -385
rect 14440 -365 14470 -335
rect 14440 -415 14470 -385
rect 14525 -365 14555 -335
rect 14525 -415 14555 -385
rect 14610 -365 14640 -335
rect 14610 -415 14640 -385
rect 14695 -365 14725 -335
rect 14695 -415 14725 -385
rect 14780 -365 14810 -335
rect 14780 -415 14810 -385
rect 14865 -365 14895 -335
rect 14865 -415 14895 -385
rect 14950 -365 14980 -335
rect 14950 -415 14980 -385
rect 15035 -365 15065 -335
rect 15035 -415 15065 -385
rect 15120 -365 15150 -335
rect 15120 -415 15150 -385
rect 15205 -365 15235 -335
rect 15205 -415 15235 -385
rect 15290 -365 15320 -335
rect 15290 -415 15320 -385
rect 15375 -365 15405 -335
rect 15375 -415 15405 -385
rect 15460 -365 15490 -335
rect 15460 -415 15490 -385
rect 15545 -365 15575 -335
rect 15545 -415 15575 -385
rect 15630 -365 15660 -335
rect 15630 -415 15660 -385
rect 15715 -365 15745 -335
rect 15715 -415 15745 -385
rect 15800 -365 15830 -335
rect 15800 -415 15830 -385
rect 15885 -365 15915 -335
rect 15885 -415 15915 -385
rect 15970 -365 16000 -335
rect 15970 -415 16000 -385
rect 16055 -365 16085 -335
rect 16055 -415 16085 -385
rect 16140 -365 16170 -335
rect 16140 -415 16170 -385
rect 16225 -365 16255 -335
rect 16225 -415 16255 -385
rect 16310 -365 16340 -335
rect 16310 -415 16340 -385
rect 16395 -365 16425 -335
rect 16395 -415 16425 -385
rect 16480 -365 16510 -335
rect 16480 -415 16510 -385
rect 16565 -365 16595 -335
rect 16565 -415 16595 -385
rect 16650 -365 16680 -335
rect 16650 -415 16680 -385
rect 16735 -365 16765 -335
rect 16735 -415 16765 -385
rect 16820 -365 16850 -335
rect 16820 -415 16850 -385
rect 16905 -365 16935 -335
rect 16905 -415 16935 -385
rect 16990 -365 17020 -335
rect 16990 -415 17020 -385
rect 17075 -365 17105 -335
rect 17075 -415 17105 -385
rect 17160 -365 17190 -335
rect 17160 -415 17190 -385
rect 17245 -365 17275 -335
rect 17245 -415 17275 -385
rect 17330 -365 17360 -335
rect 17330 -415 17360 -385
rect 17415 -365 17445 -335
rect 17415 -415 17445 -385
rect 17500 -365 17530 -335
rect 17500 -415 17530 -385
rect 17585 -365 17615 -335
rect 17585 -415 17615 -385
rect 17670 -365 17700 -335
rect 17670 -415 17700 -385
rect 17755 -365 17785 -335
rect 17755 -415 17785 -385
rect 17840 -365 17870 -335
rect 17840 -415 17870 -385
rect 17925 -365 17955 -335
rect 17925 -415 17955 -385
rect 18010 -365 18040 -335
rect 18010 -415 18040 -385
rect 18095 -365 18125 -335
rect 18095 -415 18125 -385
rect 18180 -365 18210 -335
rect 18180 -415 18210 -385
rect 18265 -365 18295 -335
rect 18265 -415 18295 -385
rect 18350 -365 18380 -335
rect 18350 -415 18380 -385
rect 18435 -365 18465 -335
rect 18435 -415 18465 -385
rect 18520 -365 18550 -335
rect 18520 -415 18550 -385
rect 18605 -365 18635 -335
rect 18605 -415 18635 -385
rect 18690 -365 18720 -335
rect 18690 -415 18720 -385
rect 18775 -365 18805 -335
rect 18775 -415 18805 -385
rect 18860 -365 18890 -335
rect 18860 -415 18890 -385
rect 18945 -365 18975 -335
rect 18945 -415 18975 -385
rect 19030 -365 19060 -335
rect 19030 -415 19060 -385
rect 19115 -365 19145 -335
rect 19115 -415 19145 -385
rect 19200 -365 19230 -335
rect 19200 -415 19230 -385
rect 19285 -365 19315 -335
rect 19285 -415 19315 -385
rect 19370 -365 19400 -335
rect 19370 -415 19400 -385
rect 19455 -365 19485 -335
rect 19455 -415 19485 -385
rect 19540 -365 19570 -335
rect 19540 -415 19570 -385
rect 19625 -365 19655 -335
rect 19625 -415 19655 -385
rect 19710 -365 19740 -335
rect 19710 -415 19740 -385
rect 19795 -365 19825 -335
rect 19795 -415 19825 -385
rect 19880 -365 19910 -335
rect 19880 -415 19910 -385
rect 19965 -365 19995 -335
rect 19965 -415 19995 -385
rect 20050 -365 20080 -335
rect 20050 -415 20080 -385
rect 20135 -365 20165 -335
rect 20135 -415 20165 -385
rect 20220 -365 20250 -335
rect 20220 -415 20250 -385
rect 20305 -365 20335 -335
rect 20305 -415 20335 -385
rect 20390 -365 20420 -335
rect 20390 -415 20420 -385
rect 20475 -365 20505 -335
rect 20475 -415 20505 -385
rect 20560 -365 20590 -335
rect 20560 -415 20590 -385
rect 20645 -365 20675 -335
rect 20645 -415 20675 -385
rect 20730 -365 20760 -335
rect 20730 -415 20760 -385
rect 20815 -365 20845 -335
rect 20815 -415 20845 -385
rect 20900 -365 20930 -335
rect 20900 -415 20930 -385
rect 20985 -365 21015 -335
rect 20985 -415 21015 -385
rect 21070 -365 21100 -335
rect 21070 -415 21100 -385
rect 21155 -365 21185 -335
rect 21155 -415 21185 -385
rect 21240 -365 21270 -335
rect 21240 -415 21270 -385
rect 21325 -365 21355 -335
rect 21325 -415 21355 -385
rect 21410 -365 21440 -335
rect 21410 -415 21440 -385
rect 21495 -365 21525 -335
rect 21495 -415 21525 -385
rect 21580 -365 21610 -335
rect 21580 -415 21610 -385
rect 21665 -365 21695 -335
rect 21665 -415 21695 -385
rect 21750 -365 21780 -335
rect 21750 -415 21780 -385
rect 21835 -365 21865 -335
rect 21835 -415 21865 -385
rect 21920 -365 21950 -335
rect 21920 -415 21950 -385
rect 22005 -365 22035 -335
rect 22005 -415 22035 -385
rect 22090 -365 22120 -335
rect 22090 -415 22120 -385
rect 22175 -365 22205 -335
rect 22175 -415 22205 -385
rect 22260 -365 22290 -335
rect 22260 -415 22290 -385
rect 22345 -365 22375 -335
rect 22345 -415 22375 -385
rect 22430 -365 22460 -335
rect 22430 -415 22460 -385
rect 22515 -365 22545 -335
rect 22515 -415 22545 -385
rect 22600 -365 22630 -335
rect 22600 -415 22630 -385
rect 22685 -365 22715 -335
rect 22685 -415 22715 -385
rect 22770 -365 22800 -335
rect 22770 -415 22800 -385
rect 22855 -365 22885 -335
rect 22855 -415 22885 -385
rect 22940 -365 22970 -335
rect 22940 -415 22970 -385
rect 23025 -365 23055 -335
rect 23025 -415 23055 -385
rect 23110 -365 23140 -335
rect 23110 -415 23140 -385
rect 23195 -365 23225 -335
rect 23195 -415 23225 -385
rect 23280 -365 23310 -335
rect 23280 -415 23310 -385
rect 23365 -365 23395 -335
rect 23365 -415 23395 -385
rect 23450 -365 23480 -335
rect 23450 -415 23480 -385
rect 23535 -365 23565 -335
rect 23535 -415 23565 -385
rect 23620 -365 23650 -335
rect 23620 -415 23650 -385
rect 23705 -365 23735 -335
rect 23705 -415 23735 -385
rect 23790 -365 23820 -335
rect 23790 -415 23820 -385
rect 23875 -365 23905 -335
rect 23875 -415 23905 -385
rect 23960 -365 23990 -335
rect 23960 -415 23990 -385
rect 24045 -365 24075 -335
rect 24045 -415 24075 -385
rect 24130 -365 24160 -335
rect 24130 -415 24160 -385
rect 24215 -365 24245 -335
rect 24215 -415 24245 -385
rect 24300 -365 24330 -335
rect 24300 -415 24330 -385
rect 24385 -365 24415 -335
rect 24385 -415 24415 -385
rect 24470 -365 24500 -335
rect 24470 -415 24500 -385
rect 24555 -365 24585 -335
rect 24555 -415 24585 -385
rect 24640 -365 24670 -335
rect 24640 -415 24670 -385
rect 24725 -365 24755 -335
rect 24725 -415 24755 -385
rect 24810 -365 24840 -335
rect 24810 -415 24840 -385
rect 24895 -365 24925 -335
rect 24895 -415 24925 -385
rect 24980 -365 25010 -335
rect 24980 -415 25010 -385
rect 25065 -365 25095 -335
rect 25065 -415 25095 -385
rect 25150 -365 25180 -335
rect 25150 -415 25180 -385
rect 25235 -365 25265 -335
rect 25235 -415 25265 -385
rect 25320 -365 25350 -335
rect 25320 -415 25350 -385
rect 25405 -365 25435 -335
rect 25405 -415 25435 -385
rect 25490 -365 25520 -335
rect 25490 -415 25520 -385
rect 25575 -365 25605 -335
rect 25575 -415 25605 -385
rect 25660 -365 25690 -335
rect 25660 -415 25690 -385
rect 25745 -365 25775 -335
rect 25745 -415 25775 -385
rect 25830 -365 25860 -335
rect 25830 -415 25860 -385
rect 25915 -365 25945 -335
rect 25915 -415 25945 -385
rect 26000 -365 26030 -335
rect 26000 -415 26030 -385
rect 26085 -365 26115 -335
rect 26085 -415 26115 -385
rect 26170 -365 26200 -335
rect 26170 -415 26200 -385
rect 26255 -365 26285 -335
rect 26255 -415 26285 -385
rect 26340 -365 26370 -335
rect 26340 -415 26370 -385
rect 26425 -365 26455 -335
rect 26425 -415 26455 -385
rect 26510 -365 26540 -335
rect 26510 -415 26540 -385
rect 26595 -365 26625 -335
rect 26595 -415 26625 -385
rect 26680 -365 26710 -335
rect 26680 -415 26710 -385
rect 26765 -365 26795 -335
rect 26765 -415 26795 -385
rect 26850 -365 26880 -335
rect 26850 -415 26880 -385
rect 26935 -365 26965 -335
rect 26935 -415 26965 -385
rect 27020 -365 27050 -335
rect 27020 -415 27050 -385
rect 27105 -365 27135 -335
rect 27105 -415 27135 -385
rect 27190 -365 27220 -335
rect 27190 -415 27220 -385
rect 27275 -365 27305 -335
rect 27275 -415 27305 -385
rect 27360 -365 27390 -335
rect 27360 -415 27390 -385
rect 27445 -365 27475 -335
rect 27445 -415 27475 -385
rect 27530 -365 27560 -335
rect 27530 -415 27560 -385
rect 27615 -365 27645 -335
rect 27615 -415 27645 -385
rect 27700 -365 27730 -335
rect 27700 -415 27730 -385
rect 27785 -365 27815 -335
rect 27785 -415 27815 -385
rect 27870 -365 27900 -335
rect 27870 -415 27900 -385
rect 27955 -365 27985 -335
rect 27955 -415 27985 -385
rect 28040 -365 28070 -335
rect 28040 -415 28070 -385
rect 28125 -365 28155 -335
rect 28125 -415 28155 -385
rect 28210 -365 28240 -335
rect 28210 -415 28240 -385
rect 28295 -365 28325 -335
rect 28295 -415 28325 -385
rect 28380 -365 28410 -335
rect 28380 -415 28410 -385
rect 28465 -365 28495 -335
rect 28465 -415 28495 -385
rect 28550 -365 28580 -335
rect 28550 -415 28580 -385
rect 28635 -365 28665 -335
rect 28635 -415 28665 -385
rect 28720 -365 28750 -335
rect 28720 -415 28750 -385
rect 28805 -365 28835 -335
rect 28805 -415 28835 -385
rect 28890 -365 28920 -335
rect 28890 -415 28920 -385
rect 28975 -365 29005 -335
rect 28975 -415 29005 -385
rect 29060 -365 29090 -335
rect 29060 -415 29090 -385
rect 29145 -365 29175 -335
rect 29145 -415 29175 -385
rect 29230 -365 29260 -335
rect 29230 -415 29260 -385
rect 29315 -365 29345 -335
rect 29315 -415 29345 -385
rect 29400 -365 29430 -335
rect 29400 -415 29430 -385
rect 29485 -365 29515 -335
rect 29485 -415 29515 -385
rect 29570 -365 29600 -335
rect 29570 -415 29600 -385
rect 29655 -365 29685 -335
rect 29655 -415 29685 -385
rect 29740 -365 29770 -335
rect 29740 -415 29770 -385
rect 29825 -365 29855 -335
rect 29825 -415 29855 -385
rect 29910 -365 29940 -335
rect 29910 -415 29940 -385
rect 29995 -365 30025 -335
rect 29995 -415 30025 -385
rect 30080 -365 30110 -335
rect 30080 -415 30110 -385
rect 30165 -365 30195 -335
rect 30165 -415 30195 -385
rect 30250 -365 30280 -335
rect 30250 -415 30280 -385
rect 30335 -365 30365 -335
rect 30335 -415 30365 -385
rect 30420 -365 30450 -335
rect 30420 -415 30450 -385
rect 30505 -365 30535 -335
rect 30505 -415 30535 -385
rect 30590 -365 30620 -335
rect 30590 -415 30620 -385
rect 30675 -365 30705 -335
rect 30675 -415 30705 -385
rect 30760 -365 30790 -335
rect 30760 -415 30790 -385
rect 30845 -365 30875 -335
rect 30845 -415 30875 -385
rect 30930 -365 30960 -335
rect 30930 -415 30960 -385
rect 31015 -365 31045 -335
rect 31015 -415 31045 -385
rect 31100 -365 31130 -335
rect 31100 -415 31130 -385
rect 31185 -365 31215 -335
rect 31185 -415 31215 -385
rect 31270 -365 31300 -335
rect 31270 -415 31300 -385
rect 31355 -365 31385 -335
rect 31355 -415 31385 -385
rect 31440 -365 31470 -335
rect 31440 -415 31470 -385
rect 31525 -365 31555 -335
rect 31525 -415 31555 -385
rect 31610 -365 31640 -335
rect 31610 -415 31640 -385
rect 31695 -365 31725 -335
rect 31695 -415 31725 -385
rect 31780 -365 31810 -335
rect 31780 -415 31810 -385
rect 31865 -365 31895 -335
rect 31865 -415 31895 -385
rect 31950 -365 31980 -335
rect 31950 -415 31980 -385
rect 32035 -365 32065 -335
rect 32035 -415 32065 -385
rect 32120 -365 32150 -335
rect 32120 -415 32150 -385
rect 32205 -365 32235 -335
rect 32205 -415 32235 -385
rect 32290 -365 32320 -335
rect 32290 -415 32320 -385
rect 32375 -365 32405 -335
rect 32375 -415 32405 -385
rect 32460 -365 32490 -335
rect 32460 -415 32490 -385
rect 32545 -365 32575 -335
rect 32545 -415 32575 -385
rect 32630 -365 32660 -335
rect 32630 -415 32660 -385
rect 32715 -365 32745 -335
rect 32715 -415 32745 -385
rect 32800 -365 32830 -335
rect 32800 -415 32830 -385
rect 32885 -365 32915 -335
rect 32885 -415 32915 -385
rect 32970 -365 33000 -335
rect 32970 -415 33000 -385
rect 33055 -365 33085 -335
rect 33055 -415 33085 -385
rect 33140 -365 33170 -335
rect 33140 -415 33170 -385
rect 33225 -365 33255 -335
rect 33225 -415 33255 -385
rect 33310 -365 33340 -335
rect 33310 -415 33340 -385
rect 33395 -365 33425 -335
rect 33395 -415 33425 -385
rect 33480 -365 33510 -335
rect 33480 -415 33510 -385
rect 33565 -365 33595 -335
rect 33565 -415 33595 -385
rect 33650 -365 33680 -335
rect 33650 -415 33680 -385
rect 33735 -365 33765 -335
rect 33735 -415 33765 -385
rect 33820 -365 33850 -335
rect 33820 -415 33850 -385
rect 33905 -365 33935 -335
rect 33905 -415 33935 -385
rect 33990 -365 34020 -335
rect 33990 -415 34020 -385
rect 34075 -365 34105 -335
rect 34075 -415 34105 -385
rect 34160 -365 34190 -335
rect 34160 -415 34190 -385
rect 34245 -365 34275 -335
rect 34245 -415 34275 -385
rect 34330 -365 34360 -335
rect 34330 -415 34360 -385
rect 34415 -365 34445 -335
rect 34415 -415 34445 -385
rect 34500 -365 34530 -335
rect 34500 -415 34530 -385
rect 34585 -365 34615 -335
rect 34585 -415 34615 -385
rect 34670 -365 34700 -335
rect 34670 -415 34700 -385
rect 34755 -365 34785 -335
rect 34755 -415 34785 -385
rect 34840 -365 34870 -335
rect 34840 -415 34870 -385
rect 34925 -365 34955 -335
rect 34925 -415 34955 -385
rect 35010 -365 35040 -335
rect 35010 -415 35040 -385
rect 35095 -365 35125 -335
rect 35095 -415 35125 -385
rect 35180 -365 35210 -335
rect 35180 -415 35210 -385
rect 35265 -365 35295 -335
rect 35265 -415 35295 -385
rect 35350 -365 35380 -335
rect 35350 -415 35380 -385
rect 35435 -365 35465 -335
rect 35435 -415 35465 -385
rect 35520 -365 35550 -335
rect 35520 -415 35550 -385
rect 35605 -365 35635 -335
rect 35605 -415 35635 -385
rect 35690 -365 35720 -335
rect 35690 -415 35720 -385
rect 35775 -365 35805 -335
rect 35775 -415 35805 -385
rect 35860 -365 35890 -335
rect 35860 -415 35890 -385
rect 35945 -365 35975 -335
rect 35945 -415 35975 -385
rect 36030 -365 36060 -335
rect 36030 -415 36060 -385
rect 36115 -365 36145 -335
rect 36115 -415 36145 -385
rect 36200 -365 36230 -335
rect 36200 -415 36230 -385
rect 36285 -365 36315 -335
rect 36285 -415 36315 -385
rect 36370 -365 36400 -335
rect 36370 -415 36400 -385
rect 36455 -365 36485 -335
rect 36455 -415 36485 -385
rect 36540 -365 36570 -335
rect 36540 -415 36570 -385
rect 36625 -365 36655 -335
rect 36625 -415 36655 -385
rect 36710 -365 36740 -335
rect 36710 -415 36740 -385
rect 36795 -365 36825 -335
rect 36795 -415 36825 -385
rect 36880 -365 36910 -335
rect 36880 -415 36910 -385
rect 36965 -365 36995 -335
rect 36965 -415 36995 -385
rect 37050 -365 37080 -335
rect 37050 -415 37080 -385
rect 37135 -365 37165 -335
rect 37135 -415 37165 -385
rect 37220 -365 37250 -335
rect 37220 -415 37250 -385
rect 37305 -365 37335 -335
rect 37305 -415 37335 -385
rect 37390 -365 37420 -335
rect 37390 -415 37420 -385
rect 37475 -365 37505 -335
rect 37475 -415 37505 -385
rect 37560 -365 37590 -335
rect 37560 -415 37590 -385
rect 37645 -365 37675 -335
rect 37645 -415 37675 -385
rect 37730 -365 37760 -335
rect 37730 -415 37760 -385
rect 37815 -365 37845 -335
rect 37815 -415 37845 -385
rect 37900 -365 37930 -335
rect 37900 -415 37930 -385
rect 37985 -365 38015 -335
rect 37985 -415 38015 -385
rect 38070 -365 38100 -335
rect 38070 -415 38100 -385
rect 38155 -365 38185 -335
rect 38155 -415 38185 -385
rect 38240 -365 38270 -335
rect 38240 -415 38270 -385
rect 38325 -365 38355 -335
rect 38325 -415 38355 -385
rect 38410 -365 38440 -335
rect 38410 -415 38440 -385
rect 38495 -365 38525 -335
rect 38495 -415 38525 -385
rect 38580 -365 38610 -335
rect 38580 -415 38610 -385
rect 38665 -365 38695 -335
rect 38665 -415 38695 -385
rect 38750 -365 38780 -335
rect 38750 -415 38780 -385
rect 38835 -365 38865 -335
rect 38835 -415 38865 -385
rect 38920 -365 38950 -335
rect 38920 -415 38950 -385
rect 39005 -365 39035 -335
rect 39005 -415 39035 -385
rect 39090 -365 39120 -335
rect 39090 -415 39120 -385
rect 39175 -365 39205 -335
rect 39175 -415 39205 -385
rect 39260 -365 39290 -335
rect 39260 -415 39290 -385
rect 39345 -365 39375 -335
rect 39345 -415 39375 -385
rect 39430 -365 39460 -335
rect 39430 -415 39460 -385
rect 39515 -365 39545 -335
rect 39515 -415 39545 -385
rect 39600 -365 39630 -335
rect 39600 -415 39630 -385
rect 39685 -365 39715 -335
rect 39685 -415 39715 -385
rect 39770 -365 39800 -335
rect 39770 -415 39800 -385
rect 39855 -365 39885 -335
rect 39855 -415 39885 -385
rect 39940 -365 39970 -335
rect 39940 -415 39970 -385
rect 40025 -365 40055 -335
rect 40025 -415 40055 -385
rect 40110 -365 40140 -335
rect 40110 -415 40140 -385
rect 40195 -365 40225 -335
rect 40195 -415 40225 -385
rect 40280 -365 40310 -335
rect 40280 -415 40310 -385
rect 40365 -365 40395 -335
rect 40365 -415 40395 -385
rect 40450 -365 40480 -335
rect 40450 -415 40480 -385
rect 40535 -365 40565 -335
rect 40535 -415 40565 -385
rect 40620 -365 40650 -335
rect 40620 -415 40650 -385
rect 40705 -365 40735 -335
rect 40705 -415 40735 -385
rect 40790 -365 40820 -335
rect 40790 -415 40820 -385
rect 40875 -365 40905 -335
rect 40875 -415 40905 -385
rect 40960 -365 40990 -335
rect 40960 -415 40990 -385
rect 41045 -365 41075 -335
rect 41045 -415 41075 -385
rect 41130 -365 41160 -335
rect 41130 -415 41160 -385
rect 41215 -365 41245 -335
rect 41215 -415 41245 -385
rect 41300 -365 41330 -335
rect 41300 -415 41330 -385
rect 41385 -365 41415 -335
rect 41385 -415 41415 -385
rect 41470 -365 41500 -335
rect 41470 -415 41500 -385
rect 41555 -365 41585 -335
rect 41555 -415 41585 -385
rect 41640 -365 41670 -335
rect 41640 -415 41670 -385
rect 41725 -365 41755 -335
rect 41725 -415 41755 -385
rect 41810 -365 41840 -335
rect 41810 -415 41840 -385
rect 41895 -365 41925 -335
rect 41895 -415 41925 -385
rect 41980 -365 42010 -335
rect 41980 -415 42010 -385
rect 42065 -365 42095 -335
rect 42065 -415 42095 -385
rect 42150 -365 42180 -335
rect 42150 -415 42180 -385
rect 42235 -365 42265 -335
rect 42235 -415 42265 -385
rect 42320 -365 42350 -335
rect 42320 -415 42350 -385
rect 42405 -365 42435 -335
rect 42405 -415 42435 -385
rect 42490 -365 42520 -335
rect 42490 -415 42520 -385
rect 42575 -365 42605 -335
rect 42575 -415 42605 -385
rect 42660 -365 42690 -335
rect 42660 -415 42690 -385
rect 42745 -365 42775 -335
rect 42745 -415 42775 -385
rect 42830 -365 42860 -335
rect 42830 -415 42860 -385
rect 42915 -365 42945 -335
rect 42915 -415 42945 -385
rect 43000 -365 43030 -335
rect 43000 -415 43030 -385
rect 43085 -365 43115 -335
rect 43085 -415 43115 -385
rect 43170 -365 43200 -335
rect 43170 -415 43200 -385
rect 43255 -365 43285 -335
rect 43255 -415 43285 -385
rect 43340 -365 43370 -335
rect 43340 -415 43370 -385
rect 43425 -365 43455 -335
rect 43425 -415 43455 -385
rect 43510 -365 43540 -335
rect 43510 -415 43540 -385
rect 43595 -365 43625 -335
rect 43595 -415 43625 -385
<< pdiffc >>
rect 15 175 45 205
rect 15 125 45 155
rect 100 175 130 205
rect 100 125 130 155
rect 225 175 255 205
rect 225 125 255 155
rect 310 175 340 205
rect 310 125 340 155
rect 395 175 425 205
rect 395 125 425 155
rect 480 175 510 205
rect 480 125 510 155
rect 565 175 595 205
rect 565 125 595 155
rect 760 175 790 205
rect 760 125 790 155
rect 845 175 875 205
rect 845 125 875 155
rect 930 175 960 205
rect 930 125 960 155
rect 1015 175 1045 205
rect 1015 125 1045 155
rect 1100 175 1130 205
rect 1100 125 1130 155
rect 1185 175 1215 205
rect 1185 125 1215 155
rect 1270 175 1300 205
rect 1270 125 1300 155
rect 1355 175 1385 205
rect 1355 125 1385 155
rect 1440 175 1470 205
rect 1440 125 1470 155
rect 1525 175 1555 205
rect 1525 125 1555 155
rect 1610 175 1640 205
rect 1610 125 1640 155
rect 1695 175 1725 205
rect 1695 125 1725 155
rect 1780 175 1810 205
rect 1780 125 1810 155
rect 1865 175 1895 205
rect 1865 125 1895 155
rect 1950 175 1980 205
rect 1950 125 1980 155
rect 2035 175 2065 205
rect 2035 125 2065 155
rect 2120 175 2150 205
rect 2120 125 2150 155
rect 2270 175 2300 205
rect 2270 125 2300 155
rect 2355 175 2385 205
rect 2355 125 2385 155
rect 2440 175 2470 205
rect 2440 125 2470 155
rect 2525 175 2555 205
rect 2525 125 2555 155
rect 2610 175 2640 205
rect 2610 125 2640 155
rect 2695 175 2725 205
rect 2695 125 2725 155
rect 2780 175 2810 205
rect 2780 125 2810 155
rect 2865 175 2895 205
rect 2865 125 2895 155
rect 2950 175 2980 205
rect 2950 125 2980 155
rect 3035 175 3065 205
rect 3035 125 3065 155
rect 3120 175 3150 205
rect 3120 125 3150 155
rect 3205 175 3235 205
rect 3205 125 3235 155
rect 3290 175 3320 205
rect 3290 125 3320 155
rect 3375 175 3405 205
rect 3375 125 3405 155
rect 3460 175 3490 205
rect 3460 125 3490 155
rect 3545 175 3575 205
rect 3545 125 3575 155
rect 3630 175 3660 205
rect 3630 125 3660 155
rect 3715 175 3745 205
rect 3715 125 3745 155
rect 3800 175 3830 205
rect 3800 125 3830 155
rect 3885 175 3915 205
rect 3885 125 3915 155
rect 3970 175 4000 205
rect 3970 125 4000 155
rect 4055 175 4085 205
rect 4055 125 4085 155
rect 4140 175 4170 205
rect 4140 125 4170 155
rect 4225 175 4255 205
rect 4225 125 4255 155
rect 4310 175 4340 205
rect 4310 125 4340 155
rect 4395 175 4425 205
rect 4395 125 4425 155
rect 4480 175 4510 205
rect 4480 125 4510 155
rect 4565 175 4595 205
rect 4565 125 4595 155
rect 4650 175 4680 205
rect 4650 125 4680 155
rect 4735 175 4765 205
rect 4735 125 4765 155
rect 4820 175 4850 205
rect 4820 125 4850 155
rect 4905 175 4935 205
rect 4905 125 4935 155
rect 4990 175 5020 205
rect 4990 125 5020 155
rect 5075 175 5105 205
rect 5075 125 5105 155
rect 5160 175 5190 205
rect 5160 125 5190 155
rect 5245 175 5275 205
rect 5245 125 5275 155
rect 5330 175 5360 205
rect 5330 125 5360 155
rect 5415 175 5445 205
rect 5415 125 5445 155
rect 5500 175 5530 205
rect 5500 125 5530 155
rect 5585 175 5615 205
rect 5585 125 5615 155
rect 5670 175 5700 205
rect 5670 125 5700 155
rect 5755 175 5785 205
rect 5755 125 5785 155
rect 5840 175 5870 205
rect 5840 125 5870 155
rect 5925 175 5955 205
rect 5925 125 5955 155
rect 6010 175 6040 205
rect 6010 125 6040 155
rect 6095 175 6125 205
rect 6095 125 6125 155
rect 6180 175 6210 205
rect 6180 125 6210 155
rect 6265 175 6295 205
rect 6265 125 6295 155
rect 6350 175 6380 205
rect 6350 125 6380 155
rect 6435 175 6465 205
rect 6435 125 6465 155
rect 6520 175 6550 205
rect 6520 125 6550 155
rect 6605 175 6635 205
rect 6605 125 6635 155
rect 6690 175 6720 205
rect 6690 125 6720 155
rect 6775 175 6805 205
rect 6775 125 6805 155
rect 6860 175 6890 205
rect 6860 125 6890 155
rect 6945 175 6975 205
rect 6945 125 6975 155
rect 7030 175 7060 205
rect 7030 125 7060 155
rect 7115 175 7145 205
rect 7115 125 7145 155
rect 7200 175 7230 205
rect 7200 125 7230 155
rect 7285 175 7315 205
rect 7285 125 7315 155
rect 7370 175 7400 205
rect 7370 125 7400 155
rect 7455 175 7485 205
rect 7455 125 7485 155
rect 7540 175 7570 205
rect 7540 125 7570 155
rect 7625 175 7655 205
rect 7625 125 7655 155
rect 7710 175 7740 205
rect 7710 125 7740 155
rect 7860 175 7890 205
rect 7860 125 7890 155
rect 7945 175 7975 205
rect 7945 125 7975 155
rect 8030 175 8060 205
rect 8030 125 8060 155
rect 8115 175 8145 205
rect 8115 125 8145 155
rect 8200 175 8230 205
rect 8200 125 8230 155
rect 8285 175 8315 205
rect 8285 125 8315 155
rect 8370 175 8400 205
rect 8370 125 8400 155
rect 8455 175 8485 205
rect 8455 125 8485 155
rect 8540 175 8570 205
rect 8540 125 8570 155
rect 8625 175 8655 205
rect 8625 125 8655 155
rect 8710 175 8740 205
rect 8710 125 8740 155
rect 8795 175 8825 205
rect 8795 125 8825 155
rect 8880 175 8910 205
rect 8880 125 8910 155
rect 8965 175 8995 205
rect 8965 125 8995 155
rect 9050 175 9080 205
rect 9050 125 9080 155
rect 9135 175 9165 205
rect 9135 125 9165 155
rect 9220 175 9250 205
rect 9220 125 9250 155
rect 9305 175 9335 205
rect 9305 125 9335 155
rect 9390 175 9420 205
rect 9390 125 9420 155
rect 9475 175 9505 205
rect 9475 125 9505 155
rect 9560 175 9590 205
rect 9560 125 9590 155
rect 9645 175 9675 205
rect 9645 125 9675 155
rect 9730 175 9760 205
rect 9730 125 9760 155
rect 9815 175 9845 205
rect 9815 125 9845 155
rect 9900 175 9930 205
rect 9900 125 9930 155
rect 9985 175 10015 205
rect 9985 125 10015 155
rect 10070 175 10100 205
rect 10070 125 10100 155
rect 10155 175 10185 205
rect 10155 125 10185 155
rect 10240 175 10270 205
rect 10240 125 10270 155
rect 10325 175 10355 205
rect 10325 125 10355 155
rect 10410 175 10440 205
rect 10410 125 10440 155
rect 10495 175 10525 205
rect 10495 125 10525 155
rect 10580 175 10610 205
rect 10580 125 10610 155
rect 10665 175 10695 205
rect 10665 125 10695 155
rect 10750 175 10780 205
rect 10750 125 10780 155
rect 10835 175 10865 205
rect 10835 125 10865 155
rect 10920 175 10950 205
rect 10920 125 10950 155
rect 11005 175 11035 205
rect 11005 125 11035 155
rect 11090 175 11120 205
rect 11090 125 11120 155
rect 11175 175 11205 205
rect 11175 125 11205 155
rect 11260 175 11290 205
rect 11260 125 11290 155
rect 11345 175 11375 205
rect 11345 125 11375 155
rect 11430 175 11460 205
rect 11430 125 11460 155
rect 11515 175 11545 205
rect 11515 125 11545 155
rect 11600 175 11630 205
rect 11600 125 11630 155
rect 11685 175 11715 205
rect 11685 125 11715 155
rect 11770 175 11800 205
rect 11770 125 11800 155
rect 11855 175 11885 205
rect 11855 125 11885 155
rect 11940 175 11970 205
rect 11940 125 11970 155
rect 12025 175 12055 205
rect 12025 125 12055 155
rect 12110 175 12140 205
rect 12110 125 12140 155
rect 12195 175 12225 205
rect 12195 125 12225 155
rect 12280 175 12310 205
rect 12280 125 12310 155
rect 12365 175 12395 205
rect 12365 125 12395 155
rect 12450 175 12480 205
rect 12450 125 12480 155
rect 12535 175 12565 205
rect 12535 125 12565 155
rect 12620 175 12650 205
rect 12620 125 12650 155
rect 12705 175 12735 205
rect 12705 125 12735 155
rect 12790 175 12820 205
rect 12790 125 12820 155
rect 12875 175 12905 205
rect 12875 125 12905 155
rect 12960 175 12990 205
rect 12960 125 12990 155
rect 13045 175 13075 205
rect 13045 125 13075 155
rect 13130 175 13160 205
rect 13130 125 13160 155
rect 13215 175 13245 205
rect 13215 125 13245 155
rect 13300 175 13330 205
rect 13300 125 13330 155
rect 13385 175 13415 205
rect 13385 125 13415 155
rect 13470 175 13500 205
rect 13470 125 13500 155
rect 13555 175 13585 205
rect 13555 125 13585 155
rect 13640 175 13670 205
rect 13640 125 13670 155
rect 13725 175 13755 205
rect 13725 125 13755 155
rect 13810 175 13840 205
rect 13810 125 13840 155
rect 13895 175 13925 205
rect 13895 125 13925 155
rect 13980 175 14010 205
rect 13980 125 14010 155
rect 14065 175 14095 205
rect 14065 125 14095 155
rect 14150 175 14180 205
rect 14150 125 14180 155
rect 14235 175 14265 205
rect 14235 125 14265 155
rect 14320 175 14350 205
rect 14320 125 14350 155
rect 14405 175 14435 205
rect 14405 125 14435 155
rect 14490 175 14520 205
rect 14490 125 14520 155
rect 14575 175 14605 205
rect 14575 125 14605 155
rect 14660 175 14690 205
rect 14660 125 14690 155
rect 14745 175 14775 205
rect 14745 125 14775 155
rect 14830 175 14860 205
rect 14830 125 14860 155
rect 14915 175 14945 205
rect 14915 125 14945 155
rect 15000 175 15030 205
rect 15000 125 15030 155
rect 15085 175 15115 205
rect 15085 125 15115 155
rect 15170 175 15200 205
rect 15170 125 15200 155
rect 15255 175 15285 205
rect 15255 125 15285 155
rect 15340 175 15370 205
rect 15340 125 15370 155
rect 15425 175 15455 205
rect 15425 125 15455 155
rect 15510 175 15540 205
rect 15510 125 15540 155
rect 15595 175 15625 205
rect 15595 125 15625 155
rect 15680 175 15710 205
rect 15680 125 15710 155
rect 15765 175 15795 205
rect 15765 125 15795 155
rect 15850 175 15880 205
rect 15850 125 15880 155
rect 15935 175 15965 205
rect 15935 125 15965 155
rect 16020 175 16050 205
rect 16020 125 16050 155
rect 16105 175 16135 205
rect 16105 125 16135 155
rect 16190 175 16220 205
rect 16190 125 16220 155
rect 16275 175 16305 205
rect 16275 125 16305 155
rect 16360 175 16390 205
rect 16360 125 16390 155
rect 16445 175 16475 205
rect 16445 125 16475 155
rect 16530 175 16560 205
rect 16530 125 16560 155
rect 16615 175 16645 205
rect 16615 125 16645 155
rect 16700 175 16730 205
rect 16700 125 16730 155
rect 16785 175 16815 205
rect 16785 125 16815 155
rect 16870 175 16900 205
rect 16870 125 16900 155
rect 16955 175 16985 205
rect 16955 125 16985 155
rect 17040 175 17070 205
rect 17040 125 17070 155
rect 17125 175 17155 205
rect 17125 125 17155 155
rect 17210 175 17240 205
rect 17210 125 17240 155
rect 17295 175 17325 205
rect 17295 125 17325 155
rect 17380 175 17410 205
rect 17380 125 17410 155
rect 17465 175 17495 205
rect 17465 125 17495 155
rect 17550 175 17580 205
rect 17550 125 17580 155
rect 17635 175 17665 205
rect 17635 125 17665 155
rect 17720 175 17750 205
rect 17720 125 17750 155
rect 17805 175 17835 205
rect 17805 125 17835 155
rect 17890 175 17920 205
rect 17890 125 17920 155
rect 17975 175 18005 205
rect 17975 125 18005 155
rect 18060 175 18090 205
rect 18060 125 18090 155
rect 18145 175 18175 205
rect 18145 125 18175 155
rect 18230 175 18260 205
rect 18230 125 18260 155
rect 18315 175 18345 205
rect 18315 125 18345 155
rect 18400 175 18430 205
rect 18400 125 18430 155
rect 18485 175 18515 205
rect 18485 125 18515 155
rect 18570 175 18600 205
rect 18570 125 18600 155
rect 18655 175 18685 205
rect 18655 125 18685 155
rect 18740 175 18770 205
rect 18740 125 18770 155
rect 18825 175 18855 205
rect 18825 125 18855 155
rect 18910 175 18940 205
rect 18910 125 18940 155
rect 18995 175 19025 205
rect 18995 125 19025 155
rect 19080 175 19110 205
rect 19080 125 19110 155
rect 19165 175 19195 205
rect 19165 125 19195 155
rect 19250 175 19280 205
rect 19250 125 19280 155
rect 19335 175 19365 205
rect 19335 125 19365 155
rect 19420 175 19450 205
rect 19420 125 19450 155
rect 19505 175 19535 205
rect 19505 125 19535 155
rect 19590 175 19620 205
rect 19590 125 19620 155
rect 19675 175 19705 205
rect 19675 125 19705 155
rect 19760 175 19790 205
rect 19760 125 19790 155
rect 19845 175 19875 205
rect 19845 125 19875 155
rect 19930 175 19960 205
rect 19930 125 19960 155
rect 20015 175 20045 205
rect 20015 125 20045 155
rect 20100 175 20130 205
rect 20100 125 20130 155
rect 20185 175 20215 205
rect 20185 125 20215 155
rect 20270 175 20300 205
rect 20270 125 20300 155
rect 20355 175 20385 205
rect 20355 125 20385 155
rect 20440 175 20470 205
rect 20440 125 20470 155
rect 20525 175 20555 205
rect 20525 125 20555 155
rect 20610 175 20640 205
rect 20610 125 20640 155
rect 20695 175 20725 205
rect 20695 125 20725 155
rect 20780 175 20810 205
rect 20780 125 20810 155
rect 20865 175 20895 205
rect 20865 125 20895 155
rect 20950 175 20980 205
rect 20950 125 20980 155
rect 21035 175 21065 205
rect 21035 125 21065 155
rect 21120 175 21150 205
rect 21120 125 21150 155
rect 21205 175 21235 205
rect 21205 125 21235 155
rect 21290 175 21320 205
rect 21290 125 21320 155
rect 21375 175 21405 205
rect 21375 125 21405 155
rect 21460 175 21490 205
rect 21460 125 21490 155
rect 21545 175 21575 205
rect 21545 125 21575 155
rect 21630 175 21660 205
rect 21630 125 21660 155
rect 21715 175 21745 205
rect 21715 125 21745 155
rect 21800 175 21830 205
rect 21800 125 21830 155
rect 21885 175 21915 205
rect 21885 125 21915 155
rect 21970 175 22000 205
rect 21970 125 22000 155
rect 22055 175 22085 205
rect 22055 125 22085 155
rect 22140 175 22170 205
rect 22140 125 22170 155
rect 22225 175 22255 205
rect 22225 125 22255 155
rect 22310 175 22340 205
rect 22310 125 22340 155
rect 22395 175 22425 205
rect 22395 125 22425 155
rect 22480 175 22510 205
rect 22480 125 22510 155
rect 22565 175 22595 205
rect 22565 125 22595 155
rect 22650 175 22680 205
rect 22650 125 22680 155
rect 22735 175 22765 205
rect 22735 125 22765 155
rect 22820 175 22850 205
rect 22820 125 22850 155
rect 22905 175 22935 205
rect 22905 125 22935 155
rect 22990 175 23020 205
rect 22990 125 23020 155
rect 23075 175 23105 205
rect 23075 125 23105 155
rect 23160 175 23190 205
rect 23160 125 23190 155
rect 23245 175 23275 205
rect 23245 125 23275 155
rect 23330 175 23360 205
rect 23330 125 23360 155
rect 23415 175 23445 205
rect 23415 125 23445 155
rect 23500 175 23530 205
rect 23500 125 23530 155
rect 23585 175 23615 205
rect 23585 125 23615 155
rect 23670 175 23700 205
rect 23670 125 23700 155
rect 23755 175 23785 205
rect 23755 125 23785 155
rect 23840 175 23870 205
rect 23840 125 23870 155
rect 23925 175 23955 205
rect 23925 125 23955 155
rect 24010 175 24040 205
rect 24010 125 24040 155
rect 24095 175 24125 205
rect 24095 125 24125 155
rect 24180 175 24210 205
rect 24180 125 24210 155
rect 24265 175 24295 205
rect 24265 125 24295 155
rect 24350 175 24380 205
rect 24350 125 24380 155
rect 24435 175 24465 205
rect 24435 125 24465 155
rect 24520 175 24550 205
rect 24520 125 24550 155
rect 24605 175 24635 205
rect 24605 125 24635 155
rect 24690 175 24720 205
rect 24690 125 24720 155
rect 24775 175 24805 205
rect 24775 125 24805 155
rect 24860 175 24890 205
rect 24860 125 24890 155
rect 24945 175 24975 205
rect 24945 125 24975 155
rect 25030 175 25060 205
rect 25030 125 25060 155
rect 25115 175 25145 205
rect 25115 125 25145 155
rect 25200 175 25230 205
rect 25200 125 25230 155
rect 25285 175 25315 205
rect 25285 125 25315 155
rect 25370 175 25400 205
rect 25370 125 25400 155
rect 25455 175 25485 205
rect 25455 125 25485 155
rect 25540 175 25570 205
rect 25540 125 25570 155
rect 25625 175 25655 205
rect 25625 125 25655 155
rect 25710 175 25740 205
rect 25710 125 25740 155
rect 25795 175 25825 205
rect 25795 125 25825 155
rect 25880 175 25910 205
rect 25880 125 25910 155
rect 25965 175 25995 205
rect 25965 125 25995 155
rect 26050 175 26080 205
rect 26050 125 26080 155
rect 26135 175 26165 205
rect 26135 125 26165 155
rect 26220 175 26250 205
rect 26220 125 26250 155
rect 26305 175 26335 205
rect 26305 125 26335 155
rect 26390 175 26420 205
rect 26390 125 26420 155
rect 26475 175 26505 205
rect 26475 125 26505 155
rect 26560 175 26590 205
rect 26560 125 26590 155
rect 26645 175 26675 205
rect 26645 125 26675 155
rect 26730 175 26760 205
rect 26730 125 26760 155
rect 26815 175 26845 205
rect 26815 125 26845 155
rect 26900 175 26930 205
rect 26900 125 26930 155
rect 26985 175 27015 205
rect 26985 125 27015 155
rect 27070 175 27100 205
rect 27070 125 27100 155
rect 27155 175 27185 205
rect 27155 125 27185 155
rect 27240 175 27270 205
rect 27240 125 27270 155
rect 27325 175 27355 205
rect 27325 125 27355 155
rect 27410 175 27440 205
rect 27410 125 27440 155
rect 27495 175 27525 205
rect 27495 125 27525 155
rect 27580 175 27610 205
rect 27580 125 27610 155
rect 27665 175 27695 205
rect 27665 125 27695 155
rect 27750 175 27780 205
rect 27750 125 27780 155
rect 27835 175 27865 205
rect 27835 125 27865 155
rect 27920 175 27950 205
rect 27920 125 27950 155
rect 28005 175 28035 205
rect 28005 125 28035 155
rect 28090 175 28120 205
rect 28090 125 28120 155
rect 28175 175 28205 205
rect 28175 125 28205 155
rect 28260 175 28290 205
rect 28260 125 28290 155
rect 28345 175 28375 205
rect 28345 125 28375 155
rect 28430 175 28460 205
rect 28430 125 28460 155
rect 28515 175 28545 205
rect 28515 125 28545 155
rect 28600 175 28630 205
rect 28600 125 28630 155
rect 28685 175 28715 205
rect 28685 125 28715 155
rect 28770 175 28800 205
rect 28770 125 28800 155
rect 28855 175 28885 205
rect 28855 125 28885 155
rect 28940 175 28970 205
rect 28940 125 28970 155
rect 29025 175 29055 205
rect 29025 125 29055 155
rect 29110 175 29140 205
rect 29110 125 29140 155
rect 29195 175 29225 205
rect 29195 125 29225 155
rect 29280 175 29310 205
rect 29280 125 29310 155
rect 29365 175 29395 205
rect 29365 125 29395 155
rect 29450 175 29480 205
rect 29450 125 29480 155
rect 29535 175 29565 205
rect 29535 125 29565 155
rect 29620 175 29650 205
rect 29620 125 29650 155
rect 75 -530 105 -500
rect 75 -580 105 -550
rect 75 -630 105 -600
rect 75 -680 105 -650
rect 160 -530 190 -500
rect 160 -580 190 -550
rect 160 -630 190 -600
rect 160 -680 190 -650
rect 245 -530 275 -500
rect 245 -580 275 -550
rect 245 -630 275 -600
rect 245 -680 275 -650
rect 330 -530 360 -500
rect 330 -580 360 -550
rect 330 -630 360 -600
rect 330 -680 360 -650
rect 415 -530 445 -500
rect 415 -580 445 -550
rect 415 -630 445 -600
rect 415 -680 445 -650
rect 500 -530 530 -500
rect 500 -580 530 -550
rect 500 -630 530 -600
rect 500 -680 530 -650
rect 585 -530 615 -500
rect 585 -580 615 -550
rect 585 -630 615 -600
rect 585 -680 615 -650
rect 670 -530 700 -500
rect 670 -580 700 -550
rect 670 -630 700 -600
rect 670 -680 700 -650
rect 755 -530 785 -500
rect 755 -580 785 -550
rect 755 -630 785 -600
rect 755 -680 785 -650
rect 840 -530 870 -500
rect 840 -580 870 -550
rect 840 -630 870 -600
rect 840 -680 870 -650
rect 925 -530 955 -500
rect 925 -580 955 -550
rect 925 -630 955 -600
rect 925 -680 955 -650
rect 1010 -530 1040 -500
rect 1010 -580 1040 -550
rect 1010 -630 1040 -600
rect 1010 -680 1040 -650
rect 1095 -530 1125 -500
rect 1095 -580 1125 -550
rect 1095 -630 1125 -600
rect 1095 -680 1125 -650
rect 1180 -530 1210 -500
rect 1180 -580 1210 -550
rect 1180 -630 1210 -600
rect 1180 -680 1210 -650
rect 1265 -530 1295 -500
rect 1265 -580 1295 -550
rect 1265 -630 1295 -600
rect 1265 -680 1295 -650
rect 1350 -530 1380 -500
rect 1350 -580 1380 -550
rect 1350 -630 1380 -600
rect 1350 -680 1380 -650
rect 1435 -530 1465 -500
rect 1435 -580 1465 -550
rect 1435 -630 1465 -600
rect 1435 -680 1465 -650
rect 1520 -530 1550 -500
rect 1520 -580 1550 -550
rect 1520 -630 1550 -600
rect 1520 -680 1550 -650
rect 1605 -530 1635 -500
rect 1605 -580 1635 -550
rect 1605 -630 1635 -600
rect 1605 -680 1635 -650
rect 1690 -530 1720 -500
rect 1690 -580 1720 -550
rect 1690 -630 1720 -600
rect 1690 -680 1720 -650
rect 1775 -530 1805 -500
rect 1775 -580 1805 -550
rect 1775 -630 1805 -600
rect 1775 -680 1805 -650
rect 1860 -530 1890 -500
rect 1860 -580 1890 -550
rect 1860 -630 1890 -600
rect 1860 -680 1890 -650
rect 1945 -530 1975 -500
rect 1945 -580 1975 -550
rect 1945 -630 1975 -600
rect 1945 -680 1975 -650
rect 2030 -530 2060 -500
rect 2030 -580 2060 -550
rect 2030 -630 2060 -600
rect 2030 -680 2060 -650
rect 2115 -530 2145 -500
rect 2115 -580 2145 -550
rect 2115 -630 2145 -600
rect 2115 -680 2145 -650
rect 2200 -530 2230 -500
rect 2200 -580 2230 -550
rect 2200 -630 2230 -600
rect 2200 -680 2230 -650
rect 2285 -530 2315 -500
rect 2285 -580 2315 -550
rect 2285 -630 2315 -600
rect 2285 -680 2315 -650
rect 2370 -530 2400 -500
rect 2370 -580 2400 -550
rect 2370 -630 2400 -600
rect 2370 -680 2400 -650
rect 2455 -530 2485 -500
rect 2455 -580 2485 -550
rect 2455 -630 2485 -600
rect 2455 -680 2485 -650
rect 2540 -530 2570 -500
rect 2540 -580 2570 -550
rect 2540 -630 2570 -600
rect 2540 -680 2570 -650
rect 2625 -530 2655 -500
rect 2625 -580 2655 -550
rect 2625 -630 2655 -600
rect 2625 -680 2655 -650
rect 2710 -530 2740 -500
rect 2710 -580 2740 -550
rect 2710 -630 2740 -600
rect 2710 -680 2740 -650
rect 2795 -530 2825 -500
rect 2795 -580 2825 -550
rect 2795 -630 2825 -600
rect 2795 -680 2825 -650
rect 2880 -530 2910 -500
rect 2880 -580 2910 -550
rect 2880 -630 2910 -600
rect 2880 -680 2910 -650
rect 2965 -530 2995 -500
rect 2965 -580 2995 -550
rect 2965 -630 2995 -600
rect 2965 -680 2995 -650
rect 3050 -530 3080 -500
rect 3050 -580 3080 -550
rect 3050 -630 3080 -600
rect 3050 -680 3080 -650
rect 3135 -530 3165 -500
rect 3135 -580 3165 -550
rect 3135 -630 3165 -600
rect 3135 -680 3165 -650
rect 3220 -530 3250 -500
rect 3220 -580 3250 -550
rect 3220 -630 3250 -600
rect 3220 -680 3250 -650
rect 3305 -530 3335 -500
rect 3305 -580 3335 -550
rect 3305 -630 3335 -600
rect 3305 -680 3335 -650
rect 3390 -530 3420 -500
rect 3390 -580 3420 -550
rect 3390 -630 3420 -600
rect 3390 -680 3420 -650
rect 3475 -530 3505 -500
rect 3475 -580 3505 -550
rect 3475 -630 3505 -600
rect 3475 -680 3505 -650
rect 3560 -530 3590 -500
rect 3560 -580 3590 -550
rect 3560 -630 3590 -600
rect 3560 -680 3590 -650
rect 3645 -530 3675 -500
rect 3645 -580 3675 -550
rect 3645 -630 3675 -600
rect 3645 -680 3675 -650
rect 3730 -530 3760 -500
rect 3730 -580 3760 -550
rect 3730 -630 3760 -600
rect 3730 -680 3760 -650
rect 3815 -530 3845 -500
rect 3815 -580 3845 -550
rect 3815 -630 3845 -600
rect 3815 -680 3845 -650
rect 3900 -530 3930 -500
rect 3900 -580 3930 -550
rect 3900 -630 3930 -600
rect 3900 -680 3930 -650
rect 3985 -530 4015 -500
rect 3985 -580 4015 -550
rect 3985 -630 4015 -600
rect 3985 -680 4015 -650
rect 4070 -530 4100 -500
rect 4070 -580 4100 -550
rect 4070 -630 4100 -600
rect 4070 -680 4100 -650
rect 4155 -530 4185 -500
rect 4155 -580 4185 -550
rect 4155 -630 4185 -600
rect 4155 -680 4185 -650
rect 4240 -530 4270 -500
rect 4240 -580 4270 -550
rect 4240 -630 4270 -600
rect 4240 -680 4270 -650
rect 4325 -530 4355 -500
rect 4325 -580 4355 -550
rect 4325 -630 4355 -600
rect 4325 -680 4355 -650
rect 4410 -530 4440 -500
rect 4410 -580 4440 -550
rect 4410 -630 4440 -600
rect 4410 -680 4440 -650
rect 4495 -530 4525 -500
rect 4495 -580 4525 -550
rect 4495 -630 4525 -600
rect 4495 -680 4525 -650
rect 4580 -530 4610 -500
rect 4580 -580 4610 -550
rect 4580 -630 4610 -600
rect 4580 -680 4610 -650
rect 4665 -530 4695 -500
rect 4665 -580 4695 -550
rect 4665 -630 4695 -600
rect 4665 -680 4695 -650
rect 4750 -530 4780 -500
rect 4750 -580 4780 -550
rect 4750 -630 4780 -600
rect 4750 -680 4780 -650
rect 4835 -530 4865 -500
rect 4835 -580 4865 -550
rect 4835 -630 4865 -600
rect 4835 -680 4865 -650
rect 4920 -530 4950 -500
rect 4920 -580 4950 -550
rect 4920 -630 4950 -600
rect 4920 -680 4950 -650
rect 5005 -530 5035 -500
rect 5005 -580 5035 -550
rect 5005 -630 5035 -600
rect 5005 -680 5035 -650
rect 5090 -530 5120 -500
rect 5090 -580 5120 -550
rect 5090 -630 5120 -600
rect 5090 -680 5120 -650
rect 5175 -530 5205 -500
rect 5175 -580 5205 -550
rect 5175 -630 5205 -600
rect 5175 -680 5205 -650
rect 5260 -530 5290 -500
rect 5260 -580 5290 -550
rect 5260 -630 5290 -600
rect 5260 -680 5290 -650
rect 5345 -530 5375 -500
rect 5345 -580 5375 -550
rect 5345 -630 5375 -600
rect 5345 -680 5375 -650
rect 5430 -530 5460 -500
rect 5430 -580 5460 -550
rect 5430 -630 5460 -600
rect 5430 -680 5460 -650
rect 5515 -530 5545 -500
rect 5515 -580 5545 -550
rect 5515 -630 5545 -600
rect 5515 -680 5545 -650
rect 5600 -530 5630 -500
rect 5600 -580 5630 -550
rect 5600 -630 5630 -600
rect 5600 -680 5630 -650
rect 5685 -530 5715 -500
rect 5685 -580 5715 -550
rect 5685 -630 5715 -600
rect 5685 -680 5715 -650
rect 5770 -530 5800 -500
rect 5770 -580 5800 -550
rect 5770 -630 5800 -600
rect 5770 -680 5800 -650
rect 5855 -530 5885 -500
rect 5855 -580 5885 -550
rect 5855 -630 5885 -600
rect 5855 -680 5885 -650
rect 5940 -530 5970 -500
rect 5940 -580 5970 -550
rect 5940 -630 5970 -600
rect 5940 -680 5970 -650
rect 6025 -530 6055 -500
rect 6025 -580 6055 -550
rect 6025 -630 6055 -600
rect 6025 -680 6055 -650
rect 6110 -530 6140 -500
rect 6110 -580 6140 -550
rect 6110 -630 6140 -600
rect 6110 -680 6140 -650
rect 6195 -530 6225 -500
rect 6195 -580 6225 -550
rect 6195 -630 6225 -600
rect 6195 -680 6225 -650
rect 6280 -530 6310 -500
rect 6280 -580 6310 -550
rect 6280 -630 6310 -600
rect 6280 -680 6310 -650
rect 6365 -530 6395 -500
rect 6365 -580 6395 -550
rect 6365 -630 6395 -600
rect 6365 -680 6395 -650
rect 6450 -530 6480 -500
rect 6450 -580 6480 -550
rect 6450 -630 6480 -600
rect 6450 -680 6480 -650
rect 6535 -530 6565 -500
rect 6535 -580 6565 -550
rect 6535 -630 6565 -600
rect 6535 -680 6565 -650
rect 6620 -530 6650 -500
rect 6620 -580 6650 -550
rect 6620 -630 6650 -600
rect 6620 -680 6650 -650
rect 6705 -530 6735 -500
rect 6705 -580 6735 -550
rect 6705 -630 6735 -600
rect 6705 -680 6735 -650
rect 6790 -530 6820 -500
rect 6790 -580 6820 -550
rect 6790 -630 6820 -600
rect 6790 -680 6820 -650
rect 6875 -530 6905 -500
rect 6875 -580 6905 -550
rect 6875 -630 6905 -600
rect 6875 -680 6905 -650
rect 6960 -530 6990 -500
rect 6960 -580 6990 -550
rect 6960 -630 6990 -600
rect 6960 -680 6990 -650
rect 7045 -530 7075 -500
rect 7045 -580 7075 -550
rect 7045 -630 7075 -600
rect 7045 -680 7075 -650
rect 7130 -530 7160 -500
rect 7130 -580 7160 -550
rect 7130 -630 7160 -600
rect 7130 -680 7160 -650
rect 7215 -530 7245 -500
rect 7215 -580 7245 -550
rect 7215 -630 7245 -600
rect 7215 -680 7245 -650
rect 7300 -530 7330 -500
rect 7300 -580 7330 -550
rect 7300 -630 7330 -600
rect 7300 -680 7330 -650
rect 7385 -530 7415 -500
rect 7385 -580 7415 -550
rect 7385 -630 7415 -600
rect 7385 -680 7415 -650
rect 7470 -530 7500 -500
rect 7470 -580 7500 -550
rect 7470 -630 7500 -600
rect 7470 -680 7500 -650
rect 7555 -530 7585 -500
rect 7555 -580 7585 -550
rect 7555 -630 7585 -600
rect 7555 -680 7585 -650
rect 7640 -530 7670 -500
rect 7640 -580 7670 -550
rect 7640 -630 7670 -600
rect 7640 -680 7670 -650
rect 7725 -530 7755 -500
rect 7725 -580 7755 -550
rect 7725 -630 7755 -600
rect 7725 -680 7755 -650
rect 7810 -530 7840 -500
rect 7810 -580 7840 -550
rect 7810 -630 7840 -600
rect 7810 -680 7840 -650
rect 7895 -530 7925 -500
rect 7895 -580 7925 -550
rect 7895 -630 7925 -600
rect 7895 -680 7925 -650
rect 7980 -530 8010 -500
rect 7980 -580 8010 -550
rect 7980 -630 8010 -600
rect 7980 -680 8010 -650
rect 8065 -530 8095 -500
rect 8065 -580 8095 -550
rect 8065 -630 8095 -600
rect 8065 -680 8095 -650
rect 8150 -530 8180 -500
rect 8150 -580 8180 -550
rect 8150 -630 8180 -600
rect 8150 -680 8180 -650
rect 8235 -530 8265 -500
rect 8235 -580 8265 -550
rect 8235 -630 8265 -600
rect 8235 -680 8265 -650
rect 8320 -530 8350 -500
rect 8320 -580 8350 -550
rect 8320 -630 8350 -600
rect 8320 -680 8350 -650
rect 8405 -530 8435 -500
rect 8405 -580 8435 -550
rect 8405 -630 8435 -600
rect 8405 -680 8435 -650
rect 8490 -530 8520 -500
rect 8490 -580 8520 -550
rect 8490 -630 8520 -600
rect 8490 -680 8520 -650
rect 8575 -530 8605 -500
rect 8575 -580 8605 -550
rect 8575 -630 8605 -600
rect 8575 -680 8605 -650
rect 8660 -530 8690 -500
rect 8660 -580 8690 -550
rect 8660 -630 8690 -600
rect 8660 -680 8690 -650
rect 8745 -530 8775 -500
rect 8745 -580 8775 -550
rect 8745 -630 8775 -600
rect 8745 -680 8775 -650
rect 8830 -530 8860 -500
rect 8830 -580 8860 -550
rect 8830 -630 8860 -600
rect 8830 -680 8860 -650
rect 8915 -530 8945 -500
rect 8915 -580 8945 -550
rect 8915 -630 8945 -600
rect 8915 -680 8945 -650
rect 9000 -530 9030 -500
rect 9000 -580 9030 -550
rect 9000 -630 9030 -600
rect 9000 -680 9030 -650
rect 9085 -530 9115 -500
rect 9085 -580 9115 -550
rect 9085 -630 9115 -600
rect 9085 -680 9115 -650
rect 9170 -530 9200 -500
rect 9170 -580 9200 -550
rect 9170 -630 9200 -600
rect 9170 -680 9200 -650
rect 9255 -530 9285 -500
rect 9255 -580 9285 -550
rect 9255 -630 9285 -600
rect 9255 -680 9285 -650
rect 9340 -530 9370 -500
rect 9340 -580 9370 -550
rect 9340 -630 9370 -600
rect 9340 -680 9370 -650
rect 9425 -530 9455 -500
rect 9425 -580 9455 -550
rect 9425 -630 9455 -600
rect 9425 -680 9455 -650
rect 9510 -530 9540 -500
rect 9510 -580 9540 -550
rect 9510 -630 9540 -600
rect 9510 -680 9540 -650
rect 9595 -530 9625 -500
rect 9595 -580 9625 -550
rect 9595 -630 9625 -600
rect 9595 -680 9625 -650
rect 9680 -530 9710 -500
rect 9680 -580 9710 -550
rect 9680 -630 9710 -600
rect 9680 -680 9710 -650
rect 9765 -530 9795 -500
rect 9765 -580 9795 -550
rect 9765 -630 9795 -600
rect 9765 -680 9795 -650
rect 9850 -530 9880 -500
rect 9850 -580 9880 -550
rect 9850 -630 9880 -600
rect 9850 -680 9880 -650
rect 9935 -530 9965 -500
rect 9935 -580 9965 -550
rect 9935 -630 9965 -600
rect 9935 -680 9965 -650
rect 10020 -530 10050 -500
rect 10020 -580 10050 -550
rect 10020 -630 10050 -600
rect 10020 -680 10050 -650
rect 10105 -530 10135 -500
rect 10105 -580 10135 -550
rect 10105 -630 10135 -600
rect 10105 -680 10135 -650
rect 10190 -530 10220 -500
rect 10190 -580 10220 -550
rect 10190 -630 10220 -600
rect 10190 -680 10220 -650
rect 10275 -530 10305 -500
rect 10275 -580 10305 -550
rect 10275 -630 10305 -600
rect 10275 -680 10305 -650
rect 10360 -530 10390 -500
rect 10360 -580 10390 -550
rect 10360 -630 10390 -600
rect 10360 -680 10390 -650
rect 10445 -530 10475 -500
rect 10445 -580 10475 -550
rect 10445 -630 10475 -600
rect 10445 -680 10475 -650
rect 10530 -530 10560 -500
rect 10530 -580 10560 -550
rect 10530 -630 10560 -600
rect 10530 -680 10560 -650
rect 10615 -530 10645 -500
rect 10615 -580 10645 -550
rect 10615 -630 10645 -600
rect 10615 -680 10645 -650
rect 10700 -530 10730 -500
rect 10700 -580 10730 -550
rect 10700 -630 10730 -600
rect 10700 -680 10730 -650
rect 10785 -530 10815 -500
rect 10785 -580 10815 -550
rect 10785 -630 10815 -600
rect 10785 -680 10815 -650
rect 10870 -530 10900 -500
rect 10870 -580 10900 -550
rect 10870 -630 10900 -600
rect 10870 -680 10900 -650
rect 10955 -530 10985 -500
rect 10955 -580 10985 -550
rect 10955 -630 10985 -600
rect 10955 -680 10985 -650
rect 11040 -530 11070 -500
rect 11040 -580 11070 -550
rect 11040 -630 11070 -600
rect 11040 -680 11070 -650
rect 11125 -530 11155 -500
rect 11125 -580 11155 -550
rect 11125 -630 11155 -600
rect 11125 -680 11155 -650
rect 11210 -530 11240 -500
rect 11210 -580 11240 -550
rect 11210 -630 11240 -600
rect 11210 -680 11240 -650
rect 11295 -530 11325 -500
rect 11295 -580 11325 -550
rect 11295 -630 11325 -600
rect 11295 -680 11325 -650
rect 11380 -530 11410 -500
rect 11380 -580 11410 -550
rect 11380 -630 11410 -600
rect 11380 -680 11410 -650
rect 11465 -530 11495 -500
rect 11465 -580 11495 -550
rect 11465 -630 11495 -600
rect 11465 -680 11495 -650
rect 11550 -530 11580 -500
rect 11550 -580 11580 -550
rect 11550 -630 11580 -600
rect 11550 -680 11580 -650
rect 11635 -530 11665 -500
rect 11635 -580 11665 -550
rect 11635 -630 11665 -600
rect 11635 -680 11665 -650
rect 11720 -530 11750 -500
rect 11720 -580 11750 -550
rect 11720 -630 11750 -600
rect 11720 -680 11750 -650
rect 11805 -530 11835 -500
rect 11805 -580 11835 -550
rect 11805 -630 11835 -600
rect 11805 -680 11835 -650
rect 11890 -530 11920 -500
rect 11890 -580 11920 -550
rect 11890 -630 11920 -600
rect 11890 -680 11920 -650
rect 11975 -530 12005 -500
rect 11975 -580 12005 -550
rect 11975 -630 12005 -600
rect 11975 -680 12005 -650
rect 12060 -530 12090 -500
rect 12060 -580 12090 -550
rect 12060 -630 12090 -600
rect 12060 -680 12090 -650
rect 12145 -530 12175 -500
rect 12145 -580 12175 -550
rect 12145 -630 12175 -600
rect 12145 -680 12175 -650
rect 12230 -530 12260 -500
rect 12230 -580 12260 -550
rect 12230 -630 12260 -600
rect 12230 -680 12260 -650
rect 12315 -530 12345 -500
rect 12315 -580 12345 -550
rect 12315 -630 12345 -600
rect 12315 -680 12345 -650
rect 12400 -530 12430 -500
rect 12400 -580 12430 -550
rect 12400 -630 12430 -600
rect 12400 -680 12430 -650
rect 12485 -530 12515 -500
rect 12485 -580 12515 -550
rect 12485 -630 12515 -600
rect 12485 -680 12515 -650
rect 12570 -530 12600 -500
rect 12570 -580 12600 -550
rect 12570 -630 12600 -600
rect 12570 -680 12600 -650
rect 12655 -530 12685 -500
rect 12655 -580 12685 -550
rect 12655 -630 12685 -600
rect 12655 -680 12685 -650
rect 12740 -530 12770 -500
rect 12740 -580 12770 -550
rect 12740 -630 12770 -600
rect 12740 -680 12770 -650
rect 12825 -530 12855 -500
rect 12825 -580 12855 -550
rect 12825 -630 12855 -600
rect 12825 -680 12855 -650
rect 12910 -530 12940 -500
rect 12910 -580 12940 -550
rect 12910 -630 12940 -600
rect 12910 -680 12940 -650
rect 12995 -530 13025 -500
rect 12995 -580 13025 -550
rect 12995 -630 13025 -600
rect 12995 -680 13025 -650
rect 13080 -530 13110 -500
rect 13080 -580 13110 -550
rect 13080 -630 13110 -600
rect 13080 -680 13110 -650
rect 13165 -530 13195 -500
rect 13165 -580 13195 -550
rect 13165 -630 13195 -600
rect 13165 -680 13195 -650
rect 13250 -530 13280 -500
rect 13250 -580 13280 -550
rect 13250 -630 13280 -600
rect 13250 -680 13280 -650
rect 13335 -530 13365 -500
rect 13335 -580 13365 -550
rect 13335 -630 13365 -600
rect 13335 -680 13365 -650
rect 13420 -530 13450 -500
rect 13420 -580 13450 -550
rect 13420 -630 13450 -600
rect 13420 -680 13450 -650
rect 13505 -530 13535 -500
rect 13505 -580 13535 -550
rect 13505 -630 13535 -600
rect 13505 -680 13535 -650
rect 13590 -530 13620 -500
rect 13590 -580 13620 -550
rect 13590 -630 13620 -600
rect 13590 -680 13620 -650
rect 13675 -530 13705 -500
rect 13675 -580 13705 -550
rect 13675 -630 13705 -600
rect 13675 -680 13705 -650
rect 13760 -530 13790 -500
rect 13760 -580 13790 -550
rect 13760 -630 13790 -600
rect 13760 -680 13790 -650
rect 13845 -530 13875 -500
rect 13845 -580 13875 -550
rect 13845 -630 13875 -600
rect 13845 -680 13875 -650
rect 13930 -530 13960 -500
rect 13930 -580 13960 -550
rect 13930 -630 13960 -600
rect 13930 -680 13960 -650
rect 14015 -530 14045 -500
rect 14015 -580 14045 -550
rect 14015 -630 14045 -600
rect 14015 -680 14045 -650
rect 14100 -530 14130 -500
rect 14100 -580 14130 -550
rect 14100 -630 14130 -600
rect 14100 -680 14130 -650
rect 14185 -530 14215 -500
rect 14185 -580 14215 -550
rect 14185 -630 14215 -600
rect 14185 -680 14215 -650
rect 14270 -530 14300 -500
rect 14270 -580 14300 -550
rect 14270 -630 14300 -600
rect 14270 -680 14300 -650
rect 14355 -530 14385 -500
rect 14355 -580 14385 -550
rect 14355 -630 14385 -600
rect 14355 -680 14385 -650
rect 14440 -530 14470 -500
rect 14440 -580 14470 -550
rect 14440 -630 14470 -600
rect 14440 -680 14470 -650
rect 14525 -530 14555 -500
rect 14525 -580 14555 -550
rect 14525 -630 14555 -600
rect 14525 -680 14555 -650
rect 14610 -530 14640 -500
rect 14610 -580 14640 -550
rect 14610 -630 14640 -600
rect 14610 -680 14640 -650
rect 14695 -530 14725 -500
rect 14695 -580 14725 -550
rect 14695 -630 14725 -600
rect 14695 -680 14725 -650
rect 14780 -530 14810 -500
rect 14780 -580 14810 -550
rect 14780 -630 14810 -600
rect 14780 -680 14810 -650
rect 14865 -530 14895 -500
rect 14865 -580 14895 -550
rect 14865 -630 14895 -600
rect 14865 -680 14895 -650
rect 14950 -530 14980 -500
rect 14950 -580 14980 -550
rect 14950 -630 14980 -600
rect 14950 -680 14980 -650
rect 15035 -530 15065 -500
rect 15035 -580 15065 -550
rect 15035 -630 15065 -600
rect 15035 -680 15065 -650
rect 15120 -530 15150 -500
rect 15120 -580 15150 -550
rect 15120 -630 15150 -600
rect 15120 -680 15150 -650
rect 15205 -530 15235 -500
rect 15205 -580 15235 -550
rect 15205 -630 15235 -600
rect 15205 -680 15235 -650
rect 15290 -530 15320 -500
rect 15290 -580 15320 -550
rect 15290 -630 15320 -600
rect 15290 -680 15320 -650
rect 15375 -530 15405 -500
rect 15375 -580 15405 -550
rect 15375 -630 15405 -600
rect 15375 -680 15405 -650
rect 15460 -530 15490 -500
rect 15460 -580 15490 -550
rect 15460 -630 15490 -600
rect 15460 -680 15490 -650
rect 15545 -530 15575 -500
rect 15545 -580 15575 -550
rect 15545 -630 15575 -600
rect 15545 -680 15575 -650
rect 15630 -530 15660 -500
rect 15630 -580 15660 -550
rect 15630 -630 15660 -600
rect 15630 -680 15660 -650
rect 15715 -530 15745 -500
rect 15715 -580 15745 -550
rect 15715 -630 15745 -600
rect 15715 -680 15745 -650
rect 15800 -530 15830 -500
rect 15800 -580 15830 -550
rect 15800 -630 15830 -600
rect 15800 -680 15830 -650
rect 15885 -530 15915 -500
rect 15885 -580 15915 -550
rect 15885 -630 15915 -600
rect 15885 -680 15915 -650
rect 15970 -530 16000 -500
rect 15970 -580 16000 -550
rect 15970 -630 16000 -600
rect 15970 -680 16000 -650
rect 16055 -530 16085 -500
rect 16055 -580 16085 -550
rect 16055 -630 16085 -600
rect 16055 -680 16085 -650
rect 16140 -530 16170 -500
rect 16140 -580 16170 -550
rect 16140 -630 16170 -600
rect 16140 -680 16170 -650
rect 16225 -530 16255 -500
rect 16225 -580 16255 -550
rect 16225 -630 16255 -600
rect 16225 -680 16255 -650
rect 16310 -530 16340 -500
rect 16310 -580 16340 -550
rect 16310 -630 16340 -600
rect 16310 -680 16340 -650
rect 16395 -530 16425 -500
rect 16395 -580 16425 -550
rect 16395 -630 16425 -600
rect 16395 -680 16425 -650
rect 16480 -530 16510 -500
rect 16480 -580 16510 -550
rect 16480 -630 16510 -600
rect 16480 -680 16510 -650
rect 16565 -530 16595 -500
rect 16565 -580 16595 -550
rect 16565 -630 16595 -600
rect 16565 -680 16595 -650
rect 16650 -530 16680 -500
rect 16650 -580 16680 -550
rect 16650 -630 16680 -600
rect 16650 -680 16680 -650
rect 16735 -530 16765 -500
rect 16735 -580 16765 -550
rect 16735 -630 16765 -600
rect 16735 -680 16765 -650
rect 16820 -530 16850 -500
rect 16820 -580 16850 -550
rect 16820 -630 16850 -600
rect 16820 -680 16850 -650
rect 16905 -530 16935 -500
rect 16905 -580 16935 -550
rect 16905 -630 16935 -600
rect 16905 -680 16935 -650
rect 16990 -530 17020 -500
rect 16990 -580 17020 -550
rect 16990 -630 17020 -600
rect 16990 -680 17020 -650
rect 17075 -530 17105 -500
rect 17075 -580 17105 -550
rect 17075 -630 17105 -600
rect 17075 -680 17105 -650
rect 17160 -530 17190 -500
rect 17160 -580 17190 -550
rect 17160 -630 17190 -600
rect 17160 -680 17190 -650
rect 17245 -530 17275 -500
rect 17245 -580 17275 -550
rect 17245 -630 17275 -600
rect 17245 -680 17275 -650
rect 17330 -530 17360 -500
rect 17330 -580 17360 -550
rect 17330 -630 17360 -600
rect 17330 -680 17360 -650
rect 17415 -530 17445 -500
rect 17415 -580 17445 -550
rect 17415 -630 17445 -600
rect 17415 -680 17445 -650
rect 17500 -530 17530 -500
rect 17500 -580 17530 -550
rect 17500 -630 17530 -600
rect 17500 -680 17530 -650
rect 17585 -530 17615 -500
rect 17585 -580 17615 -550
rect 17585 -630 17615 -600
rect 17585 -680 17615 -650
rect 17670 -530 17700 -500
rect 17670 -580 17700 -550
rect 17670 -630 17700 -600
rect 17670 -680 17700 -650
rect 17755 -530 17785 -500
rect 17755 -580 17785 -550
rect 17755 -630 17785 -600
rect 17755 -680 17785 -650
rect 17840 -530 17870 -500
rect 17840 -580 17870 -550
rect 17840 -630 17870 -600
rect 17840 -680 17870 -650
rect 17925 -530 17955 -500
rect 17925 -580 17955 -550
rect 17925 -630 17955 -600
rect 17925 -680 17955 -650
rect 18010 -530 18040 -500
rect 18010 -580 18040 -550
rect 18010 -630 18040 -600
rect 18010 -680 18040 -650
rect 18095 -530 18125 -500
rect 18095 -580 18125 -550
rect 18095 -630 18125 -600
rect 18095 -680 18125 -650
rect 18180 -530 18210 -500
rect 18180 -580 18210 -550
rect 18180 -630 18210 -600
rect 18180 -680 18210 -650
rect 18265 -530 18295 -500
rect 18265 -580 18295 -550
rect 18265 -630 18295 -600
rect 18265 -680 18295 -650
rect 18350 -530 18380 -500
rect 18350 -580 18380 -550
rect 18350 -630 18380 -600
rect 18350 -680 18380 -650
rect 18435 -530 18465 -500
rect 18435 -580 18465 -550
rect 18435 -630 18465 -600
rect 18435 -680 18465 -650
rect 18520 -530 18550 -500
rect 18520 -580 18550 -550
rect 18520 -630 18550 -600
rect 18520 -680 18550 -650
rect 18605 -530 18635 -500
rect 18605 -580 18635 -550
rect 18605 -630 18635 -600
rect 18605 -680 18635 -650
rect 18690 -530 18720 -500
rect 18690 -580 18720 -550
rect 18690 -630 18720 -600
rect 18690 -680 18720 -650
rect 18775 -530 18805 -500
rect 18775 -580 18805 -550
rect 18775 -630 18805 -600
rect 18775 -680 18805 -650
rect 18860 -530 18890 -500
rect 18860 -580 18890 -550
rect 18860 -630 18890 -600
rect 18860 -680 18890 -650
rect 18945 -530 18975 -500
rect 18945 -580 18975 -550
rect 18945 -630 18975 -600
rect 18945 -680 18975 -650
rect 19030 -530 19060 -500
rect 19030 -580 19060 -550
rect 19030 -630 19060 -600
rect 19030 -680 19060 -650
rect 19115 -530 19145 -500
rect 19115 -580 19145 -550
rect 19115 -630 19145 -600
rect 19115 -680 19145 -650
rect 19200 -530 19230 -500
rect 19200 -580 19230 -550
rect 19200 -630 19230 -600
rect 19200 -680 19230 -650
rect 19285 -530 19315 -500
rect 19285 -580 19315 -550
rect 19285 -630 19315 -600
rect 19285 -680 19315 -650
rect 19370 -530 19400 -500
rect 19370 -580 19400 -550
rect 19370 -630 19400 -600
rect 19370 -680 19400 -650
rect 19455 -530 19485 -500
rect 19455 -580 19485 -550
rect 19455 -630 19485 -600
rect 19455 -680 19485 -650
rect 19540 -530 19570 -500
rect 19540 -580 19570 -550
rect 19540 -630 19570 -600
rect 19540 -680 19570 -650
rect 19625 -530 19655 -500
rect 19625 -580 19655 -550
rect 19625 -630 19655 -600
rect 19625 -680 19655 -650
rect 19710 -530 19740 -500
rect 19710 -580 19740 -550
rect 19710 -630 19740 -600
rect 19710 -680 19740 -650
rect 19795 -530 19825 -500
rect 19795 -580 19825 -550
rect 19795 -630 19825 -600
rect 19795 -680 19825 -650
rect 19880 -530 19910 -500
rect 19880 -580 19910 -550
rect 19880 -630 19910 -600
rect 19880 -680 19910 -650
rect 19965 -530 19995 -500
rect 19965 -580 19995 -550
rect 19965 -630 19995 -600
rect 19965 -680 19995 -650
rect 20050 -530 20080 -500
rect 20050 -580 20080 -550
rect 20050 -630 20080 -600
rect 20050 -680 20080 -650
rect 20135 -530 20165 -500
rect 20135 -580 20165 -550
rect 20135 -630 20165 -600
rect 20135 -680 20165 -650
rect 20220 -530 20250 -500
rect 20220 -580 20250 -550
rect 20220 -630 20250 -600
rect 20220 -680 20250 -650
rect 20305 -530 20335 -500
rect 20305 -580 20335 -550
rect 20305 -630 20335 -600
rect 20305 -680 20335 -650
rect 20390 -530 20420 -500
rect 20390 -580 20420 -550
rect 20390 -630 20420 -600
rect 20390 -680 20420 -650
rect 20475 -530 20505 -500
rect 20475 -580 20505 -550
rect 20475 -630 20505 -600
rect 20475 -680 20505 -650
rect 20560 -530 20590 -500
rect 20560 -580 20590 -550
rect 20560 -630 20590 -600
rect 20560 -680 20590 -650
rect 20645 -530 20675 -500
rect 20645 -580 20675 -550
rect 20645 -630 20675 -600
rect 20645 -680 20675 -650
rect 20730 -530 20760 -500
rect 20730 -580 20760 -550
rect 20730 -630 20760 -600
rect 20730 -680 20760 -650
rect 20815 -530 20845 -500
rect 20815 -580 20845 -550
rect 20815 -630 20845 -600
rect 20815 -680 20845 -650
rect 20900 -530 20930 -500
rect 20900 -580 20930 -550
rect 20900 -630 20930 -600
rect 20900 -680 20930 -650
rect 20985 -530 21015 -500
rect 20985 -580 21015 -550
rect 20985 -630 21015 -600
rect 20985 -680 21015 -650
rect 21070 -530 21100 -500
rect 21070 -580 21100 -550
rect 21070 -630 21100 -600
rect 21070 -680 21100 -650
rect 21155 -530 21185 -500
rect 21155 -580 21185 -550
rect 21155 -630 21185 -600
rect 21155 -680 21185 -650
rect 21240 -530 21270 -500
rect 21240 -580 21270 -550
rect 21240 -630 21270 -600
rect 21240 -680 21270 -650
rect 21325 -530 21355 -500
rect 21325 -580 21355 -550
rect 21325 -630 21355 -600
rect 21325 -680 21355 -650
rect 21410 -530 21440 -500
rect 21410 -580 21440 -550
rect 21410 -630 21440 -600
rect 21410 -680 21440 -650
rect 21495 -530 21525 -500
rect 21495 -580 21525 -550
rect 21495 -630 21525 -600
rect 21495 -680 21525 -650
rect 21580 -530 21610 -500
rect 21580 -580 21610 -550
rect 21580 -630 21610 -600
rect 21580 -680 21610 -650
rect 21665 -530 21695 -500
rect 21665 -580 21695 -550
rect 21665 -630 21695 -600
rect 21665 -680 21695 -650
rect 21750 -530 21780 -500
rect 21750 -580 21780 -550
rect 21750 -630 21780 -600
rect 21750 -680 21780 -650
rect 21835 -530 21865 -500
rect 21835 -580 21865 -550
rect 21835 -630 21865 -600
rect 21835 -680 21865 -650
rect 21920 -530 21950 -500
rect 21920 -580 21950 -550
rect 21920 -630 21950 -600
rect 21920 -680 21950 -650
rect 22005 -530 22035 -500
rect 22005 -580 22035 -550
rect 22005 -630 22035 -600
rect 22005 -680 22035 -650
rect 22090 -530 22120 -500
rect 22090 -580 22120 -550
rect 22090 -630 22120 -600
rect 22090 -680 22120 -650
rect 22175 -530 22205 -500
rect 22175 -580 22205 -550
rect 22175 -630 22205 -600
rect 22175 -680 22205 -650
rect 22260 -530 22290 -500
rect 22260 -580 22290 -550
rect 22260 -630 22290 -600
rect 22260 -680 22290 -650
rect 22345 -530 22375 -500
rect 22345 -580 22375 -550
rect 22345 -630 22375 -600
rect 22345 -680 22375 -650
rect 22430 -530 22460 -500
rect 22430 -580 22460 -550
rect 22430 -630 22460 -600
rect 22430 -680 22460 -650
rect 22515 -530 22545 -500
rect 22515 -580 22545 -550
rect 22515 -630 22545 -600
rect 22515 -680 22545 -650
rect 22600 -530 22630 -500
rect 22600 -580 22630 -550
rect 22600 -630 22630 -600
rect 22600 -680 22630 -650
rect 22685 -530 22715 -500
rect 22685 -580 22715 -550
rect 22685 -630 22715 -600
rect 22685 -680 22715 -650
rect 22770 -530 22800 -500
rect 22770 -580 22800 -550
rect 22770 -630 22800 -600
rect 22770 -680 22800 -650
rect 22855 -530 22885 -500
rect 22855 -580 22885 -550
rect 22855 -630 22885 -600
rect 22855 -680 22885 -650
rect 22940 -530 22970 -500
rect 22940 -580 22970 -550
rect 22940 -630 22970 -600
rect 22940 -680 22970 -650
rect 23025 -530 23055 -500
rect 23025 -580 23055 -550
rect 23025 -630 23055 -600
rect 23025 -680 23055 -650
rect 23110 -530 23140 -500
rect 23110 -580 23140 -550
rect 23110 -630 23140 -600
rect 23110 -680 23140 -650
rect 23195 -530 23225 -500
rect 23195 -580 23225 -550
rect 23195 -630 23225 -600
rect 23195 -680 23225 -650
rect 23280 -530 23310 -500
rect 23280 -580 23310 -550
rect 23280 -630 23310 -600
rect 23280 -680 23310 -650
rect 23365 -530 23395 -500
rect 23365 -580 23395 -550
rect 23365 -630 23395 -600
rect 23365 -680 23395 -650
rect 23450 -530 23480 -500
rect 23450 -580 23480 -550
rect 23450 -630 23480 -600
rect 23450 -680 23480 -650
rect 23535 -530 23565 -500
rect 23535 -580 23565 -550
rect 23535 -630 23565 -600
rect 23535 -680 23565 -650
rect 23620 -530 23650 -500
rect 23620 -580 23650 -550
rect 23620 -630 23650 -600
rect 23620 -680 23650 -650
rect 23705 -530 23735 -500
rect 23705 -580 23735 -550
rect 23705 -630 23735 -600
rect 23705 -680 23735 -650
rect 23790 -530 23820 -500
rect 23790 -580 23820 -550
rect 23790 -630 23820 -600
rect 23790 -680 23820 -650
rect 23875 -530 23905 -500
rect 23875 -580 23905 -550
rect 23875 -630 23905 -600
rect 23875 -680 23905 -650
rect 23960 -530 23990 -500
rect 23960 -580 23990 -550
rect 23960 -630 23990 -600
rect 23960 -680 23990 -650
rect 24045 -530 24075 -500
rect 24045 -580 24075 -550
rect 24045 -630 24075 -600
rect 24045 -680 24075 -650
rect 24130 -530 24160 -500
rect 24130 -580 24160 -550
rect 24130 -630 24160 -600
rect 24130 -680 24160 -650
rect 24215 -530 24245 -500
rect 24215 -580 24245 -550
rect 24215 -630 24245 -600
rect 24215 -680 24245 -650
rect 24300 -530 24330 -500
rect 24300 -580 24330 -550
rect 24300 -630 24330 -600
rect 24300 -680 24330 -650
rect 24385 -530 24415 -500
rect 24385 -580 24415 -550
rect 24385 -630 24415 -600
rect 24385 -680 24415 -650
rect 24470 -530 24500 -500
rect 24470 -580 24500 -550
rect 24470 -630 24500 -600
rect 24470 -680 24500 -650
rect 24555 -530 24585 -500
rect 24555 -580 24585 -550
rect 24555 -630 24585 -600
rect 24555 -680 24585 -650
rect 24640 -530 24670 -500
rect 24640 -580 24670 -550
rect 24640 -630 24670 -600
rect 24640 -680 24670 -650
rect 24725 -530 24755 -500
rect 24725 -580 24755 -550
rect 24725 -630 24755 -600
rect 24725 -680 24755 -650
rect 24810 -530 24840 -500
rect 24810 -580 24840 -550
rect 24810 -630 24840 -600
rect 24810 -680 24840 -650
rect 24895 -530 24925 -500
rect 24895 -580 24925 -550
rect 24895 -630 24925 -600
rect 24895 -680 24925 -650
rect 24980 -530 25010 -500
rect 24980 -580 25010 -550
rect 24980 -630 25010 -600
rect 24980 -680 25010 -650
rect 25065 -530 25095 -500
rect 25065 -580 25095 -550
rect 25065 -630 25095 -600
rect 25065 -680 25095 -650
rect 25150 -530 25180 -500
rect 25150 -580 25180 -550
rect 25150 -630 25180 -600
rect 25150 -680 25180 -650
rect 25235 -530 25265 -500
rect 25235 -580 25265 -550
rect 25235 -630 25265 -600
rect 25235 -680 25265 -650
rect 25320 -530 25350 -500
rect 25320 -580 25350 -550
rect 25320 -630 25350 -600
rect 25320 -680 25350 -650
rect 25405 -530 25435 -500
rect 25405 -580 25435 -550
rect 25405 -630 25435 -600
rect 25405 -680 25435 -650
rect 25490 -530 25520 -500
rect 25490 -580 25520 -550
rect 25490 -630 25520 -600
rect 25490 -680 25520 -650
rect 25575 -530 25605 -500
rect 25575 -580 25605 -550
rect 25575 -630 25605 -600
rect 25575 -680 25605 -650
rect 25660 -530 25690 -500
rect 25660 -580 25690 -550
rect 25660 -630 25690 -600
rect 25660 -680 25690 -650
rect 25745 -530 25775 -500
rect 25745 -580 25775 -550
rect 25745 -630 25775 -600
rect 25745 -680 25775 -650
rect 25830 -530 25860 -500
rect 25830 -580 25860 -550
rect 25830 -630 25860 -600
rect 25830 -680 25860 -650
rect 25915 -530 25945 -500
rect 25915 -580 25945 -550
rect 25915 -630 25945 -600
rect 25915 -680 25945 -650
rect 26000 -530 26030 -500
rect 26000 -580 26030 -550
rect 26000 -630 26030 -600
rect 26000 -680 26030 -650
rect 26085 -530 26115 -500
rect 26085 -580 26115 -550
rect 26085 -630 26115 -600
rect 26085 -680 26115 -650
rect 26170 -530 26200 -500
rect 26170 -580 26200 -550
rect 26170 -630 26200 -600
rect 26170 -680 26200 -650
rect 26255 -530 26285 -500
rect 26255 -580 26285 -550
rect 26255 -630 26285 -600
rect 26255 -680 26285 -650
rect 26340 -530 26370 -500
rect 26340 -580 26370 -550
rect 26340 -630 26370 -600
rect 26340 -680 26370 -650
rect 26425 -530 26455 -500
rect 26425 -580 26455 -550
rect 26425 -630 26455 -600
rect 26425 -680 26455 -650
rect 26510 -530 26540 -500
rect 26510 -580 26540 -550
rect 26510 -630 26540 -600
rect 26510 -680 26540 -650
rect 26595 -530 26625 -500
rect 26595 -580 26625 -550
rect 26595 -630 26625 -600
rect 26595 -680 26625 -650
rect 26680 -530 26710 -500
rect 26680 -580 26710 -550
rect 26680 -630 26710 -600
rect 26680 -680 26710 -650
rect 26765 -530 26795 -500
rect 26765 -580 26795 -550
rect 26765 -630 26795 -600
rect 26765 -680 26795 -650
rect 26850 -530 26880 -500
rect 26850 -580 26880 -550
rect 26850 -630 26880 -600
rect 26850 -680 26880 -650
rect 26935 -530 26965 -500
rect 26935 -580 26965 -550
rect 26935 -630 26965 -600
rect 26935 -680 26965 -650
rect 27020 -530 27050 -500
rect 27020 -580 27050 -550
rect 27020 -630 27050 -600
rect 27020 -680 27050 -650
rect 27105 -530 27135 -500
rect 27105 -580 27135 -550
rect 27105 -630 27135 -600
rect 27105 -680 27135 -650
rect 27190 -530 27220 -500
rect 27190 -580 27220 -550
rect 27190 -630 27220 -600
rect 27190 -680 27220 -650
rect 27275 -530 27305 -500
rect 27275 -580 27305 -550
rect 27275 -630 27305 -600
rect 27275 -680 27305 -650
rect 27360 -530 27390 -500
rect 27360 -580 27390 -550
rect 27360 -630 27390 -600
rect 27360 -680 27390 -650
rect 27445 -530 27475 -500
rect 27445 -580 27475 -550
rect 27445 -630 27475 -600
rect 27445 -680 27475 -650
rect 27530 -530 27560 -500
rect 27530 -580 27560 -550
rect 27530 -630 27560 -600
rect 27530 -680 27560 -650
rect 27615 -530 27645 -500
rect 27615 -580 27645 -550
rect 27615 -630 27645 -600
rect 27615 -680 27645 -650
rect 27700 -530 27730 -500
rect 27700 -580 27730 -550
rect 27700 -630 27730 -600
rect 27700 -680 27730 -650
rect 27785 -530 27815 -500
rect 27785 -580 27815 -550
rect 27785 -630 27815 -600
rect 27785 -680 27815 -650
rect 27870 -530 27900 -500
rect 27870 -580 27900 -550
rect 27870 -630 27900 -600
rect 27870 -680 27900 -650
rect 27955 -530 27985 -500
rect 27955 -580 27985 -550
rect 27955 -630 27985 -600
rect 27955 -680 27985 -650
rect 28040 -530 28070 -500
rect 28040 -580 28070 -550
rect 28040 -630 28070 -600
rect 28040 -680 28070 -650
rect 28125 -530 28155 -500
rect 28125 -580 28155 -550
rect 28125 -630 28155 -600
rect 28125 -680 28155 -650
rect 28210 -530 28240 -500
rect 28210 -580 28240 -550
rect 28210 -630 28240 -600
rect 28210 -680 28240 -650
rect 28295 -530 28325 -500
rect 28295 -580 28325 -550
rect 28295 -630 28325 -600
rect 28295 -680 28325 -650
rect 28380 -530 28410 -500
rect 28380 -580 28410 -550
rect 28380 -630 28410 -600
rect 28380 -680 28410 -650
rect 28465 -530 28495 -500
rect 28465 -580 28495 -550
rect 28465 -630 28495 -600
rect 28465 -680 28495 -650
rect 28550 -530 28580 -500
rect 28550 -580 28580 -550
rect 28550 -630 28580 -600
rect 28550 -680 28580 -650
rect 28635 -530 28665 -500
rect 28635 -580 28665 -550
rect 28635 -630 28665 -600
rect 28635 -680 28665 -650
rect 28720 -530 28750 -500
rect 28720 -580 28750 -550
rect 28720 -630 28750 -600
rect 28720 -680 28750 -650
rect 28805 -530 28835 -500
rect 28805 -580 28835 -550
rect 28805 -630 28835 -600
rect 28805 -680 28835 -650
rect 28890 -530 28920 -500
rect 28890 -580 28920 -550
rect 28890 -630 28920 -600
rect 28890 -680 28920 -650
rect 28975 -530 29005 -500
rect 28975 -580 29005 -550
rect 28975 -630 29005 -600
rect 28975 -680 29005 -650
rect 29060 -530 29090 -500
rect 29060 -580 29090 -550
rect 29060 -630 29090 -600
rect 29060 -680 29090 -650
rect 29145 -530 29175 -500
rect 29145 -580 29175 -550
rect 29145 -630 29175 -600
rect 29145 -680 29175 -650
rect 29230 -530 29260 -500
rect 29230 -580 29260 -550
rect 29230 -630 29260 -600
rect 29230 -680 29260 -650
rect 29315 -530 29345 -500
rect 29315 -580 29345 -550
rect 29315 -630 29345 -600
rect 29315 -680 29345 -650
rect 29400 -530 29430 -500
rect 29400 -580 29430 -550
rect 29400 -630 29430 -600
rect 29400 -680 29430 -650
rect 29485 -530 29515 -500
rect 29485 -580 29515 -550
rect 29485 -630 29515 -600
rect 29485 -680 29515 -650
rect 29570 -530 29600 -500
rect 29570 -580 29600 -550
rect 29570 -630 29600 -600
rect 29570 -680 29600 -650
rect 29655 -530 29685 -500
rect 29655 -580 29685 -550
rect 29655 -630 29685 -600
rect 29655 -680 29685 -650
rect 29740 -530 29770 -500
rect 29740 -580 29770 -550
rect 29740 -630 29770 -600
rect 29740 -680 29770 -650
rect 29825 -530 29855 -500
rect 29825 -580 29855 -550
rect 29825 -630 29855 -600
rect 29825 -680 29855 -650
rect 29910 -530 29940 -500
rect 29910 -580 29940 -550
rect 29910 -630 29940 -600
rect 29910 -680 29940 -650
rect 29995 -530 30025 -500
rect 29995 -580 30025 -550
rect 29995 -630 30025 -600
rect 29995 -680 30025 -650
rect 30080 -530 30110 -500
rect 30080 -580 30110 -550
rect 30080 -630 30110 -600
rect 30080 -680 30110 -650
rect 30165 -530 30195 -500
rect 30165 -580 30195 -550
rect 30165 -630 30195 -600
rect 30165 -680 30195 -650
rect 30250 -530 30280 -500
rect 30250 -580 30280 -550
rect 30250 -630 30280 -600
rect 30250 -680 30280 -650
rect 30335 -530 30365 -500
rect 30335 -580 30365 -550
rect 30335 -630 30365 -600
rect 30335 -680 30365 -650
rect 30420 -530 30450 -500
rect 30420 -580 30450 -550
rect 30420 -630 30450 -600
rect 30420 -680 30450 -650
rect 30505 -530 30535 -500
rect 30505 -580 30535 -550
rect 30505 -630 30535 -600
rect 30505 -680 30535 -650
rect 30590 -530 30620 -500
rect 30590 -580 30620 -550
rect 30590 -630 30620 -600
rect 30590 -680 30620 -650
rect 30675 -530 30705 -500
rect 30675 -580 30705 -550
rect 30675 -630 30705 -600
rect 30675 -680 30705 -650
rect 30760 -530 30790 -500
rect 30760 -580 30790 -550
rect 30760 -630 30790 -600
rect 30760 -680 30790 -650
rect 30845 -530 30875 -500
rect 30845 -580 30875 -550
rect 30845 -630 30875 -600
rect 30845 -680 30875 -650
rect 30930 -530 30960 -500
rect 30930 -580 30960 -550
rect 30930 -630 30960 -600
rect 30930 -680 30960 -650
rect 31015 -530 31045 -500
rect 31015 -580 31045 -550
rect 31015 -630 31045 -600
rect 31015 -680 31045 -650
rect 31100 -530 31130 -500
rect 31100 -580 31130 -550
rect 31100 -630 31130 -600
rect 31100 -680 31130 -650
rect 31185 -530 31215 -500
rect 31185 -580 31215 -550
rect 31185 -630 31215 -600
rect 31185 -680 31215 -650
rect 31270 -530 31300 -500
rect 31270 -580 31300 -550
rect 31270 -630 31300 -600
rect 31270 -680 31300 -650
rect 31355 -530 31385 -500
rect 31355 -580 31385 -550
rect 31355 -630 31385 -600
rect 31355 -680 31385 -650
rect 31440 -530 31470 -500
rect 31440 -580 31470 -550
rect 31440 -630 31470 -600
rect 31440 -680 31470 -650
rect 31525 -530 31555 -500
rect 31525 -580 31555 -550
rect 31525 -630 31555 -600
rect 31525 -680 31555 -650
rect 31610 -530 31640 -500
rect 31610 -580 31640 -550
rect 31610 -630 31640 -600
rect 31610 -680 31640 -650
rect 31695 -530 31725 -500
rect 31695 -580 31725 -550
rect 31695 -630 31725 -600
rect 31695 -680 31725 -650
rect 31780 -530 31810 -500
rect 31780 -580 31810 -550
rect 31780 -630 31810 -600
rect 31780 -680 31810 -650
rect 31865 -530 31895 -500
rect 31865 -580 31895 -550
rect 31865 -630 31895 -600
rect 31865 -680 31895 -650
rect 31950 -530 31980 -500
rect 31950 -580 31980 -550
rect 31950 -630 31980 -600
rect 31950 -680 31980 -650
rect 32035 -530 32065 -500
rect 32035 -580 32065 -550
rect 32035 -630 32065 -600
rect 32035 -680 32065 -650
rect 32120 -530 32150 -500
rect 32120 -580 32150 -550
rect 32120 -630 32150 -600
rect 32120 -680 32150 -650
rect 32205 -530 32235 -500
rect 32205 -580 32235 -550
rect 32205 -630 32235 -600
rect 32205 -680 32235 -650
rect 32290 -530 32320 -500
rect 32290 -580 32320 -550
rect 32290 -630 32320 -600
rect 32290 -680 32320 -650
rect 32375 -530 32405 -500
rect 32375 -580 32405 -550
rect 32375 -630 32405 -600
rect 32375 -680 32405 -650
rect 32460 -530 32490 -500
rect 32460 -580 32490 -550
rect 32460 -630 32490 -600
rect 32460 -680 32490 -650
rect 32545 -530 32575 -500
rect 32545 -580 32575 -550
rect 32545 -630 32575 -600
rect 32545 -680 32575 -650
rect 32630 -530 32660 -500
rect 32630 -580 32660 -550
rect 32630 -630 32660 -600
rect 32630 -680 32660 -650
rect 32715 -530 32745 -500
rect 32715 -580 32745 -550
rect 32715 -630 32745 -600
rect 32715 -680 32745 -650
rect 32800 -530 32830 -500
rect 32800 -580 32830 -550
rect 32800 -630 32830 -600
rect 32800 -680 32830 -650
rect 32885 -530 32915 -500
rect 32885 -580 32915 -550
rect 32885 -630 32915 -600
rect 32885 -680 32915 -650
rect 32970 -530 33000 -500
rect 32970 -580 33000 -550
rect 32970 -630 33000 -600
rect 32970 -680 33000 -650
rect 33055 -530 33085 -500
rect 33055 -580 33085 -550
rect 33055 -630 33085 -600
rect 33055 -680 33085 -650
rect 33140 -530 33170 -500
rect 33140 -580 33170 -550
rect 33140 -630 33170 -600
rect 33140 -680 33170 -650
rect 33225 -530 33255 -500
rect 33225 -580 33255 -550
rect 33225 -630 33255 -600
rect 33225 -680 33255 -650
rect 33310 -530 33340 -500
rect 33310 -580 33340 -550
rect 33310 -630 33340 -600
rect 33310 -680 33340 -650
rect 33395 -530 33425 -500
rect 33395 -580 33425 -550
rect 33395 -630 33425 -600
rect 33395 -680 33425 -650
rect 33480 -530 33510 -500
rect 33480 -580 33510 -550
rect 33480 -630 33510 -600
rect 33480 -680 33510 -650
rect 33565 -530 33595 -500
rect 33565 -580 33595 -550
rect 33565 -630 33595 -600
rect 33565 -680 33595 -650
rect 33650 -530 33680 -500
rect 33650 -580 33680 -550
rect 33650 -630 33680 -600
rect 33650 -680 33680 -650
rect 33735 -530 33765 -500
rect 33735 -580 33765 -550
rect 33735 -630 33765 -600
rect 33735 -680 33765 -650
rect 33820 -530 33850 -500
rect 33820 -580 33850 -550
rect 33820 -630 33850 -600
rect 33820 -680 33850 -650
rect 33905 -530 33935 -500
rect 33905 -580 33935 -550
rect 33905 -630 33935 -600
rect 33905 -680 33935 -650
rect 33990 -530 34020 -500
rect 33990 -580 34020 -550
rect 33990 -630 34020 -600
rect 33990 -680 34020 -650
rect 34075 -530 34105 -500
rect 34075 -580 34105 -550
rect 34075 -630 34105 -600
rect 34075 -680 34105 -650
rect 34160 -530 34190 -500
rect 34160 -580 34190 -550
rect 34160 -630 34190 -600
rect 34160 -680 34190 -650
rect 34245 -530 34275 -500
rect 34245 -580 34275 -550
rect 34245 -630 34275 -600
rect 34245 -680 34275 -650
rect 34330 -530 34360 -500
rect 34330 -580 34360 -550
rect 34330 -630 34360 -600
rect 34330 -680 34360 -650
rect 34415 -530 34445 -500
rect 34415 -580 34445 -550
rect 34415 -630 34445 -600
rect 34415 -680 34445 -650
rect 34500 -530 34530 -500
rect 34500 -580 34530 -550
rect 34500 -630 34530 -600
rect 34500 -680 34530 -650
rect 34585 -530 34615 -500
rect 34585 -580 34615 -550
rect 34585 -630 34615 -600
rect 34585 -680 34615 -650
rect 34670 -530 34700 -500
rect 34670 -580 34700 -550
rect 34670 -630 34700 -600
rect 34670 -680 34700 -650
rect 34755 -530 34785 -500
rect 34755 -580 34785 -550
rect 34755 -630 34785 -600
rect 34755 -680 34785 -650
rect 34840 -530 34870 -500
rect 34840 -580 34870 -550
rect 34840 -630 34870 -600
rect 34840 -680 34870 -650
rect 34925 -530 34955 -500
rect 34925 -580 34955 -550
rect 34925 -630 34955 -600
rect 34925 -680 34955 -650
rect 35010 -530 35040 -500
rect 35010 -580 35040 -550
rect 35010 -630 35040 -600
rect 35010 -680 35040 -650
rect 35095 -530 35125 -500
rect 35095 -580 35125 -550
rect 35095 -630 35125 -600
rect 35095 -680 35125 -650
rect 35180 -530 35210 -500
rect 35180 -580 35210 -550
rect 35180 -630 35210 -600
rect 35180 -680 35210 -650
rect 35265 -530 35295 -500
rect 35265 -580 35295 -550
rect 35265 -630 35295 -600
rect 35265 -680 35295 -650
rect 35350 -530 35380 -500
rect 35350 -580 35380 -550
rect 35350 -630 35380 -600
rect 35350 -680 35380 -650
rect 35435 -530 35465 -500
rect 35435 -580 35465 -550
rect 35435 -630 35465 -600
rect 35435 -680 35465 -650
rect 35520 -530 35550 -500
rect 35520 -580 35550 -550
rect 35520 -630 35550 -600
rect 35520 -680 35550 -650
rect 35605 -530 35635 -500
rect 35605 -580 35635 -550
rect 35605 -630 35635 -600
rect 35605 -680 35635 -650
rect 35690 -530 35720 -500
rect 35690 -580 35720 -550
rect 35690 -630 35720 -600
rect 35690 -680 35720 -650
rect 35775 -530 35805 -500
rect 35775 -580 35805 -550
rect 35775 -630 35805 -600
rect 35775 -680 35805 -650
rect 35860 -530 35890 -500
rect 35860 -580 35890 -550
rect 35860 -630 35890 -600
rect 35860 -680 35890 -650
rect 35945 -530 35975 -500
rect 35945 -580 35975 -550
rect 35945 -630 35975 -600
rect 35945 -680 35975 -650
rect 36030 -530 36060 -500
rect 36030 -580 36060 -550
rect 36030 -630 36060 -600
rect 36030 -680 36060 -650
rect 36115 -530 36145 -500
rect 36115 -580 36145 -550
rect 36115 -630 36145 -600
rect 36115 -680 36145 -650
rect 36200 -530 36230 -500
rect 36200 -580 36230 -550
rect 36200 -630 36230 -600
rect 36200 -680 36230 -650
rect 36285 -530 36315 -500
rect 36285 -580 36315 -550
rect 36285 -630 36315 -600
rect 36285 -680 36315 -650
rect 36370 -530 36400 -500
rect 36370 -580 36400 -550
rect 36370 -630 36400 -600
rect 36370 -680 36400 -650
rect 36455 -530 36485 -500
rect 36455 -580 36485 -550
rect 36455 -630 36485 -600
rect 36455 -680 36485 -650
rect 36540 -530 36570 -500
rect 36540 -580 36570 -550
rect 36540 -630 36570 -600
rect 36540 -680 36570 -650
rect 36625 -530 36655 -500
rect 36625 -580 36655 -550
rect 36625 -630 36655 -600
rect 36625 -680 36655 -650
rect 36710 -530 36740 -500
rect 36710 -580 36740 -550
rect 36710 -630 36740 -600
rect 36710 -680 36740 -650
rect 36795 -530 36825 -500
rect 36795 -580 36825 -550
rect 36795 -630 36825 -600
rect 36795 -680 36825 -650
rect 36880 -530 36910 -500
rect 36880 -580 36910 -550
rect 36880 -630 36910 -600
rect 36880 -680 36910 -650
rect 36965 -530 36995 -500
rect 36965 -580 36995 -550
rect 36965 -630 36995 -600
rect 36965 -680 36995 -650
rect 37050 -530 37080 -500
rect 37050 -580 37080 -550
rect 37050 -630 37080 -600
rect 37050 -680 37080 -650
rect 37135 -530 37165 -500
rect 37135 -580 37165 -550
rect 37135 -630 37165 -600
rect 37135 -680 37165 -650
rect 37220 -530 37250 -500
rect 37220 -580 37250 -550
rect 37220 -630 37250 -600
rect 37220 -680 37250 -650
rect 37305 -530 37335 -500
rect 37305 -580 37335 -550
rect 37305 -630 37335 -600
rect 37305 -680 37335 -650
rect 37390 -530 37420 -500
rect 37390 -580 37420 -550
rect 37390 -630 37420 -600
rect 37390 -680 37420 -650
rect 37475 -530 37505 -500
rect 37475 -580 37505 -550
rect 37475 -630 37505 -600
rect 37475 -680 37505 -650
rect 37560 -530 37590 -500
rect 37560 -580 37590 -550
rect 37560 -630 37590 -600
rect 37560 -680 37590 -650
rect 37645 -530 37675 -500
rect 37645 -580 37675 -550
rect 37645 -630 37675 -600
rect 37645 -680 37675 -650
rect 37730 -530 37760 -500
rect 37730 -580 37760 -550
rect 37730 -630 37760 -600
rect 37730 -680 37760 -650
rect 37815 -530 37845 -500
rect 37815 -580 37845 -550
rect 37815 -630 37845 -600
rect 37815 -680 37845 -650
rect 37900 -530 37930 -500
rect 37900 -580 37930 -550
rect 37900 -630 37930 -600
rect 37900 -680 37930 -650
rect 37985 -530 38015 -500
rect 37985 -580 38015 -550
rect 37985 -630 38015 -600
rect 37985 -680 38015 -650
rect 38070 -530 38100 -500
rect 38070 -580 38100 -550
rect 38070 -630 38100 -600
rect 38070 -680 38100 -650
rect 38155 -530 38185 -500
rect 38155 -580 38185 -550
rect 38155 -630 38185 -600
rect 38155 -680 38185 -650
rect 38240 -530 38270 -500
rect 38240 -580 38270 -550
rect 38240 -630 38270 -600
rect 38240 -680 38270 -650
rect 38325 -530 38355 -500
rect 38325 -580 38355 -550
rect 38325 -630 38355 -600
rect 38325 -680 38355 -650
rect 38410 -530 38440 -500
rect 38410 -580 38440 -550
rect 38410 -630 38440 -600
rect 38410 -680 38440 -650
rect 38495 -530 38525 -500
rect 38495 -580 38525 -550
rect 38495 -630 38525 -600
rect 38495 -680 38525 -650
rect 38580 -530 38610 -500
rect 38580 -580 38610 -550
rect 38580 -630 38610 -600
rect 38580 -680 38610 -650
rect 38665 -530 38695 -500
rect 38665 -580 38695 -550
rect 38665 -630 38695 -600
rect 38665 -680 38695 -650
rect 38750 -530 38780 -500
rect 38750 -580 38780 -550
rect 38750 -630 38780 -600
rect 38750 -680 38780 -650
rect 38835 -530 38865 -500
rect 38835 -580 38865 -550
rect 38835 -630 38865 -600
rect 38835 -680 38865 -650
rect 38920 -530 38950 -500
rect 38920 -580 38950 -550
rect 38920 -630 38950 -600
rect 38920 -680 38950 -650
rect 39005 -530 39035 -500
rect 39005 -580 39035 -550
rect 39005 -630 39035 -600
rect 39005 -680 39035 -650
rect 39090 -530 39120 -500
rect 39090 -580 39120 -550
rect 39090 -630 39120 -600
rect 39090 -680 39120 -650
rect 39175 -530 39205 -500
rect 39175 -580 39205 -550
rect 39175 -630 39205 -600
rect 39175 -680 39205 -650
rect 39260 -530 39290 -500
rect 39260 -580 39290 -550
rect 39260 -630 39290 -600
rect 39260 -680 39290 -650
rect 39345 -530 39375 -500
rect 39345 -580 39375 -550
rect 39345 -630 39375 -600
rect 39345 -680 39375 -650
rect 39430 -530 39460 -500
rect 39430 -580 39460 -550
rect 39430 -630 39460 -600
rect 39430 -680 39460 -650
rect 39515 -530 39545 -500
rect 39515 -580 39545 -550
rect 39515 -630 39545 -600
rect 39515 -680 39545 -650
rect 39600 -530 39630 -500
rect 39600 -580 39630 -550
rect 39600 -630 39630 -600
rect 39600 -680 39630 -650
rect 39685 -530 39715 -500
rect 39685 -580 39715 -550
rect 39685 -630 39715 -600
rect 39685 -680 39715 -650
rect 39770 -530 39800 -500
rect 39770 -580 39800 -550
rect 39770 -630 39800 -600
rect 39770 -680 39800 -650
rect 39855 -530 39885 -500
rect 39855 -580 39885 -550
rect 39855 -630 39885 -600
rect 39855 -680 39885 -650
rect 39940 -530 39970 -500
rect 39940 -580 39970 -550
rect 39940 -630 39970 -600
rect 39940 -680 39970 -650
rect 40025 -530 40055 -500
rect 40025 -580 40055 -550
rect 40025 -630 40055 -600
rect 40025 -680 40055 -650
rect 40110 -530 40140 -500
rect 40110 -580 40140 -550
rect 40110 -630 40140 -600
rect 40110 -680 40140 -650
rect 40195 -530 40225 -500
rect 40195 -580 40225 -550
rect 40195 -630 40225 -600
rect 40195 -680 40225 -650
rect 40280 -530 40310 -500
rect 40280 -580 40310 -550
rect 40280 -630 40310 -600
rect 40280 -680 40310 -650
rect 40365 -530 40395 -500
rect 40365 -580 40395 -550
rect 40365 -630 40395 -600
rect 40365 -680 40395 -650
rect 40450 -530 40480 -500
rect 40450 -580 40480 -550
rect 40450 -630 40480 -600
rect 40450 -680 40480 -650
rect 40535 -530 40565 -500
rect 40535 -580 40565 -550
rect 40535 -630 40565 -600
rect 40535 -680 40565 -650
rect 40620 -530 40650 -500
rect 40620 -580 40650 -550
rect 40620 -630 40650 -600
rect 40620 -680 40650 -650
rect 40705 -530 40735 -500
rect 40705 -580 40735 -550
rect 40705 -630 40735 -600
rect 40705 -680 40735 -650
rect 40790 -530 40820 -500
rect 40790 -580 40820 -550
rect 40790 -630 40820 -600
rect 40790 -680 40820 -650
rect 40875 -530 40905 -500
rect 40875 -580 40905 -550
rect 40875 -630 40905 -600
rect 40875 -680 40905 -650
rect 40960 -530 40990 -500
rect 40960 -580 40990 -550
rect 40960 -630 40990 -600
rect 40960 -680 40990 -650
rect 41045 -530 41075 -500
rect 41045 -580 41075 -550
rect 41045 -630 41075 -600
rect 41045 -680 41075 -650
rect 41130 -530 41160 -500
rect 41130 -580 41160 -550
rect 41130 -630 41160 -600
rect 41130 -680 41160 -650
rect 41215 -530 41245 -500
rect 41215 -580 41245 -550
rect 41215 -630 41245 -600
rect 41215 -680 41245 -650
rect 41300 -530 41330 -500
rect 41300 -580 41330 -550
rect 41300 -630 41330 -600
rect 41300 -680 41330 -650
rect 41385 -530 41415 -500
rect 41385 -580 41415 -550
rect 41385 -630 41415 -600
rect 41385 -680 41415 -650
rect 41470 -530 41500 -500
rect 41470 -580 41500 -550
rect 41470 -630 41500 -600
rect 41470 -680 41500 -650
rect 41555 -530 41585 -500
rect 41555 -580 41585 -550
rect 41555 -630 41585 -600
rect 41555 -680 41585 -650
rect 41640 -530 41670 -500
rect 41640 -580 41670 -550
rect 41640 -630 41670 -600
rect 41640 -680 41670 -650
rect 41725 -530 41755 -500
rect 41725 -580 41755 -550
rect 41725 -630 41755 -600
rect 41725 -680 41755 -650
rect 41810 -530 41840 -500
rect 41810 -580 41840 -550
rect 41810 -630 41840 -600
rect 41810 -680 41840 -650
rect 41895 -530 41925 -500
rect 41895 -580 41925 -550
rect 41895 -630 41925 -600
rect 41895 -680 41925 -650
rect 41980 -530 42010 -500
rect 41980 -580 42010 -550
rect 41980 -630 42010 -600
rect 41980 -680 42010 -650
rect 42065 -530 42095 -500
rect 42065 -580 42095 -550
rect 42065 -630 42095 -600
rect 42065 -680 42095 -650
rect 42150 -530 42180 -500
rect 42150 -580 42180 -550
rect 42150 -630 42180 -600
rect 42150 -680 42180 -650
rect 42235 -530 42265 -500
rect 42235 -580 42265 -550
rect 42235 -630 42265 -600
rect 42235 -680 42265 -650
rect 42320 -530 42350 -500
rect 42320 -580 42350 -550
rect 42320 -630 42350 -600
rect 42320 -680 42350 -650
rect 42405 -530 42435 -500
rect 42405 -580 42435 -550
rect 42405 -630 42435 -600
rect 42405 -680 42435 -650
rect 42490 -530 42520 -500
rect 42490 -580 42520 -550
rect 42490 -630 42520 -600
rect 42490 -680 42520 -650
rect 42575 -530 42605 -500
rect 42575 -580 42605 -550
rect 42575 -630 42605 -600
rect 42575 -680 42605 -650
rect 42660 -530 42690 -500
rect 42660 -580 42690 -550
rect 42660 -630 42690 -600
rect 42660 -680 42690 -650
rect 42745 -530 42775 -500
rect 42745 -580 42775 -550
rect 42745 -630 42775 -600
rect 42745 -680 42775 -650
rect 42830 -530 42860 -500
rect 42830 -580 42860 -550
rect 42830 -630 42860 -600
rect 42830 -680 42860 -650
rect 42915 -530 42945 -500
rect 42915 -580 42945 -550
rect 42915 -630 42945 -600
rect 42915 -680 42945 -650
rect 43000 -530 43030 -500
rect 43000 -580 43030 -550
rect 43000 -630 43030 -600
rect 43000 -680 43030 -650
rect 43085 -530 43115 -500
rect 43085 -580 43115 -550
rect 43085 -630 43115 -600
rect 43085 -680 43115 -650
rect 43170 -530 43200 -500
rect 43170 -580 43200 -550
rect 43170 -630 43200 -600
rect 43170 -680 43200 -650
rect 43255 -530 43285 -500
rect 43255 -580 43285 -550
rect 43255 -630 43285 -600
rect 43255 -680 43285 -650
rect 43340 -530 43370 -500
rect 43340 -580 43370 -550
rect 43340 -630 43370 -600
rect 43340 -680 43370 -650
rect 43425 -530 43455 -500
rect 43425 -580 43455 -550
rect 43425 -630 43455 -600
rect 43425 -680 43455 -650
rect 43510 -530 43540 -500
rect 43510 -580 43540 -550
rect 43510 -630 43540 -600
rect 43510 -680 43540 -650
rect 43595 -530 43625 -500
rect 43595 -580 43625 -550
rect 43595 -630 43625 -600
rect 43595 -680 43625 -650
<< poly >>
rect 65 215 80 230
rect 275 215 290 230
rect 360 215 375 230
rect 445 215 460 230
rect 530 215 545 230
rect 810 215 825 230
rect 895 215 910 230
rect 980 215 995 230
rect 1065 215 1080 230
rect 1150 215 1165 230
rect 1235 215 1250 230
rect 1320 215 1335 230
rect 1405 215 1420 230
rect 1490 215 1505 230
rect 1575 215 1590 230
rect 1660 215 1675 230
rect 1745 215 1760 230
rect 1830 215 1845 230
rect 1915 215 1930 230
rect 2000 215 2015 230
rect 2085 215 2100 230
rect 2320 215 2335 230
rect 2405 215 2420 230
rect 2490 215 2505 230
rect 2575 215 2590 230
rect 2660 215 2675 230
rect 2745 215 2760 230
rect 2830 215 2845 230
rect 2915 215 2930 230
rect 3000 215 3015 230
rect 3085 215 3100 230
rect 3170 215 3185 230
rect 3255 215 3270 230
rect 3340 215 3355 230
rect 3425 215 3440 230
rect 3510 215 3525 230
rect 3595 215 3610 230
rect 3680 215 3695 230
rect 3765 215 3780 230
rect 3850 215 3865 230
rect 3935 215 3950 230
rect 4020 215 4035 230
rect 4105 215 4120 230
rect 4190 215 4205 230
rect 4275 215 4290 230
rect 4360 215 4375 230
rect 4445 215 4460 230
rect 4530 215 4545 230
rect 4615 215 4630 230
rect 4700 215 4715 230
rect 4785 215 4800 230
rect 4870 215 4885 230
rect 4955 215 4970 230
rect 5040 215 5055 230
rect 5125 215 5140 230
rect 5210 215 5225 230
rect 5295 215 5310 230
rect 5380 215 5395 230
rect 5465 215 5480 230
rect 5550 215 5565 230
rect 5635 215 5650 230
rect 5720 215 5735 230
rect 5805 215 5820 230
rect 5890 215 5905 230
rect 5975 215 5990 230
rect 6060 215 6075 230
rect 6145 215 6160 230
rect 6230 215 6245 230
rect 6315 215 6330 230
rect 6400 215 6415 230
rect 6485 215 6500 230
rect 6570 215 6585 230
rect 6655 215 6670 230
rect 6740 215 6755 230
rect 6825 215 6840 230
rect 6910 215 6925 230
rect 6995 215 7010 230
rect 7080 215 7095 230
rect 7165 215 7180 230
rect 7250 215 7265 230
rect 7335 215 7350 230
rect 7420 215 7435 230
rect 7505 215 7520 230
rect 7590 215 7605 230
rect 7675 215 7690 230
rect 7910 215 7925 230
rect 7995 215 8010 230
rect 8080 215 8095 230
rect 8165 215 8180 230
rect 8250 215 8265 230
rect 8335 215 8350 230
rect 8420 215 8435 230
rect 8505 215 8520 230
rect 8590 215 8605 230
rect 8675 215 8690 230
rect 8760 215 8775 230
rect 8845 215 8860 230
rect 8930 215 8945 230
rect 9015 215 9030 230
rect 9100 215 9115 230
rect 9185 215 9200 230
rect 9270 215 9285 230
rect 9355 215 9370 230
rect 9440 215 9455 230
rect 9525 215 9540 230
rect 9610 215 9625 230
rect 9695 215 9710 230
rect 9780 215 9795 230
rect 9865 215 9880 230
rect 9950 215 9965 230
rect 10035 215 10050 230
rect 10120 215 10135 230
rect 10205 215 10220 230
rect 10290 215 10305 230
rect 10375 215 10390 230
rect 10460 215 10475 230
rect 10545 215 10560 230
rect 10630 215 10645 230
rect 10715 215 10730 230
rect 10800 215 10815 230
rect 10885 215 10900 230
rect 10970 215 10985 230
rect 11055 215 11070 230
rect 11140 215 11155 230
rect 11225 215 11240 230
rect 11310 215 11325 230
rect 11395 215 11410 230
rect 11480 215 11495 230
rect 11565 215 11580 230
rect 11650 215 11665 230
rect 11735 215 11750 230
rect 11820 215 11835 230
rect 11905 215 11920 230
rect 11990 215 12005 230
rect 12075 215 12090 230
rect 12160 215 12175 230
rect 12245 215 12260 230
rect 12330 215 12345 230
rect 12415 215 12430 230
rect 12500 215 12515 230
rect 12585 215 12600 230
rect 12670 215 12685 230
rect 12755 215 12770 230
rect 12840 215 12855 230
rect 12925 215 12940 230
rect 13010 215 13025 230
rect 13095 215 13110 230
rect 13180 215 13195 230
rect 13265 215 13280 230
rect 13350 215 13365 230
rect 13435 215 13450 230
rect 13520 215 13535 230
rect 13605 215 13620 230
rect 13690 215 13705 230
rect 13775 215 13790 230
rect 13860 215 13875 230
rect 13945 215 13960 230
rect 14030 215 14045 230
rect 14115 215 14130 230
rect 14200 215 14215 230
rect 14285 215 14300 230
rect 14370 215 14385 230
rect 14455 215 14470 230
rect 14540 215 14555 230
rect 14625 215 14640 230
rect 14710 215 14725 230
rect 14795 215 14810 230
rect 14880 215 14895 230
rect 14965 215 14980 230
rect 15050 215 15065 230
rect 15135 215 15150 230
rect 15220 215 15235 230
rect 15305 215 15320 230
rect 15390 215 15405 230
rect 15475 215 15490 230
rect 15560 215 15575 230
rect 15645 215 15660 230
rect 15730 215 15745 230
rect 15815 215 15830 230
rect 15900 215 15915 230
rect 15985 215 16000 230
rect 16070 215 16085 230
rect 16155 215 16170 230
rect 16240 215 16255 230
rect 16325 215 16340 230
rect 16410 215 16425 230
rect 16495 215 16510 230
rect 16580 215 16595 230
rect 16665 215 16680 230
rect 16750 215 16765 230
rect 16835 215 16850 230
rect 16920 215 16935 230
rect 17005 215 17020 230
rect 17090 215 17105 230
rect 17175 215 17190 230
rect 17260 215 17275 230
rect 17345 215 17360 230
rect 17430 215 17445 230
rect 17515 215 17530 230
rect 17600 215 17615 230
rect 17685 215 17700 230
rect 17770 215 17785 230
rect 17855 215 17870 230
rect 17940 215 17955 230
rect 18025 215 18040 230
rect 18110 215 18125 230
rect 18195 215 18210 230
rect 18280 215 18295 230
rect 18365 215 18380 230
rect 18450 215 18465 230
rect 18535 215 18550 230
rect 18620 215 18635 230
rect 18705 215 18720 230
rect 18790 215 18805 230
rect 18875 215 18890 230
rect 18960 215 18975 230
rect 19045 215 19060 230
rect 19130 215 19145 230
rect 19215 215 19230 230
rect 19300 215 19315 230
rect 19385 215 19400 230
rect 19470 215 19485 230
rect 19555 215 19570 230
rect 19640 215 19655 230
rect 19725 215 19740 230
rect 19810 215 19825 230
rect 19895 215 19910 230
rect 19980 215 19995 230
rect 20065 215 20080 230
rect 20150 215 20165 230
rect 20235 215 20250 230
rect 20320 215 20335 230
rect 20405 215 20420 230
rect 20490 215 20505 230
rect 20575 215 20590 230
rect 20660 215 20675 230
rect 20745 215 20760 230
rect 20830 215 20845 230
rect 20915 215 20930 230
rect 21000 215 21015 230
rect 21085 215 21100 230
rect 21170 215 21185 230
rect 21255 215 21270 230
rect 21340 215 21355 230
rect 21425 215 21440 230
rect 21510 215 21525 230
rect 21595 215 21610 230
rect 21680 215 21695 230
rect 21765 215 21780 230
rect 21850 215 21865 230
rect 21935 215 21950 230
rect 22020 215 22035 230
rect 22105 215 22120 230
rect 22190 215 22205 230
rect 22275 215 22290 230
rect 22360 215 22375 230
rect 22445 215 22460 230
rect 22530 215 22545 230
rect 22615 215 22630 230
rect 22700 215 22715 230
rect 22785 215 22800 230
rect 22870 215 22885 230
rect 22955 215 22970 230
rect 23040 215 23055 230
rect 23125 215 23140 230
rect 23210 215 23225 230
rect 23295 215 23310 230
rect 23380 215 23395 230
rect 23465 215 23480 230
rect 23550 215 23565 230
rect 23635 215 23650 230
rect 23720 215 23735 230
rect 23805 215 23820 230
rect 23890 215 23905 230
rect 23975 215 23990 230
rect 24060 215 24075 230
rect 24145 215 24160 230
rect 24230 215 24245 230
rect 24315 215 24330 230
rect 24400 215 24415 230
rect 24485 215 24500 230
rect 24570 215 24585 230
rect 24655 215 24670 230
rect 24740 215 24755 230
rect 24825 215 24840 230
rect 24910 215 24925 230
rect 24995 215 25010 230
rect 25080 215 25095 230
rect 25165 215 25180 230
rect 25250 215 25265 230
rect 25335 215 25350 230
rect 25420 215 25435 230
rect 25505 215 25520 230
rect 25590 215 25605 230
rect 25675 215 25690 230
rect 25760 215 25775 230
rect 25845 215 25860 230
rect 25930 215 25945 230
rect 26015 215 26030 230
rect 26100 215 26115 230
rect 26185 215 26200 230
rect 26270 215 26285 230
rect 26355 215 26370 230
rect 26440 215 26455 230
rect 26525 215 26540 230
rect 26610 215 26625 230
rect 26695 215 26710 230
rect 26780 215 26795 230
rect 26865 215 26880 230
rect 26950 215 26965 230
rect 27035 215 27050 230
rect 27120 215 27135 230
rect 27205 215 27220 230
rect 27290 215 27305 230
rect 27375 215 27390 230
rect 27460 215 27475 230
rect 27545 215 27560 230
rect 27630 215 27645 230
rect 27715 215 27730 230
rect 27800 215 27815 230
rect 27885 215 27900 230
rect 27970 215 27985 230
rect 28055 215 28070 230
rect 28140 215 28155 230
rect 28225 215 28240 230
rect 28310 215 28325 230
rect 28395 215 28410 230
rect 28480 215 28495 230
rect 28565 215 28580 230
rect 28650 215 28665 230
rect 28735 215 28750 230
rect 28820 215 28835 230
rect 28905 215 28920 230
rect 28990 215 29005 230
rect 29075 215 29090 230
rect 29160 215 29175 230
rect 29245 215 29260 230
rect 29330 215 29345 230
rect 29415 215 29430 230
rect 29500 215 29515 230
rect 29585 215 29600 230
rect 65 65 80 115
rect 25 55 80 65
rect 25 15 35 55
rect 65 15 80 55
rect 275 50 290 115
rect 360 50 375 115
rect 445 50 460 115
rect 530 50 545 115
rect 810 50 825 115
rect 895 50 910 115
rect 980 50 995 115
rect 1065 50 1080 115
rect 1150 50 1165 115
rect 1235 50 1250 115
rect 1320 50 1335 115
rect 1405 50 1420 115
rect 1490 50 1505 115
rect 1575 50 1590 115
rect 1660 50 1675 115
rect 1745 50 1760 115
rect 1830 50 1845 115
rect 1915 50 1930 115
rect 2000 50 2015 115
rect 2085 50 2100 115
rect 2320 50 2335 115
rect 2405 50 2420 115
rect 2490 50 2505 115
rect 2575 50 2590 115
rect 2660 50 2675 115
rect 2745 50 2760 115
rect 2830 50 2845 115
rect 2915 50 2930 115
rect 3000 50 3015 115
rect 3085 50 3100 115
rect 3170 50 3185 115
rect 3255 50 3270 115
rect 3340 50 3355 115
rect 3425 50 3440 115
rect 3510 50 3525 115
rect 3595 50 3610 115
rect 3680 50 3695 115
rect 3765 50 3780 115
rect 3850 50 3865 115
rect 3935 50 3950 115
rect 4020 50 4035 115
rect 4105 50 4120 115
rect 4190 50 4205 115
rect 4275 50 4290 115
rect 4360 50 4375 115
rect 4445 50 4460 115
rect 4530 50 4545 115
rect 4615 50 4630 115
rect 4700 50 4715 115
rect 4785 50 4800 115
rect 4870 50 4885 115
rect 4955 50 4970 115
rect 5040 50 5055 115
rect 5125 50 5140 115
rect 5210 50 5225 115
rect 5295 50 5310 115
rect 5380 50 5395 115
rect 5465 50 5480 115
rect 5550 50 5565 115
rect 5635 50 5650 115
rect 5720 50 5735 115
rect 5805 50 5820 115
rect 5890 50 5905 115
rect 5975 50 5990 115
rect 6060 50 6075 115
rect 6145 50 6160 115
rect 6230 50 6245 115
rect 6315 50 6330 115
rect 6400 50 6415 115
rect 6485 50 6500 115
rect 6570 50 6585 115
rect 6655 50 6670 115
rect 6740 50 6755 115
rect 6825 50 6840 115
rect 6910 50 6925 115
rect 6995 50 7010 115
rect 7080 50 7095 115
rect 7165 50 7180 115
rect 7250 50 7265 115
rect 7335 50 7350 115
rect 7420 50 7435 115
rect 7505 50 7520 115
rect 7590 50 7605 115
rect 7675 50 7690 115
rect 7910 50 7925 115
rect 7995 50 8010 115
rect 8080 50 8095 115
rect 8165 50 8180 115
rect 8250 50 8265 115
rect 8335 50 8350 115
rect 8420 50 8435 115
rect 8505 50 8520 115
rect 8590 50 8605 115
rect 8675 50 8690 115
rect 8760 50 8775 115
rect 8845 50 8860 115
rect 8930 50 8945 115
rect 9015 50 9030 115
rect 9100 50 9115 115
rect 9185 50 9200 115
rect 9270 50 9285 115
rect 9355 50 9370 115
rect 9440 50 9455 115
rect 9525 50 9540 115
rect 9610 50 9625 115
rect 9695 50 9710 115
rect 9780 50 9795 115
rect 9865 50 9880 115
rect 9950 50 9965 115
rect 10035 50 10050 115
rect 10120 50 10135 115
rect 10205 50 10220 115
rect 10290 50 10305 115
rect 10375 50 10390 115
rect 10460 50 10475 115
rect 10545 50 10560 115
rect 10630 50 10645 115
rect 10715 50 10730 115
rect 10800 50 10815 115
rect 10885 50 10900 115
rect 10970 50 10985 115
rect 11055 50 11070 115
rect 11140 50 11155 115
rect 11225 50 11240 115
rect 11310 50 11325 115
rect 11395 50 11410 115
rect 11480 50 11495 115
rect 11565 50 11580 115
rect 11650 50 11665 115
rect 11735 50 11750 115
rect 11820 50 11835 115
rect 11905 50 11920 115
rect 11990 50 12005 115
rect 12075 50 12090 115
rect 12160 50 12175 115
rect 12245 50 12260 115
rect 12330 50 12345 115
rect 12415 50 12430 115
rect 12500 50 12515 115
rect 12585 50 12600 115
rect 12670 50 12685 115
rect 12755 50 12770 115
rect 12840 50 12855 115
rect 12925 50 12940 115
rect 13010 50 13025 115
rect 13095 50 13110 115
rect 13180 50 13195 115
rect 13265 50 13280 115
rect 13350 50 13365 115
rect 13435 50 13450 115
rect 13520 50 13535 115
rect 13605 50 13620 115
rect 13690 50 13705 115
rect 13775 50 13790 115
rect 13860 50 13875 115
rect 13945 50 13960 115
rect 14030 50 14045 115
rect 14115 50 14130 115
rect 14200 50 14215 115
rect 14285 50 14300 115
rect 14370 50 14385 115
rect 14455 50 14470 115
rect 14540 50 14555 115
rect 14625 50 14640 115
rect 14710 50 14725 115
rect 14795 50 14810 115
rect 14880 50 14895 115
rect 14965 50 14980 115
rect 15050 50 15065 115
rect 15135 50 15150 115
rect 15220 50 15235 115
rect 15305 50 15320 115
rect 15390 50 15405 115
rect 15475 50 15490 115
rect 15560 50 15575 115
rect 15645 50 15660 115
rect 15730 50 15745 115
rect 15815 50 15830 115
rect 15900 50 15915 115
rect 15985 50 16000 115
rect 16070 50 16085 115
rect 16155 50 16170 115
rect 16240 50 16255 115
rect 16325 50 16340 115
rect 16410 50 16425 115
rect 16495 50 16510 115
rect 16580 50 16595 115
rect 16665 50 16680 115
rect 16750 50 16765 115
rect 16835 50 16850 115
rect 16920 50 16935 115
rect 17005 50 17020 115
rect 17090 50 17105 115
rect 17175 50 17190 115
rect 17260 50 17275 115
rect 17345 50 17360 115
rect 17430 50 17445 115
rect 17515 50 17530 115
rect 17600 50 17615 115
rect 17685 50 17700 115
rect 17770 50 17785 115
rect 17855 50 17870 115
rect 17940 50 17955 115
rect 18025 50 18040 115
rect 18110 50 18125 115
rect 18195 50 18210 115
rect 18280 50 18295 115
rect 18365 50 18380 115
rect 18450 50 18465 115
rect 18535 50 18550 115
rect 18620 50 18635 115
rect 18705 50 18720 115
rect 18790 50 18805 115
rect 18875 50 18890 115
rect 18960 50 18975 115
rect 19045 50 19060 115
rect 19130 50 19145 115
rect 19215 50 19230 115
rect 19300 50 19315 115
rect 19385 50 19400 115
rect 19470 50 19485 115
rect 19555 50 19570 115
rect 19640 50 19655 115
rect 19725 50 19740 115
rect 19810 50 19825 115
rect 19895 50 19910 115
rect 19980 50 19995 115
rect 20065 50 20080 115
rect 20150 50 20165 115
rect 20235 50 20250 115
rect 20320 50 20335 115
rect 20405 50 20420 115
rect 20490 50 20505 115
rect 20575 50 20590 115
rect 20660 50 20675 115
rect 20745 50 20760 115
rect 20830 50 20845 115
rect 20915 50 20930 115
rect 21000 50 21015 115
rect 21085 50 21100 115
rect 21170 50 21185 115
rect 21255 50 21270 115
rect 21340 50 21355 115
rect 21425 50 21440 115
rect 21510 50 21525 115
rect 21595 50 21610 115
rect 21680 50 21695 115
rect 21765 50 21780 115
rect 21850 50 21865 115
rect 21935 50 21950 115
rect 22020 50 22035 115
rect 22105 50 22120 115
rect 22190 50 22205 115
rect 22275 50 22290 115
rect 22360 50 22375 115
rect 22445 50 22460 115
rect 22530 50 22545 115
rect 22615 50 22630 115
rect 22700 50 22715 115
rect 22785 50 22800 115
rect 22870 50 22885 115
rect 22955 50 22970 115
rect 23040 50 23055 115
rect 23125 50 23140 115
rect 23210 50 23225 115
rect 23295 50 23310 115
rect 23380 50 23395 115
rect 23465 50 23480 115
rect 23550 50 23565 115
rect 23635 50 23650 115
rect 23720 50 23735 115
rect 23805 50 23820 115
rect 23890 50 23905 115
rect 23975 50 23990 115
rect 24060 50 24075 115
rect 24145 50 24160 115
rect 24230 50 24245 115
rect 24315 50 24330 115
rect 24400 50 24415 115
rect 24485 50 24500 115
rect 24570 50 24585 115
rect 24655 50 24670 115
rect 24740 50 24755 115
rect 24825 50 24840 115
rect 24910 50 24925 115
rect 24995 50 25010 115
rect 25080 50 25095 115
rect 25165 50 25180 115
rect 25250 50 25265 115
rect 25335 50 25350 115
rect 25420 50 25435 115
rect 25505 50 25520 115
rect 25590 50 25605 115
rect 25675 50 25690 115
rect 25760 50 25775 115
rect 25845 50 25860 115
rect 25930 50 25945 115
rect 26015 50 26030 115
rect 26100 50 26115 115
rect 26185 50 26200 115
rect 26270 50 26285 115
rect 26355 50 26370 115
rect 26440 50 26455 115
rect 26525 50 26540 115
rect 26610 50 26625 115
rect 26695 50 26710 115
rect 26780 50 26795 115
rect 26865 50 26880 115
rect 26950 50 26965 115
rect 27035 50 27050 115
rect 27120 50 27135 115
rect 27205 50 27220 115
rect 27290 50 27305 115
rect 27375 50 27390 115
rect 27460 50 27475 115
rect 27545 50 27560 115
rect 27630 50 27645 115
rect 27715 50 27730 115
rect 27800 50 27815 115
rect 27885 50 27900 115
rect 27970 50 27985 115
rect 28055 50 28070 115
rect 28140 50 28155 115
rect 28225 50 28240 115
rect 28310 50 28325 115
rect 28395 50 28410 115
rect 28480 50 28495 115
rect 28565 50 28580 115
rect 28650 50 28665 115
rect 28735 50 28750 115
rect 28820 50 28835 115
rect 28905 50 28920 115
rect 28990 50 29005 115
rect 29075 50 29090 115
rect 29160 50 29175 115
rect 29245 50 29260 115
rect 29330 50 29345 115
rect 29415 50 29430 115
rect 29500 50 29515 115
rect 29585 50 29600 115
rect 25 5 80 15
rect 65 -20 80 5
rect 275 -20 290 0
rect 360 -20 375 0
rect 445 -20 460 0
rect 530 -20 545 0
rect 810 -20 825 0
rect 895 -20 910 0
rect 980 -20 995 0
rect 1065 -20 1080 0
rect 1150 -20 1165 0
rect 1235 -20 1250 0
rect 1320 -20 1335 0
rect 1405 -20 1420 0
rect 1490 -20 1505 0
rect 1575 -20 1590 0
rect 1660 -20 1675 0
rect 1745 -20 1760 0
rect 1830 -20 1845 0
rect 1915 -20 1930 0
rect 2000 -20 2015 0
rect 2085 -20 2100 0
rect 2320 -20 2335 0
rect 2405 -20 2420 0
rect 2490 -20 2505 0
rect 2575 -20 2590 0
rect 2660 -20 2675 0
rect 2745 -20 2760 0
rect 2830 -20 2845 0
rect 2915 -20 2930 0
rect 3000 -20 3015 0
rect 3085 -20 3100 0
rect 3170 -20 3185 0
rect 3255 -20 3270 0
rect 3340 -20 3355 0
rect 3425 -20 3440 0
rect 3510 -20 3525 0
rect 3595 -20 3610 0
rect 3680 -20 3695 0
rect 3765 -20 3780 0
rect 3850 -20 3865 0
rect 3935 -20 3950 0
rect 4020 -20 4035 0
rect 4105 -20 4120 0
rect 4190 -20 4205 0
rect 4275 -20 4290 0
rect 4360 -20 4375 0
rect 4445 -20 4460 0
rect 4530 -20 4545 0
rect 4615 -20 4630 0
rect 4700 -20 4715 0
rect 4785 -20 4800 0
rect 4870 -20 4885 0
rect 4955 -20 4970 0
rect 5040 -20 5055 0
rect 5125 -20 5140 0
rect 5210 -20 5225 0
rect 5295 -20 5310 0
rect 5380 -20 5395 0
rect 5465 -20 5480 0
rect 5550 -20 5565 0
rect 5635 -20 5650 0
rect 5720 -20 5735 0
rect 5805 -20 5820 0
rect 5890 -20 5905 0
rect 5975 -20 5990 0
rect 6060 -20 6075 0
rect 6145 -20 6160 0
rect 6230 -20 6245 0
rect 6315 -20 6330 0
rect 6400 -20 6415 0
rect 6485 -20 6500 0
rect 6570 -20 6585 0
rect 6655 -20 6670 0
rect 6740 -20 6755 0
rect 6825 -20 6840 0
rect 6910 -20 6925 0
rect 6995 -20 7010 0
rect 7080 -20 7095 0
rect 7165 -20 7180 0
rect 7250 -20 7265 0
rect 7335 -20 7350 0
rect 7420 -20 7435 0
rect 7505 -20 7520 0
rect 7590 -20 7605 0
rect 7675 -20 7690 0
rect 7910 -20 7925 0
rect 7995 -20 8010 0
rect 8080 -20 8095 0
rect 8165 -20 8180 0
rect 8250 -20 8265 0
rect 8335 -20 8350 0
rect 8420 -20 8435 0
rect 8505 -20 8520 0
rect 8590 -20 8605 0
rect 8675 -20 8690 0
rect 8760 -20 8775 0
rect 8845 -20 8860 0
rect 8930 -20 8945 0
rect 9015 -20 9030 0
rect 9100 -20 9115 0
rect 9185 -20 9200 0
rect 9270 -20 9285 0
rect 9355 -20 9370 0
rect 9440 -20 9455 0
rect 9525 -20 9540 0
rect 9610 -20 9625 0
rect 9695 -20 9710 0
rect 9780 -20 9795 0
rect 9865 -20 9880 0
rect 9950 -20 9965 0
rect 10035 -20 10050 0
rect 10120 -20 10135 0
rect 10205 -20 10220 0
rect 10290 -20 10305 0
rect 10375 -20 10390 0
rect 10460 -20 10475 0
rect 10545 -20 10560 0
rect 10630 -20 10645 0
rect 10715 -20 10730 0
rect 10800 -20 10815 0
rect 10885 -20 10900 0
rect 10970 -20 10985 0
rect 11055 -20 11070 0
rect 11140 -20 11155 0
rect 11225 -20 11240 0
rect 11310 -20 11325 0
rect 11395 -20 11410 0
rect 11480 -20 11495 0
rect 11565 -20 11580 0
rect 11650 -20 11665 0
rect 11735 -20 11750 0
rect 11820 -20 11835 0
rect 11905 -20 11920 0
rect 11990 -20 12005 0
rect 12075 -20 12090 0
rect 12160 -20 12175 0
rect 12245 -20 12260 0
rect 12330 -20 12345 0
rect 12415 -20 12430 0
rect 12500 -20 12515 0
rect 12585 -20 12600 0
rect 12670 -20 12685 0
rect 12755 -20 12770 0
rect 12840 -20 12855 0
rect 12925 -20 12940 0
rect 13010 -20 13025 0
rect 13095 -20 13110 0
rect 13180 -20 13195 0
rect 13265 -20 13280 0
rect 13350 -20 13365 0
rect 13435 -20 13450 0
rect 13520 -20 13535 0
rect 13605 -20 13620 0
rect 13690 -20 13705 0
rect 13775 -20 13790 0
rect 13860 -20 13875 0
rect 13945 -20 13960 0
rect 14030 -20 14045 0
rect 14115 -20 14130 0
rect 14200 -20 14215 0
rect 14285 -20 14300 0
rect 14370 -20 14385 0
rect 14455 -20 14470 0
rect 14540 -20 14555 0
rect 14625 -20 14640 0
rect 14710 -20 14725 0
rect 14795 -20 14810 0
rect 14880 -20 14895 0
rect 14965 -20 14980 0
rect 15050 -20 15065 0
rect 15135 -20 15150 0
rect 15220 -20 15235 0
rect 15305 -20 15320 0
rect 15390 -20 15405 0
rect 15475 -20 15490 0
rect 15560 -20 15575 0
rect 15645 -20 15660 0
rect 15730 -20 15745 0
rect 15815 -20 15830 0
rect 15900 -20 15915 0
rect 15985 -20 16000 0
rect 16070 -20 16085 0
rect 16155 -20 16170 0
rect 16240 -20 16255 0
rect 16325 -20 16340 0
rect 16410 -20 16425 0
rect 16495 -20 16510 0
rect 16580 -20 16595 0
rect 16665 -20 16680 0
rect 16750 -20 16765 0
rect 16835 -20 16850 0
rect 16920 -20 16935 0
rect 17005 -20 17020 0
rect 17090 -20 17105 0
rect 17175 -20 17190 0
rect 17260 -20 17275 0
rect 17345 -20 17360 0
rect 17430 -20 17445 0
rect 17515 -20 17530 0
rect 17600 -20 17615 0
rect 17685 -20 17700 0
rect 17770 -20 17785 0
rect 17855 -20 17870 0
rect 17940 -20 17955 0
rect 18025 -20 18040 0
rect 18110 -20 18125 0
rect 18195 -20 18210 0
rect 18280 -20 18295 0
rect 18365 -20 18380 0
rect 18450 -20 18465 0
rect 18535 -20 18550 0
rect 18620 -20 18635 0
rect 18705 -20 18720 0
rect 18790 -20 18805 0
rect 18875 -20 18890 0
rect 18960 -20 18975 0
rect 19045 -20 19060 0
rect 19130 -20 19145 0
rect 19215 -20 19230 0
rect 19300 -20 19315 0
rect 19385 -20 19400 0
rect 19470 -20 19485 0
rect 19555 -20 19570 0
rect 19640 -20 19655 0
rect 19725 -20 19740 0
rect 19810 -20 19825 0
rect 19895 -20 19910 0
rect 19980 -20 19995 0
rect 20065 -20 20080 0
rect 20150 -20 20165 0
rect 20235 -20 20250 0
rect 20320 -20 20335 0
rect 20405 -20 20420 0
rect 20490 -20 20505 0
rect 20575 -20 20590 0
rect 20660 -20 20675 0
rect 20745 -20 20760 0
rect 20830 -20 20845 0
rect 20915 -20 20930 0
rect 21000 -20 21015 0
rect 21085 -20 21100 0
rect 21170 -20 21185 0
rect 21255 -20 21270 0
rect 21340 -20 21355 0
rect 21425 -20 21440 0
rect 21510 -20 21525 0
rect 21595 -20 21610 0
rect 21680 -20 21695 0
rect 21765 -20 21780 0
rect 21850 -20 21865 0
rect 21935 -20 21950 0
rect 22020 -20 22035 0
rect 22105 -20 22120 0
rect 22190 -20 22205 0
rect 22275 -20 22290 0
rect 22360 -20 22375 0
rect 22445 -20 22460 0
rect 22530 -20 22545 0
rect 22615 -20 22630 0
rect 22700 -20 22715 0
rect 22785 -20 22800 0
rect 22870 -20 22885 0
rect 22955 -20 22970 0
rect 23040 -20 23055 0
rect 23125 -20 23140 0
rect 23210 -20 23225 0
rect 23295 -20 23310 0
rect 23380 -20 23395 0
rect 23465 -20 23480 0
rect 23550 -20 23565 0
rect 23635 -20 23650 0
rect 23720 -20 23735 0
rect 23805 -20 23820 0
rect 23890 -20 23905 0
rect 23975 -20 23990 0
rect 24060 -20 24075 0
rect 24145 -20 24160 0
rect 24230 -20 24245 0
rect 24315 -20 24330 0
rect 24400 -20 24415 0
rect 24485 -20 24500 0
rect 24570 -20 24585 0
rect 24655 -20 24670 0
rect 24740 -20 24755 0
rect 24825 -20 24840 0
rect 24910 -20 24925 0
rect 24995 -20 25010 0
rect 25080 -20 25095 0
rect 25165 -20 25180 0
rect 25250 -20 25265 0
rect 25335 -20 25350 0
rect 25420 -20 25435 0
rect 25505 -20 25520 0
rect 25590 -20 25605 0
rect 25675 -20 25690 0
rect 25760 -20 25775 0
rect 25845 -20 25860 0
rect 25930 -20 25945 0
rect 26015 -20 26030 0
rect 26100 -20 26115 0
rect 26185 -20 26200 0
rect 26270 -20 26285 0
rect 26355 -20 26370 0
rect 26440 -20 26455 0
rect 26525 -20 26540 0
rect 26610 -20 26625 0
rect 26695 -20 26710 0
rect 26780 -20 26795 0
rect 26865 -20 26880 0
rect 26950 -20 26965 0
rect 27035 -20 27050 0
rect 27120 -20 27135 0
rect 27205 -20 27220 0
rect 27290 -20 27305 0
rect 27375 -20 27390 0
rect 27460 -20 27475 0
rect 27545 -20 27560 0
rect 27630 -20 27645 0
rect 27715 -20 27730 0
rect 27800 -20 27815 0
rect 27885 -20 27900 0
rect 27970 -20 27985 0
rect 28055 -20 28070 0
rect 28140 -20 28155 0
rect 28225 -20 28240 0
rect 28310 -20 28325 0
rect 28395 -20 28410 0
rect 28480 -20 28495 0
rect 28565 -20 28580 0
rect 28650 -20 28665 0
rect 28735 -20 28750 0
rect 28820 -20 28835 0
rect 28905 -20 28920 0
rect 28990 -20 29005 0
rect 29075 -20 29090 0
rect 29160 -20 29175 0
rect 29245 -20 29260 0
rect 29330 -20 29345 0
rect 29415 -20 29430 0
rect 29500 -20 29515 0
rect 29585 -20 29600 0
rect 255 -30 310 -20
rect 255 -60 265 -30
rect 300 -60 310 -30
rect 255 -70 310 -60
rect 340 -30 395 -20
rect 340 -60 350 -30
rect 385 -60 395 -30
rect 340 -70 395 -60
rect 425 -30 480 -20
rect 425 -60 435 -30
rect 470 -60 480 -30
rect 425 -70 480 -60
rect 510 -30 565 -20
rect 510 -60 520 -30
rect 555 -60 565 -30
rect 510 -70 565 -60
rect 790 -30 845 -20
rect 790 -60 800 -30
rect 835 -60 845 -30
rect 790 -70 845 -60
rect 875 -30 930 -20
rect 875 -60 885 -30
rect 920 -60 930 -30
rect 875 -70 930 -60
rect 960 -30 1015 -20
rect 960 -60 970 -30
rect 1005 -60 1015 -30
rect 960 -70 1015 -60
rect 1045 -30 1100 -20
rect 1045 -60 1055 -30
rect 1090 -60 1100 -30
rect 1045 -70 1100 -60
rect 1130 -30 1185 -20
rect 1130 -60 1140 -30
rect 1175 -60 1185 -30
rect 1130 -70 1185 -60
rect 1215 -30 1270 -20
rect 1215 -60 1225 -30
rect 1260 -60 1270 -30
rect 1215 -70 1270 -60
rect 1300 -30 1355 -20
rect 1300 -60 1310 -30
rect 1345 -60 1355 -30
rect 1300 -70 1355 -60
rect 1385 -30 1440 -20
rect 1385 -60 1395 -30
rect 1430 -60 1440 -30
rect 1385 -70 1440 -60
rect 1470 -30 1525 -20
rect 1470 -60 1480 -30
rect 1515 -60 1525 -30
rect 1470 -70 1525 -60
rect 1555 -30 1610 -20
rect 1555 -60 1565 -30
rect 1600 -60 1610 -30
rect 1555 -70 1610 -60
rect 1640 -30 1695 -20
rect 1640 -60 1650 -30
rect 1685 -60 1695 -30
rect 1640 -70 1695 -60
rect 1725 -30 1780 -20
rect 1725 -60 1735 -30
rect 1770 -60 1780 -30
rect 1725 -70 1780 -60
rect 1810 -30 1865 -20
rect 1810 -60 1820 -30
rect 1855 -60 1865 -30
rect 1810 -70 1865 -60
rect 1895 -30 1950 -20
rect 1895 -60 1905 -30
rect 1940 -60 1950 -30
rect 1895 -70 1950 -60
rect 1980 -30 2035 -20
rect 1980 -60 1990 -30
rect 2025 -60 2035 -30
rect 1980 -70 2035 -60
rect 2065 -30 2120 -20
rect 2065 -60 2075 -30
rect 2110 -60 2120 -30
rect 2065 -70 2120 -60
rect 2300 -30 2355 -20
rect 2300 -60 2310 -30
rect 2345 -60 2355 -30
rect 2300 -70 2355 -60
rect 2385 -30 2440 -20
rect 2385 -60 2395 -30
rect 2430 -60 2440 -30
rect 2385 -70 2440 -60
rect 2470 -30 2525 -20
rect 2470 -60 2480 -30
rect 2515 -60 2525 -30
rect 2470 -70 2525 -60
rect 2555 -30 2610 -20
rect 2555 -60 2565 -30
rect 2600 -60 2610 -30
rect 2555 -70 2610 -60
rect 2640 -30 2695 -20
rect 2640 -60 2650 -30
rect 2685 -60 2695 -30
rect 2640 -70 2695 -60
rect 2725 -30 2780 -20
rect 2725 -60 2735 -30
rect 2770 -60 2780 -30
rect 2725 -70 2780 -60
rect 2810 -30 2865 -20
rect 2810 -60 2820 -30
rect 2855 -60 2865 -30
rect 2810 -70 2865 -60
rect 2895 -30 2950 -20
rect 2895 -60 2905 -30
rect 2940 -60 2950 -30
rect 2895 -70 2950 -60
rect 2980 -30 3035 -20
rect 2980 -60 2990 -30
rect 3025 -60 3035 -30
rect 2980 -70 3035 -60
rect 3065 -30 3120 -20
rect 3065 -60 3075 -30
rect 3110 -60 3120 -30
rect 3065 -70 3120 -60
rect 3150 -30 3205 -20
rect 3150 -60 3160 -30
rect 3195 -60 3205 -30
rect 3150 -70 3205 -60
rect 3235 -30 3290 -20
rect 3235 -60 3245 -30
rect 3280 -60 3290 -30
rect 3235 -70 3290 -60
rect 3320 -30 3375 -20
rect 3320 -60 3330 -30
rect 3365 -60 3375 -30
rect 3320 -70 3375 -60
rect 3405 -30 3460 -20
rect 3405 -60 3415 -30
rect 3450 -60 3460 -30
rect 3405 -70 3460 -60
rect 3490 -30 3545 -20
rect 3490 -60 3500 -30
rect 3535 -60 3545 -30
rect 3490 -70 3545 -60
rect 3575 -30 3630 -20
rect 3575 -60 3585 -30
rect 3620 -60 3630 -30
rect 3575 -70 3630 -60
rect 3660 -30 3715 -20
rect 3660 -60 3670 -30
rect 3705 -60 3715 -30
rect 3660 -70 3715 -60
rect 3745 -30 3800 -20
rect 3745 -60 3755 -30
rect 3790 -60 3800 -30
rect 3745 -70 3800 -60
rect 3830 -30 3885 -20
rect 3830 -60 3840 -30
rect 3875 -60 3885 -30
rect 3830 -70 3885 -60
rect 3915 -30 3970 -20
rect 3915 -60 3925 -30
rect 3960 -60 3970 -30
rect 3915 -70 3970 -60
rect 4000 -30 4055 -20
rect 4000 -60 4010 -30
rect 4045 -60 4055 -30
rect 4000 -70 4055 -60
rect 4085 -30 4140 -20
rect 4085 -60 4095 -30
rect 4130 -60 4140 -30
rect 4085 -70 4140 -60
rect 4170 -30 4225 -20
rect 4170 -60 4180 -30
rect 4215 -60 4225 -30
rect 4170 -70 4225 -60
rect 4255 -30 4310 -20
rect 4255 -60 4265 -30
rect 4300 -60 4310 -30
rect 4255 -70 4310 -60
rect 4340 -30 4395 -20
rect 4340 -60 4350 -30
rect 4385 -60 4395 -30
rect 4340 -70 4395 -60
rect 4425 -30 4480 -20
rect 4425 -60 4435 -30
rect 4470 -60 4480 -30
rect 4425 -70 4480 -60
rect 4510 -30 4565 -20
rect 4510 -60 4520 -30
rect 4555 -60 4565 -30
rect 4510 -70 4565 -60
rect 4595 -30 4650 -20
rect 4595 -60 4605 -30
rect 4640 -60 4650 -30
rect 4595 -70 4650 -60
rect 4680 -30 4735 -20
rect 4680 -60 4690 -30
rect 4725 -60 4735 -30
rect 4680 -70 4735 -60
rect 4765 -30 4820 -20
rect 4765 -60 4775 -30
rect 4810 -60 4820 -30
rect 4765 -70 4820 -60
rect 4850 -30 4905 -20
rect 4850 -60 4860 -30
rect 4895 -60 4905 -30
rect 4850 -70 4905 -60
rect 4935 -30 4990 -20
rect 4935 -60 4945 -30
rect 4980 -60 4990 -30
rect 4935 -70 4990 -60
rect 5020 -30 5075 -20
rect 5020 -60 5030 -30
rect 5065 -60 5075 -30
rect 5020 -70 5075 -60
rect 5105 -30 5160 -20
rect 5105 -60 5115 -30
rect 5150 -60 5160 -30
rect 5105 -70 5160 -60
rect 5190 -30 5245 -20
rect 5190 -60 5200 -30
rect 5235 -60 5245 -30
rect 5190 -70 5245 -60
rect 5275 -30 5330 -20
rect 5275 -60 5285 -30
rect 5320 -60 5330 -30
rect 5275 -70 5330 -60
rect 5360 -30 5415 -20
rect 5360 -60 5370 -30
rect 5405 -60 5415 -30
rect 5360 -70 5415 -60
rect 5445 -30 5500 -20
rect 5445 -60 5455 -30
rect 5490 -60 5500 -30
rect 5445 -70 5500 -60
rect 5530 -30 5585 -20
rect 5530 -60 5540 -30
rect 5575 -60 5585 -30
rect 5530 -70 5585 -60
rect 5615 -30 5670 -20
rect 5615 -60 5625 -30
rect 5660 -60 5670 -30
rect 5615 -70 5670 -60
rect 5700 -30 5755 -20
rect 5700 -60 5710 -30
rect 5745 -60 5755 -30
rect 5700 -70 5755 -60
rect 5785 -30 5840 -20
rect 5785 -60 5795 -30
rect 5830 -60 5840 -30
rect 5785 -70 5840 -60
rect 5870 -30 5925 -20
rect 5870 -60 5880 -30
rect 5915 -60 5925 -30
rect 5870 -70 5925 -60
rect 5955 -30 6010 -20
rect 5955 -60 5965 -30
rect 6000 -60 6010 -30
rect 5955 -70 6010 -60
rect 6040 -30 6095 -20
rect 6040 -60 6050 -30
rect 6085 -60 6095 -30
rect 6040 -70 6095 -60
rect 6125 -30 6180 -20
rect 6125 -60 6135 -30
rect 6170 -60 6180 -30
rect 6125 -70 6180 -60
rect 6210 -30 6265 -20
rect 6210 -60 6220 -30
rect 6255 -60 6265 -30
rect 6210 -70 6265 -60
rect 6295 -30 6350 -20
rect 6295 -60 6305 -30
rect 6340 -60 6350 -30
rect 6295 -70 6350 -60
rect 6380 -30 6435 -20
rect 6380 -60 6390 -30
rect 6425 -60 6435 -30
rect 6380 -70 6435 -60
rect 6465 -30 6520 -20
rect 6465 -60 6475 -30
rect 6510 -60 6520 -30
rect 6465 -70 6520 -60
rect 6550 -30 6605 -20
rect 6550 -60 6560 -30
rect 6595 -60 6605 -30
rect 6550 -70 6605 -60
rect 6635 -30 6690 -20
rect 6635 -60 6645 -30
rect 6680 -60 6690 -30
rect 6635 -70 6690 -60
rect 6720 -30 6775 -20
rect 6720 -60 6730 -30
rect 6765 -60 6775 -30
rect 6720 -70 6775 -60
rect 6805 -30 6860 -20
rect 6805 -60 6815 -30
rect 6850 -60 6860 -30
rect 6805 -70 6860 -60
rect 6890 -30 6945 -20
rect 6890 -60 6900 -30
rect 6935 -60 6945 -30
rect 6890 -70 6945 -60
rect 6975 -30 7030 -20
rect 6975 -60 6985 -30
rect 7020 -60 7030 -30
rect 6975 -70 7030 -60
rect 7060 -30 7115 -20
rect 7060 -60 7070 -30
rect 7105 -60 7115 -30
rect 7060 -70 7115 -60
rect 7145 -30 7200 -20
rect 7145 -60 7155 -30
rect 7190 -60 7200 -30
rect 7145 -70 7200 -60
rect 7230 -30 7285 -20
rect 7230 -60 7240 -30
rect 7275 -60 7285 -30
rect 7230 -70 7285 -60
rect 7315 -30 7370 -20
rect 7315 -60 7325 -30
rect 7360 -60 7370 -30
rect 7315 -70 7370 -60
rect 7400 -30 7455 -20
rect 7400 -60 7410 -30
rect 7445 -60 7455 -30
rect 7400 -70 7455 -60
rect 7485 -30 7540 -20
rect 7485 -60 7495 -30
rect 7530 -60 7540 -30
rect 7485 -70 7540 -60
rect 7570 -30 7625 -20
rect 7570 -60 7580 -30
rect 7615 -60 7625 -30
rect 7570 -70 7625 -60
rect 7655 -30 7710 -20
rect 7655 -60 7665 -30
rect 7700 -60 7710 -30
rect 7655 -70 7710 -60
rect 7890 -30 7945 -20
rect 7890 -60 7900 -30
rect 7935 -60 7945 -30
rect 7890 -70 7945 -60
rect 7975 -30 8030 -20
rect 7975 -60 7985 -30
rect 8020 -60 8030 -30
rect 7975 -70 8030 -60
rect 8060 -30 8115 -20
rect 8060 -60 8070 -30
rect 8105 -60 8115 -30
rect 8060 -70 8115 -60
rect 8145 -30 8200 -20
rect 8145 -60 8155 -30
rect 8190 -60 8200 -30
rect 8145 -70 8200 -60
rect 8230 -30 8285 -20
rect 8230 -60 8240 -30
rect 8275 -60 8285 -30
rect 8230 -70 8285 -60
rect 8315 -30 8370 -20
rect 8315 -60 8325 -30
rect 8360 -60 8370 -30
rect 8315 -70 8370 -60
rect 8400 -30 8455 -20
rect 8400 -60 8410 -30
rect 8445 -60 8455 -30
rect 8400 -70 8455 -60
rect 8485 -30 8540 -20
rect 8485 -60 8495 -30
rect 8530 -60 8540 -30
rect 8485 -70 8540 -60
rect 8570 -30 8625 -20
rect 8570 -60 8580 -30
rect 8615 -60 8625 -30
rect 8570 -70 8625 -60
rect 8655 -30 8710 -20
rect 8655 -60 8665 -30
rect 8700 -60 8710 -30
rect 8655 -70 8710 -60
rect 8740 -30 8795 -20
rect 8740 -60 8750 -30
rect 8785 -60 8795 -30
rect 8740 -70 8795 -60
rect 8825 -30 8880 -20
rect 8825 -60 8835 -30
rect 8870 -60 8880 -30
rect 8825 -70 8880 -60
rect 8910 -30 8965 -20
rect 8910 -60 8920 -30
rect 8955 -60 8965 -30
rect 8910 -70 8965 -60
rect 8995 -30 9050 -20
rect 8995 -60 9005 -30
rect 9040 -60 9050 -30
rect 8995 -70 9050 -60
rect 9080 -30 9135 -20
rect 9080 -60 9090 -30
rect 9125 -60 9135 -30
rect 9080 -70 9135 -60
rect 9165 -30 9220 -20
rect 9165 -60 9175 -30
rect 9210 -60 9220 -30
rect 9165 -70 9220 -60
rect 9250 -30 9305 -20
rect 9250 -60 9260 -30
rect 9295 -60 9305 -30
rect 9250 -70 9305 -60
rect 9335 -30 9390 -20
rect 9335 -60 9345 -30
rect 9380 -60 9390 -30
rect 9335 -70 9390 -60
rect 9420 -30 9475 -20
rect 9420 -60 9430 -30
rect 9465 -60 9475 -30
rect 9420 -70 9475 -60
rect 9505 -30 9560 -20
rect 9505 -60 9515 -30
rect 9550 -60 9560 -30
rect 9505 -70 9560 -60
rect 9590 -30 9645 -20
rect 9590 -60 9600 -30
rect 9635 -60 9645 -30
rect 9590 -70 9645 -60
rect 9675 -30 9730 -20
rect 9675 -60 9685 -30
rect 9720 -60 9730 -30
rect 9675 -70 9730 -60
rect 9760 -30 9815 -20
rect 9760 -60 9770 -30
rect 9805 -60 9815 -30
rect 9760 -70 9815 -60
rect 9845 -30 9900 -20
rect 9845 -60 9855 -30
rect 9890 -60 9900 -30
rect 9845 -70 9900 -60
rect 9930 -30 9985 -20
rect 9930 -60 9940 -30
rect 9975 -60 9985 -30
rect 9930 -70 9985 -60
rect 10015 -30 10070 -20
rect 10015 -60 10025 -30
rect 10060 -60 10070 -30
rect 10015 -70 10070 -60
rect 10100 -30 10155 -20
rect 10100 -60 10110 -30
rect 10145 -60 10155 -30
rect 10100 -70 10155 -60
rect 10185 -30 10240 -20
rect 10185 -60 10195 -30
rect 10230 -60 10240 -30
rect 10185 -70 10240 -60
rect 10270 -30 10325 -20
rect 10270 -60 10280 -30
rect 10315 -60 10325 -30
rect 10270 -70 10325 -60
rect 10355 -30 10410 -20
rect 10355 -60 10365 -30
rect 10400 -60 10410 -30
rect 10355 -70 10410 -60
rect 10440 -30 10495 -20
rect 10440 -60 10450 -30
rect 10485 -60 10495 -30
rect 10440 -70 10495 -60
rect 10525 -30 10580 -20
rect 10525 -60 10535 -30
rect 10570 -60 10580 -30
rect 10525 -70 10580 -60
rect 10610 -30 10665 -20
rect 10610 -60 10620 -30
rect 10655 -60 10665 -30
rect 10610 -70 10665 -60
rect 10695 -30 10750 -20
rect 10695 -60 10705 -30
rect 10740 -60 10750 -30
rect 10695 -70 10750 -60
rect 10780 -30 10835 -20
rect 10780 -60 10790 -30
rect 10825 -60 10835 -30
rect 10780 -70 10835 -60
rect 10865 -30 10920 -20
rect 10865 -60 10875 -30
rect 10910 -60 10920 -30
rect 10865 -70 10920 -60
rect 10950 -30 11005 -20
rect 10950 -60 10960 -30
rect 10995 -60 11005 -30
rect 10950 -70 11005 -60
rect 11035 -30 11090 -20
rect 11035 -60 11045 -30
rect 11080 -60 11090 -30
rect 11035 -70 11090 -60
rect 11120 -30 11175 -20
rect 11120 -60 11130 -30
rect 11165 -60 11175 -30
rect 11120 -70 11175 -60
rect 11205 -30 11260 -20
rect 11205 -60 11215 -30
rect 11250 -60 11260 -30
rect 11205 -70 11260 -60
rect 11290 -30 11345 -20
rect 11290 -60 11300 -30
rect 11335 -60 11345 -30
rect 11290 -70 11345 -60
rect 11375 -30 11430 -20
rect 11375 -60 11385 -30
rect 11420 -60 11430 -30
rect 11375 -70 11430 -60
rect 11460 -30 11515 -20
rect 11460 -60 11470 -30
rect 11505 -60 11515 -30
rect 11460 -70 11515 -60
rect 11545 -30 11600 -20
rect 11545 -60 11555 -30
rect 11590 -60 11600 -30
rect 11545 -70 11600 -60
rect 11630 -30 11685 -20
rect 11630 -60 11640 -30
rect 11675 -60 11685 -30
rect 11630 -70 11685 -60
rect 11715 -30 11770 -20
rect 11715 -60 11725 -30
rect 11760 -60 11770 -30
rect 11715 -70 11770 -60
rect 11800 -30 11855 -20
rect 11800 -60 11810 -30
rect 11845 -60 11855 -30
rect 11800 -70 11855 -60
rect 11885 -30 11940 -20
rect 11885 -60 11895 -30
rect 11930 -60 11940 -30
rect 11885 -70 11940 -60
rect 11970 -30 12025 -20
rect 11970 -60 11980 -30
rect 12015 -60 12025 -30
rect 11970 -70 12025 -60
rect 12055 -30 12110 -20
rect 12055 -60 12065 -30
rect 12100 -60 12110 -30
rect 12055 -70 12110 -60
rect 12140 -30 12195 -20
rect 12140 -60 12150 -30
rect 12185 -60 12195 -30
rect 12140 -70 12195 -60
rect 12225 -30 12280 -20
rect 12225 -60 12235 -30
rect 12270 -60 12280 -30
rect 12225 -70 12280 -60
rect 12310 -30 12365 -20
rect 12310 -60 12320 -30
rect 12355 -60 12365 -30
rect 12310 -70 12365 -60
rect 12395 -30 12450 -20
rect 12395 -60 12405 -30
rect 12440 -60 12450 -30
rect 12395 -70 12450 -60
rect 12480 -30 12535 -20
rect 12480 -60 12490 -30
rect 12525 -60 12535 -30
rect 12480 -70 12535 -60
rect 12565 -30 12620 -20
rect 12565 -60 12575 -30
rect 12610 -60 12620 -30
rect 12565 -70 12620 -60
rect 12650 -30 12705 -20
rect 12650 -60 12660 -30
rect 12695 -60 12705 -30
rect 12650 -70 12705 -60
rect 12735 -30 12790 -20
rect 12735 -60 12745 -30
rect 12780 -60 12790 -30
rect 12735 -70 12790 -60
rect 12820 -30 12875 -20
rect 12820 -60 12830 -30
rect 12865 -60 12875 -30
rect 12820 -70 12875 -60
rect 12905 -30 12960 -20
rect 12905 -60 12915 -30
rect 12950 -60 12960 -30
rect 12905 -70 12960 -60
rect 12990 -30 13045 -20
rect 12990 -60 13000 -30
rect 13035 -60 13045 -30
rect 12990 -70 13045 -60
rect 13075 -30 13130 -20
rect 13075 -60 13085 -30
rect 13120 -60 13130 -30
rect 13075 -70 13130 -60
rect 13160 -30 13215 -20
rect 13160 -60 13170 -30
rect 13205 -60 13215 -30
rect 13160 -70 13215 -60
rect 13245 -30 13300 -20
rect 13245 -60 13255 -30
rect 13290 -60 13300 -30
rect 13245 -70 13300 -60
rect 13330 -30 13385 -20
rect 13330 -60 13340 -30
rect 13375 -60 13385 -30
rect 13330 -70 13385 -60
rect 13415 -30 13470 -20
rect 13415 -60 13425 -30
rect 13460 -60 13470 -30
rect 13415 -70 13470 -60
rect 13500 -30 13555 -20
rect 13500 -60 13510 -30
rect 13545 -60 13555 -30
rect 13500 -70 13555 -60
rect 13585 -30 13640 -20
rect 13585 -60 13595 -30
rect 13630 -60 13640 -30
rect 13585 -70 13640 -60
rect 13670 -30 13725 -20
rect 13670 -60 13680 -30
rect 13715 -60 13725 -30
rect 13670 -70 13725 -60
rect 13755 -30 13810 -20
rect 13755 -60 13765 -30
rect 13800 -60 13810 -30
rect 13755 -70 13810 -60
rect 13840 -30 13895 -20
rect 13840 -60 13850 -30
rect 13885 -60 13895 -30
rect 13840 -70 13895 -60
rect 13925 -30 13980 -20
rect 13925 -60 13935 -30
rect 13970 -60 13980 -30
rect 13925 -70 13980 -60
rect 14010 -30 14065 -20
rect 14010 -60 14020 -30
rect 14055 -60 14065 -30
rect 14010 -70 14065 -60
rect 14095 -30 14150 -20
rect 14095 -60 14105 -30
rect 14140 -60 14150 -30
rect 14095 -70 14150 -60
rect 14180 -30 14235 -20
rect 14180 -60 14190 -30
rect 14225 -60 14235 -30
rect 14180 -70 14235 -60
rect 14265 -30 14320 -20
rect 14265 -60 14275 -30
rect 14310 -60 14320 -30
rect 14265 -70 14320 -60
rect 14350 -30 14405 -20
rect 14350 -60 14360 -30
rect 14395 -60 14405 -30
rect 14350 -70 14405 -60
rect 14435 -30 14490 -20
rect 14435 -60 14445 -30
rect 14480 -60 14490 -30
rect 14435 -70 14490 -60
rect 14520 -30 14575 -20
rect 14520 -60 14530 -30
rect 14565 -60 14575 -30
rect 14520 -70 14575 -60
rect 14605 -30 14660 -20
rect 14605 -60 14615 -30
rect 14650 -60 14660 -30
rect 14605 -70 14660 -60
rect 14690 -30 14745 -20
rect 14690 -60 14700 -30
rect 14735 -60 14745 -30
rect 14690 -70 14745 -60
rect 14775 -30 14830 -20
rect 14775 -60 14785 -30
rect 14820 -60 14830 -30
rect 14775 -70 14830 -60
rect 14860 -30 14915 -20
rect 14860 -60 14870 -30
rect 14905 -60 14915 -30
rect 14860 -70 14915 -60
rect 14945 -30 15000 -20
rect 14945 -60 14955 -30
rect 14990 -60 15000 -30
rect 14945 -70 15000 -60
rect 15030 -30 15085 -20
rect 15030 -60 15040 -30
rect 15075 -60 15085 -30
rect 15030 -70 15085 -60
rect 15115 -30 15170 -20
rect 15115 -60 15125 -30
rect 15160 -60 15170 -30
rect 15115 -70 15170 -60
rect 15200 -30 15255 -20
rect 15200 -60 15210 -30
rect 15245 -60 15255 -30
rect 15200 -70 15255 -60
rect 15285 -30 15340 -20
rect 15285 -60 15295 -30
rect 15330 -60 15340 -30
rect 15285 -70 15340 -60
rect 15370 -30 15425 -20
rect 15370 -60 15380 -30
rect 15415 -60 15425 -30
rect 15370 -70 15425 -60
rect 15455 -30 15510 -20
rect 15455 -60 15465 -30
rect 15500 -60 15510 -30
rect 15455 -70 15510 -60
rect 15540 -30 15595 -20
rect 15540 -60 15550 -30
rect 15585 -60 15595 -30
rect 15540 -70 15595 -60
rect 15625 -30 15680 -20
rect 15625 -60 15635 -30
rect 15670 -60 15680 -30
rect 15625 -70 15680 -60
rect 15710 -30 15765 -20
rect 15710 -60 15720 -30
rect 15755 -60 15765 -30
rect 15710 -70 15765 -60
rect 15795 -30 15850 -20
rect 15795 -60 15805 -30
rect 15840 -60 15850 -30
rect 15795 -70 15850 -60
rect 15880 -30 15935 -20
rect 15880 -60 15890 -30
rect 15925 -60 15935 -30
rect 15880 -70 15935 -60
rect 15965 -30 16020 -20
rect 15965 -60 15975 -30
rect 16010 -60 16020 -30
rect 15965 -70 16020 -60
rect 16050 -30 16105 -20
rect 16050 -60 16060 -30
rect 16095 -60 16105 -30
rect 16050 -70 16105 -60
rect 16135 -30 16190 -20
rect 16135 -60 16145 -30
rect 16180 -60 16190 -30
rect 16135 -70 16190 -60
rect 16220 -30 16275 -20
rect 16220 -60 16230 -30
rect 16265 -60 16275 -30
rect 16220 -70 16275 -60
rect 16305 -30 16360 -20
rect 16305 -60 16315 -30
rect 16350 -60 16360 -30
rect 16305 -70 16360 -60
rect 16390 -30 16445 -20
rect 16390 -60 16400 -30
rect 16435 -60 16445 -30
rect 16390 -70 16445 -60
rect 16475 -30 16530 -20
rect 16475 -60 16485 -30
rect 16520 -60 16530 -30
rect 16475 -70 16530 -60
rect 16560 -30 16615 -20
rect 16560 -60 16570 -30
rect 16605 -60 16615 -30
rect 16560 -70 16615 -60
rect 16645 -30 16700 -20
rect 16645 -60 16655 -30
rect 16690 -60 16700 -30
rect 16645 -70 16700 -60
rect 16730 -30 16785 -20
rect 16730 -60 16740 -30
rect 16775 -60 16785 -30
rect 16730 -70 16785 -60
rect 16815 -30 16870 -20
rect 16815 -60 16825 -30
rect 16860 -60 16870 -30
rect 16815 -70 16870 -60
rect 16900 -30 16955 -20
rect 16900 -60 16910 -30
rect 16945 -60 16955 -30
rect 16900 -70 16955 -60
rect 16985 -30 17040 -20
rect 16985 -60 16995 -30
rect 17030 -60 17040 -30
rect 16985 -70 17040 -60
rect 17070 -30 17125 -20
rect 17070 -60 17080 -30
rect 17115 -60 17125 -30
rect 17070 -70 17125 -60
rect 17155 -30 17210 -20
rect 17155 -60 17165 -30
rect 17200 -60 17210 -30
rect 17155 -70 17210 -60
rect 17240 -30 17295 -20
rect 17240 -60 17250 -30
rect 17285 -60 17295 -30
rect 17240 -70 17295 -60
rect 17325 -30 17380 -20
rect 17325 -60 17335 -30
rect 17370 -60 17380 -30
rect 17325 -70 17380 -60
rect 17410 -30 17465 -20
rect 17410 -60 17420 -30
rect 17455 -60 17465 -30
rect 17410 -70 17465 -60
rect 17495 -30 17550 -20
rect 17495 -60 17505 -30
rect 17540 -60 17550 -30
rect 17495 -70 17550 -60
rect 17580 -30 17635 -20
rect 17580 -60 17590 -30
rect 17625 -60 17635 -30
rect 17580 -70 17635 -60
rect 17665 -30 17720 -20
rect 17665 -60 17675 -30
rect 17710 -60 17720 -30
rect 17665 -70 17720 -60
rect 17750 -30 17805 -20
rect 17750 -60 17760 -30
rect 17795 -60 17805 -30
rect 17750 -70 17805 -60
rect 17835 -30 17890 -20
rect 17835 -60 17845 -30
rect 17880 -60 17890 -30
rect 17835 -70 17890 -60
rect 17920 -30 17975 -20
rect 17920 -60 17930 -30
rect 17965 -60 17975 -30
rect 17920 -70 17975 -60
rect 18005 -30 18060 -20
rect 18005 -60 18015 -30
rect 18050 -60 18060 -30
rect 18005 -70 18060 -60
rect 18090 -30 18145 -20
rect 18090 -60 18100 -30
rect 18135 -60 18145 -30
rect 18090 -70 18145 -60
rect 18175 -30 18230 -20
rect 18175 -60 18185 -30
rect 18220 -60 18230 -30
rect 18175 -70 18230 -60
rect 18260 -30 18315 -20
rect 18260 -60 18270 -30
rect 18305 -60 18315 -30
rect 18260 -70 18315 -60
rect 18345 -30 18400 -20
rect 18345 -60 18355 -30
rect 18390 -60 18400 -30
rect 18345 -70 18400 -60
rect 18430 -30 18485 -20
rect 18430 -60 18440 -30
rect 18475 -60 18485 -30
rect 18430 -70 18485 -60
rect 18515 -30 18570 -20
rect 18515 -60 18525 -30
rect 18560 -60 18570 -30
rect 18515 -70 18570 -60
rect 18600 -30 18655 -20
rect 18600 -60 18610 -30
rect 18645 -60 18655 -30
rect 18600 -70 18655 -60
rect 18685 -30 18740 -20
rect 18685 -60 18695 -30
rect 18730 -60 18740 -30
rect 18685 -70 18740 -60
rect 18770 -30 18825 -20
rect 18770 -60 18780 -30
rect 18815 -60 18825 -30
rect 18770 -70 18825 -60
rect 18855 -30 18910 -20
rect 18855 -60 18865 -30
rect 18900 -60 18910 -30
rect 18855 -70 18910 -60
rect 18940 -30 18995 -20
rect 18940 -60 18950 -30
rect 18985 -60 18995 -30
rect 18940 -70 18995 -60
rect 19025 -30 19080 -20
rect 19025 -60 19035 -30
rect 19070 -60 19080 -30
rect 19025 -70 19080 -60
rect 19110 -30 19165 -20
rect 19110 -60 19120 -30
rect 19155 -60 19165 -30
rect 19110 -70 19165 -60
rect 19195 -30 19250 -20
rect 19195 -60 19205 -30
rect 19240 -60 19250 -30
rect 19195 -70 19250 -60
rect 19280 -30 19335 -20
rect 19280 -60 19290 -30
rect 19325 -60 19335 -30
rect 19280 -70 19335 -60
rect 19365 -30 19420 -20
rect 19365 -60 19375 -30
rect 19410 -60 19420 -30
rect 19365 -70 19420 -60
rect 19450 -30 19505 -20
rect 19450 -60 19460 -30
rect 19495 -60 19505 -30
rect 19450 -70 19505 -60
rect 19535 -30 19590 -20
rect 19535 -60 19545 -30
rect 19580 -60 19590 -30
rect 19535 -70 19590 -60
rect 19620 -30 19675 -20
rect 19620 -60 19630 -30
rect 19665 -60 19675 -30
rect 19620 -70 19675 -60
rect 19705 -30 19760 -20
rect 19705 -60 19715 -30
rect 19750 -60 19760 -30
rect 19705 -70 19760 -60
rect 19790 -30 19845 -20
rect 19790 -60 19800 -30
rect 19835 -60 19845 -30
rect 19790 -70 19845 -60
rect 19875 -30 19930 -20
rect 19875 -60 19885 -30
rect 19920 -60 19930 -30
rect 19875 -70 19930 -60
rect 19960 -30 20015 -20
rect 19960 -60 19970 -30
rect 20005 -60 20015 -30
rect 19960 -70 20015 -60
rect 20045 -30 20100 -20
rect 20045 -60 20055 -30
rect 20090 -60 20100 -30
rect 20045 -70 20100 -60
rect 20130 -30 20185 -20
rect 20130 -60 20140 -30
rect 20175 -60 20185 -30
rect 20130 -70 20185 -60
rect 20215 -30 20270 -20
rect 20215 -60 20225 -30
rect 20260 -60 20270 -30
rect 20215 -70 20270 -60
rect 20300 -30 20355 -20
rect 20300 -60 20310 -30
rect 20345 -60 20355 -30
rect 20300 -70 20355 -60
rect 20385 -30 20440 -20
rect 20385 -60 20395 -30
rect 20430 -60 20440 -30
rect 20385 -70 20440 -60
rect 20470 -30 20525 -20
rect 20470 -60 20480 -30
rect 20515 -60 20525 -30
rect 20470 -70 20525 -60
rect 20555 -30 20610 -20
rect 20555 -60 20565 -30
rect 20600 -60 20610 -30
rect 20555 -70 20610 -60
rect 20640 -30 20695 -20
rect 20640 -60 20650 -30
rect 20685 -60 20695 -30
rect 20640 -70 20695 -60
rect 20725 -30 20780 -20
rect 20725 -60 20735 -30
rect 20770 -60 20780 -30
rect 20725 -70 20780 -60
rect 20810 -30 20865 -20
rect 20810 -60 20820 -30
rect 20855 -60 20865 -30
rect 20810 -70 20865 -60
rect 20895 -30 20950 -20
rect 20895 -60 20905 -30
rect 20940 -60 20950 -30
rect 20895 -70 20950 -60
rect 20980 -30 21035 -20
rect 20980 -60 20990 -30
rect 21025 -60 21035 -30
rect 20980 -70 21035 -60
rect 21065 -30 21120 -20
rect 21065 -60 21075 -30
rect 21110 -60 21120 -30
rect 21065 -70 21120 -60
rect 21150 -30 21205 -20
rect 21150 -60 21160 -30
rect 21195 -60 21205 -30
rect 21150 -70 21205 -60
rect 21235 -30 21290 -20
rect 21235 -60 21245 -30
rect 21280 -60 21290 -30
rect 21235 -70 21290 -60
rect 21320 -30 21375 -20
rect 21320 -60 21330 -30
rect 21365 -60 21375 -30
rect 21320 -70 21375 -60
rect 21405 -30 21460 -20
rect 21405 -60 21415 -30
rect 21450 -60 21460 -30
rect 21405 -70 21460 -60
rect 21490 -30 21545 -20
rect 21490 -60 21500 -30
rect 21535 -60 21545 -30
rect 21490 -70 21545 -60
rect 21575 -30 21630 -20
rect 21575 -60 21585 -30
rect 21620 -60 21630 -30
rect 21575 -70 21630 -60
rect 21660 -30 21715 -20
rect 21660 -60 21670 -30
rect 21705 -60 21715 -30
rect 21660 -70 21715 -60
rect 21745 -30 21800 -20
rect 21745 -60 21755 -30
rect 21790 -60 21800 -30
rect 21745 -70 21800 -60
rect 21830 -30 21885 -20
rect 21830 -60 21840 -30
rect 21875 -60 21885 -30
rect 21830 -70 21885 -60
rect 21915 -30 21970 -20
rect 21915 -60 21925 -30
rect 21960 -60 21970 -30
rect 21915 -70 21970 -60
rect 22000 -30 22055 -20
rect 22000 -60 22010 -30
rect 22045 -60 22055 -30
rect 22000 -70 22055 -60
rect 22085 -30 22140 -20
rect 22085 -60 22095 -30
rect 22130 -60 22140 -30
rect 22085 -70 22140 -60
rect 22170 -30 22225 -20
rect 22170 -60 22180 -30
rect 22215 -60 22225 -30
rect 22170 -70 22225 -60
rect 22255 -30 22310 -20
rect 22255 -60 22265 -30
rect 22300 -60 22310 -30
rect 22255 -70 22310 -60
rect 22340 -30 22395 -20
rect 22340 -60 22350 -30
rect 22385 -60 22395 -30
rect 22340 -70 22395 -60
rect 22425 -30 22480 -20
rect 22425 -60 22435 -30
rect 22470 -60 22480 -30
rect 22425 -70 22480 -60
rect 22510 -30 22565 -20
rect 22510 -60 22520 -30
rect 22555 -60 22565 -30
rect 22510 -70 22565 -60
rect 22595 -30 22650 -20
rect 22595 -60 22605 -30
rect 22640 -60 22650 -30
rect 22595 -70 22650 -60
rect 22680 -30 22735 -20
rect 22680 -60 22690 -30
rect 22725 -60 22735 -30
rect 22680 -70 22735 -60
rect 22765 -30 22820 -20
rect 22765 -60 22775 -30
rect 22810 -60 22820 -30
rect 22765 -70 22820 -60
rect 22850 -30 22905 -20
rect 22850 -60 22860 -30
rect 22895 -60 22905 -30
rect 22850 -70 22905 -60
rect 22935 -30 22990 -20
rect 22935 -60 22945 -30
rect 22980 -60 22990 -30
rect 22935 -70 22990 -60
rect 23020 -30 23075 -20
rect 23020 -60 23030 -30
rect 23065 -60 23075 -30
rect 23020 -70 23075 -60
rect 23105 -30 23160 -20
rect 23105 -60 23115 -30
rect 23150 -60 23160 -30
rect 23105 -70 23160 -60
rect 23190 -30 23245 -20
rect 23190 -60 23200 -30
rect 23235 -60 23245 -30
rect 23190 -70 23245 -60
rect 23275 -30 23330 -20
rect 23275 -60 23285 -30
rect 23320 -60 23330 -30
rect 23275 -70 23330 -60
rect 23360 -30 23415 -20
rect 23360 -60 23370 -30
rect 23405 -60 23415 -30
rect 23360 -70 23415 -60
rect 23445 -30 23500 -20
rect 23445 -60 23455 -30
rect 23490 -60 23500 -30
rect 23445 -70 23500 -60
rect 23530 -30 23585 -20
rect 23530 -60 23540 -30
rect 23575 -60 23585 -30
rect 23530 -70 23585 -60
rect 23615 -30 23670 -20
rect 23615 -60 23625 -30
rect 23660 -60 23670 -30
rect 23615 -70 23670 -60
rect 23700 -30 23755 -20
rect 23700 -60 23710 -30
rect 23745 -60 23755 -30
rect 23700 -70 23755 -60
rect 23785 -30 23840 -20
rect 23785 -60 23795 -30
rect 23830 -60 23840 -30
rect 23785 -70 23840 -60
rect 23870 -30 23925 -20
rect 23870 -60 23880 -30
rect 23915 -60 23925 -30
rect 23870 -70 23925 -60
rect 23955 -30 24010 -20
rect 23955 -60 23965 -30
rect 24000 -60 24010 -30
rect 23955 -70 24010 -60
rect 24040 -30 24095 -20
rect 24040 -60 24050 -30
rect 24085 -60 24095 -30
rect 24040 -70 24095 -60
rect 24125 -30 24180 -20
rect 24125 -60 24135 -30
rect 24170 -60 24180 -30
rect 24125 -70 24180 -60
rect 24210 -30 24265 -20
rect 24210 -60 24220 -30
rect 24255 -60 24265 -30
rect 24210 -70 24265 -60
rect 24295 -30 24350 -20
rect 24295 -60 24305 -30
rect 24340 -60 24350 -30
rect 24295 -70 24350 -60
rect 24380 -30 24435 -20
rect 24380 -60 24390 -30
rect 24425 -60 24435 -30
rect 24380 -70 24435 -60
rect 24465 -30 24520 -20
rect 24465 -60 24475 -30
rect 24510 -60 24520 -30
rect 24465 -70 24520 -60
rect 24550 -30 24605 -20
rect 24550 -60 24560 -30
rect 24595 -60 24605 -30
rect 24550 -70 24605 -60
rect 24635 -30 24690 -20
rect 24635 -60 24645 -30
rect 24680 -60 24690 -30
rect 24635 -70 24690 -60
rect 24720 -30 24775 -20
rect 24720 -60 24730 -30
rect 24765 -60 24775 -30
rect 24720 -70 24775 -60
rect 24805 -30 24860 -20
rect 24805 -60 24815 -30
rect 24850 -60 24860 -30
rect 24805 -70 24860 -60
rect 24890 -30 24945 -20
rect 24890 -60 24900 -30
rect 24935 -60 24945 -30
rect 24890 -70 24945 -60
rect 24975 -30 25030 -20
rect 24975 -60 24985 -30
rect 25020 -60 25030 -30
rect 24975 -70 25030 -60
rect 25060 -30 25115 -20
rect 25060 -60 25070 -30
rect 25105 -60 25115 -30
rect 25060 -70 25115 -60
rect 25145 -30 25200 -20
rect 25145 -60 25155 -30
rect 25190 -60 25200 -30
rect 25145 -70 25200 -60
rect 25230 -30 25285 -20
rect 25230 -60 25240 -30
rect 25275 -60 25285 -30
rect 25230 -70 25285 -60
rect 25315 -30 25370 -20
rect 25315 -60 25325 -30
rect 25360 -60 25370 -30
rect 25315 -70 25370 -60
rect 25400 -30 25455 -20
rect 25400 -60 25410 -30
rect 25445 -60 25455 -30
rect 25400 -70 25455 -60
rect 25485 -30 25540 -20
rect 25485 -60 25495 -30
rect 25530 -60 25540 -30
rect 25485 -70 25540 -60
rect 25570 -30 25625 -20
rect 25570 -60 25580 -30
rect 25615 -60 25625 -30
rect 25570 -70 25625 -60
rect 25655 -30 25710 -20
rect 25655 -60 25665 -30
rect 25700 -60 25710 -30
rect 25655 -70 25710 -60
rect 25740 -30 25795 -20
rect 25740 -60 25750 -30
rect 25785 -60 25795 -30
rect 25740 -70 25795 -60
rect 25825 -30 25880 -20
rect 25825 -60 25835 -30
rect 25870 -60 25880 -30
rect 25825 -70 25880 -60
rect 25910 -30 25965 -20
rect 25910 -60 25920 -30
rect 25955 -60 25965 -30
rect 25910 -70 25965 -60
rect 25995 -30 26050 -20
rect 25995 -60 26005 -30
rect 26040 -60 26050 -30
rect 25995 -70 26050 -60
rect 26080 -30 26135 -20
rect 26080 -60 26090 -30
rect 26125 -60 26135 -30
rect 26080 -70 26135 -60
rect 26165 -30 26220 -20
rect 26165 -60 26175 -30
rect 26210 -60 26220 -30
rect 26165 -70 26220 -60
rect 26250 -30 26305 -20
rect 26250 -60 26260 -30
rect 26295 -60 26305 -30
rect 26250 -70 26305 -60
rect 26335 -30 26390 -20
rect 26335 -60 26345 -30
rect 26380 -60 26390 -30
rect 26335 -70 26390 -60
rect 26420 -30 26475 -20
rect 26420 -60 26430 -30
rect 26465 -60 26475 -30
rect 26420 -70 26475 -60
rect 26505 -30 26560 -20
rect 26505 -60 26515 -30
rect 26550 -60 26560 -30
rect 26505 -70 26560 -60
rect 26590 -30 26645 -20
rect 26590 -60 26600 -30
rect 26635 -60 26645 -30
rect 26590 -70 26645 -60
rect 26675 -30 26730 -20
rect 26675 -60 26685 -30
rect 26720 -60 26730 -30
rect 26675 -70 26730 -60
rect 26760 -30 26815 -20
rect 26760 -60 26770 -30
rect 26805 -60 26815 -30
rect 26760 -70 26815 -60
rect 26845 -30 26900 -20
rect 26845 -60 26855 -30
rect 26890 -60 26900 -30
rect 26845 -70 26900 -60
rect 26930 -30 26985 -20
rect 26930 -60 26940 -30
rect 26975 -60 26985 -30
rect 26930 -70 26985 -60
rect 27015 -30 27070 -20
rect 27015 -60 27025 -30
rect 27060 -60 27070 -30
rect 27015 -70 27070 -60
rect 27100 -30 27155 -20
rect 27100 -60 27110 -30
rect 27145 -60 27155 -30
rect 27100 -70 27155 -60
rect 27185 -30 27240 -20
rect 27185 -60 27195 -30
rect 27230 -60 27240 -30
rect 27185 -70 27240 -60
rect 27270 -30 27325 -20
rect 27270 -60 27280 -30
rect 27315 -60 27325 -30
rect 27270 -70 27325 -60
rect 27355 -30 27410 -20
rect 27355 -60 27365 -30
rect 27400 -60 27410 -30
rect 27355 -70 27410 -60
rect 27440 -30 27495 -20
rect 27440 -60 27450 -30
rect 27485 -60 27495 -30
rect 27440 -70 27495 -60
rect 27525 -30 27580 -20
rect 27525 -60 27535 -30
rect 27570 -60 27580 -30
rect 27525 -70 27580 -60
rect 27610 -30 27665 -20
rect 27610 -60 27620 -30
rect 27655 -60 27665 -30
rect 27610 -70 27665 -60
rect 27695 -30 27750 -20
rect 27695 -60 27705 -30
rect 27740 -60 27750 -30
rect 27695 -70 27750 -60
rect 27780 -30 27835 -20
rect 27780 -60 27790 -30
rect 27825 -60 27835 -30
rect 27780 -70 27835 -60
rect 27865 -30 27920 -20
rect 27865 -60 27875 -30
rect 27910 -60 27920 -30
rect 27865 -70 27920 -60
rect 27950 -30 28005 -20
rect 27950 -60 27960 -30
rect 27995 -60 28005 -30
rect 27950 -70 28005 -60
rect 28035 -30 28090 -20
rect 28035 -60 28045 -30
rect 28080 -60 28090 -30
rect 28035 -70 28090 -60
rect 28120 -30 28175 -20
rect 28120 -60 28130 -30
rect 28165 -60 28175 -30
rect 28120 -70 28175 -60
rect 28205 -30 28260 -20
rect 28205 -60 28215 -30
rect 28250 -60 28260 -30
rect 28205 -70 28260 -60
rect 28290 -30 28345 -20
rect 28290 -60 28300 -30
rect 28335 -60 28345 -30
rect 28290 -70 28345 -60
rect 28375 -30 28430 -20
rect 28375 -60 28385 -30
rect 28420 -60 28430 -30
rect 28375 -70 28430 -60
rect 28460 -30 28515 -20
rect 28460 -60 28470 -30
rect 28505 -60 28515 -30
rect 28460 -70 28515 -60
rect 28545 -30 28600 -20
rect 28545 -60 28555 -30
rect 28590 -60 28600 -30
rect 28545 -70 28600 -60
rect 28630 -30 28685 -20
rect 28630 -60 28640 -30
rect 28675 -60 28685 -30
rect 28630 -70 28685 -60
rect 28715 -30 28770 -20
rect 28715 -60 28725 -30
rect 28760 -60 28770 -30
rect 28715 -70 28770 -60
rect 28800 -30 28855 -20
rect 28800 -60 28810 -30
rect 28845 -60 28855 -30
rect 28800 -70 28855 -60
rect 28885 -30 28940 -20
rect 28885 -60 28895 -30
rect 28930 -60 28940 -30
rect 28885 -70 28940 -60
rect 28970 -30 29025 -20
rect 28970 -60 28980 -30
rect 29015 -60 29025 -30
rect 28970 -70 29025 -60
rect 29055 -30 29110 -20
rect 29055 -60 29065 -30
rect 29100 -60 29110 -30
rect 29055 -70 29110 -60
rect 29140 -30 29195 -20
rect 29140 -60 29150 -30
rect 29185 -60 29195 -30
rect 29140 -70 29195 -60
rect 29225 -30 29280 -20
rect 29225 -60 29235 -30
rect 29270 -60 29280 -30
rect 29225 -70 29280 -60
rect 29310 -30 29365 -20
rect 29310 -60 29320 -30
rect 29355 -60 29365 -30
rect 29310 -70 29365 -60
rect 29395 -30 29450 -20
rect 29395 -60 29405 -30
rect 29440 -60 29450 -30
rect 29395 -70 29450 -60
rect 29480 -30 29535 -20
rect 29480 -60 29490 -30
rect 29525 -60 29535 -30
rect 29480 -70 29535 -60
rect 29565 -30 29620 -20
rect 29565 -60 29575 -30
rect 29610 -60 29620 -30
rect 29565 -70 29620 -60
rect 65 -85 80 -70
rect 105 -265 160 -255
rect 105 -295 115 -265
rect 150 -295 160 -265
rect 105 -305 160 -295
rect 190 -265 245 -255
rect 190 -295 200 -265
rect 235 -295 245 -265
rect 190 -305 245 -295
rect 275 -265 330 -255
rect 275 -295 285 -265
rect 320 -295 330 -265
rect 275 -305 330 -295
rect 360 -265 415 -255
rect 360 -295 370 -265
rect 405 -295 415 -265
rect 360 -305 415 -295
rect 445 -265 500 -255
rect 445 -295 455 -265
rect 490 -295 500 -265
rect 445 -305 500 -295
rect 530 -265 585 -255
rect 530 -295 540 -265
rect 575 -295 585 -265
rect 530 -305 585 -295
rect 615 -265 670 -255
rect 615 -295 625 -265
rect 660 -295 670 -265
rect 615 -305 670 -295
rect 700 -265 755 -255
rect 700 -295 710 -265
rect 745 -295 755 -265
rect 700 -305 755 -295
rect 785 -265 840 -255
rect 785 -295 795 -265
rect 830 -295 840 -265
rect 785 -305 840 -295
rect 870 -265 925 -255
rect 870 -295 880 -265
rect 915 -295 925 -265
rect 870 -305 925 -295
rect 955 -265 1010 -255
rect 955 -295 965 -265
rect 1000 -295 1010 -265
rect 955 -305 1010 -295
rect 1040 -265 1095 -255
rect 1040 -295 1050 -265
rect 1085 -295 1095 -265
rect 1040 -305 1095 -295
rect 1125 -265 1180 -255
rect 1125 -295 1135 -265
rect 1170 -295 1180 -265
rect 1125 -305 1180 -295
rect 1210 -265 1265 -255
rect 1210 -295 1220 -265
rect 1255 -295 1265 -265
rect 1210 -305 1265 -295
rect 1295 -265 1350 -255
rect 1295 -295 1305 -265
rect 1340 -295 1350 -265
rect 1295 -305 1350 -295
rect 1380 -265 1435 -255
rect 1380 -295 1390 -265
rect 1425 -295 1435 -265
rect 1380 -305 1435 -295
rect 1465 -265 1520 -255
rect 1465 -295 1475 -265
rect 1510 -295 1520 -265
rect 1465 -305 1520 -295
rect 1550 -265 1605 -255
rect 1550 -295 1560 -265
rect 1595 -295 1605 -265
rect 1550 -305 1605 -295
rect 1635 -265 1690 -255
rect 1635 -295 1645 -265
rect 1680 -295 1690 -265
rect 1635 -305 1690 -295
rect 1720 -265 1775 -255
rect 1720 -295 1730 -265
rect 1765 -295 1775 -265
rect 1720 -305 1775 -295
rect 1805 -265 1860 -255
rect 1805 -295 1815 -265
rect 1850 -295 1860 -265
rect 1805 -305 1860 -295
rect 1890 -265 1945 -255
rect 1890 -295 1900 -265
rect 1935 -295 1945 -265
rect 1890 -305 1945 -295
rect 1975 -265 2030 -255
rect 1975 -295 1985 -265
rect 2020 -295 2030 -265
rect 1975 -305 2030 -295
rect 2060 -265 2115 -255
rect 2060 -295 2070 -265
rect 2105 -295 2115 -265
rect 2060 -305 2115 -295
rect 2145 -265 2200 -255
rect 2145 -295 2155 -265
rect 2190 -295 2200 -265
rect 2145 -305 2200 -295
rect 2230 -265 2285 -255
rect 2230 -295 2240 -265
rect 2275 -295 2285 -265
rect 2230 -305 2285 -295
rect 2315 -265 2370 -255
rect 2315 -295 2325 -265
rect 2360 -295 2370 -265
rect 2315 -305 2370 -295
rect 2400 -265 2455 -255
rect 2400 -295 2410 -265
rect 2445 -295 2455 -265
rect 2400 -305 2455 -295
rect 2485 -265 2540 -255
rect 2485 -295 2495 -265
rect 2530 -295 2540 -265
rect 2485 -305 2540 -295
rect 2570 -265 2625 -255
rect 2570 -295 2580 -265
rect 2615 -295 2625 -265
rect 2570 -305 2625 -295
rect 2655 -265 2710 -255
rect 2655 -295 2665 -265
rect 2700 -295 2710 -265
rect 2655 -305 2710 -295
rect 2740 -265 2795 -255
rect 2740 -295 2750 -265
rect 2785 -295 2795 -265
rect 2740 -305 2795 -295
rect 2825 -265 2880 -255
rect 2825 -295 2835 -265
rect 2870 -295 2880 -265
rect 2825 -305 2880 -295
rect 2910 -265 2965 -255
rect 2910 -295 2920 -265
rect 2955 -295 2965 -265
rect 2910 -305 2965 -295
rect 2995 -265 3050 -255
rect 2995 -295 3005 -265
rect 3040 -295 3050 -265
rect 2995 -305 3050 -295
rect 3080 -265 3135 -255
rect 3080 -295 3090 -265
rect 3125 -295 3135 -265
rect 3080 -305 3135 -295
rect 3165 -265 3220 -255
rect 3165 -295 3175 -265
rect 3210 -295 3220 -265
rect 3165 -305 3220 -295
rect 3250 -265 3305 -255
rect 3250 -295 3260 -265
rect 3295 -295 3305 -265
rect 3250 -305 3305 -295
rect 3335 -265 3390 -255
rect 3335 -295 3345 -265
rect 3380 -295 3390 -265
rect 3335 -305 3390 -295
rect 3420 -265 3475 -255
rect 3420 -295 3430 -265
rect 3465 -295 3475 -265
rect 3420 -305 3475 -295
rect 3505 -265 3560 -255
rect 3505 -295 3515 -265
rect 3550 -295 3560 -265
rect 3505 -305 3560 -295
rect 3590 -265 3645 -255
rect 3590 -295 3600 -265
rect 3635 -295 3645 -265
rect 3590 -305 3645 -295
rect 3675 -265 3730 -255
rect 3675 -295 3685 -265
rect 3720 -295 3730 -265
rect 3675 -305 3730 -295
rect 3760 -265 3815 -255
rect 3760 -295 3770 -265
rect 3805 -295 3815 -265
rect 3760 -305 3815 -295
rect 3845 -265 3900 -255
rect 3845 -295 3855 -265
rect 3890 -295 3900 -265
rect 3845 -305 3900 -295
rect 3930 -265 3985 -255
rect 3930 -295 3940 -265
rect 3975 -295 3985 -265
rect 3930 -305 3985 -295
rect 4015 -265 4070 -255
rect 4015 -295 4025 -265
rect 4060 -295 4070 -265
rect 4015 -305 4070 -295
rect 4100 -265 4155 -255
rect 4100 -295 4110 -265
rect 4145 -295 4155 -265
rect 4100 -305 4155 -295
rect 4185 -265 4240 -255
rect 4185 -295 4195 -265
rect 4230 -295 4240 -265
rect 4185 -305 4240 -295
rect 4270 -265 4325 -255
rect 4270 -295 4280 -265
rect 4315 -295 4325 -265
rect 4270 -305 4325 -295
rect 4355 -265 4410 -255
rect 4355 -295 4365 -265
rect 4400 -295 4410 -265
rect 4355 -305 4410 -295
rect 4440 -265 4495 -255
rect 4440 -295 4450 -265
rect 4485 -295 4495 -265
rect 4440 -305 4495 -295
rect 4525 -265 4580 -255
rect 4525 -295 4535 -265
rect 4570 -295 4580 -265
rect 4525 -305 4580 -295
rect 4610 -265 4665 -255
rect 4610 -295 4620 -265
rect 4655 -295 4665 -265
rect 4610 -305 4665 -295
rect 4695 -265 4750 -255
rect 4695 -295 4705 -265
rect 4740 -295 4750 -265
rect 4695 -305 4750 -295
rect 4780 -265 4835 -255
rect 4780 -295 4790 -265
rect 4825 -295 4835 -265
rect 4780 -305 4835 -295
rect 4865 -265 4920 -255
rect 4865 -295 4875 -265
rect 4910 -295 4920 -265
rect 4865 -305 4920 -295
rect 4950 -265 5005 -255
rect 4950 -295 4960 -265
rect 4995 -295 5005 -265
rect 4950 -305 5005 -295
rect 5035 -265 5090 -255
rect 5035 -295 5045 -265
rect 5080 -295 5090 -265
rect 5035 -305 5090 -295
rect 5120 -265 5175 -255
rect 5120 -295 5130 -265
rect 5165 -295 5175 -265
rect 5120 -305 5175 -295
rect 5205 -265 5260 -255
rect 5205 -295 5215 -265
rect 5250 -295 5260 -265
rect 5205 -305 5260 -295
rect 5290 -265 5345 -255
rect 5290 -295 5300 -265
rect 5335 -295 5345 -265
rect 5290 -305 5345 -295
rect 5375 -265 5430 -255
rect 5375 -295 5385 -265
rect 5420 -295 5430 -265
rect 5375 -305 5430 -295
rect 5460 -265 5515 -255
rect 5460 -295 5470 -265
rect 5505 -295 5515 -265
rect 5460 -305 5515 -295
rect 5545 -265 5600 -255
rect 5545 -295 5555 -265
rect 5590 -295 5600 -265
rect 5545 -305 5600 -295
rect 5630 -265 5685 -255
rect 5630 -295 5640 -265
rect 5675 -295 5685 -265
rect 5630 -305 5685 -295
rect 5715 -265 5770 -255
rect 5715 -295 5725 -265
rect 5760 -295 5770 -265
rect 5715 -305 5770 -295
rect 5800 -265 5855 -255
rect 5800 -295 5810 -265
rect 5845 -295 5855 -265
rect 5800 -305 5855 -295
rect 5885 -265 5940 -255
rect 5885 -295 5895 -265
rect 5930 -295 5940 -265
rect 5885 -305 5940 -295
rect 5970 -265 6025 -255
rect 5970 -295 5980 -265
rect 6015 -295 6025 -265
rect 5970 -305 6025 -295
rect 6055 -265 6110 -255
rect 6055 -295 6065 -265
rect 6100 -295 6110 -265
rect 6055 -305 6110 -295
rect 6140 -265 6195 -255
rect 6140 -295 6150 -265
rect 6185 -295 6195 -265
rect 6140 -305 6195 -295
rect 6225 -265 6280 -255
rect 6225 -295 6235 -265
rect 6270 -295 6280 -265
rect 6225 -305 6280 -295
rect 6310 -265 6365 -255
rect 6310 -295 6320 -265
rect 6355 -295 6365 -265
rect 6310 -305 6365 -295
rect 6395 -265 6450 -255
rect 6395 -295 6405 -265
rect 6440 -295 6450 -265
rect 6395 -305 6450 -295
rect 6480 -265 6535 -255
rect 6480 -295 6490 -265
rect 6525 -295 6535 -265
rect 6480 -305 6535 -295
rect 6565 -265 6620 -255
rect 6565 -295 6575 -265
rect 6610 -295 6620 -265
rect 6565 -305 6620 -295
rect 6650 -265 6705 -255
rect 6650 -295 6660 -265
rect 6695 -295 6705 -265
rect 6650 -305 6705 -295
rect 6735 -265 6790 -255
rect 6735 -295 6745 -265
rect 6780 -295 6790 -265
rect 6735 -305 6790 -295
rect 6820 -265 6875 -255
rect 6820 -295 6830 -265
rect 6865 -295 6875 -265
rect 6820 -305 6875 -295
rect 6905 -265 6960 -255
rect 6905 -295 6915 -265
rect 6950 -295 6960 -265
rect 6905 -305 6960 -295
rect 6990 -265 7045 -255
rect 6990 -295 7000 -265
rect 7035 -295 7045 -265
rect 6990 -305 7045 -295
rect 7075 -265 7130 -255
rect 7075 -295 7085 -265
rect 7120 -295 7130 -265
rect 7075 -305 7130 -295
rect 7160 -265 7215 -255
rect 7160 -295 7170 -265
rect 7205 -295 7215 -265
rect 7160 -305 7215 -295
rect 7245 -265 7300 -255
rect 7245 -295 7255 -265
rect 7290 -295 7300 -265
rect 7245 -305 7300 -295
rect 7330 -265 7385 -255
rect 7330 -295 7340 -265
rect 7375 -295 7385 -265
rect 7330 -305 7385 -295
rect 7415 -265 7470 -255
rect 7415 -295 7425 -265
rect 7460 -295 7470 -265
rect 7415 -305 7470 -295
rect 7500 -265 7555 -255
rect 7500 -295 7510 -265
rect 7545 -295 7555 -265
rect 7500 -305 7555 -295
rect 7585 -265 7640 -255
rect 7585 -295 7595 -265
rect 7630 -295 7640 -265
rect 7585 -305 7640 -295
rect 7670 -265 7725 -255
rect 7670 -295 7680 -265
rect 7715 -295 7725 -265
rect 7670 -305 7725 -295
rect 7755 -265 7810 -255
rect 7755 -295 7765 -265
rect 7800 -295 7810 -265
rect 7755 -305 7810 -295
rect 7840 -265 7895 -255
rect 7840 -295 7850 -265
rect 7885 -295 7895 -265
rect 7840 -305 7895 -295
rect 7925 -265 7980 -255
rect 7925 -295 7935 -265
rect 7970 -295 7980 -265
rect 7925 -305 7980 -295
rect 8010 -265 8065 -255
rect 8010 -295 8020 -265
rect 8055 -295 8065 -265
rect 8010 -305 8065 -295
rect 8095 -265 8150 -255
rect 8095 -295 8105 -265
rect 8140 -295 8150 -265
rect 8095 -305 8150 -295
rect 8180 -265 8235 -255
rect 8180 -295 8190 -265
rect 8225 -295 8235 -265
rect 8180 -305 8235 -295
rect 8265 -265 8320 -255
rect 8265 -295 8275 -265
rect 8310 -295 8320 -265
rect 8265 -305 8320 -295
rect 8350 -265 8405 -255
rect 8350 -295 8360 -265
rect 8395 -295 8405 -265
rect 8350 -305 8405 -295
rect 8435 -265 8490 -255
rect 8435 -295 8445 -265
rect 8480 -295 8490 -265
rect 8435 -305 8490 -295
rect 8520 -265 8575 -255
rect 8520 -295 8530 -265
rect 8565 -295 8575 -265
rect 8520 -305 8575 -295
rect 8605 -265 8660 -255
rect 8605 -295 8615 -265
rect 8650 -295 8660 -265
rect 8605 -305 8660 -295
rect 8690 -265 8745 -255
rect 8690 -295 8700 -265
rect 8735 -295 8745 -265
rect 8690 -305 8745 -295
rect 8775 -265 8830 -255
rect 8775 -295 8785 -265
rect 8820 -295 8830 -265
rect 8775 -305 8830 -295
rect 8860 -265 8915 -255
rect 8860 -295 8870 -265
rect 8905 -295 8915 -265
rect 8860 -305 8915 -295
rect 8945 -265 9000 -255
rect 8945 -295 8955 -265
rect 8990 -295 9000 -265
rect 8945 -305 9000 -295
rect 9030 -265 9085 -255
rect 9030 -295 9040 -265
rect 9075 -295 9085 -265
rect 9030 -305 9085 -295
rect 9115 -265 9170 -255
rect 9115 -295 9125 -265
rect 9160 -295 9170 -265
rect 9115 -305 9170 -295
rect 9200 -265 9255 -255
rect 9200 -295 9210 -265
rect 9245 -295 9255 -265
rect 9200 -305 9255 -295
rect 9285 -265 9340 -255
rect 9285 -295 9295 -265
rect 9330 -295 9340 -265
rect 9285 -305 9340 -295
rect 9370 -265 9425 -255
rect 9370 -295 9380 -265
rect 9415 -295 9425 -265
rect 9370 -305 9425 -295
rect 9455 -265 9510 -255
rect 9455 -295 9465 -265
rect 9500 -295 9510 -265
rect 9455 -305 9510 -295
rect 9540 -265 9595 -255
rect 9540 -295 9550 -265
rect 9585 -295 9595 -265
rect 9540 -305 9595 -295
rect 9625 -265 9680 -255
rect 9625 -295 9635 -265
rect 9670 -295 9680 -265
rect 9625 -305 9680 -295
rect 9710 -265 9765 -255
rect 9710 -295 9720 -265
rect 9755 -295 9765 -265
rect 9710 -305 9765 -295
rect 9795 -265 9850 -255
rect 9795 -295 9805 -265
rect 9840 -295 9850 -265
rect 9795 -305 9850 -295
rect 9880 -265 9935 -255
rect 9880 -295 9890 -265
rect 9925 -295 9935 -265
rect 9880 -305 9935 -295
rect 9965 -265 10020 -255
rect 9965 -295 9975 -265
rect 10010 -295 10020 -265
rect 9965 -305 10020 -295
rect 10050 -265 10105 -255
rect 10050 -295 10060 -265
rect 10095 -295 10105 -265
rect 10050 -305 10105 -295
rect 10135 -265 10190 -255
rect 10135 -295 10145 -265
rect 10180 -295 10190 -265
rect 10135 -305 10190 -295
rect 10220 -265 10275 -255
rect 10220 -295 10230 -265
rect 10265 -295 10275 -265
rect 10220 -305 10275 -295
rect 10305 -265 10360 -255
rect 10305 -295 10315 -265
rect 10350 -295 10360 -265
rect 10305 -305 10360 -295
rect 10390 -265 10445 -255
rect 10390 -295 10400 -265
rect 10435 -295 10445 -265
rect 10390 -305 10445 -295
rect 10475 -265 10530 -255
rect 10475 -295 10485 -265
rect 10520 -295 10530 -265
rect 10475 -305 10530 -295
rect 10560 -265 10615 -255
rect 10560 -295 10570 -265
rect 10605 -295 10615 -265
rect 10560 -305 10615 -295
rect 10645 -265 10700 -255
rect 10645 -295 10655 -265
rect 10690 -295 10700 -265
rect 10645 -305 10700 -295
rect 10730 -265 10785 -255
rect 10730 -295 10740 -265
rect 10775 -295 10785 -265
rect 10730 -305 10785 -295
rect 10815 -265 10870 -255
rect 10815 -295 10825 -265
rect 10860 -295 10870 -265
rect 10815 -305 10870 -295
rect 10900 -265 10955 -255
rect 10900 -295 10910 -265
rect 10945 -295 10955 -265
rect 10900 -305 10955 -295
rect 10985 -265 11040 -255
rect 10985 -295 10995 -265
rect 11030 -295 11040 -265
rect 10985 -305 11040 -295
rect 11070 -265 11125 -255
rect 11070 -295 11080 -265
rect 11115 -295 11125 -265
rect 11070 -305 11125 -295
rect 11155 -265 11210 -255
rect 11155 -295 11165 -265
rect 11200 -295 11210 -265
rect 11155 -305 11210 -295
rect 11240 -265 11295 -255
rect 11240 -295 11250 -265
rect 11285 -295 11295 -265
rect 11240 -305 11295 -295
rect 11325 -265 11380 -255
rect 11325 -295 11335 -265
rect 11370 -295 11380 -265
rect 11325 -305 11380 -295
rect 11410 -265 11465 -255
rect 11410 -295 11420 -265
rect 11455 -295 11465 -265
rect 11410 -305 11465 -295
rect 11495 -265 11550 -255
rect 11495 -295 11505 -265
rect 11540 -295 11550 -265
rect 11495 -305 11550 -295
rect 11580 -265 11635 -255
rect 11580 -295 11590 -265
rect 11625 -295 11635 -265
rect 11580 -305 11635 -295
rect 11665 -265 11720 -255
rect 11665 -295 11675 -265
rect 11710 -295 11720 -265
rect 11665 -305 11720 -295
rect 11750 -265 11805 -255
rect 11750 -295 11760 -265
rect 11795 -295 11805 -265
rect 11750 -305 11805 -295
rect 11835 -265 11890 -255
rect 11835 -295 11845 -265
rect 11880 -295 11890 -265
rect 11835 -305 11890 -295
rect 11920 -265 11975 -255
rect 11920 -295 11930 -265
rect 11965 -295 11975 -265
rect 11920 -305 11975 -295
rect 12005 -265 12060 -255
rect 12005 -295 12015 -265
rect 12050 -295 12060 -265
rect 12005 -305 12060 -295
rect 12090 -265 12145 -255
rect 12090 -295 12100 -265
rect 12135 -295 12145 -265
rect 12090 -305 12145 -295
rect 12175 -265 12230 -255
rect 12175 -295 12185 -265
rect 12220 -295 12230 -265
rect 12175 -305 12230 -295
rect 12260 -265 12315 -255
rect 12260 -295 12270 -265
rect 12305 -295 12315 -265
rect 12260 -305 12315 -295
rect 12345 -265 12400 -255
rect 12345 -295 12355 -265
rect 12390 -295 12400 -265
rect 12345 -305 12400 -295
rect 12430 -265 12485 -255
rect 12430 -295 12440 -265
rect 12475 -295 12485 -265
rect 12430 -305 12485 -295
rect 12515 -265 12570 -255
rect 12515 -295 12525 -265
rect 12560 -295 12570 -265
rect 12515 -305 12570 -295
rect 12600 -265 12655 -255
rect 12600 -295 12610 -265
rect 12645 -295 12655 -265
rect 12600 -305 12655 -295
rect 12685 -265 12740 -255
rect 12685 -295 12695 -265
rect 12730 -295 12740 -265
rect 12685 -305 12740 -295
rect 12770 -265 12825 -255
rect 12770 -295 12780 -265
rect 12815 -295 12825 -265
rect 12770 -305 12825 -295
rect 12855 -265 12910 -255
rect 12855 -295 12865 -265
rect 12900 -295 12910 -265
rect 12855 -305 12910 -295
rect 12940 -265 12995 -255
rect 12940 -295 12950 -265
rect 12985 -295 12995 -265
rect 12940 -305 12995 -295
rect 13025 -265 13080 -255
rect 13025 -295 13035 -265
rect 13070 -295 13080 -265
rect 13025 -305 13080 -295
rect 13110 -265 13165 -255
rect 13110 -295 13120 -265
rect 13155 -295 13165 -265
rect 13110 -305 13165 -295
rect 13195 -265 13250 -255
rect 13195 -295 13205 -265
rect 13240 -295 13250 -265
rect 13195 -305 13250 -295
rect 13280 -265 13335 -255
rect 13280 -295 13290 -265
rect 13325 -295 13335 -265
rect 13280 -305 13335 -295
rect 13365 -265 13420 -255
rect 13365 -295 13375 -265
rect 13410 -295 13420 -265
rect 13365 -305 13420 -295
rect 13450 -265 13505 -255
rect 13450 -295 13460 -265
rect 13495 -295 13505 -265
rect 13450 -305 13505 -295
rect 13535 -265 13590 -255
rect 13535 -295 13545 -265
rect 13580 -295 13590 -265
rect 13535 -305 13590 -295
rect 13620 -265 13675 -255
rect 13620 -295 13630 -265
rect 13665 -295 13675 -265
rect 13620 -305 13675 -295
rect 13705 -265 13760 -255
rect 13705 -295 13715 -265
rect 13750 -295 13760 -265
rect 13705 -305 13760 -295
rect 13790 -265 13845 -255
rect 13790 -295 13800 -265
rect 13835 -295 13845 -265
rect 13790 -305 13845 -295
rect 13875 -265 13930 -255
rect 13875 -295 13885 -265
rect 13920 -295 13930 -265
rect 13875 -305 13930 -295
rect 13960 -265 14015 -255
rect 13960 -295 13970 -265
rect 14005 -295 14015 -265
rect 13960 -305 14015 -295
rect 14045 -265 14100 -255
rect 14045 -295 14055 -265
rect 14090 -295 14100 -265
rect 14045 -305 14100 -295
rect 14130 -265 14185 -255
rect 14130 -295 14140 -265
rect 14175 -295 14185 -265
rect 14130 -305 14185 -295
rect 14215 -265 14270 -255
rect 14215 -295 14225 -265
rect 14260 -295 14270 -265
rect 14215 -305 14270 -295
rect 14300 -265 14355 -255
rect 14300 -295 14310 -265
rect 14345 -295 14355 -265
rect 14300 -305 14355 -295
rect 14385 -265 14440 -255
rect 14385 -295 14395 -265
rect 14430 -295 14440 -265
rect 14385 -305 14440 -295
rect 14470 -265 14525 -255
rect 14470 -295 14480 -265
rect 14515 -295 14525 -265
rect 14470 -305 14525 -295
rect 14555 -265 14610 -255
rect 14555 -295 14565 -265
rect 14600 -295 14610 -265
rect 14555 -305 14610 -295
rect 14640 -265 14695 -255
rect 14640 -295 14650 -265
rect 14685 -295 14695 -265
rect 14640 -305 14695 -295
rect 14725 -265 14780 -255
rect 14725 -295 14735 -265
rect 14770 -295 14780 -265
rect 14725 -305 14780 -295
rect 14810 -265 14865 -255
rect 14810 -295 14820 -265
rect 14855 -295 14865 -265
rect 14810 -305 14865 -295
rect 14895 -265 14950 -255
rect 14895 -295 14905 -265
rect 14940 -295 14950 -265
rect 14895 -305 14950 -295
rect 14980 -265 15035 -255
rect 14980 -295 14990 -265
rect 15025 -295 15035 -265
rect 14980 -305 15035 -295
rect 15065 -265 15120 -255
rect 15065 -295 15075 -265
rect 15110 -295 15120 -265
rect 15065 -305 15120 -295
rect 15150 -265 15205 -255
rect 15150 -295 15160 -265
rect 15195 -295 15205 -265
rect 15150 -305 15205 -295
rect 15235 -265 15290 -255
rect 15235 -295 15245 -265
rect 15280 -295 15290 -265
rect 15235 -305 15290 -295
rect 15320 -265 15375 -255
rect 15320 -295 15330 -265
rect 15365 -295 15375 -265
rect 15320 -305 15375 -295
rect 15405 -265 15460 -255
rect 15405 -295 15415 -265
rect 15450 -295 15460 -265
rect 15405 -305 15460 -295
rect 15490 -265 15545 -255
rect 15490 -295 15500 -265
rect 15535 -295 15545 -265
rect 15490 -305 15545 -295
rect 15575 -265 15630 -255
rect 15575 -295 15585 -265
rect 15620 -295 15630 -265
rect 15575 -305 15630 -295
rect 15660 -265 15715 -255
rect 15660 -295 15670 -265
rect 15705 -295 15715 -265
rect 15660 -305 15715 -295
rect 15745 -265 15800 -255
rect 15745 -295 15755 -265
rect 15790 -295 15800 -265
rect 15745 -305 15800 -295
rect 15830 -265 15885 -255
rect 15830 -295 15840 -265
rect 15875 -295 15885 -265
rect 15830 -305 15885 -295
rect 15915 -265 15970 -255
rect 15915 -295 15925 -265
rect 15960 -295 15970 -265
rect 15915 -305 15970 -295
rect 16000 -265 16055 -255
rect 16000 -295 16010 -265
rect 16045 -295 16055 -265
rect 16000 -305 16055 -295
rect 16085 -265 16140 -255
rect 16085 -295 16095 -265
rect 16130 -295 16140 -265
rect 16085 -305 16140 -295
rect 16170 -265 16225 -255
rect 16170 -295 16180 -265
rect 16215 -295 16225 -265
rect 16170 -305 16225 -295
rect 16255 -265 16310 -255
rect 16255 -295 16265 -265
rect 16300 -295 16310 -265
rect 16255 -305 16310 -295
rect 16340 -265 16395 -255
rect 16340 -295 16350 -265
rect 16385 -295 16395 -265
rect 16340 -305 16395 -295
rect 16425 -265 16480 -255
rect 16425 -295 16435 -265
rect 16470 -295 16480 -265
rect 16425 -305 16480 -295
rect 16510 -265 16565 -255
rect 16510 -295 16520 -265
rect 16555 -295 16565 -265
rect 16510 -305 16565 -295
rect 16595 -265 16650 -255
rect 16595 -295 16605 -265
rect 16640 -295 16650 -265
rect 16595 -305 16650 -295
rect 16680 -265 16735 -255
rect 16680 -295 16690 -265
rect 16725 -295 16735 -265
rect 16680 -305 16735 -295
rect 16765 -265 16820 -255
rect 16765 -295 16775 -265
rect 16810 -295 16820 -265
rect 16765 -305 16820 -295
rect 16850 -265 16905 -255
rect 16850 -295 16860 -265
rect 16895 -295 16905 -265
rect 16850 -305 16905 -295
rect 16935 -265 16990 -255
rect 16935 -295 16945 -265
rect 16980 -295 16990 -265
rect 16935 -305 16990 -295
rect 17020 -265 17075 -255
rect 17020 -295 17030 -265
rect 17065 -295 17075 -265
rect 17020 -305 17075 -295
rect 17105 -265 17160 -255
rect 17105 -295 17115 -265
rect 17150 -295 17160 -265
rect 17105 -305 17160 -295
rect 17190 -265 17245 -255
rect 17190 -295 17200 -265
rect 17235 -295 17245 -265
rect 17190 -305 17245 -295
rect 17275 -265 17330 -255
rect 17275 -295 17285 -265
rect 17320 -295 17330 -265
rect 17275 -305 17330 -295
rect 17360 -265 17415 -255
rect 17360 -295 17370 -265
rect 17405 -295 17415 -265
rect 17360 -305 17415 -295
rect 17445 -265 17500 -255
rect 17445 -295 17455 -265
rect 17490 -295 17500 -265
rect 17445 -305 17500 -295
rect 17530 -265 17585 -255
rect 17530 -295 17540 -265
rect 17575 -295 17585 -265
rect 17530 -305 17585 -295
rect 17615 -265 17670 -255
rect 17615 -295 17625 -265
rect 17660 -295 17670 -265
rect 17615 -305 17670 -295
rect 17700 -265 17755 -255
rect 17700 -295 17710 -265
rect 17745 -295 17755 -265
rect 17700 -305 17755 -295
rect 17785 -265 17840 -255
rect 17785 -295 17795 -265
rect 17830 -295 17840 -265
rect 17785 -305 17840 -295
rect 17870 -265 17925 -255
rect 17870 -295 17880 -265
rect 17915 -295 17925 -265
rect 17870 -305 17925 -295
rect 17955 -265 18010 -255
rect 17955 -295 17965 -265
rect 18000 -295 18010 -265
rect 17955 -305 18010 -295
rect 18040 -265 18095 -255
rect 18040 -295 18050 -265
rect 18085 -295 18095 -265
rect 18040 -305 18095 -295
rect 18125 -265 18180 -255
rect 18125 -295 18135 -265
rect 18170 -295 18180 -265
rect 18125 -305 18180 -295
rect 18210 -265 18265 -255
rect 18210 -295 18220 -265
rect 18255 -295 18265 -265
rect 18210 -305 18265 -295
rect 18295 -265 18350 -255
rect 18295 -295 18305 -265
rect 18340 -295 18350 -265
rect 18295 -305 18350 -295
rect 18380 -265 18435 -255
rect 18380 -295 18390 -265
rect 18425 -295 18435 -265
rect 18380 -305 18435 -295
rect 18465 -265 18520 -255
rect 18465 -295 18475 -265
rect 18510 -295 18520 -265
rect 18465 -305 18520 -295
rect 18550 -265 18605 -255
rect 18550 -295 18560 -265
rect 18595 -295 18605 -265
rect 18550 -305 18605 -295
rect 18635 -265 18690 -255
rect 18635 -295 18645 -265
rect 18680 -295 18690 -265
rect 18635 -305 18690 -295
rect 18720 -265 18775 -255
rect 18720 -295 18730 -265
rect 18765 -295 18775 -265
rect 18720 -305 18775 -295
rect 18805 -265 18860 -255
rect 18805 -295 18815 -265
rect 18850 -295 18860 -265
rect 18805 -305 18860 -295
rect 18890 -265 18945 -255
rect 18890 -295 18900 -265
rect 18935 -295 18945 -265
rect 18890 -305 18945 -295
rect 18975 -265 19030 -255
rect 18975 -295 18985 -265
rect 19020 -295 19030 -265
rect 18975 -305 19030 -295
rect 19060 -265 19115 -255
rect 19060 -295 19070 -265
rect 19105 -295 19115 -265
rect 19060 -305 19115 -295
rect 19145 -265 19200 -255
rect 19145 -295 19155 -265
rect 19190 -295 19200 -265
rect 19145 -305 19200 -295
rect 19230 -265 19285 -255
rect 19230 -295 19240 -265
rect 19275 -295 19285 -265
rect 19230 -305 19285 -295
rect 19315 -265 19370 -255
rect 19315 -295 19325 -265
rect 19360 -295 19370 -265
rect 19315 -305 19370 -295
rect 19400 -265 19455 -255
rect 19400 -295 19410 -265
rect 19445 -295 19455 -265
rect 19400 -305 19455 -295
rect 19485 -265 19540 -255
rect 19485 -295 19495 -265
rect 19530 -295 19540 -265
rect 19485 -305 19540 -295
rect 19570 -265 19625 -255
rect 19570 -295 19580 -265
rect 19615 -295 19625 -265
rect 19570 -305 19625 -295
rect 19655 -265 19710 -255
rect 19655 -295 19665 -265
rect 19700 -295 19710 -265
rect 19655 -305 19710 -295
rect 19740 -265 19795 -255
rect 19740 -295 19750 -265
rect 19785 -295 19795 -265
rect 19740 -305 19795 -295
rect 19825 -265 19880 -255
rect 19825 -295 19835 -265
rect 19870 -295 19880 -265
rect 19825 -305 19880 -295
rect 19910 -265 19965 -255
rect 19910 -295 19920 -265
rect 19955 -295 19965 -265
rect 19910 -305 19965 -295
rect 19995 -265 20050 -255
rect 19995 -295 20005 -265
rect 20040 -295 20050 -265
rect 19995 -305 20050 -295
rect 20080 -265 20135 -255
rect 20080 -295 20090 -265
rect 20125 -295 20135 -265
rect 20080 -305 20135 -295
rect 20165 -265 20220 -255
rect 20165 -295 20175 -265
rect 20210 -295 20220 -265
rect 20165 -305 20220 -295
rect 20250 -265 20305 -255
rect 20250 -295 20260 -265
rect 20295 -295 20305 -265
rect 20250 -305 20305 -295
rect 20335 -265 20390 -255
rect 20335 -295 20345 -265
rect 20380 -295 20390 -265
rect 20335 -305 20390 -295
rect 20420 -265 20475 -255
rect 20420 -295 20430 -265
rect 20465 -295 20475 -265
rect 20420 -305 20475 -295
rect 20505 -265 20560 -255
rect 20505 -295 20515 -265
rect 20550 -295 20560 -265
rect 20505 -305 20560 -295
rect 20590 -265 20645 -255
rect 20590 -295 20600 -265
rect 20635 -295 20645 -265
rect 20590 -305 20645 -295
rect 20675 -265 20730 -255
rect 20675 -295 20685 -265
rect 20720 -295 20730 -265
rect 20675 -305 20730 -295
rect 20760 -265 20815 -255
rect 20760 -295 20770 -265
rect 20805 -295 20815 -265
rect 20760 -305 20815 -295
rect 20845 -265 20900 -255
rect 20845 -295 20855 -265
rect 20890 -295 20900 -265
rect 20845 -305 20900 -295
rect 20930 -265 20985 -255
rect 20930 -295 20940 -265
rect 20975 -295 20985 -265
rect 20930 -305 20985 -295
rect 21015 -265 21070 -255
rect 21015 -295 21025 -265
rect 21060 -295 21070 -265
rect 21015 -305 21070 -295
rect 21100 -265 21155 -255
rect 21100 -295 21110 -265
rect 21145 -295 21155 -265
rect 21100 -305 21155 -295
rect 21185 -265 21240 -255
rect 21185 -295 21195 -265
rect 21230 -295 21240 -265
rect 21185 -305 21240 -295
rect 21270 -265 21325 -255
rect 21270 -295 21280 -265
rect 21315 -295 21325 -265
rect 21270 -305 21325 -295
rect 21355 -265 21410 -255
rect 21355 -295 21365 -265
rect 21400 -295 21410 -265
rect 21355 -305 21410 -295
rect 21440 -265 21495 -255
rect 21440 -295 21450 -265
rect 21485 -295 21495 -265
rect 21440 -305 21495 -295
rect 21525 -265 21580 -255
rect 21525 -295 21535 -265
rect 21570 -295 21580 -265
rect 21525 -305 21580 -295
rect 21610 -265 21665 -255
rect 21610 -295 21620 -265
rect 21655 -295 21665 -265
rect 21610 -305 21665 -295
rect 21695 -265 21750 -255
rect 21695 -295 21705 -265
rect 21740 -295 21750 -265
rect 21695 -305 21750 -295
rect 21780 -265 21835 -255
rect 21780 -295 21790 -265
rect 21825 -295 21835 -265
rect 21780 -305 21835 -295
rect 21865 -265 21920 -255
rect 21865 -295 21875 -265
rect 21910 -295 21920 -265
rect 21865 -305 21920 -295
rect 21950 -265 22005 -255
rect 21950 -295 21960 -265
rect 21995 -295 22005 -265
rect 21950 -305 22005 -295
rect 22035 -265 22090 -255
rect 22035 -295 22045 -265
rect 22080 -295 22090 -265
rect 22035 -305 22090 -295
rect 22120 -265 22175 -255
rect 22120 -295 22130 -265
rect 22165 -295 22175 -265
rect 22120 -305 22175 -295
rect 22205 -265 22260 -255
rect 22205 -295 22215 -265
rect 22250 -295 22260 -265
rect 22205 -305 22260 -295
rect 22290 -265 22345 -255
rect 22290 -295 22300 -265
rect 22335 -295 22345 -265
rect 22290 -305 22345 -295
rect 22375 -265 22430 -255
rect 22375 -295 22385 -265
rect 22420 -295 22430 -265
rect 22375 -305 22430 -295
rect 22460 -265 22515 -255
rect 22460 -295 22470 -265
rect 22505 -295 22515 -265
rect 22460 -305 22515 -295
rect 22545 -265 22600 -255
rect 22545 -295 22555 -265
rect 22590 -295 22600 -265
rect 22545 -305 22600 -295
rect 22630 -265 22685 -255
rect 22630 -295 22640 -265
rect 22675 -295 22685 -265
rect 22630 -305 22685 -295
rect 22715 -265 22770 -255
rect 22715 -295 22725 -265
rect 22760 -295 22770 -265
rect 22715 -305 22770 -295
rect 22800 -265 22855 -255
rect 22800 -295 22810 -265
rect 22845 -295 22855 -265
rect 22800 -305 22855 -295
rect 22885 -265 22940 -255
rect 22885 -295 22895 -265
rect 22930 -295 22940 -265
rect 22885 -305 22940 -295
rect 22970 -265 23025 -255
rect 22970 -295 22980 -265
rect 23015 -295 23025 -265
rect 22970 -305 23025 -295
rect 23055 -265 23110 -255
rect 23055 -295 23065 -265
rect 23100 -295 23110 -265
rect 23055 -305 23110 -295
rect 23140 -265 23195 -255
rect 23140 -295 23150 -265
rect 23185 -295 23195 -265
rect 23140 -305 23195 -295
rect 23225 -265 23280 -255
rect 23225 -295 23235 -265
rect 23270 -295 23280 -265
rect 23225 -305 23280 -295
rect 23310 -265 23365 -255
rect 23310 -295 23320 -265
rect 23355 -295 23365 -265
rect 23310 -305 23365 -295
rect 23395 -265 23450 -255
rect 23395 -295 23405 -265
rect 23440 -295 23450 -265
rect 23395 -305 23450 -295
rect 23480 -265 23535 -255
rect 23480 -295 23490 -265
rect 23525 -295 23535 -265
rect 23480 -305 23535 -295
rect 23565 -265 23620 -255
rect 23565 -295 23575 -265
rect 23610 -295 23620 -265
rect 23565 -305 23620 -295
rect 23650 -265 23705 -255
rect 23650 -295 23660 -265
rect 23695 -295 23705 -265
rect 23650 -305 23705 -295
rect 23735 -265 23790 -255
rect 23735 -295 23745 -265
rect 23780 -295 23790 -265
rect 23735 -305 23790 -295
rect 23820 -265 23875 -255
rect 23820 -295 23830 -265
rect 23865 -295 23875 -265
rect 23820 -305 23875 -295
rect 23905 -265 23960 -255
rect 23905 -295 23915 -265
rect 23950 -295 23960 -265
rect 23905 -305 23960 -295
rect 23990 -265 24045 -255
rect 23990 -295 24000 -265
rect 24035 -295 24045 -265
rect 23990 -305 24045 -295
rect 24075 -265 24130 -255
rect 24075 -295 24085 -265
rect 24120 -295 24130 -265
rect 24075 -305 24130 -295
rect 24160 -265 24215 -255
rect 24160 -295 24170 -265
rect 24205 -295 24215 -265
rect 24160 -305 24215 -295
rect 24245 -265 24300 -255
rect 24245 -295 24255 -265
rect 24290 -295 24300 -265
rect 24245 -305 24300 -295
rect 24330 -265 24385 -255
rect 24330 -295 24340 -265
rect 24375 -295 24385 -265
rect 24330 -305 24385 -295
rect 24415 -265 24470 -255
rect 24415 -295 24425 -265
rect 24460 -295 24470 -265
rect 24415 -305 24470 -295
rect 24500 -265 24555 -255
rect 24500 -295 24510 -265
rect 24545 -295 24555 -265
rect 24500 -305 24555 -295
rect 24585 -265 24640 -255
rect 24585 -295 24595 -265
rect 24630 -295 24640 -265
rect 24585 -305 24640 -295
rect 24670 -265 24725 -255
rect 24670 -295 24680 -265
rect 24715 -295 24725 -265
rect 24670 -305 24725 -295
rect 24755 -265 24810 -255
rect 24755 -295 24765 -265
rect 24800 -295 24810 -265
rect 24755 -305 24810 -295
rect 24840 -265 24895 -255
rect 24840 -295 24850 -265
rect 24885 -295 24895 -265
rect 24840 -305 24895 -295
rect 24925 -265 24980 -255
rect 24925 -295 24935 -265
rect 24970 -295 24980 -265
rect 24925 -305 24980 -295
rect 25010 -265 25065 -255
rect 25010 -295 25020 -265
rect 25055 -295 25065 -265
rect 25010 -305 25065 -295
rect 25095 -265 25150 -255
rect 25095 -295 25105 -265
rect 25140 -295 25150 -265
rect 25095 -305 25150 -295
rect 25180 -265 25235 -255
rect 25180 -295 25190 -265
rect 25225 -295 25235 -265
rect 25180 -305 25235 -295
rect 25265 -265 25320 -255
rect 25265 -295 25275 -265
rect 25310 -295 25320 -265
rect 25265 -305 25320 -295
rect 25350 -265 25405 -255
rect 25350 -295 25360 -265
rect 25395 -295 25405 -265
rect 25350 -305 25405 -295
rect 25435 -265 25490 -255
rect 25435 -295 25445 -265
rect 25480 -295 25490 -265
rect 25435 -305 25490 -295
rect 25520 -265 25575 -255
rect 25520 -295 25530 -265
rect 25565 -295 25575 -265
rect 25520 -305 25575 -295
rect 25605 -265 25660 -255
rect 25605 -295 25615 -265
rect 25650 -295 25660 -265
rect 25605 -305 25660 -295
rect 25690 -265 25745 -255
rect 25690 -295 25700 -265
rect 25735 -295 25745 -265
rect 25690 -305 25745 -295
rect 25775 -265 25830 -255
rect 25775 -295 25785 -265
rect 25820 -295 25830 -265
rect 25775 -305 25830 -295
rect 25860 -265 25915 -255
rect 25860 -295 25870 -265
rect 25905 -295 25915 -265
rect 25860 -305 25915 -295
rect 25945 -265 26000 -255
rect 25945 -295 25955 -265
rect 25990 -295 26000 -265
rect 25945 -305 26000 -295
rect 26030 -265 26085 -255
rect 26030 -295 26040 -265
rect 26075 -295 26085 -265
rect 26030 -305 26085 -295
rect 26115 -265 26170 -255
rect 26115 -295 26125 -265
rect 26160 -295 26170 -265
rect 26115 -305 26170 -295
rect 26200 -265 26255 -255
rect 26200 -295 26210 -265
rect 26245 -295 26255 -265
rect 26200 -305 26255 -295
rect 26285 -265 26340 -255
rect 26285 -295 26295 -265
rect 26330 -295 26340 -265
rect 26285 -305 26340 -295
rect 26370 -265 26425 -255
rect 26370 -295 26380 -265
rect 26415 -295 26425 -265
rect 26370 -305 26425 -295
rect 26455 -265 26510 -255
rect 26455 -295 26465 -265
rect 26500 -295 26510 -265
rect 26455 -305 26510 -295
rect 26540 -265 26595 -255
rect 26540 -295 26550 -265
rect 26585 -295 26595 -265
rect 26540 -305 26595 -295
rect 26625 -265 26680 -255
rect 26625 -295 26635 -265
rect 26670 -295 26680 -265
rect 26625 -305 26680 -295
rect 26710 -265 26765 -255
rect 26710 -295 26720 -265
rect 26755 -295 26765 -265
rect 26710 -305 26765 -295
rect 26795 -265 26850 -255
rect 26795 -295 26805 -265
rect 26840 -295 26850 -265
rect 26795 -305 26850 -295
rect 26880 -265 26935 -255
rect 26880 -295 26890 -265
rect 26925 -295 26935 -265
rect 26880 -305 26935 -295
rect 26965 -265 27020 -255
rect 26965 -295 26975 -265
rect 27010 -295 27020 -265
rect 26965 -305 27020 -295
rect 27050 -265 27105 -255
rect 27050 -295 27060 -265
rect 27095 -295 27105 -265
rect 27050 -305 27105 -295
rect 27135 -265 27190 -255
rect 27135 -295 27145 -265
rect 27180 -295 27190 -265
rect 27135 -305 27190 -295
rect 27220 -265 27275 -255
rect 27220 -295 27230 -265
rect 27265 -295 27275 -265
rect 27220 -305 27275 -295
rect 27305 -265 27360 -255
rect 27305 -295 27315 -265
rect 27350 -295 27360 -265
rect 27305 -305 27360 -295
rect 27390 -265 27445 -255
rect 27390 -295 27400 -265
rect 27435 -295 27445 -265
rect 27390 -305 27445 -295
rect 27475 -265 27530 -255
rect 27475 -295 27485 -265
rect 27520 -295 27530 -265
rect 27475 -305 27530 -295
rect 27560 -265 27615 -255
rect 27560 -295 27570 -265
rect 27605 -295 27615 -265
rect 27560 -305 27615 -295
rect 27645 -265 27700 -255
rect 27645 -295 27655 -265
rect 27690 -295 27700 -265
rect 27645 -305 27700 -295
rect 27730 -265 27785 -255
rect 27730 -295 27740 -265
rect 27775 -295 27785 -265
rect 27730 -305 27785 -295
rect 27815 -265 27870 -255
rect 27815 -295 27825 -265
rect 27860 -295 27870 -265
rect 27815 -305 27870 -295
rect 27900 -265 27955 -255
rect 27900 -295 27910 -265
rect 27945 -295 27955 -265
rect 27900 -305 27955 -295
rect 27985 -265 28040 -255
rect 27985 -295 27995 -265
rect 28030 -295 28040 -265
rect 27985 -305 28040 -295
rect 28070 -265 28125 -255
rect 28070 -295 28080 -265
rect 28115 -295 28125 -265
rect 28070 -305 28125 -295
rect 28155 -265 28210 -255
rect 28155 -295 28165 -265
rect 28200 -295 28210 -265
rect 28155 -305 28210 -295
rect 28240 -265 28295 -255
rect 28240 -295 28250 -265
rect 28285 -295 28295 -265
rect 28240 -305 28295 -295
rect 28325 -265 28380 -255
rect 28325 -295 28335 -265
rect 28370 -295 28380 -265
rect 28325 -305 28380 -295
rect 28410 -265 28465 -255
rect 28410 -295 28420 -265
rect 28455 -295 28465 -265
rect 28410 -305 28465 -295
rect 28495 -265 28550 -255
rect 28495 -295 28505 -265
rect 28540 -295 28550 -265
rect 28495 -305 28550 -295
rect 28580 -265 28635 -255
rect 28580 -295 28590 -265
rect 28625 -295 28635 -265
rect 28580 -305 28635 -295
rect 28665 -265 28720 -255
rect 28665 -295 28675 -265
rect 28710 -295 28720 -265
rect 28665 -305 28720 -295
rect 28750 -265 28805 -255
rect 28750 -295 28760 -265
rect 28795 -295 28805 -265
rect 28750 -305 28805 -295
rect 28835 -265 28890 -255
rect 28835 -295 28845 -265
rect 28880 -295 28890 -265
rect 28835 -305 28890 -295
rect 28920 -265 28975 -255
rect 28920 -295 28930 -265
rect 28965 -295 28975 -265
rect 28920 -305 28975 -295
rect 29005 -265 29060 -255
rect 29005 -295 29015 -265
rect 29050 -295 29060 -265
rect 29005 -305 29060 -295
rect 29090 -265 29145 -255
rect 29090 -295 29100 -265
rect 29135 -295 29145 -265
rect 29090 -305 29145 -295
rect 29175 -265 29230 -255
rect 29175 -295 29185 -265
rect 29220 -295 29230 -265
rect 29175 -305 29230 -295
rect 29260 -265 29315 -255
rect 29260 -295 29270 -265
rect 29305 -295 29315 -265
rect 29260 -305 29315 -295
rect 29345 -265 29400 -255
rect 29345 -295 29355 -265
rect 29390 -295 29400 -265
rect 29345 -305 29400 -295
rect 29430 -265 29485 -255
rect 29430 -295 29440 -265
rect 29475 -295 29485 -265
rect 29430 -305 29485 -295
rect 29515 -265 29570 -255
rect 29515 -295 29525 -265
rect 29560 -295 29570 -265
rect 29515 -305 29570 -295
rect 29600 -265 29655 -255
rect 29600 -295 29610 -265
rect 29645 -295 29655 -265
rect 29600 -305 29655 -295
rect 29685 -265 29740 -255
rect 29685 -295 29695 -265
rect 29730 -295 29740 -265
rect 29685 -305 29740 -295
rect 29770 -265 29825 -255
rect 29770 -295 29780 -265
rect 29815 -295 29825 -265
rect 29770 -305 29825 -295
rect 29855 -265 29910 -255
rect 29855 -295 29865 -265
rect 29900 -295 29910 -265
rect 29855 -305 29910 -295
rect 29940 -265 29995 -255
rect 29940 -295 29950 -265
rect 29985 -295 29995 -265
rect 29940 -305 29995 -295
rect 30025 -265 30080 -255
rect 30025 -295 30035 -265
rect 30070 -295 30080 -265
rect 30025 -305 30080 -295
rect 30110 -265 30165 -255
rect 30110 -295 30120 -265
rect 30155 -295 30165 -265
rect 30110 -305 30165 -295
rect 30195 -265 30250 -255
rect 30195 -295 30205 -265
rect 30240 -295 30250 -265
rect 30195 -305 30250 -295
rect 30280 -265 30335 -255
rect 30280 -295 30290 -265
rect 30325 -295 30335 -265
rect 30280 -305 30335 -295
rect 30365 -265 30420 -255
rect 30365 -295 30375 -265
rect 30410 -295 30420 -265
rect 30365 -305 30420 -295
rect 30450 -265 30505 -255
rect 30450 -295 30460 -265
rect 30495 -295 30505 -265
rect 30450 -305 30505 -295
rect 30535 -265 30590 -255
rect 30535 -295 30545 -265
rect 30580 -295 30590 -265
rect 30535 -305 30590 -295
rect 30620 -265 30675 -255
rect 30620 -295 30630 -265
rect 30665 -295 30675 -265
rect 30620 -305 30675 -295
rect 30705 -265 30760 -255
rect 30705 -295 30715 -265
rect 30750 -295 30760 -265
rect 30705 -305 30760 -295
rect 30790 -265 30845 -255
rect 30790 -295 30800 -265
rect 30835 -295 30845 -265
rect 30790 -305 30845 -295
rect 30875 -265 30930 -255
rect 30875 -295 30885 -265
rect 30920 -295 30930 -265
rect 30875 -305 30930 -295
rect 30960 -265 31015 -255
rect 30960 -295 30970 -265
rect 31005 -295 31015 -265
rect 30960 -305 31015 -295
rect 31045 -265 31100 -255
rect 31045 -295 31055 -265
rect 31090 -295 31100 -265
rect 31045 -305 31100 -295
rect 31130 -265 31185 -255
rect 31130 -295 31140 -265
rect 31175 -295 31185 -265
rect 31130 -305 31185 -295
rect 31215 -265 31270 -255
rect 31215 -295 31225 -265
rect 31260 -295 31270 -265
rect 31215 -305 31270 -295
rect 31300 -265 31355 -255
rect 31300 -295 31310 -265
rect 31345 -295 31355 -265
rect 31300 -305 31355 -295
rect 31385 -265 31440 -255
rect 31385 -295 31395 -265
rect 31430 -295 31440 -265
rect 31385 -305 31440 -295
rect 31470 -265 31525 -255
rect 31470 -295 31480 -265
rect 31515 -295 31525 -265
rect 31470 -305 31525 -295
rect 31555 -265 31610 -255
rect 31555 -295 31565 -265
rect 31600 -295 31610 -265
rect 31555 -305 31610 -295
rect 31640 -265 31695 -255
rect 31640 -295 31650 -265
rect 31685 -295 31695 -265
rect 31640 -305 31695 -295
rect 31725 -265 31780 -255
rect 31725 -295 31735 -265
rect 31770 -295 31780 -265
rect 31725 -305 31780 -295
rect 31810 -265 31865 -255
rect 31810 -295 31820 -265
rect 31855 -295 31865 -265
rect 31810 -305 31865 -295
rect 31895 -265 31950 -255
rect 31895 -295 31905 -265
rect 31940 -295 31950 -265
rect 31895 -305 31950 -295
rect 31980 -265 32035 -255
rect 31980 -295 31990 -265
rect 32025 -295 32035 -265
rect 31980 -305 32035 -295
rect 32065 -265 32120 -255
rect 32065 -295 32075 -265
rect 32110 -295 32120 -265
rect 32065 -305 32120 -295
rect 32150 -265 32205 -255
rect 32150 -295 32160 -265
rect 32195 -295 32205 -265
rect 32150 -305 32205 -295
rect 32235 -265 32290 -255
rect 32235 -295 32245 -265
rect 32280 -295 32290 -265
rect 32235 -305 32290 -295
rect 32320 -265 32375 -255
rect 32320 -295 32330 -265
rect 32365 -295 32375 -265
rect 32320 -305 32375 -295
rect 32405 -265 32460 -255
rect 32405 -295 32415 -265
rect 32450 -295 32460 -265
rect 32405 -305 32460 -295
rect 32490 -265 32545 -255
rect 32490 -295 32500 -265
rect 32535 -295 32545 -265
rect 32490 -305 32545 -295
rect 32575 -265 32630 -255
rect 32575 -295 32585 -265
rect 32620 -295 32630 -265
rect 32575 -305 32630 -295
rect 32660 -265 32715 -255
rect 32660 -295 32670 -265
rect 32705 -295 32715 -265
rect 32660 -305 32715 -295
rect 32745 -265 32800 -255
rect 32745 -295 32755 -265
rect 32790 -295 32800 -265
rect 32745 -305 32800 -295
rect 32830 -265 32885 -255
rect 32830 -295 32840 -265
rect 32875 -295 32885 -265
rect 32830 -305 32885 -295
rect 32915 -265 32970 -255
rect 32915 -295 32925 -265
rect 32960 -295 32970 -265
rect 32915 -305 32970 -295
rect 33000 -265 33055 -255
rect 33000 -295 33010 -265
rect 33045 -295 33055 -265
rect 33000 -305 33055 -295
rect 33085 -265 33140 -255
rect 33085 -295 33095 -265
rect 33130 -295 33140 -265
rect 33085 -305 33140 -295
rect 33170 -265 33225 -255
rect 33170 -295 33180 -265
rect 33215 -295 33225 -265
rect 33170 -305 33225 -295
rect 33255 -265 33310 -255
rect 33255 -295 33265 -265
rect 33300 -295 33310 -265
rect 33255 -305 33310 -295
rect 33340 -265 33395 -255
rect 33340 -295 33350 -265
rect 33385 -295 33395 -265
rect 33340 -305 33395 -295
rect 33425 -265 33480 -255
rect 33425 -295 33435 -265
rect 33470 -295 33480 -265
rect 33425 -305 33480 -295
rect 33510 -265 33565 -255
rect 33510 -295 33520 -265
rect 33555 -295 33565 -265
rect 33510 -305 33565 -295
rect 33595 -265 33650 -255
rect 33595 -295 33605 -265
rect 33640 -295 33650 -265
rect 33595 -305 33650 -295
rect 33680 -265 33735 -255
rect 33680 -295 33690 -265
rect 33725 -295 33735 -265
rect 33680 -305 33735 -295
rect 33765 -265 33820 -255
rect 33765 -295 33775 -265
rect 33810 -295 33820 -265
rect 33765 -305 33820 -295
rect 33850 -265 33905 -255
rect 33850 -295 33860 -265
rect 33895 -295 33905 -265
rect 33850 -305 33905 -295
rect 33935 -265 33990 -255
rect 33935 -295 33945 -265
rect 33980 -295 33990 -265
rect 33935 -305 33990 -295
rect 34020 -265 34075 -255
rect 34020 -295 34030 -265
rect 34065 -295 34075 -265
rect 34020 -305 34075 -295
rect 34105 -265 34160 -255
rect 34105 -295 34115 -265
rect 34150 -295 34160 -265
rect 34105 -305 34160 -295
rect 34190 -265 34245 -255
rect 34190 -295 34200 -265
rect 34235 -295 34245 -265
rect 34190 -305 34245 -295
rect 34275 -265 34330 -255
rect 34275 -295 34285 -265
rect 34320 -295 34330 -265
rect 34275 -305 34330 -295
rect 34360 -265 34415 -255
rect 34360 -295 34370 -265
rect 34405 -295 34415 -265
rect 34360 -305 34415 -295
rect 34445 -265 34500 -255
rect 34445 -295 34455 -265
rect 34490 -295 34500 -265
rect 34445 -305 34500 -295
rect 34530 -265 34585 -255
rect 34530 -295 34540 -265
rect 34575 -295 34585 -265
rect 34530 -305 34585 -295
rect 34615 -265 34670 -255
rect 34615 -295 34625 -265
rect 34660 -295 34670 -265
rect 34615 -305 34670 -295
rect 34700 -265 34755 -255
rect 34700 -295 34710 -265
rect 34745 -295 34755 -265
rect 34700 -305 34755 -295
rect 34785 -265 34840 -255
rect 34785 -295 34795 -265
rect 34830 -295 34840 -265
rect 34785 -305 34840 -295
rect 34870 -265 34925 -255
rect 34870 -295 34880 -265
rect 34915 -295 34925 -265
rect 34870 -305 34925 -295
rect 34955 -265 35010 -255
rect 34955 -295 34965 -265
rect 35000 -295 35010 -265
rect 34955 -305 35010 -295
rect 35040 -265 35095 -255
rect 35040 -295 35050 -265
rect 35085 -295 35095 -265
rect 35040 -305 35095 -295
rect 35125 -265 35180 -255
rect 35125 -295 35135 -265
rect 35170 -295 35180 -265
rect 35125 -305 35180 -295
rect 35210 -265 35265 -255
rect 35210 -295 35220 -265
rect 35255 -295 35265 -265
rect 35210 -305 35265 -295
rect 35295 -265 35350 -255
rect 35295 -295 35305 -265
rect 35340 -295 35350 -265
rect 35295 -305 35350 -295
rect 35380 -265 35435 -255
rect 35380 -295 35390 -265
rect 35425 -295 35435 -265
rect 35380 -305 35435 -295
rect 35465 -265 35520 -255
rect 35465 -295 35475 -265
rect 35510 -295 35520 -265
rect 35465 -305 35520 -295
rect 35550 -265 35605 -255
rect 35550 -295 35560 -265
rect 35595 -295 35605 -265
rect 35550 -305 35605 -295
rect 35635 -265 35690 -255
rect 35635 -295 35645 -265
rect 35680 -295 35690 -265
rect 35635 -305 35690 -295
rect 35720 -265 35775 -255
rect 35720 -295 35730 -265
rect 35765 -295 35775 -265
rect 35720 -305 35775 -295
rect 35805 -265 35860 -255
rect 35805 -295 35815 -265
rect 35850 -295 35860 -265
rect 35805 -305 35860 -295
rect 35890 -265 35945 -255
rect 35890 -295 35900 -265
rect 35935 -295 35945 -265
rect 35890 -305 35945 -295
rect 35975 -265 36030 -255
rect 35975 -295 35985 -265
rect 36020 -295 36030 -265
rect 35975 -305 36030 -295
rect 36060 -265 36115 -255
rect 36060 -295 36070 -265
rect 36105 -295 36115 -265
rect 36060 -305 36115 -295
rect 36145 -265 36200 -255
rect 36145 -295 36155 -265
rect 36190 -295 36200 -265
rect 36145 -305 36200 -295
rect 36230 -265 36285 -255
rect 36230 -295 36240 -265
rect 36275 -295 36285 -265
rect 36230 -305 36285 -295
rect 36315 -265 36370 -255
rect 36315 -295 36325 -265
rect 36360 -295 36370 -265
rect 36315 -305 36370 -295
rect 36400 -265 36455 -255
rect 36400 -295 36410 -265
rect 36445 -295 36455 -265
rect 36400 -305 36455 -295
rect 36485 -265 36540 -255
rect 36485 -295 36495 -265
rect 36530 -295 36540 -265
rect 36485 -305 36540 -295
rect 36570 -265 36625 -255
rect 36570 -295 36580 -265
rect 36615 -295 36625 -265
rect 36570 -305 36625 -295
rect 36655 -265 36710 -255
rect 36655 -295 36665 -265
rect 36700 -295 36710 -265
rect 36655 -305 36710 -295
rect 36740 -265 36795 -255
rect 36740 -295 36750 -265
rect 36785 -295 36795 -265
rect 36740 -305 36795 -295
rect 36825 -265 36880 -255
rect 36825 -295 36835 -265
rect 36870 -295 36880 -265
rect 36825 -305 36880 -295
rect 36910 -265 36965 -255
rect 36910 -295 36920 -265
rect 36955 -295 36965 -265
rect 36910 -305 36965 -295
rect 36995 -265 37050 -255
rect 36995 -295 37005 -265
rect 37040 -295 37050 -265
rect 36995 -305 37050 -295
rect 37080 -265 37135 -255
rect 37080 -295 37090 -265
rect 37125 -295 37135 -265
rect 37080 -305 37135 -295
rect 37165 -265 37220 -255
rect 37165 -295 37175 -265
rect 37210 -295 37220 -265
rect 37165 -305 37220 -295
rect 37250 -265 37305 -255
rect 37250 -295 37260 -265
rect 37295 -295 37305 -265
rect 37250 -305 37305 -295
rect 37335 -265 37390 -255
rect 37335 -295 37345 -265
rect 37380 -295 37390 -265
rect 37335 -305 37390 -295
rect 37420 -265 37475 -255
rect 37420 -295 37430 -265
rect 37465 -295 37475 -265
rect 37420 -305 37475 -295
rect 37505 -265 37560 -255
rect 37505 -295 37515 -265
rect 37550 -295 37560 -265
rect 37505 -305 37560 -295
rect 37590 -265 37645 -255
rect 37590 -295 37600 -265
rect 37635 -295 37645 -265
rect 37590 -305 37645 -295
rect 37675 -265 37730 -255
rect 37675 -295 37685 -265
rect 37720 -295 37730 -265
rect 37675 -305 37730 -295
rect 37760 -265 37815 -255
rect 37760 -295 37770 -265
rect 37805 -295 37815 -265
rect 37760 -305 37815 -295
rect 37845 -265 37900 -255
rect 37845 -295 37855 -265
rect 37890 -295 37900 -265
rect 37845 -305 37900 -295
rect 37930 -265 37985 -255
rect 37930 -295 37940 -265
rect 37975 -295 37985 -265
rect 37930 -305 37985 -295
rect 38015 -265 38070 -255
rect 38015 -295 38025 -265
rect 38060 -295 38070 -265
rect 38015 -305 38070 -295
rect 38100 -265 38155 -255
rect 38100 -295 38110 -265
rect 38145 -295 38155 -265
rect 38100 -305 38155 -295
rect 38185 -265 38240 -255
rect 38185 -295 38195 -265
rect 38230 -295 38240 -265
rect 38185 -305 38240 -295
rect 38270 -265 38325 -255
rect 38270 -295 38280 -265
rect 38315 -295 38325 -265
rect 38270 -305 38325 -295
rect 38355 -265 38410 -255
rect 38355 -295 38365 -265
rect 38400 -295 38410 -265
rect 38355 -305 38410 -295
rect 38440 -265 38495 -255
rect 38440 -295 38450 -265
rect 38485 -295 38495 -265
rect 38440 -305 38495 -295
rect 38525 -265 38580 -255
rect 38525 -295 38535 -265
rect 38570 -295 38580 -265
rect 38525 -305 38580 -295
rect 38610 -265 38665 -255
rect 38610 -295 38620 -265
rect 38655 -295 38665 -265
rect 38610 -305 38665 -295
rect 38695 -265 38750 -255
rect 38695 -295 38705 -265
rect 38740 -295 38750 -265
rect 38695 -305 38750 -295
rect 38780 -265 38835 -255
rect 38780 -295 38790 -265
rect 38825 -295 38835 -265
rect 38780 -305 38835 -295
rect 38865 -265 38920 -255
rect 38865 -295 38875 -265
rect 38910 -295 38920 -265
rect 38865 -305 38920 -295
rect 38950 -265 39005 -255
rect 38950 -295 38960 -265
rect 38995 -295 39005 -265
rect 38950 -305 39005 -295
rect 39035 -265 39090 -255
rect 39035 -295 39045 -265
rect 39080 -295 39090 -265
rect 39035 -305 39090 -295
rect 39120 -265 39175 -255
rect 39120 -295 39130 -265
rect 39165 -295 39175 -265
rect 39120 -305 39175 -295
rect 39205 -265 39260 -255
rect 39205 -295 39215 -265
rect 39250 -295 39260 -265
rect 39205 -305 39260 -295
rect 39290 -265 39345 -255
rect 39290 -295 39300 -265
rect 39335 -295 39345 -265
rect 39290 -305 39345 -295
rect 39375 -265 39430 -255
rect 39375 -295 39385 -265
rect 39420 -295 39430 -265
rect 39375 -305 39430 -295
rect 39460 -265 39515 -255
rect 39460 -295 39470 -265
rect 39505 -295 39515 -265
rect 39460 -305 39515 -295
rect 39545 -265 39600 -255
rect 39545 -295 39555 -265
rect 39590 -295 39600 -265
rect 39545 -305 39600 -295
rect 39630 -265 39685 -255
rect 39630 -295 39640 -265
rect 39675 -295 39685 -265
rect 39630 -305 39685 -295
rect 39715 -265 39770 -255
rect 39715 -295 39725 -265
rect 39760 -295 39770 -265
rect 39715 -305 39770 -295
rect 39800 -265 39855 -255
rect 39800 -295 39810 -265
rect 39845 -295 39855 -265
rect 39800 -305 39855 -295
rect 39885 -265 39940 -255
rect 39885 -295 39895 -265
rect 39930 -295 39940 -265
rect 39885 -305 39940 -295
rect 39970 -265 40025 -255
rect 39970 -295 39980 -265
rect 40015 -295 40025 -265
rect 39970 -305 40025 -295
rect 40055 -265 40110 -255
rect 40055 -295 40065 -265
rect 40100 -295 40110 -265
rect 40055 -305 40110 -295
rect 40140 -265 40195 -255
rect 40140 -295 40150 -265
rect 40185 -295 40195 -265
rect 40140 -305 40195 -295
rect 40225 -265 40280 -255
rect 40225 -295 40235 -265
rect 40270 -295 40280 -265
rect 40225 -305 40280 -295
rect 40310 -265 40365 -255
rect 40310 -295 40320 -265
rect 40355 -295 40365 -265
rect 40310 -305 40365 -295
rect 40395 -265 40450 -255
rect 40395 -295 40405 -265
rect 40440 -295 40450 -265
rect 40395 -305 40450 -295
rect 40480 -265 40535 -255
rect 40480 -295 40490 -265
rect 40525 -295 40535 -265
rect 40480 -305 40535 -295
rect 40565 -265 40620 -255
rect 40565 -295 40575 -265
rect 40610 -295 40620 -265
rect 40565 -305 40620 -295
rect 40650 -265 40705 -255
rect 40650 -295 40660 -265
rect 40695 -295 40705 -265
rect 40650 -305 40705 -295
rect 40735 -265 40790 -255
rect 40735 -295 40745 -265
rect 40780 -295 40790 -265
rect 40735 -305 40790 -295
rect 40820 -265 40875 -255
rect 40820 -295 40830 -265
rect 40865 -295 40875 -265
rect 40820 -305 40875 -295
rect 40905 -265 40960 -255
rect 40905 -295 40915 -265
rect 40950 -295 40960 -265
rect 40905 -305 40960 -295
rect 40990 -265 41045 -255
rect 40990 -295 41000 -265
rect 41035 -295 41045 -265
rect 40990 -305 41045 -295
rect 41075 -265 41130 -255
rect 41075 -295 41085 -265
rect 41120 -295 41130 -265
rect 41075 -305 41130 -295
rect 41160 -265 41215 -255
rect 41160 -295 41170 -265
rect 41205 -295 41215 -265
rect 41160 -305 41215 -295
rect 41245 -265 41300 -255
rect 41245 -295 41255 -265
rect 41290 -295 41300 -265
rect 41245 -305 41300 -295
rect 41330 -265 41385 -255
rect 41330 -295 41340 -265
rect 41375 -295 41385 -265
rect 41330 -305 41385 -295
rect 41415 -265 41470 -255
rect 41415 -295 41425 -265
rect 41460 -295 41470 -265
rect 41415 -305 41470 -295
rect 41500 -265 41555 -255
rect 41500 -295 41510 -265
rect 41545 -295 41555 -265
rect 41500 -305 41555 -295
rect 41585 -265 41640 -255
rect 41585 -295 41595 -265
rect 41630 -295 41640 -265
rect 41585 -305 41640 -295
rect 41670 -265 41725 -255
rect 41670 -295 41680 -265
rect 41715 -295 41725 -265
rect 41670 -305 41725 -295
rect 41755 -265 41810 -255
rect 41755 -295 41765 -265
rect 41800 -295 41810 -265
rect 41755 -305 41810 -295
rect 41840 -265 41895 -255
rect 41840 -295 41850 -265
rect 41885 -295 41895 -265
rect 41840 -305 41895 -295
rect 41925 -265 41980 -255
rect 41925 -295 41935 -265
rect 41970 -295 41980 -265
rect 41925 -305 41980 -295
rect 42010 -265 42065 -255
rect 42010 -295 42020 -265
rect 42055 -295 42065 -265
rect 42010 -305 42065 -295
rect 42095 -265 42150 -255
rect 42095 -295 42105 -265
rect 42140 -295 42150 -265
rect 42095 -305 42150 -295
rect 42180 -265 42235 -255
rect 42180 -295 42190 -265
rect 42225 -295 42235 -265
rect 42180 -305 42235 -295
rect 42265 -265 42320 -255
rect 42265 -295 42275 -265
rect 42310 -295 42320 -265
rect 42265 -305 42320 -295
rect 42350 -265 42405 -255
rect 42350 -295 42360 -265
rect 42395 -295 42405 -265
rect 42350 -305 42405 -295
rect 42435 -265 42490 -255
rect 42435 -295 42445 -265
rect 42480 -295 42490 -265
rect 42435 -305 42490 -295
rect 42520 -265 42575 -255
rect 42520 -295 42530 -265
rect 42565 -295 42575 -265
rect 42520 -305 42575 -295
rect 42605 -265 42660 -255
rect 42605 -295 42615 -265
rect 42650 -295 42660 -265
rect 42605 -305 42660 -295
rect 42690 -265 42745 -255
rect 42690 -295 42700 -265
rect 42735 -295 42745 -265
rect 42690 -305 42745 -295
rect 42775 -265 42830 -255
rect 42775 -295 42785 -265
rect 42820 -295 42830 -265
rect 42775 -305 42830 -295
rect 42860 -265 42915 -255
rect 42860 -295 42870 -265
rect 42905 -295 42915 -265
rect 42860 -305 42915 -295
rect 42945 -265 43000 -255
rect 42945 -295 42955 -265
rect 42990 -295 43000 -265
rect 42945 -305 43000 -295
rect 43030 -265 43085 -255
rect 43030 -295 43040 -265
rect 43075 -295 43085 -265
rect 43030 -305 43085 -295
rect 43115 -265 43170 -255
rect 43115 -295 43125 -265
rect 43160 -295 43170 -265
rect 43115 -305 43170 -295
rect 43200 -265 43255 -255
rect 43200 -295 43210 -265
rect 43245 -295 43255 -265
rect 43200 -305 43255 -295
rect 43285 -265 43340 -255
rect 43285 -295 43295 -265
rect 43330 -295 43340 -265
rect 43285 -305 43340 -295
rect 43370 -265 43425 -255
rect 43370 -295 43380 -265
rect 43415 -295 43425 -265
rect 43370 -305 43425 -295
rect 43455 -265 43510 -255
rect 43455 -295 43465 -265
rect 43500 -295 43510 -265
rect 43455 -305 43510 -295
rect 43540 -265 43595 -255
rect 43540 -295 43550 -265
rect 43585 -295 43595 -265
rect 43540 -305 43595 -295
rect 125 -325 140 -305
rect 210 -325 225 -305
rect 295 -325 310 -305
rect 380 -325 395 -305
rect 465 -325 480 -305
rect 550 -325 565 -305
rect 635 -325 650 -305
rect 720 -325 735 -305
rect 805 -325 820 -305
rect 890 -325 905 -305
rect 975 -325 990 -305
rect 1060 -325 1075 -305
rect 1145 -325 1160 -305
rect 1230 -325 1245 -305
rect 1315 -325 1330 -305
rect 1400 -325 1415 -305
rect 1485 -325 1500 -305
rect 1570 -325 1585 -305
rect 1655 -325 1670 -305
rect 1740 -325 1755 -305
rect 1825 -325 1840 -305
rect 1910 -325 1925 -305
rect 1995 -325 2010 -305
rect 2080 -325 2095 -305
rect 2165 -325 2180 -305
rect 2250 -325 2265 -305
rect 2335 -325 2350 -305
rect 2420 -325 2435 -305
rect 2505 -325 2520 -305
rect 2590 -325 2605 -305
rect 2675 -325 2690 -305
rect 2760 -325 2775 -305
rect 2845 -325 2860 -305
rect 2930 -325 2945 -305
rect 3015 -325 3030 -305
rect 3100 -325 3115 -305
rect 3185 -325 3200 -305
rect 3270 -325 3285 -305
rect 3355 -325 3370 -305
rect 3440 -325 3455 -305
rect 3525 -325 3540 -305
rect 3610 -325 3625 -305
rect 3695 -325 3710 -305
rect 3780 -325 3795 -305
rect 3865 -325 3880 -305
rect 3950 -325 3965 -305
rect 4035 -325 4050 -305
rect 4120 -325 4135 -305
rect 4205 -325 4220 -305
rect 4290 -325 4305 -305
rect 4375 -325 4390 -305
rect 4460 -325 4475 -305
rect 4545 -325 4560 -305
rect 4630 -325 4645 -305
rect 4715 -325 4730 -305
rect 4800 -325 4815 -305
rect 4885 -325 4900 -305
rect 4970 -325 4985 -305
rect 5055 -325 5070 -305
rect 5140 -325 5155 -305
rect 5225 -325 5240 -305
rect 5310 -325 5325 -305
rect 5395 -325 5410 -305
rect 5480 -325 5495 -305
rect 5565 -325 5580 -305
rect 5650 -325 5665 -305
rect 5735 -325 5750 -305
rect 5820 -325 5835 -305
rect 5905 -325 5920 -305
rect 5990 -325 6005 -305
rect 6075 -325 6090 -305
rect 6160 -325 6175 -305
rect 6245 -325 6260 -305
rect 6330 -325 6345 -305
rect 6415 -325 6430 -305
rect 6500 -325 6515 -305
rect 6585 -325 6600 -305
rect 6670 -325 6685 -305
rect 6755 -325 6770 -305
rect 6840 -325 6855 -305
rect 6925 -325 6940 -305
rect 7010 -325 7025 -305
rect 7095 -325 7110 -305
rect 7180 -325 7195 -305
rect 7265 -325 7280 -305
rect 7350 -325 7365 -305
rect 7435 -325 7450 -305
rect 7520 -325 7535 -305
rect 7605 -325 7620 -305
rect 7690 -325 7705 -305
rect 7775 -325 7790 -305
rect 7860 -325 7875 -305
rect 7945 -325 7960 -305
rect 8030 -325 8045 -305
rect 8115 -325 8130 -305
rect 8200 -325 8215 -305
rect 8285 -325 8300 -305
rect 8370 -325 8385 -305
rect 8455 -325 8470 -305
rect 8540 -325 8555 -305
rect 8625 -325 8640 -305
rect 8710 -325 8725 -305
rect 8795 -325 8810 -305
rect 8880 -325 8895 -305
rect 8965 -325 8980 -305
rect 9050 -325 9065 -305
rect 9135 -325 9150 -305
rect 9220 -325 9235 -305
rect 9305 -325 9320 -305
rect 9390 -325 9405 -305
rect 9475 -325 9490 -305
rect 9560 -325 9575 -305
rect 9645 -325 9660 -305
rect 9730 -325 9745 -305
rect 9815 -325 9830 -305
rect 9900 -325 9915 -305
rect 9985 -325 10000 -305
rect 10070 -325 10085 -305
rect 10155 -325 10170 -305
rect 10240 -325 10255 -305
rect 10325 -325 10340 -305
rect 10410 -325 10425 -305
rect 10495 -325 10510 -305
rect 10580 -325 10595 -305
rect 10665 -325 10680 -305
rect 10750 -325 10765 -305
rect 10835 -325 10850 -305
rect 10920 -325 10935 -305
rect 11005 -325 11020 -305
rect 11090 -325 11105 -305
rect 11175 -325 11190 -305
rect 11260 -325 11275 -305
rect 11345 -325 11360 -305
rect 11430 -325 11445 -305
rect 11515 -325 11530 -305
rect 11600 -325 11615 -305
rect 11685 -325 11700 -305
rect 11770 -325 11785 -305
rect 11855 -325 11870 -305
rect 11940 -325 11955 -305
rect 12025 -325 12040 -305
rect 12110 -325 12125 -305
rect 12195 -325 12210 -305
rect 12280 -325 12295 -305
rect 12365 -325 12380 -305
rect 12450 -325 12465 -305
rect 12535 -325 12550 -305
rect 12620 -325 12635 -305
rect 12705 -325 12720 -305
rect 12790 -325 12805 -305
rect 12875 -325 12890 -305
rect 12960 -325 12975 -305
rect 13045 -325 13060 -305
rect 13130 -325 13145 -305
rect 13215 -325 13230 -305
rect 13300 -325 13315 -305
rect 13385 -325 13400 -305
rect 13470 -325 13485 -305
rect 13555 -325 13570 -305
rect 13640 -325 13655 -305
rect 13725 -325 13740 -305
rect 13810 -325 13825 -305
rect 13895 -325 13910 -305
rect 13980 -325 13995 -305
rect 14065 -325 14080 -305
rect 14150 -325 14165 -305
rect 14235 -325 14250 -305
rect 14320 -325 14335 -305
rect 14405 -325 14420 -305
rect 14490 -325 14505 -305
rect 14575 -325 14590 -305
rect 14660 -325 14675 -305
rect 14745 -325 14760 -305
rect 14830 -325 14845 -305
rect 14915 -325 14930 -305
rect 15000 -325 15015 -305
rect 15085 -325 15100 -305
rect 15170 -325 15185 -305
rect 15255 -325 15270 -305
rect 15340 -325 15355 -305
rect 15425 -325 15440 -305
rect 15510 -325 15525 -305
rect 15595 -325 15610 -305
rect 15680 -325 15695 -305
rect 15765 -325 15780 -305
rect 15850 -325 15865 -305
rect 15935 -325 15950 -305
rect 16020 -325 16035 -305
rect 16105 -325 16120 -305
rect 16190 -325 16205 -305
rect 16275 -325 16290 -305
rect 16360 -325 16375 -305
rect 16445 -325 16460 -305
rect 16530 -325 16545 -305
rect 16615 -325 16630 -305
rect 16700 -325 16715 -305
rect 16785 -325 16800 -305
rect 16870 -325 16885 -305
rect 16955 -325 16970 -305
rect 17040 -325 17055 -305
rect 17125 -325 17140 -305
rect 17210 -325 17225 -305
rect 17295 -325 17310 -305
rect 17380 -325 17395 -305
rect 17465 -325 17480 -305
rect 17550 -325 17565 -305
rect 17635 -325 17650 -305
rect 17720 -325 17735 -305
rect 17805 -325 17820 -305
rect 17890 -325 17905 -305
rect 17975 -325 17990 -305
rect 18060 -325 18075 -305
rect 18145 -325 18160 -305
rect 18230 -325 18245 -305
rect 18315 -325 18330 -305
rect 18400 -325 18415 -305
rect 18485 -325 18500 -305
rect 18570 -325 18585 -305
rect 18655 -325 18670 -305
rect 18740 -325 18755 -305
rect 18825 -325 18840 -305
rect 18910 -325 18925 -305
rect 18995 -325 19010 -305
rect 19080 -325 19095 -305
rect 19165 -325 19180 -305
rect 19250 -325 19265 -305
rect 19335 -325 19350 -305
rect 19420 -325 19435 -305
rect 19505 -325 19520 -305
rect 19590 -325 19605 -305
rect 19675 -325 19690 -305
rect 19760 -325 19775 -305
rect 19845 -325 19860 -305
rect 19930 -325 19945 -305
rect 20015 -325 20030 -305
rect 20100 -325 20115 -305
rect 20185 -325 20200 -305
rect 20270 -325 20285 -305
rect 20355 -325 20370 -305
rect 20440 -325 20455 -305
rect 20525 -325 20540 -305
rect 20610 -325 20625 -305
rect 20695 -325 20710 -305
rect 20780 -325 20795 -305
rect 20865 -325 20880 -305
rect 20950 -325 20965 -305
rect 21035 -325 21050 -305
rect 21120 -325 21135 -305
rect 21205 -325 21220 -305
rect 21290 -325 21305 -305
rect 21375 -325 21390 -305
rect 21460 -325 21475 -305
rect 21545 -325 21560 -305
rect 21630 -325 21645 -305
rect 21715 -325 21730 -305
rect 21800 -325 21815 -305
rect 21885 -325 21900 -305
rect 21970 -325 21985 -305
rect 22055 -325 22070 -305
rect 22140 -325 22155 -305
rect 22225 -325 22240 -305
rect 22310 -325 22325 -305
rect 22395 -325 22410 -305
rect 22480 -325 22495 -305
rect 22565 -325 22580 -305
rect 22650 -325 22665 -305
rect 22735 -325 22750 -305
rect 22820 -325 22835 -305
rect 22905 -325 22920 -305
rect 22990 -325 23005 -305
rect 23075 -325 23090 -305
rect 23160 -325 23175 -305
rect 23245 -325 23260 -305
rect 23330 -325 23345 -305
rect 23415 -325 23430 -305
rect 23500 -325 23515 -305
rect 23585 -325 23600 -305
rect 23670 -325 23685 -305
rect 23755 -325 23770 -305
rect 23840 -325 23855 -305
rect 23925 -325 23940 -305
rect 24010 -325 24025 -305
rect 24095 -325 24110 -305
rect 24180 -325 24195 -305
rect 24265 -325 24280 -305
rect 24350 -325 24365 -305
rect 24435 -325 24450 -305
rect 24520 -325 24535 -305
rect 24605 -325 24620 -305
rect 24690 -325 24705 -305
rect 24775 -325 24790 -305
rect 24860 -325 24875 -305
rect 24945 -325 24960 -305
rect 25030 -325 25045 -305
rect 25115 -325 25130 -305
rect 25200 -325 25215 -305
rect 25285 -325 25300 -305
rect 25370 -325 25385 -305
rect 25455 -325 25470 -305
rect 25540 -325 25555 -305
rect 25625 -325 25640 -305
rect 25710 -325 25725 -305
rect 25795 -325 25810 -305
rect 25880 -325 25895 -305
rect 25965 -325 25980 -305
rect 26050 -325 26065 -305
rect 26135 -325 26150 -305
rect 26220 -325 26235 -305
rect 26305 -325 26320 -305
rect 26390 -325 26405 -305
rect 26475 -325 26490 -305
rect 26560 -325 26575 -305
rect 26645 -325 26660 -305
rect 26730 -325 26745 -305
rect 26815 -325 26830 -305
rect 26900 -325 26915 -305
rect 26985 -325 27000 -305
rect 27070 -325 27085 -305
rect 27155 -325 27170 -305
rect 27240 -325 27255 -305
rect 27325 -325 27340 -305
rect 27410 -325 27425 -305
rect 27495 -325 27510 -305
rect 27580 -325 27595 -305
rect 27665 -325 27680 -305
rect 27750 -325 27765 -305
rect 27835 -325 27850 -305
rect 27920 -325 27935 -305
rect 28005 -325 28020 -305
rect 28090 -325 28105 -305
rect 28175 -325 28190 -305
rect 28260 -325 28275 -305
rect 28345 -325 28360 -305
rect 28430 -325 28445 -305
rect 28515 -325 28530 -305
rect 28600 -325 28615 -305
rect 28685 -325 28700 -305
rect 28770 -325 28785 -305
rect 28855 -325 28870 -305
rect 28940 -325 28955 -305
rect 29025 -325 29040 -305
rect 29110 -325 29125 -305
rect 29195 -325 29210 -305
rect 29280 -325 29295 -305
rect 29365 -325 29380 -305
rect 29450 -325 29465 -305
rect 29535 -325 29550 -305
rect 29620 -325 29635 -305
rect 29705 -325 29720 -305
rect 29790 -325 29805 -305
rect 29875 -325 29890 -305
rect 29960 -325 29975 -305
rect 30045 -325 30060 -305
rect 30130 -325 30145 -305
rect 30215 -325 30230 -305
rect 30300 -325 30315 -305
rect 30385 -325 30400 -305
rect 30470 -325 30485 -305
rect 30555 -325 30570 -305
rect 30640 -325 30655 -305
rect 30725 -325 30740 -305
rect 30810 -325 30825 -305
rect 30895 -325 30910 -305
rect 30980 -325 30995 -305
rect 31065 -325 31080 -305
rect 31150 -325 31165 -305
rect 31235 -325 31250 -305
rect 31320 -325 31335 -305
rect 31405 -325 31420 -305
rect 31490 -325 31505 -305
rect 31575 -325 31590 -305
rect 31660 -325 31675 -305
rect 31745 -325 31760 -305
rect 31830 -325 31845 -305
rect 31915 -325 31930 -305
rect 32000 -325 32015 -305
rect 32085 -325 32100 -305
rect 32170 -325 32185 -305
rect 32255 -325 32270 -305
rect 32340 -325 32355 -305
rect 32425 -325 32440 -305
rect 32510 -325 32525 -305
rect 32595 -325 32610 -305
rect 32680 -325 32695 -305
rect 32765 -325 32780 -305
rect 32850 -325 32865 -305
rect 32935 -325 32950 -305
rect 33020 -325 33035 -305
rect 33105 -325 33120 -305
rect 33190 -325 33205 -305
rect 33275 -325 33290 -305
rect 33360 -325 33375 -305
rect 33445 -325 33460 -305
rect 33530 -325 33545 -305
rect 33615 -325 33630 -305
rect 33700 -325 33715 -305
rect 33785 -325 33800 -305
rect 33870 -325 33885 -305
rect 33955 -325 33970 -305
rect 34040 -325 34055 -305
rect 34125 -325 34140 -305
rect 34210 -325 34225 -305
rect 34295 -325 34310 -305
rect 34380 -325 34395 -305
rect 34465 -325 34480 -305
rect 34550 -325 34565 -305
rect 34635 -325 34650 -305
rect 34720 -325 34735 -305
rect 34805 -325 34820 -305
rect 34890 -325 34905 -305
rect 34975 -325 34990 -305
rect 35060 -325 35075 -305
rect 35145 -325 35160 -305
rect 35230 -325 35245 -305
rect 35315 -325 35330 -305
rect 35400 -325 35415 -305
rect 35485 -325 35500 -305
rect 35570 -325 35585 -305
rect 35655 -325 35670 -305
rect 35740 -325 35755 -305
rect 35825 -325 35840 -305
rect 35910 -325 35925 -305
rect 35995 -325 36010 -305
rect 36080 -325 36095 -305
rect 36165 -325 36180 -305
rect 36250 -325 36265 -305
rect 36335 -325 36350 -305
rect 36420 -325 36435 -305
rect 36505 -325 36520 -305
rect 36590 -325 36605 -305
rect 36675 -325 36690 -305
rect 36760 -325 36775 -305
rect 36845 -325 36860 -305
rect 36930 -325 36945 -305
rect 37015 -325 37030 -305
rect 37100 -325 37115 -305
rect 37185 -325 37200 -305
rect 37270 -325 37285 -305
rect 37355 -325 37370 -305
rect 37440 -325 37455 -305
rect 37525 -325 37540 -305
rect 37610 -325 37625 -305
rect 37695 -325 37710 -305
rect 37780 -325 37795 -305
rect 37865 -325 37880 -305
rect 37950 -325 37965 -305
rect 38035 -325 38050 -305
rect 38120 -325 38135 -305
rect 38205 -325 38220 -305
rect 38290 -325 38305 -305
rect 38375 -325 38390 -305
rect 38460 -325 38475 -305
rect 38545 -325 38560 -305
rect 38630 -325 38645 -305
rect 38715 -325 38730 -305
rect 38800 -325 38815 -305
rect 38885 -325 38900 -305
rect 38970 -325 38985 -305
rect 39055 -325 39070 -305
rect 39140 -325 39155 -305
rect 39225 -325 39240 -305
rect 39310 -325 39325 -305
rect 39395 -325 39410 -305
rect 39480 -325 39495 -305
rect 39565 -325 39580 -305
rect 39650 -325 39665 -305
rect 39735 -325 39750 -305
rect 39820 -325 39835 -305
rect 39905 -325 39920 -305
rect 39990 -325 40005 -305
rect 40075 -325 40090 -305
rect 40160 -325 40175 -305
rect 40245 -325 40260 -305
rect 40330 -325 40345 -305
rect 40415 -325 40430 -305
rect 40500 -325 40515 -305
rect 40585 -325 40600 -305
rect 40670 -325 40685 -305
rect 40755 -325 40770 -305
rect 40840 -325 40855 -305
rect 40925 -325 40940 -305
rect 41010 -325 41025 -305
rect 41095 -325 41110 -305
rect 41180 -325 41195 -305
rect 41265 -325 41280 -305
rect 41350 -325 41365 -305
rect 41435 -325 41450 -305
rect 41520 -325 41535 -305
rect 41605 -325 41620 -305
rect 41690 -325 41705 -305
rect 41775 -325 41790 -305
rect 41860 -325 41875 -305
rect 41945 -325 41960 -305
rect 42030 -325 42045 -305
rect 42115 -325 42130 -305
rect 42200 -325 42215 -305
rect 42285 -325 42300 -305
rect 42370 -325 42385 -305
rect 42455 -325 42470 -305
rect 42540 -325 42555 -305
rect 42625 -325 42640 -305
rect 42710 -325 42725 -305
rect 42795 -325 42810 -305
rect 42880 -325 42895 -305
rect 42965 -325 42980 -305
rect 43050 -325 43065 -305
rect 43135 -325 43150 -305
rect 43220 -325 43235 -305
rect 43305 -325 43320 -305
rect 43390 -325 43405 -305
rect 43475 -325 43490 -305
rect 43560 -325 43575 -305
rect 125 -490 140 -425
rect 210 -490 225 -425
rect 295 -490 310 -425
rect 380 -490 395 -425
rect 465 -490 480 -425
rect 550 -490 565 -425
rect 635 -490 650 -425
rect 720 -490 735 -425
rect 805 -490 820 -425
rect 890 -490 905 -425
rect 975 -490 990 -425
rect 1060 -490 1075 -425
rect 1145 -490 1160 -425
rect 1230 -490 1245 -425
rect 1315 -490 1330 -425
rect 1400 -490 1415 -425
rect 1485 -490 1500 -425
rect 1570 -490 1585 -425
rect 1655 -490 1670 -425
rect 1740 -490 1755 -425
rect 1825 -490 1840 -425
rect 1910 -490 1925 -425
rect 1995 -490 2010 -425
rect 2080 -490 2095 -425
rect 2165 -490 2180 -425
rect 2250 -490 2265 -425
rect 2335 -490 2350 -425
rect 2420 -490 2435 -425
rect 2505 -490 2520 -425
rect 2590 -490 2605 -425
rect 2675 -490 2690 -425
rect 2760 -490 2775 -425
rect 2845 -490 2860 -425
rect 2930 -490 2945 -425
rect 3015 -490 3030 -425
rect 3100 -490 3115 -425
rect 3185 -490 3200 -425
rect 3270 -490 3285 -425
rect 3355 -490 3370 -425
rect 3440 -490 3455 -425
rect 3525 -490 3540 -425
rect 3610 -490 3625 -425
rect 3695 -490 3710 -425
rect 3780 -490 3795 -425
rect 3865 -490 3880 -425
rect 3950 -490 3965 -425
rect 4035 -490 4050 -425
rect 4120 -490 4135 -425
rect 4205 -490 4220 -425
rect 4290 -490 4305 -425
rect 4375 -490 4390 -425
rect 4460 -490 4475 -425
rect 4545 -490 4560 -425
rect 4630 -490 4645 -425
rect 4715 -490 4730 -425
rect 4800 -490 4815 -425
rect 4885 -490 4900 -425
rect 4970 -490 4985 -425
rect 5055 -490 5070 -425
rect 5140 -490 5155 -425
rect 5225 -490 5240 -425
rect 5310 -490 5325 -425
rect 5395 -490 5410 -425
rect 5480 -490 5495 -425
rect 5565 -490 5580 -425
rect 5650 -490 5665 -425
rect 5735 -490 5750 -425
rect 5820 -490 5835 -425
rect 5905 -490 5920 -425
rect 5990 -490 6005 -425
rect 6075 -490 6090 -425
rect 6160 -490 6175 -425
rect 6245 -490 6260 -425
rect 6330 -490 6345 -425
rect 6415 -490 6430 -425
rect 6500 -490 6515 -425
rect 6585 -490 6600 -425
rect 6670 -490 6685 -425
rect 6755 -490 6770 -425
rect 6840 -490 6855 -425
rect 6925 -490 6940 -425
rect 7010 -490 7025 -425
rect 7095 -490 7110 -425
rect 7180 -490 7195 -425
rect 7265 -490 7280 -425
rect 7350 -490 7365 -425
rect 7435 -490 7450 -425
rect 7520 -490 7535 -425
rect 7605 -490 7620 -425
rect 7690 -490 7705 -425
rect 7775 -490 7790 -425
rect 7860 -490 7875 -425
rect 7945 -490 7960 -425
rect 8030 -490 8045 -425
rect 8115 -490 8130 -425
rect 8200 -490 8215 -425
rect 8285 -490 8300 -425
rect 8370 -490 8385 -425
rect 8455 -490 8470 -425
rect 8540 -490 8555 -425
rect 8625 -490 8640 -425
rect 8710 -490 8725 -425
rect 8795 -490 8810 -425
rect 8880 -490 8895 -425
rect 8965 -490 8980 -425
rect 9050 -490 9065 -425
rect 9135 -490 9150 -425
rect 9220 -490 9235 -425
rect 9305 -490 9320 -425
rect 9390 -490 9405 -425
rect 9475 -490 9490 -425
rect 9560 -490 9575 -425
rect 9645 -490 9660 -425
rect 9730 -490 9745 -425
rect 9815 -490 9830 -425
rect 9900 -490 9915 -425
rect 9985 -490 10000 -425
rect 10070 -490 10085 -425
rect 10155 -490 10170 -425
rect 10240 -490 10255 -425
rect 10325 -490 10340 -425
rect 10410 -490 10425 -425
rect 10495 -490 10510 -425
rect 10580 -490 10595 -425
rect 10665 -490 10680 -425
rect 10750 -490 10765 -425
rect 10835 -490 10850 -425
rect 10920 -490 10935 -425
rect 11005 -490 11020 -425
rect 11090 -490 11105 -425
rect 11175 -490 11190 -425
rect 11260 -490 11275 -425
rect 11345 -490 11360 -425
rect 11430 -490 11445 -425
rect 11515 -490 11530 -425
rect 11600 -490 11615 -425
rect 11685 -490 11700 -425
rect 11770 -490 11785 -425
rect 11855 -490 11870 -425
rect 11940 -490 11955 -425
rect 12025 -490 12040 -425
rect 12110 -490 12125 -425
rect 12195 -490 12210 -425
rect 12280 -490 12295 -425
rect 12365 -490 12380 -425
rect 12450 -490 12465 -425
rect 12535 -490 12550 -425
rect 12620 -490 12635 -425
rect 12705 -490 12720 -425
rect 12790 -490 12805 -425
rect 12875 -490 12890 -425
rect 12960 -490 12975 -425
rect 13045 -490 13060 -425
rect 13130 -490 13145 -425
rect 13215 -490 13230 -425
rect 13300 -490 13315 -425
rect 13385 -490 13400 -425
rect 13470 -490 13485 -425
rect 13555 -490 13570 -425
rect 13640 -490 13655 -425
rect 13725 -490 13740 -425
rect 13810 -490 13825 -425
rect 13895 -490 13910 -425
rect 13980 -490 13995 -425
rect 14065 -490 14080 -425
rect 14150 -490 14165 -425
rect 14235 -490 14250 -425
rect 14320 -490 14335 -425
rect 14405 -490 14420 -425
rect 14490 -490 14505 -425
rect 14575 -490 14590 -425
rect 14660 -490 14675 -425
rect 14745 -490 14760 -425
rect 14830 -490 14845 -425
rect 14915 -490 14930 -425
rect 15000 -490 15015 -425
rect 15085 -490 15100 -425
rect 15170 -490 15185 -425
rect 15255 -490 15270 -425
rect 15340 -490 15355 -425
rect 15425 -490 15440 -425
rect 15510 -490 15525 -425
rect 15595 -490 15610 -425
rect 15680 -490 15695 -425
rect 15765 -490 15780 -425
rect 15850 -490 15865 -425
rect 15935 -490 15950 -425
rect 16020 -490 16035 -425
rect 16105 -490 16120 -425
rect 16190 -490 16205 -425
rect 16275 -490 16290 -425
rect 16360 -490 16375 -425
rect 16445 -490 16460 -425
rect 16530 -490 16545 -425
rect 16615 -490 16630 -425
rect 16700 -490 16715 -425
rect 16785 -490 16800 -425
rect 16870 -490 16885 -425
rect 16955 -490 16970 -425
rect 17040 -490 17055 -425
rect 17125 -490 17140 -425
rect 17210 -490 17225 -425
rect 17295 -490 17310 -425
rect 17380 -490 17395 -425
rect 17465 -490 17480 -425
rect 17550 -490 17565 -425
rect 17635 -490 17650 -425
rect 17720 -490 17735 -425
rect 17805 -490 17820 -425
rect 17890 -490 17905 -425
rect 17975 -490 17990 -425
rect 18060 -490 18075 -425
rect 18145 -490 18160 -425
rect 18230 -490 18245 -425
rect 18315 -490 18330 -425
rect 18400 -490 18415 -425
rect 18485 -490 18500 -425
rect 18570 -490 18585 -425
rect 18655 -490 18670 -425
rect 18740 -490 18755 -425
rect 18825 -490 18840 -425
rect 18910 -490 18925 -425
rect 18995 -490 19010 -425
rect 19080 -490 19095 -425
rect 19165 -490 19180 -425
rect 19250 -490 19265 -425
rect 19335 -490 19350 -425
rect 19420 -490 19435 -425
rect 19505 -490 19520 -425
rect 19590 -490 19605 -425
rect 19675 -490 19690 -425
rect 19760 -490 19775 -425
rect 19845 -490 19860 -425
rect 19930 -490 19945 -425
rect 20015 -490 20030 -425
rect 20100 -490 20115 -425
rect 20185 -490 20200 -425
rect 20270 -490 20285 -425
rect 20355 -490 20370 -425
rect 20440 -490 20455 -425
rect 20525 -490 20540 -425
rect 20610 -490 20625 -425
rect 20695 -490 20710 -425
rect 20780 -490 20795 -425
rect 20865 -490 20880 -425
rect 20950 -490 20965 -425
rect 21035 -490 21050 -425
rect 21120 -490 21135 -425
rect 21205 -490 21220 -425
rect 21290 -490 21305 -425
rect 21375 -490 21390 -425
rect 21460 -490 21475 -425
rect 21545 -490 21560 -425
rect 21630 -490 21645 -425
rect 21715 -490 21730 -425
rect 21800 -490 21815 -425
rect 21885 -490 21900 -425
rect 21970 -490 21985 -425
rect 22055 -490 22070 -425
rect 22140 -490 22155 -425
rect 22225 -490 22240 -425
rect 22310 -490 22325 -425
rect 22395 -490 22410 -425
rect 22480 -490 22495 -425
rect 22565 -490 22580 -425
rect 22650 -490 22665 -425
rect 22735 -490 22750 -425
rect 22820 -490 22835 -425
rect 22905 -490 22920 -425
rect 22990 -490 23005 -425
rect 23075 -490 23090 -425
rect 23160 -490 23175 -425
rect 23245 -490 23260 -425
rect 23330 -490 23345 -425
rect 23415 -490 23430 -425
rect 23500 -490 23515 -425
rect 23585 -490 23600 -425
rect 23670 -490 23685 -425
rect 23755 -490 23770 -425
rect 23840 -490 23855 -425
rect 23925 -490 23940 -425
rect 24010 -490 24025 -425
rect 24095 -490 24110 -425
rect 24180 -490 24195 -425
rect 24265 -490 24280 -425
rect 24350 -490 24365 -425
rect 24435 -490 24450 -425
rect 24520 -490 24535 -425
rect 24605 -490 24620 -425
rect 24690 -490 24705 -425
rect 24775 -490 24790 -425
rect 24860 -490 24875 -425
rect 24945 -490 24960 -425
rect 25030 -490 25045 -425
rect 25115 -490 25130 -425
rect 25200 -490 25215 -425
rect 25285 -490 25300 -425
rect 25370 -490 25385 -425
rect 25455 -490 25470 -425
rect 25540 -490 25555 -425
rect 25625 -490 25640 -425
rect 25710 -490 25725 -425
rect 25795 -490 25810 -425
rect 25880 -490 25895 -425
rect 25965 -490 25980 -425
rect 26050 -490 26065 -425
rect 26135 -490 26150 -425
rect 26220 -490 26235 -425
rect 26305 -490 26320 -425
rect 26390 -490 26405 -425
rect 26475 -490 26490 -425
rect 26560 -490 26575 -425
rect 26645 -490 26660 -425
rect 26730 -490 26745 -425
rect 26815 -490 26830 -425
rect 26900 -490 26915 -425
rect 26985 -490 27000 -425
rect 27070 -490 27085 -425
rect 27155 -490 27170 -425
rect 27240 -490 27255 -425
rect 27325 -490 27340 -425
rect 27410 -490 27425 -425
rect 27495 -490 27510 -425
rect 27580 -490 27595 -425
rect 27665 -490 27680 -425
rect 27750 -490 27765 -425
rect 27835 -490 27850 -425
rect 27920 -490 27935 -425
rect 28005 -490 28020 -425
rect 28090 -490 28105 -425
rect 28175 -490 28190 -425
rect 28260 -490 28275 -425
rect 28345 -490 28360 -425
rect 28430 -490 28445 -425
rect 28515 -490 28530 -425
rect 28600 -490 28615 -425
rect 28685 -490 28700 -425
rect 28770 -490 28785 -425
rect 28855 -490 28870 -425
rect 28940 -490 28955 -425
rect 29025 -490 29040 -425
rect 29110 -490 29125 -425
rect 29195 -490 29210 -425
rect 29280 -490 29295 -425
rect 29365 -490 29380 -425
rect 29450 -490 29465 -425
rect 29535 -490 29550 -425
rect 29620 -490 29635 -425
rect 29705 -490 29720 -425
rect 29790 -490 29805 -425
rect 29875 -490 29890 -425
rect 29960 -490 29975 -425
rect 30045 -490 30060 -425
rect 30130 -490 30145 -425
rect 30215 -490 30230 -425
rect 30300 -490 30315 -425
rect 30385 -490 30400 -425
rect 30470 -490 30485 -425
rect 30555 -490 30570 -425
rect 30640 -490 30655 -425
rect 30725 -490 30740 -425
rect 30810 -490 30825 -425
rect 30895 -490 30910 -425
rect 30980 -490 30995 -425
rect 31065 -490 31080 -425
rect 31150 -490 31165 -425
rect 31235 -490 31250 -425
rect 31320 -490 31335 -425
rect 31405 -490 31420 -425
rect 31490 -490 31505 -425
rect 31575 -490 31590 -425
rect 31660 -490 31675 -425
rect 31745 -490 31760 -425
rect 31830 -490 31845 -425
rect 31915 -490 31930 -425
rect 32000 -490 32015 -425
rect 32085 -490 32100 -425
rect 32170 -490 32185 -425
rect 32255 -490 32270 -425
rect 32340 -490 32355 -425
rect 32425 -490 32440 -425
rect 32510 -490 32525 -425
rect 32595 -490 32610 -425
rect 32680 -490 32695 -425
rect 32765 -490 32780 -425
rect 32850 -490 32865 -425
rect 32935 -490 32950 -425
rect 33020 -490 33035 -425
rect 33105 -490 33120 -425
rect 33190 -490 33205 -425
rect 33275 -490 33290 -425
rect 33360 -490 33375 -425
rect 33445 -490 33460 -425
rect 33530 -490 33545 -425
rect 33615 -490 33630 -425
rect 33700 -490 33715 -425
rect 33785 -490 33800 -425
rect 33870 -490 33885 -425
rect 33955 -490 33970 -425
rect 34040 -490 34055 -425
rect 34125 -490 34140 -425
rect 34210 -490 34225 -425
rect 34295 -490 34310 -425
rect 34380 -490 34395 -425
rect 34465 -490 34480 -425
rect 34550 -490 34565 -425
rect 34635 -490 34650 -425
rect 34720 -490 34735 -425
rect 34805 -490 34820 -425
rect 34890 -490 34905 -425
rect 34975 -490 34990 -425
rect 35060 -490 35075 -425
rect 35145 -490 35160 -425
rect 35230 -490 35245 -425
rect 35315 -490 35330 -425
rect 35400 -490 35415 -425
rect 35485 -490 35500 -425
rect 35570 -490 35585 -425
rect 35655 -490 35670 -425
rect 35740 -490 35755 -425
rect 35825 -490 35840 -425
rect 35910 -490 35925 -425
rect 35995 -490 36010 -425
rect 36080 -490 36095 -425
rect 36165 -490 36180 -425
rect 36250 -490 36265 -425
rect 36335 -490 36350 -425
rect 36420 -490 36435 -425
rect 36505 -490 36520 -425
rect 36590 -490 36605 -425
rect 36675 -490 36690 -425
rect 36760 -490 36775 -425
rect 36845 -490 36860 -425
rect 36930 -490 36945 -425
rect 37015 -490 37030 -425
rect 37100 -490 37115 -425
rect 37185 -490 37200 -425
rect 37270 -490 37285 -425
rect 37355 -490 37370 -425
rect 37440 -490 37455 -425
rect 37525 -490 37540 -425
rect 37610 -490 37625 -425
rect 37695 -490 37710 -425
rect 37780 -490 37795 -425
rect 37865 -490 37880 -425
rect 37950 -490 37965 -425
rect 38035 -490 38050 -425
rect 38120 -490 38135 -425
rect 38205 -490 38220 -425
rect 38290 -490 38305 -425
rect 38375 -490 38390 -425
rect 38460 -490 38475 -425
rect 38545 -490 38560 -425
rect 38630 -490 38645 -425
rect 38715 -490 38730 -425
rect 38800 -490 38815 -425
rect 38885 -490 38900 -425
rect 38970 -490 38985 -425
rect 39055 -490 39070 -425
rect 39140 -490 39155 -425
rect 39225 -490 39240 -425
rect 39310 -490 39325 -425
rect 39395 -490 39410 -425
rect 39480 -490 39495 -425
rect 39565 -490 39580 -425
rect 39650 -490 39665 -425
rect 39735 -490 39750 -425
rect 39820 -490 39835 -425
rect 39905 -490 39920 -425
rect 39990 -490 40005 -425
rect 40075 -490 40090 -425
rect 40160 -490 40175 -425
rect 40245 -490 40260 -425
rect 40330 -490 40345 -425
rect 40415 -490 40430 -425
rect 40500 -490 40515 -425
rect 40585 -490 40600 -425
rect 40670 -490 40685 -425
rect 40755 -490 40770 -425
rect 40840 -490 40855 -425
rect 40925 -490 40940 -425
rect 41010 -490 41025 -425
rect 41095 -490 41110 -425
rect 41180 -490 41195 -425
rect 41265 -490 41280 -425
rect 41350 -490 41365 -425
rect 41435 -490 41450 -425
rect 41520 -490 41535 -425
rect 41605 -490 41620 -425
rect 41690 -490 41705 -425
rect 41775 -490 41790 -425
rect 41860 -490 41875 -425
rect 41945 -490 41960 -425
rect 42030 -490 42045 -425
rect 42115 -490 42130 -425
rect 42200 -490 42215 -425
rect 42285 -490 42300 -425
rect 42370 -490 42385 -425
rect 42455 -490 42470 -425
rect 42540 -490 42555 -425
rect 42625 -490 42640 -425
rect 42710 -490 42725 -425
rect 42795 -490 42810 -425
rect 42880 -490 42895 -425
rect 42965 -490 42980 -425
rect 43050 -490 43065 -425
rect 43135 -490 43150 -425
rect 43220 -490 43235 -425
rect 43305 -490 43320 -425
rect 43390 -490 43405 -425
rect 43475 -490 43490 -425
rect 43560 -490 43575 -425
rect 125 -705 140 -690
rect 210 -705 225 -690
rect 295 -705 310 -690
rect 380 -705 395 -690
rect 465 -705 480 -690
rect 550 -705 565 -690
rect 635 -705 650 -690
rect 720 -705 735 -690
rect 805 -705 820 -690
rect 890 -705 905 -690
rect 975 -705 990 -690
rect 1060 -705 1075 -690
rect 1145 -705 1160 -690
rect 1230 -705 1245 -690
rect 1315 -705 1330 -690
rect 1400 -705 1415 -690
rect 1485 -705 1500 -690
rect 1570 -705 1585 -690
rect 1655 -705 1670 -690
rect 1740 -705 1755 -690
rect 1825 -705 1840 -690
rect 1910 -705 1925 -690
rect 1995 -705 2010 -690
rect 2080 -705 2095 -690
rect 2165 -705 2180 -690
rect 2250 -705 2265 -690
rect 2335 -705 2350 -690
rect 2420 -705 2435 -690
rect 2505 -705 2520 -690
rect 2590 -705 2605 -690
rect 2675 -705 2690 -690
rect 2760 -705 2775 -690
rect 2845 -705 2860 -690
rect 2930 -705 2945 -690
rect 3015 -705 3030 -690
rect 3100 -705 3115 -690
rect 3185 -705 3200 -690
rect 3270 -705 3285 -690
rect 3355 -705 3370 -690
rect 3440 -705 3455 -690
rect 3525 -705 3540 -690
rect 3610 -705 3625 -690
rect 3695 -705 3710 -690
rect 3780 -705 3795 -690
rect 3865 -705 3880 -690
rect 3950 -705 3965 -690
rect 4035 -705 4050 -690
rect 4120 -705 4135 -690
rect 4205 -705 4220 -690
rect 4290 -705 4305 -690
rect 4375 -705 4390 -690
rect 4460 -705 4475 -690
rect 4545 -705 4560 -690
rect 4630 -705 4645 -690
rect 4715 -705 4730 -690
rect 4800 -705 4815 -690
rect 4885 -705 4900 -690
rect 4970 -705 4985 -690
rect 5055 -705 5070 -690
rect 5140 -705 5155 -690
rect 5225 -705 5240 -690
rect 5310 -705 5325 -690
rect 5395 -705 5410 -690
rect 5480 -705 5495 -690
rect 5565 -705 5580 -690
rect 5650 -705 5665 -690
rect 5735 -705 5750 -690
rect 5820 -705 5835 -690
rect 5905 -705 5920 -690
rect 5990 -705 6005 -690
rect 6075 -705 6090 -690
rect 6160 -705 6175 -690
rect 6245 -705 6260 -690
rect 6330 -705 6345 -690
rect 6415 -705 6430 -690
rect 6500 -705 6515 -690
rect 6585 -705 6600 -690
rect 6670 -705 6685 -690
rect 6755 -705 6770 -690
rect 6840 -705 6855 -690
rect 6925 -705 6940 -690
rect 7010 -705 7025 -690
rect 7095 -705 7110 -690
rect 7180 -705 7195 -690
rect 7265 -705 7280 -690
rect 7350 -705 7365 -690
rect 7435 -705 7450 -690
rect 7520 -705 7535 -690
rect 7605 -705 7620 -690
rect 7690 -705 7705 -690
rect 7775 -705 7790 -690
rect 7860 -705 7875 -690
rect 7945 -705 7960 -690
rect 8030 -705 8045 -690
rect 8115 -705 8130 -690
rect 8200 -705 8215 -690
rect 8285 -705 8300 -690
rect 8370 -705 8385 -690
rect 8455 -705 8470 -690
rect 8540 -705 8555 -690
rect 8625 -705 8640 -690
rect 8710 -705 8725 -690
rect 8795 -705 8810 -690
rect 8880 -705 8895 -690
rect 8965 -705 8980 -690
rect 9050 -705 9065 -690
rect 9135 -705 9150 -690
rect 9220 -705 9235 -690
rect 9305 -705 9320 -690
rect 9390 -705 9405 -690
rect 9475 -705 9490 -690
rect 9560 -705 9575 -690
rect 9645 -705 9660 -690
rect 9730 -705 9745 -690
rect 9815 -705 9830 -690
rect 9900 -705 9915 -690
rect 9985 -705 10000 -690
rect 10070 -705 10085 -690
rect 10155 -705 10170 -690
rect 10240 -705 10255 -690
rect 10325 -705 10340 -690
rect 10410 -705 10425 -690
rect 10495 -705 10510 -690
rect 10580 -705 10595 -690
rect 10665 -705 10680 -690
rect 10750 -705 10765 -690
rect 10835 -705 10850 -690
rect 10920 -705 10935 -690
rect 11005 -705 11020 -690
rect 11090 -705 11105 -690
rect 11175 -705 11190 -690
rect 11260 -705 11275 -690
rect 11345 -705 11360 -690
rect 11430 -705 11445 -690
rect 11515 -705 11530 -690
rect 11600 -705 11615 -690
rect 11685 -705 11700 -690
rect 11770 -705 11785 -690
rect 11855 -705 11870 -690
rect 11940 -705 11955 -690
rect 12025 -705 12040 -690
rect 12110 -705 12125 -690
rect 12195 -705 12210 -690
rect 12280 -705 12295 -690
rect 12365 -705 12380 -690
rect 12450 -705 12465 -690
rect 12535 -705 12550 -690
rect 12620 -705 12635 -690
rect 12705 -705 12720 -690
rect 12790 -705 12805 -690
rect 12875 -705 12890 -690
rect 12960 -705 12975 -690
rect 13045 -705 13060 -690
rect 13130 -705 13145 -690
rect 13215 -705 13230 -690
rect 13300 -705 13315 -690
rect 13385 -705 13400 -690
rect 13470 -705 13485 -690
rect 13555 -705 13570 -690
rect 13640 -705 13655 -690
rect 13725 -705 13740 -690
rect 13810 -705 13825 -690
rect 13895 -705 13910 -690
rect 13980 -705 13995 -690
rect 14065 -705 14080 -690
rect 14150 -705 14165 -690
rect 14235 -705 14250 -690
rect 14320 -705 14335 -690
rect 14405 -705 14420 -690
rect 14490 -705 14505 -690
rect 14575 -705 14590 -690
rect 14660 -705 14675 -690
rect 14745 -705 14760 -690
rect 14830 -705 14845 -690
rect 14915 -705 14930 -690
rect 15000 -705 15015 -690
rect 15085 -705 15100 -690
rect 15170 -705 15185 -690
rect 15255 -705 15270 -690
rect 15340 -705 15355 -690
rect 15425 -705 15440 -690
rect 15510 -705 15525 -690
rect 15595 -705 15610 -690
rect 15680 -705 15695 -690
rect 15765 -705 15780 -690
rect 15850 -705 15865 -690
rect 15935 -705 15950 -690
rect 16020 -705 16035 -690
rect 16105 -705 16120 -690
rect 16190 -705 16205 -690
rect 16275 -705 16290 -690
rect 16360 -705 16375 -690
rect 16445 -705 16460 -690
rect 16530 -705 16545 -690
rect 16615 -705 16630 -690
rect 16700 -705 16715 -690
rect 16785 -705 16800 -690
rect 16870 -705 16885 -690
rect 16955 -705 16970 -690
rect 17040 -705 17055 -690
rect 17125 -705 17140 -690
rect 17210 -705 17225 -690
rect 17295 -705 17310 -690
rect 17380 -705 17395 -690
rect 17465 -705 17480 -690
rect 17550 -705 17565 -690
rect 17635 -705 17650 -690
rect 17720 -705 17735 -690
rect 17805 -705 17820 -690
rect 17890 -705 17905 -690
rect 17975 -705 17990 -690
rect 18060 -705 18075 -690
rect 18145 -705 18160 -690
rect 18230 -705 18245 -690
rect 18315 -705 18330 -690
rect 18400 -705 18415 -690
rect 18485 -705 18500 -690
rect 18570 -705 18585 -690
rect 18655 -705 18670 -690
rect 18740 -705 18755 -690
rect 18825 -705 18840 -690
rect 18910 -705 18925 -690
rect 18995 -705 19010 -690
rect 19080 -705 19095 -690
rect 19165 -705 19180 -690
rect 19250 -705 19265 -690
rect 19335 -705 19350 -690
rect 19420 -705 19435 -690
rect 19505 -705 19520 -690
rect 19590 -705 19605 -690
rect 19675 -705 19690 -690
rect 19760 -705 19775 -690
rect 19845 -705 19860 -690
rect 19930 -705 19945 -690
rect 20015 -705 20030 -690
rect 20100 -705 20115 -690
rect 20185 -705 20200 -690
rect 20270 -705 20285 -690
rect 20355 -705 20370 -690
rect 20440 -705 20455 -690
rect 20525 -705 20540 -690
rect 20610 -705 20625 -690
rect 20695 -705 20710 -690
rect 20780 -705 20795 -690
rect 20865 -705 20880 -690
rect 20950 -705 20965 -690
rect 21035 -705 21050 -690
rect 21120 -705 21135 -690
rect 21205 -705 21220 -690
rect 21290 -705 21305 -690
rect 21375 -705 21390 -690
rect 21460 -705 21475 -690
rect 21545 -705 21560 -690
rect 21630 -705 21645 -690
rect 21715 -705 21730 -690
rect 21800 -705 21815 -690
rect 21885 -705 21900 -690
rect 21970 -705 21985 -690
rect 22055 -705 22070 -690
rect 22140 -705 22155 -690
rect 22225 -705 22240 -690
rect 22310 -705 22325 -690
rect 22395 -705 22410 -690
rect 22480 -705 22495 -690
rect 22565 -705 22580 -690
rect 22650 -705 22665 -690
rect 22735 -705 22750 -690
rect 22820 -705 22835 -690
rect 22905 -705 22920 -690
rect 22990 -705 23005 -690
rect 23075 -705 23090 -690
rect 23160 -705 23175 -690
rect 23245 -705 23260 -690
rect 23330 -705 23345 -690
rect 23415 -705 23430 -690
rect 23500 -705 23515 -690
rect 23585 -705 23600 -690
rect 23670 -705 23685 -690
rect 23755 -705 23770 -690
rect 23840 -705 23855 -690
rect 23925 -705 23940 -690
rect 24010 -705 24025 -690
rect 24095 -705 24110 -690
rect 24180 -705 24195 -690
rect 24265 -705 24280 -690
rect 24350 -705 24365 -690
rect 24435 -705 24450 -690
rect 24520 -705 24535 -690
rect 24605 -705 24620 -690
rect 24690 -705 24705 -690
rect 24775 -705 24790 -690
rect 24860 -705 24875 -690
rect 24945 -705 24960 -690
rect 25030 -705 25045 -690
rect 25115 -705 25130 -690
rect 25200 -705 25215 -690
rect 25285 -705 25300 -690
rect 25370 -705 25385 -690
rect 25455 -705 25470 -690
rect 25540 -705 25555 -690
rect 25625 -705 25640 -690
rect 25710 -705 25725 -690
rect 25795 -705 25810 -690
rect 25880 -705 25895 -690
rect 25965 -705 25980 -690
rect 26050 -705 26065 -690
rect 26135 -705 26150 -690
rect 26220 -705 26235 -690
rect 26305 -705 26320 -690
rect 26390 -705 26405 -690
rect 26475 -705 26490 -690
rect 26560 -705 26575 -690
rect 26645 -705 26660 -690
rect 26730 -705 26745 -690
rect 26815 -705 26830 -690
rect 26900 -705 26915 -690
rect 26985 -705 27000 -690
rect 27070 -705 27085 -690
rect 27155 -705 27170 -690
rect 27240 -705 27255 -690
rect 27325 -705 27340 -690
rect 27410 -705 27425 -690
rect 27495 -705 27510 -690
rect 27580 -705 27595 -690
rect 27665 -705 27680 -690
rect 27750 -705 27765 -690
rect 27835 -705 27850 -690
rect 27920 -705 27935 -690
rect 28005 -705 28020 -690
rect 28090 -705 28105 -690
rect 28175 -705 28190 -690
rect 28260 -705 28275 -690
rect 28345 -705 28360 -690
rect 28430 -705 28445 -690
rect 28515 -705 28530 -690
rect 28600 -705 28615 -690
rect 28685 -705 28700 -690
rect 28770 -705 28785 -690
rect 28855 -705 28870 -690
rect 28940 -705 28955 -690
rect 29025 -705 29040 -690
rect 29110 -705 29125 -690
rect 29195 -705 29210 -690
rect 29280 -705 29295 -690
rect 29365 -705 29380 -690
rect 29450 -705 29465 -690
rect 29535 -705 29550 -690
rect 29620 -705 29635 -690
rect 29705 -705 29720 -690
rect 29790 -705 29805 -690
rect 29875 -705 29890 -690
rect 29960 -705 29975 -690
rect 30045 -705 30060 -690
rect 30130 -705 30145 -690
rect 30215 -705 30230 -690
rect 30300 -705 30315 -690
rect 30385 -705 30400 -690
rect 30470 -705 30485 -690
rect 30555 -705 30570 -690
rect 30640 -705 30655 -690
rect 30725 -705 30740 -690
rect 30810 -705 30825 -690
rect 30895 -705 30910 -690
rect 30980 -705 30995 -690
rect 31065 -705 31080 -690
rect 31150 -705 31165 -690
rect 31235 -705 31250 -690
rect 31320 -705 31335 -690
rect 31405 -705 31420 -690
rect 31490 -705 31505 -690
rect 31575 -705 31590 -690
rect 31660 -705 31675 -690
rect 31745 -705 31760 -690
rect 31830 -705 31845 -690
rect 31915 -705 31930 -690
rect 32000 -705 32015 -690
rect 32085 -705 32100 -690
rect 32170 -705 32185 -690
rect 32255 -705 32270 -690
rect 32340 -705 32355 -690
rect 32425 -705 32440 -690
rect 32510 -705 32525 -690
rect 32595 -705 32610 -690
rect 32680 -705 32695 -690
rect 32765 -705 32780 -690
rect 32850 -705 32865 -690
rect 32935 -705 32950 -690
rect 33020 -705 33035 -690
rect 33105 -705 33120 -690
rect 33190 -705 33205 -690
rect 33275 -705 33290 -690
rect 33360 -705 33375 -690
rect 33445 -705 33460 -690
rect 33530 -705 33545 -690
rect 33615 -705 33630 -690
rect 33700 -705 33715 -690
rect 33785 -705 33800 -690
rect 33870 -705 33885 -690
rect 33955 -705 33970 -690
rect 34040 -705 34055 -690
rect 34125 -705 34140 -690
rect 34210 -705 34225 -690
rect 34295 -705 34310 -690
rect 34380 -705 34395 -690
rect 34465 -705 34480 -690
rect 34550 -705 34565 -690
rect 34635 -705 34650 -690
rect 34720 -705 34735 -690
rect 34805 -705 34820 -690
rect 34890 -705 34905 -690
rect 34975 -705 34990 -690
rect 35060 -705 35075 -690
rect 35145 -705 35160 -690
rect 35230 -705 35245 -690
rect 35315 -705 35330 -690
rect 35400 -705 35415 -690
rect 35485 -705 35500 -690
rect 35570 -705 35585 -690
rect 35655 -705 35670 -690
rect 35740 -705 35755 -690
rect 35825 -705 35840 -690
rect 35910 -705 35925 -690
rect 35995 -705 36010 -690
rect 36080 -705 36095 -690
rect 36165 -705 36180 -690
rect 36250 -705 36265 -690
rect 36335 -705 36350 -690
rect 36420 -705 36435 -690
rect 36505 -705 36520 -690
rect 36590 -705 36605 -690
rect 36675 -705 36690 -690
rect 36760 -705 36775 -690
rect 36845 -705 36860 -690
rect 36930 -705 36945 -690
rect 37015 -705 37030 -690
rect 37100 -705 37115 -690
rect 37185 -705 37200 -690
rect 37270 -705 37285 -690
rect 37355 -705 37370 -690
rect 37440 -705 37455 -690
rect 37525 -705 37540 -690
rect 37610 -705 37625 -690
rect 37695 -705 37710 -690
rect 37780 -705 37795 -690
rect 37865 -705 37880 -690
rect 37950 -705 37965 -690
rect 38035 -705 38050 -690
rect 38120 -705 38135 -690
rect 38205 -705 38220 -690
rect 38290 -705 38305 -690
rect 38375 -705 38390 -690
rect 38460 -705 38475 -690
rect 38545 -705 38560 -690
rect 38630 -705 38645 -690
rect 38715 -705 38730 -690
rect 38800 -705 38815 -690
rect 38885 -705 38900 -690
rect 38970 -705 38985 -690
rect 39055 -705 39070 -690
rect 39140 -705 39155 -690
rect 39225 -705 39240 -690
rect 39310 -705 39325 -690
rect 39395 -705 39410 -690
rect 39480 -705 39495 -690
rect 39565 -705 39580 -690
rect 39650 -705 39665 -690
rect 39735 -705 39750 -690
rect 39820 -705 39835 -690
rect 39905 -705 39920 -690
rect 39990 -705 40005 -690
rect 40075 -705 40090 -690
rect 40160 -705 40175 -690
rect 40245 -705 40260 -690
rect 40330 -705 40345 -690
rect 40415 -705 40430 -690
rect 40500 -705 40515 -690
rect 40585 -705 40600 -690
rect 40670 -705 40685 -690
rect 40755 -705 40770 -690
rect 40840 -705 40855 -690
rect 40925 -705 40940 -690
rect 41010 -705 41025 -690
rect 41095 -705 41110 -690
rect 41180 -705 41195 -690
rect 41265 -705 41280 -690
rect 41350 -705 41365 -690
rect 41435 -705 41450 -690
rect 41520 -705 41535 -690
rect 41605 -705 41620 -690
rect 41690 -705 41705 -690
rect 41775 -705 41790 -690
rect 41860 -705 41875 -690
rect 41945 -705 41960 -690
rect 42030 -705 42045 -690
rect 42115 -705 42130 -690
rect 42200 -705 42215 -690
rect 42285 -705 42300 -690
rect 42370 -705 42385 -690
rect 42455 -705 42470 -690
rect 42540 -705 42555 -690
rect 42625 -705 42640 -690
rect 42710 -705 42725 -690
rect 42795 -705 42810 -690
rect 42880 -705 42895 -690
rect 42965 -705 42980 -690
rect 43050 -705 43065 -690
rect 43135 -705 43150 -690
rect 43220 -705 43235 -690
rect 43305 -705 43320 -690
rect 43390 -705 43405 -690
rect 43475 -705 43490 -690
rect 43560 -705 43575 -690
<< polycont >>
rect 35 15 65 55
rect 265 -60 300 -30
rect 350 -60 385 -30
rect 435 -60 470 -30
rect 520 -60 555 -30
rect 800 -60 835 -30
rect 885 -60 920 -30
rect 970 -60 1005 -30
rect 1055 -60 1090 -30
rect 1140 -60 1175 -30
rect 1225 -60 1260 -30
rect 1310 -60 1345 -30
rect 1395 -60 1430 -30
rect 1480 -60 1515 -30
rect 1565 -60 1600 -30
rect 1650 -60 1685 -30
rect 1735 -60 1770 -30
rect 1820 -60 1855 -30
rect 1905 -60 1940 -30
rect 1990 -60 2025 -30
rect 2075 -60 2110 -30
rect 2310 -60 2345 -30
rect 2395 -60 2430 -30
rect 2480 -60 2515 -30
rect 2565 -60 2600 -30
rect 2650 -60 2685 -30
rect 2735 -60 2770 -30
rect 2820 -60 2855 -30
rect 2905 -60 2940 -30
rect 2990 -60 3025 -30
rect 3075 -60 3110 -30
rect 3160 -60 3195 -30
rect 3245 -60 3280 -30
rect 3330 -60 3365 -30
rect 3415 -60 3450 -30
rect 3500 -60 3535 -30
rect 3585 -60 3620 -30
rect 3670 -60 3705 -30
rect 3755 -60 3790 -30
rect 3840 -60 3875 -30
rect 3925 -60 3960 -30
rect 4010 -60 4045 -30
rect 4095 -60 4130 -30
rect 4180 -60 4215 -30
rect 4265 -60 4300 -30
rect 4350 -60 4385 -30
rect 4435 -60 4470 -30
rect 4520 -60 4555 -30
rect 4605 -60 4640 -30
rect 4690 -60 4725 -30
rect 4775 -60 4810 -30
rect 4860 -60 4895 -30
rect 4945 -60 4980 -30
rect 5030 -60 5065 -30
rect 5115 -60 5150 -30
rect 5200 -60 5235 -30
rect 5285 -60 5320 -30
rect 5370 -60 5405 -30
rect 5455 -60 5490 -30
rect 5540 -60 5575 -30
rect 5625 -60 5660 -30
rect 5710 -60 5745 -30
rect 5795 -60 5830 -30
rect 5880 -60 5915 -30
rect 5965 -60 6000 -30
rect 6050 -60 6085 -30
rect 6135 -60 6170 -30
rect 6220 -60 6255 -30
rect 6305 -60 6340 -30
rect 6390 -60 6425 -30
rect 6475 -60 6510 -30
rect 6560 -60 6595 -30
rect 6645 -60 6680 -30
rect 6730 -60 6765 -30
rect 6815 -60 6850 -30
rect 6900 -60 6935 -30
rect 6985 -60 7020 -30
rect 7070 -60 7105 -30
rect 7155 -60 7190 -30
rect 7240 -60 7275 -30
rect 7325 -60 7360 -30
rect 7410 -60 7445 -30
rect 7495 -60 7530 -30
rect 7580 -60 7615 -30
rect 7665 -60 7700 -30
rect 7900 -60 7935 -30
rect 7985 -60 8020 -30
rect 8070 -60 8105 -30
rect 8155 -60 8190 -30
rect 8240 -60 8275 -30
rect 8325 -60 8360 -30
rect 8410 -60 8445 -30
rect 8495 -60 8530 -30
rect 8580 -60 8615 -30
rect 8665 -60 8700 -30
rect 8750 -60 8785 -30
rect 8835 -60 8870 -30
rect 8920 -60 8955 -30
rect 9005 -60 9040 -30
rect 9090 -60 9125 -30
rect 9175 -60 9210 -30
rect 9260 -60 9295 -30
rect 9345 -60 9380 -30
rect 9430 -60 9465 -30
rect 9515 -60 9550 -30
rect 9600 -60 9635 -30
rect 9685 -60 9720 -30
rect 9770 -60 9805 -30
rect 9855 -60 9890 -30
rect 9940 -60 9975 -30
rect 10025 -60 10060 -30
rect 10110 -60 10145 -30
rect 10195 -60 10230 -30
rect 10280 -60 10315 -30
rect 10365 -60 10400 -30
rect 10450 -60 10485 -30
rect 10535 -60 10570 -30
rect 10620 -60 10655 -30
rect 10705 -60 10740 -30
rect 10790 -60 10825 -30
rect 10875 -60 10910 -30
rect 10960 -60 10995 -30
rect 11045 -60 11080 -30
rect 11130 -60 11165 -30
rect 11215 -60 11250 -30
rect 11300 -60 11335 -30
rect 11385 -60 11420 -30
rect 11470 -60 11505 -30
rect 11555 -60 11590 -30
rect 11640 -60 11675 -30
rect 11725 -60 11760 -30
rect 11810 -60 11845 -30
rect 11895 -60 11930 -30
rect 11980 -60 12015 -30
rect 12065 -60 12100 -30
rect 12150 -60 12185 -30
rect 12235 -60 12270 -30
rect 12320 -60 12355 -30
rect 12405 -60 12440 -30
rect 12490 -60 12525 -30
rect 12575 -60 12610 -30
rect 12660 -60 12695 -30
rect 12745 -60 12780 -30
rect 12830 -60 12865 -30
rect 12915 -60 12950 -30
rect 13000 -60 13035 -30
rect 13085 -60 13120 -30
rect 13170 -60 13205 -30
rect 13255 -60 13290 -30
rect 13340 -60 13375 -30
rect 13425 -60 13460 -30
rect 13510 -60 13545 -30
rect 13595 -60 13630 -30
rect 13680 -60 13715 -30
rect 13765 -60 13800 -30
rect 13850 -60 13885 -30
rect 13935 -60 13970 -30
rect 14020 -60 14055 -30
rect 14105 -60 14140 -30
rect 14190 -60 14225 -30
rect 14275 -60 14310 -30
rect 14360 -60 14395 -30
rect 14445 -60 14480 -30
rect 14530 -60 14565 -30
rect 14615 -60 14650 -30
rect 14700 -60 14735 -30
rect 14785 -60 14820 -30
rect 14870 -60 14905 -30
rect 14955 -60 14990 -30
rect 15040 -60 15075 -30
rect 15125 -60 15160 -30
rect 15210 -60 15245 -30
rect 15295 -60 15330 -30
rect 15380 -60 15415 -30
rect 15465 -60 15500 -30
rect 15550 -60 15585 -30
rect 15635 -60 15670 -30
rect 15720 -60 15755 -30
rect 15805 -60 15840 -30
rect 15890 -60 15925 -30
rect 15975 -60 16010 -30
rect 16060 -60 16095 -30
rect 16145 -60 16180 -30
rect 16230 -60 16265 -30
rect 16315 -60 16350 -30
rect 16400 -60 16435 -30
rect 16485 -60 16520 -30
rect 16570 -60 16605 -30
rect 16655 -60 16690 -30
rect 16740 -60 16775 -30
rect 16825 -60 16860 -30
rect 16910 -60 16945 -30
rect 16995 -60 17030 -30
rect 17080 -60 17115 -30
rect 17165 -60 17200 -30
rect 17250 -60 17285 -30
rect 17335 -60 17370 -30
rect 17420 -60 17455 -30
rect 17505 -60 17540 -30
rect 17590 -60 17625 -30
rect 17675 -60 17710 -30
rect 17760 -60 17795 -30
rect 17845 -60 17880 -30
rect 17930 -60 17965 -30
rect 18015 -60 18050 -30
rect 18100 -60 18135 -30
rect 18185 -60 18220 -30
rect 18270 -60 18305 -30
rect 18355 -60 18390 -30
rect 18440 -60 18475 -30
rect 18525 -60 18560 -30
rect 18610 -60 18645 -30
rect 18695 -60 18730 -30
rect 18780 -60 18815 -30
rect 18865 -60 18900 -30
rect 18950 -60 18985 -30
rect 19035 -60 19070 -30
rect 19120 -60 19155 -30
rect 19205 -60 19240 -30
rect 19290 -60 19325 -30
rect 19375 -60 19410 -30
rect 19460 -60 19495 -30
rect 19545 -60 19580 -30
rect 19630 -60 19665 -30
rect 19715 -60 19750 -30
rect 19800 -60 19835 -30
rect 19885 -60 19920 -30
rect 19970 -60 20005 -30
rect 20055 -60 20090 -30
rect 20140 -60 20175 -30
rect 20225 -60 20260 -30
rect 20310 -60 20345 -30
rect 20395 -60 20430 -30
rect 20480 -60 20515 -30
rect 20565 -60 20600 -30
rect 20650 -60 20685 -30
rect 20735 -60 20770 -30
rect 20820 -60 20855 -30
rect 20905 -60 20940 -30
rect 20990 -60 21025 -30
rect 21075 -60 21110 -30
rect 21160 -60 21195 -30
rect 21245 -60 21280 -30
rect 21330 -60 21365 -30
rect 21415 -60 21450 -30
rect 21500 -60 21535 -30
rect 21585 -60 21620 -30
rect 21670 -60 21705 -30
rect 21755 -60 21790 -30
rect 21840 -60 21875 -30
rect 21925 -60 21960 -30
rect 22010 -60 22045 -30
rect 22095 -60 22130 -30
rect 22180 -60 22215 -30
rect 22265 -60 22300 -30
rect 22350 -60 22385 -30
rect 22435 -60 22470 -30
rect 22520 -60 22555 -30
rect 22605 -60 22640 -30
rect 22690 -60 22725 -30
rect 22775 -60 22810 -30
rect 22860 -60 22895 -30
rect 22945 -60 22980 -30
rect 23030 -60 23065 -30
rect 23115 -60 23150 -30
rect 23200 -60 23235 -30
rect 23285 -60 23320 -30
rect 23370 -60 23405 -30
rect 23455 -60 23490 -30
rect 23540 -60 23575 -30
rect 23625 -60 23660 -30
rect 23710 -60 23745 -30
rect 23795 -60 23830 -30
rect 23880 -60 23915 -30
rect 23965 -60 24000 -30
rect 24050 -60 24085 -30
rect 24135 -60 24170 -30
rect 24220 -60 24255 -30
rect 24305 -60 24340 -30
rect 24390 -60 24425 -30
rect 24475 -60 24510 -30
rect 24560 -60 24595 -30
rect 24645 -60 24680 -30
rect 24730 -60 24765 -30
rect 24815 -60 24850 -30
rect 24900 -60 24935 -30
rect 24985 -60 25020 -30
rect 25070 -60 25105 -30
rect 25155 -60 25190 -30
rect 25240 -60 25275 -30
rect 25325 -60 25360 -30
rect 25410 -60 25445 -30
rect 25495 -60 25530 -30
rect 25580 -60 25615 -30
rect 25665 -60 25700 -30
rect 25750 -60 25785 -30
rect 25835 -60 25870 -30
rect 25920 -60 25955 -30
rect 26005 -60 26040 -30
rect 26090 -60 26125 -30
rect 26175 -60 26210 -30
rect 26260 -60 26295 -30
rect 26345 -60 26380 -30
rect 26430 -60 26465 -30
rect 26515 -60 26550 -30
rect 26600 -60 26635 -30
rect 26685 -60 26720 -30
rect 26770 -60 26805 -30
rect 26855 -60 26890 -30
rect 26940 -60 26975 -30
rect 27025 -60 27060 -30
rect 27110 -60 27145 -30
rect 27195 -60 27230 -30
rect 27280 -60 27315 -30
rect 27365 -60 27400 -30
rect 27450 -60 27485 -30
rect 27535 -60 27570 -30
rect 27620 -60 27655 -30
rect 27705 -60 27740 -30
rect 27790 -60 27825 -30
rect 27875 -60 27910 -30
rect 27960 -60 27995 -30
rect 28045 -60 28080 -30
rect 28130 -60 28165 -30
rect 28215 -60 28250 -30
rect 28300 -60 28335 -30
rect 28385 -60 28420 -30
rect 28470 -60 28505 -30
rect 28555 -60 28590 -30
rect 28640 -60 28675 -30
rect 28725 -60 28760 -30
rect 28810 -60 28845 -30
rect 28895 -60 28930 -30
rect 28980 -60 29015 -30
rect 29065 -60 29100 -30
rect 29150 -60 29185 -30
rect 29235 -60 29270 -30
rect 29320 -60 29355 -30
rect 29405 -60 29440 -30
rect 29490 -60 29525 -30
rect 29575 -60 29610 -30
rect 115 -295 150 -265
rect 200 -295 235 -265
rect 285 -295 320 -265
rect 370 -295 405 -265
rect 455 -295 490 -265
rect 540 -295 575 -265
rect 625 -295 660 -265
rect 710 -295 745 -265
rect 795 -295 830 -265
rect 880 -295 915 -265
rect 965 -295 1000 -265
rect 1050 -295 1085 -265
rect 1135 -295 1170 -265
rect 1220 -295 1255 -265
rect 1305 -295 1340 -265
rect 1390 -295 1425 -265
rect 1475 -295 1510 -265
rect 1560 -295 1595 -265
rect 1645 -295 1680 -265
rect 1730 -295 1765 -265
rect 1815 -295 1850 -265
rect 1900 -295 1935 -265
rect 1985 -295 2020 -265
rect 2070 -295 2105 -265
rect 2155 -295 2190 -265
rect 2240 -295 2275 -265
rect 2325 -295 2360 -265
rect 2410 -295 2445 -265
rect 2495 -295 2530 -265
rect 2580 -295 2615 -265
rect 2665 -295 2700 -265
rect 2750 -295 2785 -265
rect 2835 -295 2870 -265
rect 2920 -295 2955 -265
rect 3005 -295 3040 -265
rect 3090 -295 3125 -265
rect 3175 -295 3210 -265
rect 3260 -295 3295 -265
rect 3345 -295 3380 -265
rect 3430 -295 3465 -265
rect 3515 -295 3550 -265
rect 3600 -295 3635 -265
rect 3685 -295 3720 -265
rect 3770 -295 3805 -265
rect 3855 -295 3890 -265
rect 3940 -295 3975 -265
rect 4025 -295 4060 -265
rect 4110 -295 4145 -265
rect 4195 -295 4230 -265
rect 4280 -295 4315 -265
rect 4365 -295 4400 -265
rect 4450 -295 4485 -265
rect 4535 -295 4570 -265
rect 4620 -295 4655 -265
rect 4705 -295 4740 -265
rect 4790 -295 4825 -265
rect 4875 -295 4910 -265
rect 4960 -295 4995 -265
rect 5045 -295 5080 -265
rect 5130 -295 5165 -265
rect 5215 -295 5250 -265
rect 5300 -295 5335 -265
rect 5385 -295 5420 -265
rect 5470 -295 5505 -265
rect 5555 -295 5590 -265
rect 5640 -295 5675 -265
rect 5725 -295 5760 -265
rect 5810 -295 5845 -265
rect 5895 -295 5930 -265
rect 5980 -295 6015 -265
rect 6065 -295 6100 -265
rect 6150 -295 6185 -265
rect 6235 -295 6270 -265
rect 6320 -295 6355 -265
rect 6405 -295 6440 -265
rect 6490 -295 6525 -265
rect 6575 -295 6610 -265
rect 6660 -295 6695 -265
rect 6745 -295 6780 -265
rect 6830 -295 6865 -265
rect 6915 -295 6950 -265
rect 7000 -295 7035 -265
rect 7085 -295 7120 -265
rect 7170 -295 7205 -265
rect 7255 -295 7290 -265
rect 7340 -295 7375 -265
rect 7425 -295 7460 -265
rect 7510 -295 7545 -265
rect 7595 -295 7630 -265
rect 7680 -295 7715 -265
rect 7765 -295 7800 -265
rect 7850 -295 7885 -265
rect 7935 -295 7970 -265
rect 8020 -295 8055 -265
rect 8105 -295 8140 -265
rect 8190 -295 8225 -265
rect 8275 -295 8310 -265
rect 8360 -295 8395 -265
rect 8445 -295 8480 -265
rect 8530 -295 8565 -265
rect 8615 -295 8650 -265
rect 8700 -295 8735 -265
rect 8785 -295 8820 -265
rect 8870 -295 8905 -265
rect 8955 -295 8990 -265
rect 9040 -295 9075 -265
rect 9125 -295 9160 -265
rect 9210 -295 9245 -265
rect 9295 -295 9330 -265
rect 9380 -295 9415 -265
rect 9465 -295 9500 -265
rect 9550 -295 9585 -265
rect 9635 -295 9670 -265
rect 9720 -295 9755 -265
rect 9805 -295 9840 -265
rect 9890 -295 9925 -265
rect 9975 -295 10010 -265
rect 10060 -295 10095 -265
rect 10145 -295 10180 -265
rect 10230 -295 10265 -265
rect 10315 -295 10350 -265
rect 10400 -295 10435 -265
rect 10485 -295 10520 -265
rect 10570 -295 10605 -265
rect 10655 -295 10690 -265
rect 10740 -295 10775 -265
rect 10825 -295 10860 -265
rect 10910 -295 10945 -265
rect 10995 -295 11030 -265
rect 11080 -295 11115 -265
rect 11165 -295 11200 -265
rect 11250 -295 11285 -265
rect 11335 -295 11370 -265
rect 11420 -295 11455 -265
rect 11505 -295 11540 -265
rect 11590 -295 11625 -265
rect 11675 -295 11710 -265
rect 11760 -295 11795 -265
rect 11845 -295 11880 -265
rect 11930 -295 11965 -265
rect 12015 -295 12050 -265
rect 12100 -295 12135 -265
rect 12185 -295 12220 -265
rect 12270 -295 12305 -265
rect 12355 -295 12390 -265
rect 12440 -295 12475 -265
rect 12525 -295 12560 -265
rect 12610 -295 12645 -265
rect 12695 -295 12730 -265
rect 12780 -295 12815 -265
rect 12865 -295 12900 -265
rect 12950 -295 12985 -265
rect 13035 -295 13070 -265
rect 13120 -295 13155 -265
rect 13205 -295 13240 -265
rect 13290 -295 13325 -265
rect 13375 -295 13410 -265
rect 13460 -295 13495 -265
rect 13545 -295 13580 -265
rect 13630 -295 13665 -265
rect 13715 -295 13750 -265
rect 13800 -295 13835 -265
rect 13885 -295 13920 -265
rect 13970 -295 14005 -265
rect 14055 -295 14090 -265
rect 14140 -295 14175 -265
rect 14225 -295 14260 -265
rect 14310 -295 14345 -265
rect 14395 -295 14430 -265
rect 14480 -295 14515 -265
rect 14565 -295 14600 -265
rect 14650 -295 14685 -265
rect 14735 -295 14770 -265
rect 14820 -295 14855 -265
rect 14905 -295 14940 -265
rect 14990 -295 15025 -265
rect 15075 -295 15110 -265
rect 15160 -295 15195 -265
rect 15245 -295 15280 -265
rect 15330 -295 15365 -265
rect 15415 -295 15450 -265
rect 15500 -295 15535 -265
rect 15585 -295 15620 -265
rect 15670 -295 15705 -265
rect 15755 -295 15790 -265
rect 15840 -295 15875 -265
rect 15925 -295 15960 -265
rect 16010 -295 16045 -265
rect 16095 -295 16130 -265
rect 16180 -295 16215 -265
rect 16265 -295 16300 -265
rect 16350 -295 16385 -265
rect 16435 -295 16470 -265
rect 16520 -295 16555 -265
rect 16605 -295 16640 -265
rect 16690 -295 16725 -265
rect 16775 -295 16810 -265
rect 16860 -295 16895 -265
rect 16945 -295 16980 -265
rect 17030 -295 17065 -265
rect 17115 -295 17150 -265
rect 17200 -295 17235 -265
rect 17285 -295 17320 -265
rect 17370 -295 17405 -265
rect 17455 -295 17490 -265
rect 17540 -295 17575 -265
rect 17625 -295 17660 -265
rect 17710 -295 17745 -265
rect 17795 -295 17830 -265
rect 17880 -295 17915 -265
rect 17965 -295 18000 -265
rect 18050 -295 18085 -265
rect 18135 -295 18170 -265
rect 18220 -295 18255 -265
rect 18305 -295 18340 -265
rect 18390 -295 18425 -265
rect 18475 -295 18510 -265
rect 18560 -295 18595 -265
rect 18645 -295 18680 -265
rect 18730 -295 18765 -265
rect 18815 -295 18850 -265
rect 18900 -295 18935 -265
rect 18985 -295 19020 -265
rect 19070 -295 19105 -265
rect 19155 -295 19190 -265
rect 19240 -295 19275 -265
rect 19325 -295 19360 -265
rect 19410 -295 19445 -265
rect 19495 -295 19530 -265
rect 19580 -295 19615 -265
rect 19665 -295 19700 -265
rect 19750 -295 19785 -265
rect 19835 -295 19870 -265
rect 19920 -295 19955 -265
rect 20005 -295 20040 -265
rect 20090 -295 20125 -265
rect 20175 -295 20210 -265
rect 20260 -295 20295 -265
rect 20345 -295 20380 -265
rect 20430 -295 20465 -265
rect 20515 -295 20550 -265
rect 20600 -295 20635 -265
rect 20685 -295 20720 -265
rect 20770 -295 20805 -265
rect 20855 -295 20890 -265
rect 20940 -295 20975 -265
rect 21025 -295 21060 -265
rect 21110 -295 21145 -265
rect 21195 -295 21230 -265
rect 21280 -295 21315 -265
rect 21365 -295 21400 -265
rect 21450 -295 21485 -265
rect 21535 -295 21570 -265
rect 21620 -295 21655 -265
rect 21705 -295 21740 -265
rect 21790 -295 21825 -265
rect 21875 -295 21910 -265
rect 21960 -295 21995 -265
rect 22045 -295 22080 -265
rect 22130 -295 22165 -265
rect 22215 -295 22250 -265
rect 22300 -295 22335 -265
rect 22385 -295 22420 -265
rect 22470 -295 22505 -265
rect 22555 -295 22590 -265
rect 22640 -295 22675 -265
rect 22725 -295 22760 -265
rect 22810 -295 22845 -265
rect 22895 -295 22930 -265
rect 22980 -295 23015 -265
rect 23065 -295 23100 -265
rect 23150 -295 23185 -265
rect 23235 -295 23270 -265
rect 23320 -295 23355 -265
rect 23405 -295 23440 -265
rect 23490 -295 23525 -265
rect 23575 -295 23610 -265
rect 23660 -295 23695 -265
rect 23745 -295 23780 -265
rect 23830 -295 23865 -265
rect 23915 -295 23950 -265
rect 24000 -295 24035 -265
rect 24085 -295 24120 -265
rect 24170 -295 24205 -265
rect 24255 -295 24290 -265
rect 24340 -295 24375 -265
rect 24425 -295 24460 -265
rect 24510 -295 24545 -265
rect 24595 -295 24630 -265
rect 24680 -295 24715 -265
rect 24765 -295 24800 -265
rect 24850 -295 24885 -265
rect 24935 -295 24970 -265
rect 25020 -295 25055 -265
rect 25105 -295 25140 -265
rect 25190 -295 25225 -265
rect 25275 -295 25310 -265
rect 25360 -295 25395 -265
rect 25445 -295 25480 -265
rect 25530 -295 25565 -265
rect 25615 -295 25650 -265
rect 25700 -295 25735 -265
rect 25785 -295 25820 -265
rect 25870 -295 25905 -265
rect 25955 -295 25990 -265
rect 26040 -295 26075 -265
rect 26125 -295 26160 -265
rect 26210 -295 26245 -265
rect 26295 -295 26330 -265
rect 26380 -295 26415 -265
rect 26465 -295 26500 -265
rect 26550 -295 26585 -265
rect 26635 -295 26670 -265
rect 26720 -295 26755 -265
rect 26805 -295 26840 -265
rect 26890 -295 26925 -265
rect 26975 -295 27010 -265
rect 27060 -295 27095 -265
rect 27145 -295 27180 -265
rect 27230 -295 27265 -265
rect 27315 -295 27350 -265
rect 27400 -295 27435 -265
rect 27485 -295 27520 -265
rect 27570 -295 27605 -265
rect 27655 -295 27690 -265
rect 27740 -295 27775 -265
rect 27825 -295 27860 -265
rect 27910 -295 27945 -265
rect 27995 -295 28030 -265
rect 28080 -295 28115 -265
rect 28165 -295 28200 -265
rect 28250 -295 28285 -265
rect 28335 -295 28370 -265
rect 28420 -295 28455 -265
rect 28505 -295 28540 -265
rect 28590 -295 28625 -265
rect 28675 -295 28710 -265
rect 28760 -295 28795 -265
rect 28845 -295 28880 -265
rect 28930 -295 28965 -265
rect 29015 -295 29050 -265
rect 29100 -295 29135 -265
rect 29185 -295 29220 -265
rect 29270 -295 29305 -265
rect 29355 -295 29390 -265
rect 29440 -295 29475 -265
rect 29525 -295 29560 -265
rect 29610 -295 29645 -265
rect 29695 -295 29730 -265
rect 29780 -295 29815 -265
rect 29865 -295 29900 -265
rect 29950 -295 29985 -265
rect 30035 -295 30070 -265
rect 30120 -295 30155 -265
rect 30205 -295 30240 -265
rect 30290 -295 30325 -265
rect 30375 -295 30410 -265
rect 30460 -295 30495 -265
rect 30545 -295 30580 -265
rect 30630 -295 30665 -265
rect 30715 -295 30750 -265
rect 30800 -295 30835 -265
rect 30885 -295 30920 -265
rect 30970 -295 31005 -265
rect 31055 -295 31090 -265
rect 31140 -295 31175 -265
rect 31225 -295 31260 -265
rect 31310 -295 31345 -265
rect 31395 -295 31430 -265
rect 31480 -295 31515 -265
rect 31565 -295 31600 -265
rect 31650 -295 31685 -265
rect 31735 -295 31770 -265
rect 31820 -295 31855 -265
rect 31905 -295 31940 -265
rect 31990 -295 32025 -265
rect 32075 -295 32110 -265
rect 32160 -295 32195 -265
rect 32245 -295 32280 -265
rect 32330 -295 32365 -265
rect 32415 -295 32450 -265
rect 32500 -295 32535 -265
rect 32585 -295 32620 -265
rect 32670 -295 32705 -265
rect 32755 -295 32790 -265
rect 32840 -295 32875 -265
rect 32925 -295 32960 -265
rect 33010 -295 33045 -265
rect 33095 -295 33130 -265
rect 33180 -295 33215 -265
rect 33265 -295 33300 -265
rect 33350 -295 33385 -265
rect 33435 -295 33470 -265
rect 33520 -295 33555 -265
rect 33605 -295 33640 -265
rect 33690 -295 33725 -265
rect 33775 -295 33810 -265
rect 33860 -295 33895 -265
rect 33945 -295 33980 -265
rect 34030 -295 34065 -265
rect 34115 -295 34150 -265
rect 34200 -295 34235 -265
rect 34285 -295 34320 -265
rect 34370 -295 34405 -265
rect 34455 -295 34490 -265
rect 34540 -295 34575 -265
rect 34625 -295 34660 -265
rect 34710 -295 34745 -265
rect 34795 -295 34830 -265
rect 34880 -295 34915 -265
rect 34965 -295 35000 -265
rect 35050 -295 35085 -265
rect 35135 -295 35170 -265
rect 35220 -295 35255 -265
rect 35305 -295 35340 -265
rect 35390 -295 35425 -265
rect 35475 -295 35510 -265
rect 35560 -295 35595 -265
rect 35645 -295 35680 -265
rect 35730 -295 35765 -265
rect 35815 -295 35850 -265
rect 35900 -295 35935 -265
rect 35985 -295 36020 -265
rect 36070 -295 36105 -265
rect 36155 -295 36190 -265
rect 36240 -295 36275 -265
rect 36325 -295 36360 -265
rect 36410 -295 36445 -265
rect 36495 -295 36530 -265
rect 36580 -295 36615 -265
rect 36665 -295 36700 -265
rect 36750 -295 36785 -265
rect 36835 -295 36870 -265
rect 36920 -295 36955 -265
rect 37005 -295 37040 -265
rect 37090 -295 37125 -265
rect 37175 -295 37210 -265
rect 37260 -295 37295 -265
rect 37345 -295 37380 -265
rect 37430 -295 37465 -265
rect 37515 -295 37550 -265
rect 37600 -295 37635 -265
rect 37685 -295 37720 -265
rect 37770 -295 37805 -265
rect 37855 -295 37890 -265
rect 37940 -295 37975 -265
rect 38025 -295 38060 -265
rect 38110 -295 38145 -265
rect 38195 -295 38230 -265
rect 38280 -295 38315 -265
rect 38365 -295 38400 -265
rect 38450 -295 38485 -265
rect 38535 -295 38570 -265
rect 38620 -295 38655 -265
rect 38705 -295 38740 -265
rect 38790 -295 38825 -265
rect 38875 -295 38910 -265
rect 38960 -295 38995 -265
rect 39045 -295 39080 -265
rect 39130 -295 39165 -265
rect 39215 -295 39250 -265
rect 39300 -295 39335 -265
rect 39385 -295 39420 -265
rect 39470 -295 39505 -265
rect 39555 -295 39590 -265
rect 39640 -295 39675 -265
rect 39725 -295 39760 -265
rect 39810 -295 39845 -265
rect 39895 -295 39930 -265
rect 39980 -295 40015 -265
rect 40065 -295 40100 -265
rect 40150 -295 40185 -265
rect 40235 -295 40270 -265
rect 40320 -295 40355 -265
rect 40405 -295 40440 -265
rect 40490 -295 40525 -265
rect 40575 -295 40610 -265
rect 40660 -295 40695 -265
rect 40745 -295 40780 -265
rect 40830 -295 40865 -265
rect 40915 -295 40950 -265
rect 41000 -295 41035 -265
rect 41085 -295 41120 -265
rect 41170 -295 41205 -265
rect 41255 -295 41290 -265
rect 41340 -295 41375 -265
rect 41425 -295 41460 -265
rect 41510 -295 41545 -265
rect 41595 -295 41630 -265
rect 41680 -295 41715 -265
rect 41765 -295 41800 -265
rect 41850 -295 41885 -265
rect 41935 -295 41970 -265
rect 42020 -295 42055 -265
rect 42105 -295 42140 -265
rect 42190 -295 42225 -265
rect 42275 -295 42310 -265
rect 42360 -295 42395 -265
rect 42445 -295 42480 -265
rect 42530 -295 42565 -265
rect 42615 -295 42650 -265
rect 42700 -295 42735 -265
rect 42785 -295 42820 -265
rect 42870 -295 42905 -265
rect 42955 -295 42990 -265
rect 43040 -295 43075 -265
rect 43125 -295 43160 -265
rect 43210 -295 43245 -265
rect 43295 -295 43330 -265
rect 43380 -295 43415 -265
rect 43465 -295 43500 -265
rect 43550 -295 43585 -265
<< locali >>
rect 5 205 55 215
rect 5 175 15 205
rect 45 175 55 205
rect 5 155 55 175
rect 5 125 15 155
rect 45 125 55 155
rect 5 115 55 125
rect 90 205 140 215
rect 90 175 100 205
rect 130 175 140 205
rect 90 155 140 175
rect 90 125 100 155
rect 130 125 140 155
rect 90 115 140 125
rect 215 205 265 215
rect 215 175 225 205
rect 255 175 265 205
rect 215 155 265 175
rect 215 125 225 155
rect 255 125 265 155
rect 215 115 265 125
rect 300 205 350 215
rect 300 175 310 205
rect 340 175 350 205
rect 300 155 350 175
rect 300 125 310 155
rect 340 125 350 155
rect 300 115 350 125
rect 385 205 435 215
rect 385 175 395 205
rect 425 175 435 205
rect 385 155 435 175
rect 385 125 395 155
rect 425 125 435 155
rect 385 115 435 125
rect 470 205 520 215
rect 470 175 480 205
rect 510 175 520 205
rect 470 155 520 175
rect 470 125 480 155
rect 510 125 520 155
rect 470 115 520 125
rect 555 205 605 215
rect 555 175 565 205
rect 595 175 605 205
rect 555 155 605 175
rect 555 125 565 155
rect 595 125 605 155
rect 555 115 605 125
rect 750 205 800 215
rect 750 175 760 205
rect 790 175 800 205
rect 750 155 800 175
rect 750 125 760 155
rect 790 125 800 155
rect 750 115 800 125
rect 835 205 885 215
rect 835 175 845 205
rect 875 175 885 205
rect 835 155 885 175
rect 835 125 845 155
rect 875 125 885 155
rect 835 115 885 125
rect 920 205 970 215
rect 920 175 930 205
rect 960 175 970 205
rect 920 155 970 175
rect 920 125 930 155
rect 960 125 970 155
rect 920 115 970 125
rect 1005 205 1055 215
rect 1005 175 1015 205
rect 1045 175 1055 205
rect 1005 155 1055 175
rect 1005 125 1015 155
rect 1045 125 1055 155
rect 1005 115 1055 125
rect 1090 205 1140 215
rect 1090 175 1100 205
rect 1130 175 1140 205
rect 1090 155 1140 175
rect 1090 125 1100 155
rect 1130 125 1140 155
rect 1090 115 1140 125
rect 1175 205 1225 215
rect 1175 175 1185 205
rect 1215 175 1225 205
rect 1175 155 1225 175
rect 1175 125 1185 155
rect 1215 125 1225 155
rect 1175 115 1225 125
rect 1260 205 1310 215
rect 1260 175 1270 205
rect 1300 175 1310 205
rect 1260 155 1310 175
rect 1260 125 1270 155
rect 1300 125 1310 155
rect 1260 115 1310 125
rect 1345 205 1395 215
rect 1345 175 1355 205
rect 1385 175 1395 205
rect 1345 155 1395 175
rect 1345 125 1355 155
rect 1385 125 1395 155
rect 1345 115 1395 125
rect 1430 205 1480 215
rect 1430 175 1440 205
rect 1470 175 1480 205
rect 1430 155 1480 175
rect 1430 125 1440 155
rect 1470 125 1480 155
rect 1430 115 1480 125
rect 1515 205 1565 215
rect 1515 175 1525 205
rect 1555 175 1565 205
rect 1515 155 1565 175
rect 1515 125 1525 155
rect 1555 125 1565 155
rect 1515 115 1565 125
rect 1600 205 1650 215
rect 1600 175 1610 205
rect 1640 175 1650 205
rect 1600 155 1650 175
rect 1600 125 1610 155
rect 1640 125 1650 155
rect 1600 115 1650 125
rect 1685 205 1735 215
rect 1685 175 1695 205
rect 1725 175 1735 205
rect 1685 155 1735 175
rect 1685 125 1695 155
rect 1725 125 1735 155
rect 1685 115 1735 125
rect 1770 205 1820 215
rect 1770 175 1780 205
rect 1810 175 1820 205
rect 1770 155 1820 175
rect 1770 125 1780 155
rect 1810 125 1820 155
rect 1770 115 1820 125
rect 1855 205 1905 215
rect 1855 175 1865 205
rect 1895 175 1905 205
rect 1855 155 1905 175
rect 1855 125 1865 155
rect 1895 125 1905 155
rect 1855 115 1905 125
rect 1940 205 1990 215
rect 1940 175 1950 205
rect 1980 175 1990 205
rect 1940 155 1990 175
rect 1940 125 1950 155
rect 1980 125 1990 155
rect 1940 115 1990 125
rect 2025 205 2075 215
rect 2025 175 2035 205
rect 2065 175 2075 205
rect 2025 155 2075 175
rect 2025 125 2035 155
rect 2065 125 2075 155
rect 2025 115 2075 125
rect 2110 205 2160 215
rect 2110 175 2120 205
rect 2150 175 2160 205
rect 2110 155 2160 175
rect 2110 125 2120 155
rect 2150 125 2160 155
rect 2110 115 2160 125
rect 2260 205 2310 215
rect 2260 175 2270 205
rect 2300 175 2310 205
rect 2260 155 2310 175
rect 2260 125 2270 155
rect 2300 125 2310 155
rect 2260 115 2310 125
rect 2345 205 2395 215
rect 2345 175 2355 205
rect 2385 175 2395 205
rect 2345 155 2395 175
rect 2345 125 2355 155
rect 2385 125 2395 155
rect 2345 115 2395 125
rect 2430 205 2480 215
rect 2430 175 2440 205
rect 2470 175 2480 205
rect 2430 155 2480 175
rect 2430 125 2440 155
rect 2470 125 2480 155
rect 2430 115 2480 125
rect 2515 205 2565 215
rect 2515 175 2525 205
rect 2555 175 2565 205
rect 2515 155 2565 175
rect 2515 125 2525 155
rect 2555 125 2565 155
rect 2515 115 2565 125
rect 2600 205 2650 215
rect 2600 175 2610 205
rect 2640 175 2650 205
rect 2600 155 2650 175
rect 2600 125 2610 155
rect 2640 125 2650 155
rect 2600 115 2650 125
rect 2685 205 2735 215
rect 2685 175 2695 205
rect 2725 175 2735 205
rect 2685 155 2735 175
rect 2685 125 2695 155
rect 2725 125 2735 155
rect 2685 115 2735 125
rect 2770 205 2820 215
rect 2770 175 2780 205
rect 2810 175 2820 205
rect 2770 155 2820 175
rect 2770 125 2780 155
rect 2810 125 2820 155
rect 2770 115 2820 125
rect 2855 205 2905 215
rect 2855 175 2865 205
rect 2895 175 2905 205
rect 2855 155 2905 175
rect 2855 125 2865 155
rect 2895 125 2905 155
rect 2855 115 2905 125
rect 2940 205 2990 215
rect 2940 175 2950 205
rect 2980 175 2990 205
rect 2940 155 2990 175
rect 2940 125 2950 155
rect 2980 125 2990 155
rect 2940 115 2990 125
rect 3025 205 3075 215
rect 3025 175 3035 205
rect 3065 175 3075 205
rect 3025 155 3075 175
rect 3025 125 3035 155
rect 3065 125 3075 155
rect 3025 115 3075 125
rect 3110 205 3160 215
rect 3110 175 3120 205
rect 3150 175 3160 205
rect 3110 155 3160 175
rect 3110 125 3120 155
rect 3150 125 3160 155
rect 3110 115 3160 125
rect 3195 205 3245 215
rect 3195 175 3205 205
rect 3235 175 3245 205
rect 3195 155 3245 175
rect 3195 125 3205 155
rect 3235 125 3245 155
rect 3195 115 3245 125
rect 3280 205 3330 215
rect 3280 175 3290 205
rect 3320 175 3330 205
rect 3280 155 3330 175
rect 3280 125 3290 155
rect 3320 125 3330 155
rect 3280 115 3330 125
rect 3365 205 3415 215
rect 3365 175 3375 205
rect 3405 175 3415 205
rect 3365 155 3415 175
rect 3365 125 3375 155
rect 3405 125 3415 155
rect 3365 115 3415 125
rect 3450 205 3500 215
rect 3450 175 3460 205
rect 3490 175 3500 205
rect 3450 155 3500 175
rect 3450 125 3460 155
rect 3490 125 3500 155
rect 3450 115 3500 125
rect 3535 205 3585 215
rect 3535 175 3545 205
rect 3575 175 3585 205
rect 3535 155 3585 175
rect 3535 125 3545 155
rect 3575 125 3585 155
rect 3535 115 3585 125
rect 3620 205 3670 215
rect 3620 175 3630 205
rect 3660 175 3670 205
rect 3620 155 3670 175
rect 3620 125 3630 155
rect 3660 125 3670 155
rect 3620 115 3670 125
rect 3705 205 3755 215
rect 3705 175 3715 205
rect 3745 175 3755 205
rect 3705 155 3755 175
rect 3705 125 3715 155
rect 3745 125 3755 155
rect 3705 115 3755 125
rect 3790 205 3840 215
rect 3790 175 3800 205
rect 3830 175 3840 205
rect 3790 155 3840 175
rect 3790 125 3800 155
rect 3830 125 3840 155
rect 3790 115 3840 125
rect 3875 205 3925 215
rect 3875 175 3885 205
rect 3915 175 3925 205
rect 3875 155 3925 175
rect 3875 125 3885 155
rect 3915 125 3925 155
rect 3875 115 3925 125
rect 3960 205 4010 215
rect 3960 175 3970 205
rect 4000 175 4010 205
rect 3960 155 4010 175
rect 3960 125 3970 155
rect 4000 125 4010 155
rect 3960 115 4010 125
rect 4045 205 4095 215
rect 4045 175 4055 205
rect 4085 175 4095 205
rect 4045 155 4095 175
rect 4045 125 4055 155
rect 4085 125 4095 155
rect 4045 115 4095 125
rect 4130 205 4180 215
rect 4130 175 4140 205
rect 4170 175 4180 205
rect 4130 155 4180 175
rect 4130 125 4140 155
rect 4170 125 4180 155
rect 4130 115 4180 125
rect 4215 205 4265 215
rect 4215 175 4225 205
rect 4255 175 4265 205
rect 4215 155 4265 175
rect 4215 125 4225 155
rect 4255 125 4265 155
rect 4215 115 4265 125
rect 4300 205 4350 215
rect 4300 175 4310 205
rect 4340 175 4350 205
rect 4300 155 4350 175
rect 4300 125 4310 155
rect 4340 125 4350 155
rect 4300 115 4350 125
rect 4385 205 4435 215
rect 4385 175 4395 205
rect 4425 175 4435 205
rect 4385 155 4435 175
rect 4385 125 4395 155
rect 4425 125 4435 155
rect 4385 115 4435 125
rect 4470 205 4520 215
rect 4470 175 4480 205
rect 4510 175 4520 205
rect 4470 155 4520 175
rect 4470 125 4480 155
rect 4510 125 4520 155
rect 4470 115 4520 125
rect 4555 205 4605 215
rect 4555 175 4565 205
rect 4595 175 4605 205
rect 4555 155 4605 175
rect 4555 125 4565 155
rect 4595 125 4605 155
rect 4555 115 4605 125
rect 4640 205 4690 215
rect 4640 175 4650 205
rect 4680 175 4690 205
rect 4640 155 4690 175
rect 4640 125 4650 155
rect 4680 125 4690 155
rect 4640 115 4690 125
rect 4725 205 4775 215
rect 4725 175 4735 205
rect 4765 175 4775 205
rect 4725 155 4775 175
rect 4725 125 4735 155
rect 4765 125 4775 155
rect 4725 115 4775 125
rect 4810 205 4860 215
rect 4810 175 4820 205
rect 4850 175 4860 205
rect 4810 155 4860 175
rect 4810 125 4820 155
rect 4850 125 4860 155
rect 4810 115 4860 125
rect 4895 205 4945 215
rect 4895 175 4905 205
rect 4935 175 4945 205
rect 4895 155 4945 175
rect 4895 125 4905 155
rect 4935 125 4945 155
rect 4895 115 4945 125
rect 4980 205 5030 215
rect 4980 175 4990 205
rect 5020 175 5030 205
rect 4980 155 5030 175
rect 4980 125 4990 155
rect 5020 125 5030 155
rect 4980 115 5030 125
rect 5065 205 5115 215
rect 5065 175 5075 205
rect 5105 175 5115 205
rect 5065 155 5115 175
rect 5065 125 5075 155
rect 5105 125 5115 155
rect 5065 115 5115 125
rect 5150 205 5200 215
rect 5150 175 5160 205
rect 5190 175 5200 205
rect 5150 155 5200 175
rect 5150 125 5160 155
rect 5190 125 5200 155
rect 5150 115 5200 125
rect 5235 205 5285 215
rect 5235 175 5245 205
rect 5275 175 5285 205
rect 5235 155 5285 175
rect 5235 125 5245 155
rect 5275 125 5285 155
rect 5235 115 5285 125
rect 5320 205 5370 215
rect 5320 175 5330 205
rect 5360 175 5370 205
rect 5320 155 5370 175
rect 5320 125 5330 155
rect 5360 125 5370 155
rect 5320 115 5370 125
rect 5405 205 5455 215
rect 5405 175 5415 205
rect 5445 175 5455 205
rect 5405 155 5455 175
rect 5405 125 5415 155
rect 5445 125 5455 155
rect 5405 115 5455 125
rect 5490 205 5540 215
rect 5490 175 5500 205
rect 5530 175 5540 205
rect 5490 155 5540 175
rect 5490 125 5500 155
rect 5530 125 5540 155
rect 5490 115 5540 125
rect 5575 205 5625 215
rect 5575 175 5585 205
rect 5615 175 5625 205
rect 5575 155 5625 175
rect 5575 125 5585 155
rect 5615 125 5625 155
rect 5575 115 5625 125
rect 5660 205 5710 215
rect 5660 175 5670 205
rect 5700 175 5710 205
rect 5660 155 5710 175
rect 5660 125 5670 155
rect 5700 125 5710 155
rect 5660 115 5710 125
rect 5745 205 5795 215
rect 5745 175 5755 205
rect 5785 175 5795 205
rect 5745 155 5795 175
rect 5745 125 5755 155
rect 5785 125 5795 155
rect 5745 115 5795 125
rect 5830 205 5880 215
rect 5830 175 5840 205
rect 5870 175 5880 205
rect 5830 155 5880 175
rect 5830 125 5840 155
rect 5870 125 5880 155
rect 5830 115 5880 125
rect 5915 205 5965 215
rect 5915 175 5925 205
rect 5955 175 5965 205
rect 5915 155 5965 175
rect 5915 125 5925 155
rect 5955 125 5965 155
rect 5915 115 5965 125
rect 6000 205 6050 215
rect 6000 175 6010 205
rect 6040 175 6050 205
rect 6000 155 6050 175
rect 6000 125 6010 155
rect 6040 125 6050 155
rect 6000 115 6050 125
rect 6085 205 6135 215
rect 6085 175 6095 205
rect 6125 175 6135 205
rect 6085 155 6135 175
rect 6085 125 6095 155
rect 6125 125 6135 155
rect 6085 115 6135 125
rect 6170 205 6220 215
rect 6170 175 6180 205
rect 6210 175 6220 205
rect 6170 155 6220 175
rect 6170 125 6180 155
rect 6210 125 6220 155
rect 6170 115 6220 125
rect 6255 205 6305 215
rect 6255 175 6265 205
rect 6295 175 6305 205
rect 6255 155 6305 175
rect 6255 125 6265 155
rect 6295 125 6305 155
rect 6255 115 6305 125
rect 6340 205 6390 215
rect 6340 175 6350 205
rect 6380 175 6390 205
rect 6340 155 6390 175
rect 6340 125 6350 155
rect 6380 125 6390 155
rect 6340 115 6390 125
rect 6425 205 6475 215
rect 6425 175 6435 205
rect 6465 175 6475 205
rect 6425 155 6475 175
rect 6425 125 6435 155
rect 6465 125 6475 155
rect 6425 115 6475 125
rect 6510 205 6560 215
rect 6510 175 6520 205
rect 6550 175 6560 205
rect 6510 155 6560 175
rect 6510 125 6520 155
rect 6550 125 6560 155
rect 6510 115 6560 125
rect 6595 205 6645 215
rect 6595 175 6605 205
rect 6635 175 6645 205
rect 6595 155 6645 175
rect 6595 125 6605 155
rect 6635 125 6645 155
rect 6595 115 6645 125
rect 6680 205 6730 215
rect 6680 175 6690 205
rect 6720 175 6730 205
rect 6680 155 6730 175
rect 6680 125 6690 155
rect 6720 125 6730 155
rect 6680 115 6730 125
rect 6765 205 6815 215
rect 6765 175 6775 205
rect 6805 175 6815 205
rect 6765 155 6815 175
rect 6765 125 6775 155
rect 6805 125 6815 155
rect 6765 115 6815 125
rect 6850 205 6900 215
rect 6850 175 6860 205
rect 6890 175 6900 205
rect 6850 155 6900 175
rect 6850 125 6860 155
rect 6890 125 6900 155
rect 6850 115 6900 125
rect 6935 205 6985 215
rect 6935 175 6945 205
rect 6975 175 6985 205
rect 6935 155 6985 175
rect 6935 125 6945 155
rect 6975 125 6985 155
rect 6935 115 6985 125
rect 7020 205 7070 215
rect 7020 175 7030 205
rect 7060 175 7070 205
rect 7020 155 7070 175
rect 7020 125 7030 155
rect 7060 125 7070 155
rect 7020 115 7070 125
rect 7105 205 7155 215
rect 7105 175 7115 205
rect 7145 175 7155 205
rect 7105 155 7155 175
rect 7105 125 7115 155
rect 7145 125 7155 155
rect 7105 115 7155 125
rect 7190 205 7240 215
rect 7190 175 7200 205
rect 7230 175 7240 205
rect 7190 155 7240 175
rect 7190 125 7200 155
rect 7230 125 7240 155
rect 7190 115 7240 125
rect 7275 205 7325 215
rect 7275 175 7285 205
rect 7315 175 7325 205
rect 7275 155 7325 175
rect 7275 125 7285 155
rect 7315 125 7325 155
rect 7275 115 7325 125
rect 7360 205 7410 215
rect 7360 175 7370 205
rect 7400 175 7410 205
rect 7360 155 7410 175
rect 7360 125 7370 155
rect 7400 125 7410 155
rect 7360 115 7410 125
rect 7445 205 7495 215
rect 7445 175 7455 205
rect 7485 175 7495 205
rect 7445 155 7495 175
rect 7445 125 7455 155
rect 7485 125 7495 155
rect 7445 115 7495 125
rect 7530 205 7580 215
rect 7530 175 7540 205
rect 7570 175 7580 205
rect 7530 155 7580 175
rect 7530 125 7540 155
rect 7570 125 7580 155
rect 7530 115 7580 125
rect 7615 205 7665 215
rect 7615 175 7625 205
rect 7655 175 7665 205
rect 7615 155 7665 175
rect 7615 125 7625 155
rect 7655 125 7665 155
rect 7615 115 7665 125
rect 7700 205 7750 215
rect 7700 175 7710 205
rect 7740 175 7750 205
rect 7700 155 7750 175
rect 7700 125 7710 155
rect 7740 125 7750 155
rect 7700 115 7750 125
rect 7850 205 7900 215
rect 7850 175 7860 205
rect 7890 175 7900 205
rect 7850 155 7900 175
rect 7850 125 7860 155
rect 7890 125 7900 155
rect 7850 115 7900 125
rect 7935 205 7985 215
rect 7935 175 7945 205
rect 7975 175 7985 205
rect 7935 155 7985 175
rect 7935 125 7945 155
rect 7975 125 7985 155
rect 7935 115 7985 125
rect 8020 205 8070 215
rect 8020 175 8030 205
rect 8060 175 8070 205
rect 8020 155 8070 175
rect 8020 125 8030 155
rect 8060 125 8070 155
rect 8020 115 8070 125
rect 8105 205 8155 215
rect 8105 175 8115 205
rect 8145 175 8155 205
rect 8105 155 8155 175
rect 8105 125 8115 155
rect 8145 125 8155 155
rect 8105 115 8155 125
rect 8190 205 8240 215
rect 8190 175 8200 205
rect 8230 175 8240 205
rect 8190 155 8240 175
rect 8190 125 8200 155
rect 8230 125 8240 155
rect 8190 115 8240 125
rect 8275 205 8325 215
rect 8275 175 8285 205
rect 8315 175 8325 205
rect 8275 155 8325 175
rect 8275 125 8285 155
rect 8315 125 8325 155
rect 8275 115 8325 125
rect 8360 205 8410 215
rect 8360 175 8370 205
rect 8400 175 8410 205
rect 8360 155 8410 175
rect 8360 125 8370 155
rect 8400 125 8410 155
rect 8360 115 8410 125
rect 8445 205 8495 215
rect 8445 175 8455 205
rect 8485 175 8495 205
rect 8445 155 8495 175
rect 8445 125 8455 155
rect 8485 125 8495 155
rect 8445 115 8495 125
rect 8530 205 8580 215
rect 8530 175 8540 205
rect 8570 175 8580 205
rect 8530 155 8580 175
rect 8530 125 8540 155
rect 8570 125 8580 155
rect 8530 115 8580 125
rect 8615 205 8665 215
rect 8615 175 8625 205
rect 8655 175 8665 205
rect 8615 155 8665 175
rect 8615 125 8625 155
rect 8655 125 8665 155
rect 8615 115 8665 125
rect 8700 205 8750 215
rect 8700 175 8710 205
rect 8740 175 8750 205
rect 8700 155 8750 175
rect 8700 125 8710 155
rect 8740 125 8750 155
rect 8700 115 8750 125
rect 8785 205 8835 215
rect 8785 175 8795 205
rect 8825 175 8835 205
rect 8785 155 8835 175
rect 8785 125 8795 155
rect 8825 125 8835 155
rect 8785 115 8835 125
rect 8870 205 8920 215
rect 8870 175 8880 205
rect 8910 175 8920 205
rect 8870 155 8920 175
rect 8870 125 8880 155
rect 8910 125 8920 155
rect 8870 115 8920 125
rect 8955 205 9005 215
rect 8955 175 8965 205
rect 8995 175 9005 205
rect 8955 155 9005 175
rect 8955 125 8965 155
rect 8995 125 9005 155
rect 8955 115 9005 125
rect 9040 205 9090 215
rect 9040 175 9050 205
rect 9080 175 9090 205
rect 9040 155 9090 175
rect 9040 125 9050 155
rect 9080 125 9090 155
rect 9040 115 9090 125
rect 9125 205 9175 215
rect 9125 175 9135 205
rect 9165 175 9175 205
rect 9125 155 9175 175
rect 9125 125 9135 155
rect 9165 125 9175 155
rect 9125 115 9175 125
rect 9210 205 9260 215
rect 9210 175 9220 205
rect 9250 175 9260 205
rect 9210 155 9260 175
rect 9210 125 9220 155
rect 9250 125 9260 155
rect 9210 115 9260 125
rect 9295 205 9345 215
rect 9295 175 9305 205
rect 9335 175 9345 205
rect 9295 155 9345 175
rect 9295 125 9305 155
rect 9335 125 9345 155
rect 9295 115 9345 125
rect 9380 205 9430 215
rect 9380 175 9390 205
rect 9420 175 9430 205
rect 9380 155 9430 175
rect 9380 125 9390 155
rect 9420 125 9430 155
rect 9380 115 9430 125
rect 9465 205 9515 215
rect 9465 175 9475 205
rect 9505 175 9515 205
rect 9465 155 9515 175
rect 9465 125 9475 155
rect 9505 125 9515 155
rect 9465 115 9515 125
rect 9550 205 9600 215
rect 9550 175 9560 205
rect 9590 175 9600 205
rect 9550 155 9600 175
rect 9550 125 9560 155
rect 9590 125 9600 155
rect 9550 115 9600 125
rect 9635 205 9685 215
rect 9635 175 9645 205
rect 9675 175 9685 205
rect 9635 155 9685 175
rect 9635 125 9645 155
rect 9675 125 9685 155
rect 9635 115 9685 125
rect 9720 205 9770 215
rect 9720 175 9730 205
rect 9760 175 9770 205
rect 9720 155 9770 175
rect 9720 125 9730 155
rect 9760 125 9770 155
rect 9720 115 9770 125
rect 9805 205 9855 215
rect 9805 175 9815 205
rect 9845 175 9855 205
rect 9805 155 9855 175
rect 9805 125 9815 155
rect 9845 125 9855 155
rect 9805 115 9855 125
rect 9890 205 9940 215
rect 9890 175 9900 205
rect 9930 175 9940 205
rect 9890 155 9940 175
rect 9890 125 9900 155
rect 9930 125 9940 155
rect 9890 115 9940 125
rect 9975 205 10025 215
rect 9975 175 9985 205
rect 10015 175 10025 205
rect 9975 155 10025 175
rect 9975 125 9985 155
rect 10015 125 10025 155
rect 9975 115 10025 125
rect 10060 205 10110 215
rect 10060 175 10070 205
rect 10100 175 10110 205
rect 10060 155 10110 175
rect 10060 125 10070 155
rect 10100 125 10110 155
rect 10060 115 10110 125
rect 10145 205 10195 215
rect 10145 175 10155 205
rect 10185 175 10195 205
rect 10145 155 10195 175
rect 10145 125 10155 155
rect 10185 125 10195 155
rect 10145 115 10195 125
rect 10230 205 10280 215
rect 10230 175 10240 205
rect 10270 175 10280 205
rect 10230 155 10280 175
rect 10230 125 10240 155
rect 10270 125 10280 155
rect 10230 115 10280 125
rect 10315 205 10365 215
rect 10315 175 10325 205
rect 10355 175 10365 205
rect 10315 155 10365 175
rect 10315 125 10325 155
rect 10355 125 10365 155
rect 10315 115 10365 125
rect 10400 205 10450 215
rect 10400 175 10410 205
rect 10440 175 10450 205
rect 10400 155 10450 175
rect 10400 125 10410 155
rect 10440 125 10450 155
rect 10400 115 10450 125
rect 10485 205 10535 215
rect 10485 175 10495 205
rect 10525 175 10535 205
rect 10485 155 10535 175
rect 10485 125 10495 155
rect 10525 125 10535 155
rect 10485 115 10535 125
rect 10570 205 10620 215
rect 10570 175 10580 205
rect 10610 175 10620 205
rect 10570 155 10620 175
rect 10570 125 10580 155
rect 10610 125 10620 155
rect 10570 115 10620 125
rect 10655 205 10705 215
rect 10655 175 10665 205
rect 10695 175 10705 205
rect 10655 155 10705 175
rect 10655 125 10665 155
rect 10695 125 10705 155
rect 10655 115 10705 125
rect 10740 205 10790 215
rect 10740 175 10750 205
rect 10780 175 10790 205
rect 10740 155 10790 175
rect 10740 125 10750 155
rect 10780 125 10790 155
rect 10740 115 10790 125
rect 10825 205 10875 215
rect 10825 175 10835 205
rect 10865 175 10875 205
rect 10825 155 10875 175
rect 10825 125 10835 155
rect 10865 125 10875 155
rect 10825 115 10875 125
rect 10910 205 10960 215
rect 10910 175 10920 205
rect 10950 175 10960 205
rect 10910 155 10960 175
rect 10910 125 10920 155
rect 10950 125 10960 155
rect 10910 115 10960 125
rect 10995 205 11045 215
rect 10995 175 11005 205
rect 11035 175 11045 205
rect 10995 155 11045 175
rect 10995 125 11005 155
rect 11035 125 11045 155
rect 10995 115 11045 125
rect 11080 205 11130 215
rect 11080 175 11090 205
rect 11120 175 11130 205
rect 11080 155 11130 175
rect 11080 125 11090 155
rect 11120 125 11130 155
rect 11080 115 11130 125
rect 11165 205 11215 215
rect 11165 175 11175 205
rect 11205 175 11215 205
rect 11165 155 11215 175
rect 11165 125 11175 155
rect 11205 125 11215 155
rect 11165 115 11215 125
rect 11250 205 11300 215
rect 11250 175 11260 205
rect 11290 175 11300 205
rect 11250 155 11300 175
rect 11250 125 11260 155
rect 11290 125 11300 155
rect 11250 115 11300 125
rect 11335 205 11385 215
rect 11335 175 11345 205
rect 11375 175 11385 205
rect 11335 155 11385 175
rect 11335 125 11345 155
rect 11375 125 11385 155
rect 11335 115 11385 125
rect 11420 205 11470 215
rect 11420 175 11430 205
rect 11460 175 11470 205
rect 11420 155 11470 175
rect 11420 125 11430 155
rect 11460 125 11470 155
rect 11420 115 11470 125
rect 11505 205 11555 215
rect 11505 175 11515 205
rect 11545 175 11555 205
rect 11505 155 11555 175
rect 11505 125 11515 155
rect 11545 125 11555 155
rect 11505 115 11555 125
rect 11590 205 11640 215
rect 11590 175 11600 205
rect 11630 175 11640 205
rect 11590 155 11640 175
rect 11590 125 11600 155
rect 11630 125 11640 155
rect 11590 115 11640 125
rect 11675 205 11725 215
rect 11675 175 11685 205
rect 11715 175 11725 205
rect 11675 155 11725 175
rect 11675 125 11685 155
rect 11715 125 11725 155
rect 11675 115 11725 125
rect 11760 205 11810 215
rect 11760 175 11770 205
rect 11800 175 11810 205
rect 11760 155 11810 175
rect 11760 125 11770 155
rect 11800 125 11810 155
rect 11760 115 11810 125
rect 11845 205 11895 215
rect 11845 175 11855 205
rect 11885 175 11895 205
rect 11845 155 11895 175
rect 11845 125 11855 155
rect 11885 125 11895 155
rect 11845 115 11895 125
rect 11930 205 11980 215
rect 11930 175 11940 205
rect 11970 175 11980 205
rect 11930 155 11980 175
rect 11930 125 11940 155
rect 11970 125 11980 155
rect 11930 115 11980 125
rect 12015 205 12065 215
rect 12015 175 12025 205
rect 12055 175 12065 205
rect 12015 155 12065 175
rect 12015 125 12025 155
rect 12055 125 12065 155
rect 12015 115 12065 125
rect 12100 205 12150 215
rect 12100 175 12110 205
rect 12140 175 12150 205
rect 12100 155 12150 175
rect 12100 125 12110 155
rect 12140 125 12150 155
rect 12100 115 12150 125
rect 12185 205 12235 215
rect 12185 175 12195 205
rect 12225 175 12235 205
rect 12185 155 12235 175
rect 12185 125 12195 155
rect 12225 125 12235 155
rect 12185 115 12235 125
rect 12270 205 12320 215
rect 12270 175 12280 205
rect 12310 175 12320 205
rect 12270 155 12320 175
rect 12270 125 12280 155
rect 12310 125 12320 155
rect 12270 115 12320 125
rect 12355 205 12405 215
rect 12355 175 12365 205
rect 12395 175 12405 205
rect 12355 155 12405 175
rect 12355 125 12365 155
rect 12395 125 12405 155
rect 12355 115 12405 125
rect 12440 205 12490 215
rect 12440 175 12450 205
rect 12480 175 12490 205
rect 12440 155 12490 175
rect 12440 125 12450 155
rect 12480 125 12490 155
rect 12440 115 12490 125
rect 12525 205 12575 215
rect 12525 175 12535 205
rect 12565 175 12575 205
rect 12525 155 12575 175
rect 12525 125 12535 155
rect 12565 125 12575 155
rect 12525 115 12575 125
rect 12610 205 12660 215
rect 12610 175 12620 205
rect 12650 175 12660 205
rect 12610 155 12660 175
rect 12610 125 12620 155
rect 12650 125 12660 155
rect 12610 115 12660 125
rect 12695 205 12745 215
rect 12695 175 12705 205
rect 12735 175 12745 205
rect 12695 155 12745 175
rect 12695 125 12705 155
rect 12735 125 12745 155
rect 12695 115 12745 125
rect 12780 205 12830 215
rect 12780 175 12790 205
rect 12820 175 12830 205
rect 12780 155 12830 175
rect 12780 125 12790 155
rect 12820 125 12830 155
rect 12780 115 12830 125
rect 12865 205 12915 215
rect 12865 175 12875 205
rect 12905 175 12915 205
rect 12865 155 12915 175
rect 12865 125 12875 155
rect 12905 125 12915 155
rect 12865 115 12915 125
rect 12950 205 13000 215
rect 12950 175 12960 205
rect 12990 175 13000 205
rect 12950 155 13000 175
rect 12950 125 12960 155
rect 12990 125 13000 155
rect 12950 115 13000 125
rect 13035 205 13085 215
rect 13035 175 13045 205
rect 13075 175 13085 205
rect 13035 155 13085 175
rect 13035 125 13045 155
rect 13075 125 13085 155
rect 13035 115 13085 125
rect 13120 205 13170 215
rect 13120 175 13130 205
rect 13160 175 13170 205
rect 13120 155 13170 175
rect 13120 125 13130 155
rect 13160 125 13170 155
rect 13120 115 13170 125
rect 13205 205 13255 215
rect 13205 175 13215 205
rect 13245 175 13255 205
rect 13205 155 13255 175
rect 13205 125 13215 155
rect 13245 125 13255 155
rect 13205 115 13255 125
rect 13290 205 13340 215
rect 13290 175 13300 205
rect 13330 175 13340 205
rect 13290 155 13340 175
rect 13290 125 13300 155
rect 13330 125 13340 155
rect 13290 115 13340 125
rect 13375 205 13425 215
rect 13375 175 13385 205
rect 13415 175 13425 205
rect 13375 155 13425 175
rect 13375 125 13385 155
rect 13415 125 13425 155
rect 13375 115 13425 125
rect 13460 205 13510 215
rect 13460 175 13470 205
rect 13500 175 13510 205
rect 13460 155 13510 175
rect 13460 125 13470 155
rect 13500 125 13510 155
rect 13460 115 13510 125
rect 13545 205 13595 215
rect 13545 175 13555 205
rect 13585 175 13595 205
rect 13545 155 13595 175
rect 13545 125 13555 155
rect 13585 125 13595 155
rect 13545 115 13595 125
rect 13630 205 13680 215
rect 13630 175 13640 205
rect 13670 175 13680 205
rect 13630 155 13680 175
rect 13630 125 13640 155
rect 13670 125 13680 155
rect 13630 115 13680 125
rect 13715 205 13765 215
rect 13715 175 13725 205
rect 13755 175 13765 205
rect 13715 155 13765 175
rect 13715 125 13725 155
rect 13755 125 13765 155
rect 13715 115 13765 125
rect 13800 205 13850 215
rect 13800 175 13810 205
rect 13840 175 13850 205
rect 13800 155 13850 175
rect 13800 125 13810 155
rect 13840 125 13850 155
rect 13800 115 13850 125
rect 13885 205 13935 215
rect 13885 175 13895 205
rect 13925 175 13935 205
rect 13885 155 13935 175
rect 13885 125 13895 155
rect 13925 125 13935 155
rect 13885 115 13935 125
rect 13970 205 14020 215
rect 13970 175 13980 205
rect 14010 175 14020 205
rect 13970 155 14020 175
rect 13970 125 13980 155
rect 14010 125 14020 155
rect 13970 115 14020 125
rect 14055 205 14105 215
rect 14055 175 14065 205
rect 14095 175 14105 205
rect 14055 155 14105 175
rect 14055 125 14065 155
rect 14095 125 14105 155
rect 14055 115 14105 125
rect 14140 205 14190 215
rect 14140 175 14150 205
rect 14180 175 14190 205
rect 14140 155 14190 175
rect 14140 125 14150 155
rect 14180 125 14190 155
rect 14140 115 14190 125
rect 14225 205 14275 215
rect 14225 175 14235 205
rect 14265 175 14275 205
rect 14225 155 14275 175
rect 14225 125 14235 155
rect 14265 125 14275 155
rect 14225 115 14275 125
rect 14310 205 14360 215
rect 14310 175 14320 205
rect 14350 175 14360 205
rect 14310 155 14360 175
rect 14310 125 14320 155
rect 14350 125 14360 155
rect 14310 115 14360 125
rect 14395 205 14445 215
rect 14395 175 14405 205
rect 14435 175 14445 205
rect 14395 155 14445 175
rect 14395 125 14405 155
rect 14435 125 14445 155
rect 14395 115 14445 125
rect 14480 205 14530 215
rect 14480 175 14490 205
rect 14520 175 14530 205
rect 14480 155 14530 175
rect 14480 125 14490 155
rect 14520 125 14530 155
rect 14480 115 14530 125
rect 14565 205 14615 215
rect 14565 175 14575 205
rect 14605 175 14615 205
rect 14565 155 14615 175
rect 14565 125 14575 155
rect 14605 125 14615 155
rect 14565 115 14615 125
rect 14650 205 14700 215
rect 14650 175 14660 205
rect 14690 175 14700 205
rect 14650 155 14700 175
rect 14650 125 14660 155
rect 14690 125 14700 155
rect 14650 115 14700 125
rect 14735 205 14785 215
rect 14735 175 14745 205
rect 14775 175 14785 205
rect 14735 155 14785 175
rect 14735 125 14745 155
rect 14775 125 14785 155
rect 14735 115 14785 125
rect 14820 205 14870 215
rect 14820 175 14830 205
rect 14860 175 14870 205
rect 14820 155 14870 175
rect 14820 125 14830 155
rect 14860 125 14870 155
rect 14820 115 14870 125
rect 14905 205 14955 215
rect 14905 175 14915 205
rect 14945 175 14955 205
rect 14905 155 14955 175
rect 14905 125 14915 155
rect 14945 125 14955 155
rect 14905 115 14955 125
rect 14990 205 15040 215
rect 14990 175 15000 205
rect 15030 175 15040 205
rect 14990 155 15040 175
rect 14990 125 15000 155
rect 15030 125 15040 155
rect 14990 115 15040 125
rect 15075 205 15125 215
rect 15075 175 15085 205
rect 15115 175 15125 205
rect 15075 155 15125 175
rect 15075 125 15085 155
rect 15115 125 15125 155
rect 15075 115 15125 125
rect 15160 205 15210 215
rect 15160 175 15170 205
rect 15200 175 15210 205
rect 15160 155 15210 175
rect 15160 125 15170 155
rect 15200 125 15210 155
rect 15160 115 15210 125
rect 15245 205 15295 215
rect 15245 175 15255 205
rect 15285 175 15295 205
rect 15245 155 15295 175
rect 15245 125 15255 155
rect 15285 125 15295 155
rect 15245 115 15295 125
rect 15330 205 15380 215
rect 15330 175 15340 205
rect 15370 175 15380 205
rect 15330 155 15380 175
rect 15330 125 15340 155
rect 15370 125 15380 155
rect 15330 115 15380 125
rect 15415 205 15465 215
rect 15415 175 15425 205
rect 15455 175 15465 205
rect 15415 155 15465 175
rect 15415 125 15425 155
rect 15455 125 15465 155
rect 15415 115 15465 125
rect 15500 205 15550 215
rect 15500 175 15510 205
rect 15540 175 15550 205
rect 15500 155 15550 175
rect 15500 125 15510 155
rect 15540 125 15550 155
rect 15500 115 15550 125
rect 15585 205 15635 215
rect 15585 175 15595 205
rect 15625 175 15635 205
rect 15585 155 15635 175
rect 15585 125 15595 155
rect 15625 125 15635 155
rect 15585 115 15635 125
rect 15670 205 15720 215
rect 15670 175 15680 205
rect 15710 175 15720 205
rect 15670 155 15720 175
rect 15670 125 15680 155
rect 15710 125 15720 155
rect 15670 115 15720 125
rect 15755 205 15805 215
rect 15755 175 15765 205
rect 15795 175 15805 205
rect 15755 155 15805 175
rect 15755 125 15765 155
rect 15795 125 15805 155
rect 15755 115 15805 125
rect 15840 205 15890 215
rect 15840 175 15850 205
rect 15880 175 15890 205
rect 15840 155 15890 175
rect 15840 125 15850 155
rect 15880 125 15890 155
rect 15840 115 15890 125
rect 15925 205 15975 215
rect 15925 175 15935 205
rect 15965 175 15975 205
rect 15925 155 15975 175
rect 15925 125 15935 155
rect 15965 125 15975 155
rect 15925 115 15975 125
rect 16010 205 16060 215
rect 16010 175 16020 205
rect 16050 175 16060 205
rect 16010 155 16060 175
rect 16010 125 16020 155
rect 16050 125 16060 155
rect 16010 115 16060 125
rect 16095 205 16145 215
rect 16095 175 16105 205
rect 16135 175 16145 205
rect 16095 155 16145 175
rect 16095 125 16105 155
rect 16135 125 16145 155
rect 16095 115 16145 125
rect 16180 205 16230 215
rect 16180 175 16190 205
rect 16220 175 16230 205
rect 16180 155 16230 175
rect 16180 125 16190 155
rect 16220 125 16230 155
rect 16180 115 16230 125
rect 16265 205 16315 215
rect 16265 175 16275 205
rect 16305 175 16315 205
rect 16265 155 16315 175
rect 16265 125 16275 155
rect 16305 125 16315 155
rect 16265 115 16315 125
rect 16350 205 16400 215
rect 16350 175 16360 205
rect 16390 175 16400 205
rect 16350 155 16400 175
rect 16350 125 16360 155
rect 16390 125 16400 155
rect 16350 115 16400 125
rect 16435 205 16485 215
rect 16435 175 16445 205
rect 16475 175 16485 205
rect 16435 155 16485 175
rect 16435 125 16445 155
rect 16475 125 16485 155
rect 16435 115 16485 125
rect 16520 205 16570 215
rect 16520 175 16530 205
rect 16560 175 16570 205
rect 16520 155 16570 175
rect 16520 125 16530 155
rect 16560 125 16570 155
rect 16520 115 16570 125
rect 16605 205 16655 215
rect 16605 175 16615 205
rect 16645 175 16655 205
rect 16605 155 16655 175
rect 16605 125 16615 155
rect 16645 125 16655 155
rect 16605 115 16655 125
rect 16690 205 16740 215
rect 16690 175 16700 205
rect 16730 175 16740 205
rect 16690 155 16740 175
rect 16690 125 16700 155
rect 16730 125 16740 155
rect 16690 115 16740 125
rect 16775 205 16825 215
rect 16775 175 16785 205
rect 16815 175 16825 205
rect 16775 155 16825 175
rect 16775 125 16785 155
rect 16815 125 16825 155
rect 16775 115 16825 125
rect 16860 205 16910 215
rect 16860 175 16870 205
rect 16900 175 16910 205
rect 16860 155 16910 175
rect 16860 125 16870 155
rect 16900 125 16910 155
rect 16860 115 16910 125
rect 16945 205 16995 215
rect 16945 175 16955 205
rect 16985 175 16995 205
rect 16945 155 16995 175
rect 16945 125 16955 155
rect 16985 125 16995 155
rect 16945 115 16995 125
rect 17030 205 17080 215
rect 17030 175 17040 205
rect 17070 175 17080 205
rect 17030 155 17080 175
rect 17030 125 17040 155
rect 17070 125 17080 155
rect 17030 115 17080 125
rect 17115 205 17165 215
rect 17115 175 17125 205
rect 17155 175 17165 205
rect 17115 155 17165 175
rect 17115 125 17125 155
rect 17155 125 17165 155
rect 17115 115 17165 125
rect 17200 205 17250 215
rect 17200 175 17210 205
rect 17240 175 17250 205
rect 17200 155 17250 175
rect 17200 125 17210 155
rect 17240 125 17250 155
rect 17200 115 17250 125
rect 17285 205 17335 215
rect 17285 175 17295 205
rect 17325 175 17335 205
rect 17285 155 17335 175
rect 17285 125 17295 155
rect 17325 125 17335 155
rect 17285 115 17335 125
rect 17370 205 17420 215
rect 17370 175 17380 205
rect 17410 175 17420 205
rect 17370 155 17420 175
rect 17370 125 17380 155
rect 17410 125 17420 155
rect 17370 115 17420 125
rect 17455 205 17505 215
rect 17455 175 17465 205
rect 17495 175 17505 205
rect 17455 155 17505 175
rect 17455 125 17465 155
rect 17495 125 17505 155
rect 17455 115 17505 125
rect 17540 205 17590 215
rect 17540 175 17550 205
rect 17580 175 17590 205
rect 17540 155 17590 175
rect 17540 125 17550 155
rect 17580 125 17590 155
rect 17540 115 17590 125
rect 17625 205 17675 215
rect 17625 175 17635 205
rect 17665 175 17675 205
rect 17625 155 17675 175
rect 17625 125 17635 155
rect 17665 125 17675 155
rect 17625 115 17675 125
rect 17710 205 17760 215
rect 17710 175 17720 205
rect 17750 175 17760 205
rect 17710 155 17760 175
rect 17710 125 17720 155
rect 17750 125 17760 155
rect 17710 115 17760 125
rect 17795 205 17845 215
rect 17795 175 17805 205
rect 17835 175 17845 205
rect 17795 155 17845 175
rect 17795 125 17805 155
rect 17835 125 17845 155
rect 17795 115 17845 125
rect 17880 205 17930 215
rect 17880 175 17890 205
rect 17920 175 17930 205
rect 17880 155 17930 175
rect 17880 125 17890 155
rect 17920 125 17930 155
rect 17880 115 17930 125
rect 17965 205 18015 215
rect 17965 175 17975 205
rect 18005 175 18015 205
rect 17965 155 18015 175
rect 17965 125 17975 155
rect 18005 125 18015 155
rect 17965 115 18015 125
rect 18050 205 18100 215
rect 18050 175 18060 205
rect 18090 175 18100 205
rect 18050 155 18100 175
rect 18050 125 18060 155
rect 18090 125 18100 155
rect 18050 115 18100 125
rect 18135 205 18185 215
rect 18135 175 18145 205
rect 18175 175 18185 205
rect 18135 155 18185 175
rect 18135 125 18145 155
rect 18175 125 18185 155
rect 18135 115 18185 125
rect 18220 205 18270 215
rect 18220 175 18230 205
rect 18260 175 18270 205
rect 18220 155 18270 175
rect 18220 125 18230 155
rect 18260 125 18270 155
rect 18220 115 18270 125
rect 18305 205 18355 215
rect 18305 175 18315 205
rect 18345 175 18355 205
rect 18305 155 18355 175
rect 18305 125 18315 155
rect 18345 125 18355 155
rect 18305 115 18355 125
rect 18390 205 18440 215
rect 18390 175 18400 205
rect 18430 175 18440 205
rect 18390 155 18440 175
rect 18390 125 18400 155
rect 18430 125 18440 155
rect 18390 115 18440 125
rect 18475 205 18525 215
rect 18475 175 18485 205
rect 18515 175 18525 205
rect 18475 155 18525 175
rect 18475 125 18485 155
rect 18515 125 18525 155
rect 18475 115 18525 125
rect 18560 205 18610 215
rect 18560 175 18570 205
rect 18600 175 18610 205
rect 18560 155 18610 175
rect 18560 125 18570 155
rect 18600 125 18610 155
rect 18560 115 18610 125
rect 18645 205 18695 215
rect 18645 175 18655 205
rect 18685 175 18695 205
rect 18645 155 18695 175
rect 18645 125 18655 155
rect 18685 125 18695 155
rect 18645 115 18695 125
rect 18730 205 18780 215
rect 18730 175 18740 205
rect 18770 175 18780 205
rect 18730 155 18780 175
rect 18730 125 18740 155
rect 18770 125 18780 155
rect 18730 115 18780 125
rect 18815 205 18865 215
rect 18815 175 18825 205
rect 18855 175 18865 205
rect 18815 155 18865 175
rect 18815 125 18825 155
rect 18855 125 18865 155
rect 18815 115 18865 125
rect 18900 205 18950 215
rect 18900 175 18910 205
rect 18940 175 18950 205
rect 18900 155 18950 175
rect 18900 125 18910 155
rect 18940 125 18950 155
rect 18900 115 18950 125
rect 18985 205 19035 215
rect 18985 175 18995 205
rect 19025 175 19035 205
rect 18985 155 19035 175
rect 18985 125 18995 155
rect 19025 125 19035 155
rect 18985 115 19035 125
rect 19070 205 19120 215
rect 19070 175 19080 205
rect 19110 175 19120 205
rect 19070 155 19120 175
rect 19070 125 19080 155
rect 19110 125 19120 155
rect 19070 115 19120 125
rect 19155 205 19205 215
rect 19155 175 19165 205
rect 19195 175 19205 205
rect 19155 155 19205 175
rect 19155 125 19165 155
rect 19195 125 19205 155
rect 19155 115 19205 125
rect 19240 205 19290 215
rect 19240 175 19250 205
rect 19280 175 19290 205
rect 19240 155 19290 175
rect 19240 125 19250 155
rect 19280 125 19290 155
rect 19240 115 19290 125
rect 19325 205 19375 215
rect 19325 175 19335 205
rect 19365 175 19375 205
rect 19325 155 19375 175
rect 19325 125 19335 155
rect 19365 125 19375 155
rect 19325 115 19375 125
rect 19410 205 19460 215
rect 19410 175 19420 205
rect 19450 175 19460 205
rect 19410 155 19460 175
rect 19410 125 19420 155
rect 19450 125 19460 155
rect 19410 115 19460 125
rect 19495 205 19545 215
rect 19495 175 19505 205
rect 19535 175 19545 205
rect 19495 155 19545 175
rect 19495 125 19505 155
rect 19535 125 19545 155
rect 19495 115 19545 125
rect 19580 205 19630 215
rect 19580 175 19590 205
rect 19620 175 19630 205
rect 19580 155 19630 175
rect 19580 125 19590 155
rect 19620 125 19630 155
rect 19580 115 19630 125
rect 19665 205 19715 215
rect 19665 175 19675 205
rect 19705 175 19715 205
rect 19665 155 19715 175
rect 19665 125 19675 155
rect 19705 125 19715 155
rect 19665 115 19715 125
rect 19750 205 19800 215
rect 19750 175 19760 205
rect 19790 175 19800 205
rect 19750 155 19800 175
rect 19750 125 19760 155
rect 19790 125 19800 155
rect 19750 115 19800 125
rect 19835 205 19885 215
rect 19835 175 19845 205
rect 19875 175 19885 205
rect 19835 155 19885 175
rect 19835 125 19845 155
rect 19875 125 19885 155
rect 19835 115 19885 125
rect 19920 205 19970 215
rect 19920 175 19930 205
rect 19960 175 19970 205
rect 19920 155 19970 175
rect 19920 125 19930 155
rect 19960 125 19970 155
rect 19920 115 19970 125
rect 20005 205 20055 215
rect 20005 175 20015 205
rect 20045 175 20055 205
rect 20005 155 20055 175
rect 20005 125 20015 155
rect 20045 125 20055 155
rect 20005 115 20055 125
rect 20090 205 20140 215
rect 20090 175 20100 205
rect 20130 175 20140 205
rect 20090 155 20140 175
rect 20090 125 20100 155
rect 20130 125 20140 155
rect 20090 115 20140 125
rect 20175 205 20225 215
rect 20175 175 20185 205
rect 20215 175 20225 205
rect 20175 155 20225 175
rect 20175 125 20185 155
rect 20215 125 20225 155
rect 20175 115 20225 125
rect 20260 205 20310 215
rect 20260 175 20270 205
rect 20300 175 20310 205
rect 20260 155 20310 175
rect 20260 125 20270 155
rect 20300 125 20310 155
rect 20260 115 20310 125
rect 20345 205 20395 215
rect 20345 175 20355 205
rect 20385 175 20395 205
rect 20345 155 20395 175
rect 20345 125 20355 155
rect 20385 125 20395 155
rect 20345 115 20395 125
rect 20430 205 20480 215
rect 20430 175 20440 205
rect 20470 175 20480 205
rect 20430 155 20480 175
rect 20430 125 20440 155
rect 20470 125 20480 155
rect 20430 115 20480 125
rect 20515 205 20565 215
rect 20515 175 20525 205
rect 20555 175 20565 205
rect 20515 155 20565 175
rect 20515 125 20525 155
rect 20555 125 20565 155
rect 20515 115 20565 125
rect 20600 205 20650 215
rect 20600 175 20610 205
rect 20640 175 20650 205
rect 20600 155 20650 175
rect 20600 125 20610 155
rect 20640 125 20650 155
rect 20600 115 20650 125
rect 20685 205 20735 215
rect 20685 175 20695 205
rect 20725 175 20735 205
rect 20685 155 20735 175
rect 20685 125 20695 155
rect 20725 125 20735 155
rect 20685 115 20735 125
rect 20770 205 20820 215
rect 20770 175 20780 205
rect 20810 175 20820 205
rect 20770 155 20820 175
rect 20770 125 20780 155
rect 20810 125 20820 155
rect 20770 115 20820 125
rect 20855 205 20905 215
rect 20855 175 20865 205
rect 20895 175 20905 205
rect 20855 155 20905 175
rect 20855 125 20865 155
rect 20895 125 20905 155
rect 20855 115 20905 125
rect 20940 205 20990 215
rect 20940 175 20950 205
rect 20980 175 20990 205
rect 20940 155 20990 175
rect 20940 125 20950 155
rect 20980 125 20990 155
rect 20940 115 20990 125
rect 21025 205 21075 215
rect 21025 175 21035 205
rect 21065 175 21075 205
rect 21025 155 21075 175
rect 21025 125 21035 155
rect 21065 125 21075 155
rect 21025 115 21075 125
rect 21110 205 21160 215
rect 21110 175 21120 205
rect 21150 175 21160 205
rect 21110 155 21160 175
rect 21110 125 21120 155
rect 21150 125 21160 155
rect 21110 115 21160 125
rect 21195 205 21245 215
rect 21195 175 21205 205
rect 21235 175 21245 205
rect 21195 155 21245 175
rect 21195 125 21205 155
rect 21235 125 21245 155
rect 21195 115 21245 125
rect 21280 205 21330 215
rect 21280 175 21290 205
rect 21320 175 21330 205
rect 21280 155 21330 175
rect 21280 125 21290 155
rect 21320 125 21330 155
rect 21280 115 21330 125
rect 21365 205 21415 215
rect 21365 175 21375 205
rect 21405 175 21415 205
rect 21365 155 21415 175
rect 21365 125 21375 155
rect 21405 125 21415 155
rect 21365 115 21415 125
rect 21450 205 21500 215
rect 21450 175 21460 205
rect 21490 175 21500 205
rect 21450 155 21500 175
rect 21450 125 21460 155
rect 21490 125 21500 155
rect 21450 115 21500 125
rect 21535 205 21585 215
rect 21535 175 21545 205
rect 21575 175 21585 205
rect 21535 155 21585 175
rect 21535 125 21545 155
rect 21575 125 21585 155
rect 21535 115 21585 125
rect 21620 205 21670 215
rect 21620 175 21630 205
rect 21660 175 21670 205
rect 21620 155 21670 175
rect 21620 125 21630 155
rect 21660 125 21670 155
rect 21620 115 21670 125
rect 21705 205 21755 215
rect 21705 175 21715 205
rect 21745 175 21755 205
rect 21705 155 21755 175
rect 21705 125 21715 155
rect 21745 125 21755 155
rect 21705 115 21755 125
rect 21790 205 21840 215
rect 21790 175 21800 205
rect 21830 175 21840 205
rect 21790 155 21840 175
rect 21790 125 21800 155
rect 21830 125 21840 155
rect 21790 115 21840 125
rect 21875 205 21925 215
rect 21875 175 21885 205
rect 21915 175 21925 205
rect 21875 155 21925 175
rect 21875 125 21885 155
rect 21915 125 21925 155
rect 21875 115 21925 125
rect 21960 205 22010 215
rect 21960 175 21970 205
rect 22000 175 22010 205
rect 21960 155 22010 175
rect 21960 125 21970 155
rect 22000 125 22010 155
rect 21960 115 22010 125
rect 22045 205 22095 215
rect 22045 175 22055 205
rect 22085 175 22095 205
rect 22045 155 22095 175
rect 22045 125 22055 155
rect 22085 125 22095 155
rect 22045 115 22095 125
rect 22130 205 22180 215
rect 22130 175 22140 205
rect 22170 175 22180 205
rect 22130 155 22180 175
rect 22130 125 22140 155
rect 22170 125 22180 155
rect 22130 115 22180 125
rect 22215 205 22265 215
rect 22215 175 22225 205
rect 22255 175 22265 205
rect 22215 155 22265 175
rect 22215 125 22225 155
rect 22255 125 22265 155
rect 22215 115 22265 125
rect 22300 205 22350 215
rect 22300 175 22310 205
rect 22340 175 22350 205
rect 22300 155 22350 175
rect 22300 125 22310 155
rect 22340 125 22350 155
rect 22300 115 22350 125
rect 22385 205 22435 215
rect 22385 175 22395 205
rect 22425 175 22435 205
rect 22385 155 22435 175
rect 22385 125 22395 155
rect 22425 125 22435 155
rect 22385 115 22435 125
rect 22470 205 22520 215
rect 22470 175 22480 205
rect 22510 175 22520 205
rect 22470 155 22520 175
rect 22470 125 22480 155
rect 22510 125 22520 155
rect 22470 115 22520 125
rect 22555 205 22605 215
rect 22555 175 22565 205
rect 22595 175 22605 205
rect 22555 155 22605 175
rect 22555 125 22565 155
rect 22595 125 22605 155
rect 22555 115 22605 125
rect 22640 205 22690 215
rect 22640 175 22650 205
rect 22680 175 22690 205
rect 22640 155 22690 175
rect 22640 125 22650 155
rect 22680 125 22690 155
rect 22640 115 22690 125
rect 22725 205 22775 215
rect 22725 175 22735 205
rect 22765 175 22775 205
rect 22725 155 22775 175
rect 22725 125 22735 155
rect 22765 125 22775 155
rect 22725 115 22775 125
rect 22810 205 22860 215
rect 22810 175 22820 205
rect 22850 175 22860 205
rect 22810 155 22860 175
rect 22810 125 22820 155
rect 22850 125 22860 155
rect 22810 115 22860 125
rect 22895 205 22945 215
rect 22895 175 22905 205
rect 22935 175 22945 205
rect 22895 155 22945 175
rect 22895 125 22905 155
rect 22935 125 22945 155
rect 22895 115 22945 125
rect 22980 205 23030 215
rect 22980 175 22990 205
rect 23020 175 23030 205
rect 22980 155 23030 175
rect 22980 125 22990 155
rect 23020 125 23030 155
rect 22980 115 23030 125
rect 23065 205 23115 215
rect 23065 175 23075 205
rect 23105 175 23115 205
rect 23065 155 23115 175
rect 23065 125 23075 155
rect 23105 125 23115 155
rect 23065 115 23115 125
rect 23150 205 23200 215
rect 23150 175 23160 205
rect 23190 175 23200 205
rect 23150 155 23200 175
rect 23150 125 23160 155
rect 23190 125 23200 155
rect 23150 115 23200 125
rect 23235 205 23285 215
rect 23235 175 23245 205
rect 23275 175 23285 205
rect 23235 155 23285 175
rect 23235 125 23245 155
rect 23275 125 23285 155
rect 23235 115 23285 125
rect 23320 205 23370 215
rect 23320 175 23330 205
rect 23360 175 23370 205
rect 23320 155 23370 175
rect 23320 125 23330 155
rect 23360 125 23370 155
rect 23320 115 23370 125
rect 23405 205 23455 215
rect 23405 175 23415 205
rect 23445 175 23455 205
rect 23405 155 23455 175
rect 23405 125 23415 155
rect 23445 125 23455 155
rect 23405 115 23455 125
rect 23490 205 23540 215
rect 23490 175 23500 205
rect 23530 175 23540 205
rect 23490 155 23540 175
rect 23490 125 23500 155
rect 23530 125 23540 155
rect 23490 115 23540 125
rect 23575 205 23625 215
rect 23575 175 23585 205
rect 23615 175 23625 205
rect 23575 155 23625 175
rect 23575 125 23585 155
rect 23615 125 23625 155
rect 23575 115 23625 125
rect 23660 205 23710 215
rect 23660 175 23670 205
rect 23700 175 23710 205
rect 23660 155 23710 175
rect 23660 125 23670 155
rect 23700 125 23710 155
rect 23660 115 23710 125
rect 23745 205 23795 215
rect 23745 175 23755 205
rect 23785 175 23795 205
rect 23745 155 23795 175
rect 23745 125 23755 155
rect 23785 125 23795 155
rect 23745 115 23795 125
rect 23830 205 23880 215
rect 23830 175 23840 205
rect 23870 175 23880 205
rect 23830 155 23880 175
rect 23830 125 23840 155
rect 23870 125 23880 155
rect 23830 115 23880 125
rect 23915 205 23965 215
rect 23915 175 23925 205
rect 23955 175 23965 205
rect 23915 155 23965 175
rect 23915 125 23925 155
rect 23955 125 23965 155
rect 23915 115 23965 125
rect 24000 205 24050 215
rect 24000 175 24010 205
rect 24040 175 24050 205
rect 24000 155 24050 175
rect 24000 125 24010 155
rect 24040 125 24050 155
rect 24000 115 24050 125
rect 24085 205 24135 215
rect 24085 175 24095 205
rect 24125 175 24135 205
rect 24085 155 24135 175
rect 24085 125 24095 155
rect 24125 125 24135 155
rect 24085 115 24135 125
rect 24170 205 24220 215
rect 24170 175 24180 205
rect 24210 175 24220 205
rect 24170 155 24220 175
rect 24170 125 24180 155
rect 24210 125 24220 155
rect 24170 115 24220 125
rect 24255 205 24305 215
rect 24255 175 24265 205
rect 24295 175 24305 205
rect 24255 155 24305 175
rect 24255 125 24265 155
rect 24295 125 24305 155
rect 24255 115 24305 125
rect 24340 205 24390 215
rect 24340 175 24350 205
rect 24380 175 24390 205
rect 24340 155 24390 175
rect 24340 125 24350 155
rect 24380 125 24390 155
rect 24340 115 24390 125
rect 24425 205 24475 215
rect 24425 175 24435 205
rect 24465 175 24475 205
rect 24425 155 24475 175
rect 24425 125 24435 155
rect 24465 125 24475 155
rect 24425 115 24475 125
rect 24510 205 24560 215
rect 24510 175 24520 205
rect 24550 175 24560 205
rect 24510 155 24560 175
rect 24510 125 24520 155
rect 24550 125 24560 155
rect 24510 115 24560 125
rect 24595 205 24645 215
rect 24595 175 24605 205
rect 24635 175 24645 205
rect 24595 155 24645 175
rect 24595 125 24605 155
rect 24635 125 24645 155
rect 24595 115 24645 125
rect 24680 205 24730 215
rect 24680 175 24690 205
rect 24720 175 24730 205
rect 24680 155 24730 175
rect 24680 125 24690 155
rect 24720 125 24730 155
rect 24680 115 24730 125
rect 24765 205 24815 215
rect 24765 175 24775 205
rect 24805 175 24815 205
rect 24765 155 24815 175
rect 24765 125 24775 155
rect 24805 125 24815 155
rect 24765 115 24815 125
rect 24850 205 24900 215
rect 24850 175 24860 205
rect 24890 175 24900 205
rect 24850 155 24900 175
rect 24850 125 24860 155
rect 24890 125 24900 155
rect 24850 115 24900 125
rect 24935 205 24985 215
rect 24935 175 24945 205
rect 24975 175 24985 205
rect 24935 155 24985 175
rect 24935 125 24945 155
rect 24975 125 24985 155
rect 24935 115 24985 125
rect 25020 205 25070 215
rect 25020 175 25030 205
rect 25060 175 25070 205
rect 25020 155 25070 175
rect 25020 125 25030 155
rect 25060 125 25070 155
rect 25020 115 25070 125
rect 25105 205 25155 215
rect 25105 175 25115 205
rect 25145 175 25155 205
rect 25105 155 25155 175
rect 25105 125 25115 155
rect 25145 125 25155 155
rect 25105 115 25155 125
rect 25190 205 25240 215
rect 25190 175 25200 205
rect 25230 175 25240 205
rect 25190 155 25240 175
rect 25190 125 25200 155
rect 25230 125 25240 155
rect 25190 115 25240 125
rect 25275 205 25325 215
rect 25275 175 25285 205
rect 25315 175 25325 205
rect 25275 155 25325 175
rect 25275 125 25285 155
rect 25315 125 25325 155
rect 25275 115 25325 125
rect 25360 205 25410 215
rect 25360 175 25370 205
rect 25400 175 25410 205
rect 25360 155 25410 175
rect 25360 125 25370 155
rect 25400 125 25410 155
rect 25360 115 25410 125
rect 25445 205 25495 215
rect 25445 175 25455 205
rect 25485 175 25495 205
rect 25445 155 25495 175
rect 25445 125 25455 155
rect 25485 125 25495 155
rect 25445 115 25495 125
rect 25530 205 25580 215
rect 25530 175 25540 205
rect 25570 175 25580 205
rect 25530 155 25580 175
rect 25530 125 25540 155
rect 25570 125 25580 155
rect 25530 115 25580 125
rect 25615 205 25665 215
rect 25615 175 25625 205
rect 25655 175 25665 205
rect 25615 155 25665 175
rect 25615 125 25625 155
rect 25655 125 25665 155
rect 25615 115 25665 125
rect 25700 205 25750 215
rect 25700 175 25710 205
rect 25740 175 25750 205
rect 25700 155 25750 175
rect 25700 125 25710 155
rect 25740 125 25750 155
rect 25700 115 25750 125
rect 25785 205 25835 215
rect 25785 175 25795 205
rect 25825 175 25835 205
rect 25785 155 25835 175
rect 25785 125 25795 155
rect 25825 125 25835 155
rect 25785 115 25835 125
rect 25870 205 25920 215
rect 25870 175 25880 205
rect 25910 175 25920 205
rect 25870 155 25920 175
rect 25870 125 25880 155
rect 25910 125 25920 155
rect 25870 115 25920 125
rect 25955 205 26005 215
rect 25955 175 25965 205
rect 25995 175 26005 205
rect 25955 155 26005 175
rect 25955 125 25965 155
rect 25995 125 26005 155
rect 25955 115 26005 125
rect 26040 205 26090 215
rect 26040 175 26050 205
rect 26080 175 26090 205
rect 26040 155 26090 175
rect 26040 125 26050 155
rect 26080 125 26090 155
rect 26040 115 26090 125
rect 26125 205 26175 215
rect 26125 175 26135 205
rect 26165 175 26175 205
rect 26125 155 26175 175
rect 26125 125 26135 155
rect 26165 125 26175 155
rect 26125 115 26175 125
rect 26210 205 26260 215
rect 26210 175 26220 205
rect 26250 175 26260 205
rect 26210 155 26260 175
rect 26210 125 26220 155
rect 26250 125 26260 155
rect 26210 115 26260 125
rect 26295 205 26345 215
rect 26295 175 26305 205
rect 26335 175 26345 205
rect 26295 155 26345 175
rect 26295 125 26305 155
rect 26335 125 26345 155
rect 26295 115 26345 125
rect 26380 205 26430 215
rect 26380 175 26390 205
rect 26420 175 26430 205
rect 26380 155 26430 175
rect 26380 125 26390 155
rect 26420 125 26430 155
rect 26380 115 26430 125
rect 26465 205 26515 215
rect 26465 175 26475 205
rect 26505 175 26515 205
rect 26465 155 26515 175
rect 26465 125 26475 155
rect 26505 125 26515 155
rect 26465 115 26515 125
rect 26550 205 26600 215
rect 26550 175 26560 205
rect 26590 175 26600 205
rect 26550 155 26600 175
rect 26550 125 26560 155
rect 26590 125 26600 155
rect 26550 115 26600 125
rect 26635 205 26685 215
rect 26635 175 26645 205
rect 26675 175 26685 205
rect 26635 155 26685 175
rect 26635 125 26645 155
rect 26675 125 26685 155
rect 26635 115 26685 125
rect 26720 205 26770 215
rect 26720 175 26730 205
rect 26760 175 26770 205
rect 26720 155 26770 175
rect 26720 125 26730 155
rect 26760 125 26770 155
rect 26720 115 26770 125
rect 26805 205 26855 215
rect 26805 175 26815 205
rect 26845 175 26855 205
rect 26805 155 26855 175
rect 26805 125 26815 155
rect 26845 125 26855 155
rect 26805 115 26855 125
rect 26890 205 26940 215
rect 26890 175 26900 205
rect 26930 175 26940 205
rect 26890 155 26940 175
rect 26890 125 26900 155
rect 26930 125 26940 155
rect 26890 115 26940 125
rect 26975 205 27025 215
rect 26975 175 26985 205
rect 27015 175 27025 205
rect 26975 155 27025 175
rect 26975 125 26985 155
rect 27015 125 27025 155
rect 26975 115 27025 125
rect 27060 205 27110 215
rect 27060 175 27070 205
rect 27100 175 27110 205
rect 27060 155 27110 175
rect 27060 125 27070 155
rect 27100 125 27110 155
rect 27060 115 27110 125
rect 27145 205 27195 215
rect 27145 175 27155 205
rect 27185 175 27195 205
rect 27145 155 27195 175
rect 27145 125 27155 155
rect 27185 125 27195 155
rect 27145 115 27195 125
rect 27230 205 27280 215
rect 27230 175 27240 205
rect 27270 175 27280 205
rect 27230 155 27280 175
rect 27230 125 27240 155
rect 27270 125 27280 155
rect 27230 115 27280 125
rect 27315 205 27365 215
rect 27315 175 27325 205
rect 27355 175 27365 205
rect 27315 155 27365 175
rect 27315 125 27325 155
rect 27355 125 27365 155
rect 27315 115 27365 125
rect 27400 205 27450 215
rect 27400 175 27410 205
rect 27440 175 27450 205
rect 27400 155 27450 175
rect 27400 125 27410 155
rect 27440 125 27450 155
rect 27400 115 27450 125
rect 27485 205 27535 215
rect 27485 175 27495 205
rect 27525 175 27535 205
rect 27485 155 27535 175
rect 27485 125 27495 155
rect 27525 125 27535 155
rect 27485 115 27535 125
rect 27570 205 27620 215
rect 27570 175 27580 205
rect 27610 175 27620 205
rect 27570 155 27620 175
rect 27570 125 27580 155
rect 27610 125 27620 155
rect 27570 115 27620 125
rect 27655 205 27705 215
rect 27655 175 27665 205
rect 27695 175 27705 205
rect 27655 155 27705 175
rect 27655 125 27665 155
rect 27695 125 27705 155
rect 27655 115 27705 125
rect 27740 205 27790 215
rect 27740 175 27750 205
rect 27780 175 27790 205
rect 27740 155 27790 175
rect 27740 125 27750 155
rect 27780 125 27790 155
rect 27740 115 27790 125
rect 27825 205 27875 215
rect 27825 175 27835 205
rect 27865 175 27875 205
rect 27825 155 27875 175
rect 27825 125 27835 155
rect 27865 125 27875 155
rect 27825 115 27875 125
rect 27910 205 27960 215
rect 27910 175 27920 205
rect 27950 175 27960 205
rect 27910 155 27960 175
rect 27910 125 27920 155
rect 27950 125 27960 155
rect 27910 115 27960 125
rect 27995 205 28045 215
rect 27995 175 28005 205
rect 28035 175 28045 205
rect 27995 155 28045 175
rect 27995 125 28005 155
rect 28035 125 28045 155
rect 27995 115 28045 125
rect 28080 205 28130 215
rect 28080 175 28090 205
rect 28120 175 28130 205
rect 28080 155 28130 175
rect 28080 125 28090 155
rect 28120 125 28130 155
rect 28080 115 28130 125
rect 28165 205 28215 215
rect 28165 175 28175 205
rect 28205 175 28215 205
rect 28165 155 28215 175
rect 28165 125 28175 155
rect 28205 125 28215 155
rect 28165 115 28215 125
rect 28250 205 28300 215
rect 28250 175 28260 205
rect 28290 175 28300 205
rect 28250 155 28300 175
rect 28250 125 28260 155
rect 28290 125 28300 155
rect 28250 115 28300 125
rect 28335 205 28385 215
rect 28335 175 28345 205
rect 28375 175 28385 205
rect 28335 155 28385 175
rect 28335 125 28345 155
rect 28375 125 28385 155
rect 28335 115 28385 125
rect 28420 205 28470 215
rect 28420 175 28430 205
rect 28460 175 28470 205
rect 28420 155 28470 175
rect 28420 125 28430 155
rect 28460 125 28470 155
rect 28420 115 28470 125
rect 28505 205 28555 215
rect 28505 175 28515 205
rect 28545 175 28555 205
rect 28505 155 28555 175
rect 28505 125 28515 155
rect 28545 125 28555 155
rect 28505 115 28555 125
rect 28590 205 28640 215
rect 28590 175 28600 205
rect 28630 175 28640 205
rect 28590 155 28640 175
rect 28590 125 28600 155
rect 28630 125 28640 155
rect 28590 115 28640 125
rect 28675 205 28725 215
rect 28675 175 28685 205
rect 28715 175 28725 205
rect 28675 155 28725 175
rect 28675 125 28685 155
rect 28715 125 28725 155
rect 28675 115 28725 125
rect 28760 205 28810 215
rect 28760 175 28770 205
rect 28800 175 28810 205
rect 28760 155 28810 175
rect 28760 125 28770 155
rect 28800 125 28810 155
rect 28760 115 28810 125
rect 28845 205 28895 215
rect 28845 175 28855 205
rect 28885 175 28895 205
rect 28845 155 28895 175
rect 28845 125 28855 155
rect 28885 125 28895 155
rect 28845 115 28895 125
rect 28930 205 28980 215
rect 28930 175 28940 205
rect 28970 175 28980 205
rect 28930 155 28980 175
rect 28930 125 28940 155
rect 28970 125 28980 155
rect 28930 115 28980 125
rect 29015 205 29065 215
rect 29015 175 29025 205
rect 29055 175 29065 205
rect 29015 155 29065 175
rect 29015 125 29025 155
rect 29055 125 29065 155
rect 29015 115 29065 125
rect 29100 205 29150 215
rect 29100 175 29110 205
rect 29140 175 29150 205
rect 29100 155 29150 175
rect 29100 125 29110 155
rect 29140 125 29150 155
rect 29100 115 29150 125
rect 29185 205 29235 215
rect 29185 175 29195 205
rect 29225 175 29235 205
rect 29185 155 29235 175
rect 29185 125 29195 155
rect 29225 125 29235 155
rect 29185 115 29235 125
rect 29270 205 29320 215
rect 29270 175 29280 205
rect 29310 175 29320 205
rect 29270 155 29320 175
rect 29270 125 29280 155
rect 29310 125 29320 155
rect 29270 115 29320 125
rect 29355 205 29405 215
rect 29355 175 29365 205
rect 29395 175 29405 205
rect 29355 155 29405 175
rect 29355 125 29365 155
rect 29395 125 29405 155
rect 29355 115 29405 125
rect 29440 205 29490 215
rect 29440 175 29450 205
rect 29480 175 29490 205
rect 29440 155 29490 175
rect 29440 125 29450 155
rect 29480 125 29490 155
rect 29440 115 29490 125
rect 29525 205 29575 215
rect 29525 175 29535 205
rect 29565 175 29575 205
rect 29525 155 29575 175
rect 29525 125 29535 155
rect 29565 125 29575 155
rect 29525 115 29575 125
rect 29610 205 29660 215
rect 29610 175 29620 205
rect 29650 175 29660 205
rect 29610 155 29660 175
rect 29610 125 29620 155
rect 29650 125 29660 155
rect 29610 115 29660 125
rect 25 55 75 65
rect 25 15 35 55
rect 65 15 75 55
rect 25 5 75 15
rect 215 40 265 50
rect 215 10 225 40
rect 255 10 265 40
rect 215 0 265 10
rect 300 40 350 50
rect 300 10 310 40
rect 340 10 350 40
rect 300 0 350 10
rect 385 40 435 50
rect 385 10 395 40
rect 425 10 435 40
rect 385 0 435 10
rect 470 40 520 50
rect 470 10 480 40
rect 510 10 520 40
rect 470 0 520 10
rect 555 40 605 50
rect 555 10 565 40
rect 595 10 605 40
rect 555 0 605 10
rect 750 40 800 50
rect 750 10 760 40
rect 790 10 800 40
rect 750 0 800 10
rect 835 40 885 50
rect 835 10 845 40
rect 875 10 885 40
rect 835 0 885 10
rect 920 40 970 50
rect 920 10 930 40
rect 960 10 970 40
rect 920 0 970 10
rect 1005 40 1055 50
rect 1005 10 1015 40
rect 1045 10 1055 40
rect 1005 0 1055 10
rect 1090 40 1140 50
rect 1090 10 1100 40
rect 1130 10 1140 40
rect 1090 0 1140 10
rect 1175 40 1225 50
rect 1175 10 1185 40
rect 1215 10 1225 40
rect 1175 0 1225 10
rect 1260 40 1310 50
rect 1260 10 1270 40
rect 1300 10 1310 40
rect 1260 0 1310 10
rect 1345 40 1395 50
rect 1345 10 1355 40
rect 1385 10 1395 40
rect 1345 0 1395 10
rect 1430 40 1480 50
rect 1430 10 1440 40
rect 1470 10 1480 40
rect 1430 0 1480 10
rect 1515 40 1565 50
rect 1515 10 1525 40
rect 1555 10 1565 40
rect 1515 0 1565 10
rect 1600 40 1650 50
rect 1600 10 1610 40
rect 1640 10 1650 40
rect 1600 0 1650 10
rect 1685 40 1735 50
rect 1685 10 1695 40
rect 1725 10 1735 40
rect 1685 0 1735 10
rect 1770 40 1820 50
rect 1770 10 1780 40
rect 1810 10 1820 40
rect 1770 0 1820 10
rect 1855 40 1905 50
rect 1855 10 1865 40
rect 1895 10 1905 40
rect 1855 0 1905 10
rect 1940 40 1990 50
rect 1940 10 1950 40
rect 1980 10 1990 40
rect 1940 0 1990 10
rect 2025 40 2075 50
rect 2025 10 2035 40
rect 2065 10 2075 40
rect 2025 0 2075 10
rect 2110 40 2160 50
rect 2110 10 2120 40
rect 2150 10 2160 40
rect 2110 0 2160 10
rect 2260 40 2310 50
rect 2260 10 2270 40
rect 2300 10 2310 40
rect 2260 0 2310 10
rect 2345 40 2395 50
rect 2345 10 2355 40
rect 2385 10 2395 40
rect 2345 0 2395 10
rect 2430 40 2480 50
rect 2430 10 2440 40
rect 2470 10 2480 40
rect 2430 0 2480 10
rect 2515 40 2565 50
rect 2515 10 2525 40
rect 2555 10 2565 40
rect 2515 0 2565 10
rect 2600 40 2650 50
rect 2600 10 2610 40
rect 2640 10 2650 40
rect 2600 0 2650 10
rect 2685 40 2735 50
rect 2685 10 2695 40
rect 2725 10 2735 40
rect 2685 0 2735 10
rect 2770 40 2820 50
rect 2770 10 2780 40
rect 2810 10 2820 40
rect 2770 0 2820 10
rect 2855 40 2905 50
rect 2855 10 2865 40
rect 2895 10 2905 40
rect 2855 0 2905 10
rect 2940 40 2990 50
rect 2940 10 2950 40
rect 2980 10 2990 40
rect 2940 0 2990 10
rect 3025 40 3075 50
rect 3025 10 3035 40
rect 3065 10 3075 40
rect 3025 0 3075 10
rect 3110 40 3160 50
rect 3110 10 3120 40
rect 3150 10 3160 40
rect 3110 0 3160 10
rect 3195 40 3245 50
rect 3195 10 3205 40
rect 3235 10 3245 40
rect 3195 0 3245 10
rect 3280 40 3330 50
rect 3280 10 3290 40
rect 3320 10 3330 40
rect 3280 0 3330 10
rect 3365 40 3415 50
rect 3365 10 3375 40
rect 3405 10 3415 40
rect 3365 0 3415 10
rect 3450 40 3500 50
rect 3450 10 3460 40
rect 3490 10 3500 40
rect 3450 0 3500 10
rect 3535 40 3585 50
rect 3535 10 3545 40
rect 3575 10 3585 40
rect 3535 0 3585 10
rect 3620 40 3670 50
rect 3620 10 3630 40
rect 3660 10 3670 40
rect 3620 0 3670 10
rect 3705 40 3755 50
rect 3705 10 3715 40
rect 3745 10 3755 40
rect 3705 0 3755 10
rect 3790 40 3840 50
rect 3790 10 3800 40
rect 3830 10 3840 40
rect 3790 0 3840 10
rect 3875 40 3925 50
rect 3875 10 3885 40
rect 3915 10 3925 40
rect 3875 0 3925 10
rect 3960 40 4010 50
rect 3960 10 3970 40
rect 4000 10 4010 40
rect 3960 0 4010 10
rect 4045 40 4095 50
rect 4045 10 4055 40
rect 4085 10 4095 40
rect 4045 0 4095 10
rect 4130 40 4180 50
rect 4130 10 4140 40
rect 4170 10 4180 40
rect 4130 0 4180 10
rect 4215 40 4265 50
rect 4215 10 4225 40
rect 4255 10 4265 40
rect 4215 0 4265 10
rect 4300 40 4350 50
rect 4300 10 4310 40
rect 4340 10 4350 40
rect 4300 0 4350 10
rect 4385 40 4435 50
rect 4385 10 4395 40
rect 4425 10 4435 40
rect 4385 0 4435 10
rect 4470 40 4520 50
rect 4470 10 4480 40
rect 4510 10 4520 40
rect 4470 0 4520 10
rect 4555 40 4605 50
rect 4555 10 4565 40
rect 4595 10 4605 40
rect 4555 0 4605 10
rect 4640 40 4690 50
rect 4640 10 4650 40
rect 4680 10 4690 40
rect 4640 0 4690 10
rect 4725 40 4775 50
rect 4725 10 4735 40
rect 4765 10 4775 40
rect 4725 0 4775 10
rect 4810 40 4860 50
rect 4810 10 4820 40
rect 4850 10 4860 40
rect 4810 0 4860 10
rect 4895 40 4945 50
rect 4895 10 4905 40
rect 4935 10 4945 40
rect 4895 0 4945 10
rect 4980 40 5030 50
rect 4980 10 4990 40
rect 5020 10 5030 40
rect 4980 0 5030 10
rect 5065 40 5115 50
rect 5065 10 5075 40
rect 5105 10 5115 40
rect 5065 0 5115 10
rect 5150 40 5200 50
rect 5150 10 5160 40
rect 5190 10 5200 40
rect 5150 0 5200 10
rect 5235 40 5285 50
rect 5235 10 5245 40
rect 5275 10 5285 40
rect 5235 0 5285 10
rect 5320 40 5370 50
rect 5320 10 5330 40
rect 5360 10 5370 40
rect 5320 0 5370 10
rect 5405 40 5455 50
rect 5405 10 5415 40
rect 5445 10 5455 40
rect 5405 0 5455 10
rect 5490 40 5540 50
rect 5490 10 5500 40
rect 5530 10 5540 40
rect 5490 0 5540 10
rect 5575 40 5625 50
rect 5575 10 5585 40
rect 5615 10 5625 40
rect 5575 0 5625 10
rect 5660 40 5710 50
rect 5660 10 5670 40
rect 5700 10 5710 40
rect 5660 0 5710 10
rect 5745 40 5795 50
rect 5745 10 5755 40
rect 5785 10 5795 40
rect 5745 0 5795 10
rect 5830 40 5880 50
rect 5830 10 5840 40
rect 5870 10 5880 40
rect 5830 0 5880 10
rect 5915 40 5965 50
rect 5915 10 5925 40
rect 5955 10 5965 40
rect 5915 0 5965 10
rect 6000 40 6050 50
rect 6000 10 6010 40
rect 6040 10 6050 40
rect 6000 0 6050 10
rect 6085 40 6135 50
rect 6085 10 6095 40
rect 6125 10 6135 40
rect 6085 0 6135 10
rect 6170 40 6220 50
rect 6170 10 6180 40
rect 6210 10 6220 40
rect 6170 0 6220 10
rect 6255 40 6305 50
rect 6255 10 6265 40
rect 6295 10 6305 40
rect 6255 0 6305 10
rect 6340 40 6390 50
rect 6340 10 6350 40
rect 6380 10 6390 40
rect 6340 0 6390 10
rect 6425 40 6475 50
rect 6425 10 6435 40
rect 6465 10 6475 40
rect 6425 0 6475 10
rect 6510 40 6560 50
rect 6510 10 6520 40
rect 6550 10 6560 40
rect 6510 0 6560 10
rect 6595 40 6645 50
rect 6595 10 6605 40
rect 6635 10 6645 40
rect 6595 0 6645 10
rect 6680 40 6730 50
rect 6680 10 6690 40
rect 6720 10 6730 40
rect 6680 0 6730 10
rect 6765 40 6815 50
rect 6765 10 6775 40
rect 6805 10 6815 40
rect 6765 0 6815 10
rect 6850 40 6900 50
rect 6850 10 6860 40
rect 6890 10 6900 40
rect 6850 0 6900 10
rect 6935 40 6985 50
rect 6935 10 6945 40
rect 6975 10 6985 40
rect 6935 0 6985 10
rect 7020 40 7070 50
rect 7020 10 7030 40
rect 7060 10 7070 40
rect 7020 0 7070 10
rect 7105 40 7155 50
rect 7105 10 7115 40
rect 7145 10 7155 40
rect 7105 0 7155 10
rect 7190 40 7240 50
rect 7190 10 7200 40
rect 7230 10 7240 40
rect 7190 0 7240 10
rect 7275 40 7325 50
rect 7275 10 7285 40
rect 7315 10 7325 40
rect 7275 0 7325 10
rect 7360 40 7410 50
rect 7360 10 7370 40
rect 7400 10 7410 40
rect 7360 0 7410 10
rect 7445 40 7495 50
rect 7445 10 7455 40
rect 7485 10 7495 40
rect 7445 0 7495 10
rect 7530 40 7580 50
rect 7530 10 7540 40
rect 7570 10 7580 40
rect 7530 0 7580 10
rect 7615 40 7665 50
rect 7615 10 7625 40
rect 7655 10 7665 40
rect 7615 0 7665 10
rect 7700 40 7750 50
rect 7700 10 7710 40
rect 7740 10 7750 40
rect 7700 0 7750 10
rect 7850 40 7900 50
rect 7850 10 7860 40
rect 7890 10 7900 40
rect 7850 0 7900 10
rect 7935 40 7985 50
rect 7935 10 7945 40
rect 7975 10 7985 40
rect 7935 0 7985 10
rect 8020 40 8070 50
rect 8020 10 8030 40
rect 8060 10 8070 40
rect 8020 0 8070 10
rect 8105 40 8155 50
rect 8105 10 8115 40
rect 8145 10 8155 40
rect 8105 0 8155 10
rect 8190 40 8240 50
rect 8190 10 8200 40
rect 8230 10 8240 40
rect 8190 0 8240 10
rect 8275 40 8325 50
rect 8275 10 8285 40
rect 8315 10 8325 40
rect 8275 0 8325 10
rect 8360 40 8410 50
rect 8360 10 8370 40
rect 8400 10 8410 40
rect 8360 0 8410 10
rect 8445 40 8495 50
rect 8445 10 8455 40
rect 8485 10 8495 40
rect 8445 0 8495 10
rect 8530 40 8580 50
rect 8530 10 8540 40
rect 8570 10 8580 40
rect 8530 0 8580 10
rect 8615 40 8665 50
rect 8615 10 8625 40
rect 8655 10 8665 40
rect 8615 0 8665 10
rect 8700 40 8750 50
rect 8700 10 8710 40
rect 8740 10 8750 40
rect 8700 0 8750 10
rect 8785 40 8835 50
rect 8785 10 8795 40
rect 8825 10 8835 40
rect 8785 0 8835 10
rect 8870 40 8920 50
rect 8870 10 8880 40
rect 8910 10 8920 40
rect 8870 0 8920 10
rect 8955 40 9005 50
rect 8955 10 8965 40
rect 8995 10 9005 40
rect 8955 0 9005 10
rect 9040 40 9090 50
rect 9040 10 9050 40
rect 9080 10 9090 40
rect 9040 0 9090 10
rect 9125 40 9175 50
rect 9125 10 9135 40
rect 9165 10 9175 40
rect 9125 0 9175 10
rect 9210 40 9260 50
rect 9210 10 9220 40
rect 9250 10 9260 40
rect 9210 0 9260 10
rect 9295 40 9345 50
rect 9295 10 9305 40
rect 9335 10 9345 40
rect 9295 0 9345 10
rect 9380 40 9430 50
rect 9380 10 9390 40
rect 9420 10 9430 40
rect 9380 0 9430 10
rect 9465 40 9515 50
rect 9465 10 9475 40
rect 9505 10 9515 40
rect 9465 0 9515 10
rect 9550 40 9600 50
rect 9550 10 9560 40
rect 9590 10 9600 40
rect 9550 0 9600 10
rect 9635 40 9685 50
rect 9635 10 9645 40
rect 9675 10 9685 40
rect 9635 0 9685 10
rect 9720 40 9770 50
rect 9720 10 9730 40
rect 9760 10 9770 40
rect 9720 0 9770 10
rect 9805 40 9855 50
rect 9805 10 9815 40
rect 9845 10 9855 40
rect 9805 0 9855 10
rect 9890 40 9940 50
rect 9890 10 9900 40
rect 9930 10 9940 40
rect 9890 0 9940 10
rect 9975 40 10025 50
rect 9975 10 9985 40
rect 10015 10 10025 40
rect 9975 0 10025 10
rect 10060 40 10110 50
rect 10060 10 10070 40
rect 10100 10 10110 40
rect 10060 0 10110 10
rect 10145 40 10195 50
rect 10145 10 10155 40
rect 10185 10 10195 40
rect 10145 0 10195 10
rect 10230 40 10280 50
rect 10230 10 10240 40
rect 10270 10 10280 40
rect 10230 0 10280 10
rect 10315 40 10365 50
rect 10315 10 10325 40
rect 10355 10 10365 40
rect 10315 0 10365 10
rect 10400 40 10450 50
rect 10400 10 10410 40
rect 10440 10 10450 40
rect 10400 0 10450 10
rect 10485 40 10535 50
rect 10485 10 10495 40
rect 10525 10 10535 40
rect 10485 0 10535 10
rect 10570 40 10620 50
rect 10570 10 10580 40
rect 10610 10 10620 40
rect 10570 0 10620 10
rect 10655 40 10705 50
rect 10655 10 10665 40
rect 10695 10 10705 40
rect 10655 0 10705 10
rect 10740 40 10790 50
rect 10740 10 10750 40
rect 10780 10 10790 40
rect 10740 0 10790 10
rect 10825 40 10875 50
rect 10825 10 10835 40
rect 10865 10 10875 40
rect 10825 0 10875 10
rect 10910 40 10960 50
rect 10910 10 10920 40
rect 10950 10 10960 40
rect 10910 0 10960 10
rect 10995 40 11045 50
rect 10995 10 11005 40
rect 11035 10 11045 40
rect 10995 0 11045 10
rect 11080 40 11130 50
rect 11080 10 11090 40
rect 11120 10 11130 40
rect 11080 0 11130 10
rect 11165 40 11215 50
rect 11165 10 11175 40
rect 11205 10 11215 40
rect 11165 0 11215 10
rect 11250 40 11300 50
rect 11250 10 11260 40
rect 11290 10 11300 40
rect 11250 0 11300 10
rect 11335 40 11385 50
rect 11335 10 11345 40
rect 11375 10 11385 40
rect 11335 0 11385 10
rect 11420 40 11470 50
rect 11420 10 11430 40
rect 11460 10 11470 40
rect 11420 0 11470 10
rect 11505 40 11555 50
rect 11505 10 11515 40
rect 11545 10 11555 40
rect 11505 0 11555 10
rect 11590 40 11640 50
rect 11590 10 11600 40
rect 11630 10 11640 40
rect 11590 0 11640 10
rect 11675 40 11725 50
rect 11675 10 11685 40
rect 11715 10 11725 40
rect 11675 0 11725 10
rect 11760 40 11810 50
rect 11760 10 11770 40
rect 11800 10 11810 40
rect 11760 0 11810 10
rect 11845 40 11895 50
rect 11845 10 11855 40
rect 11885 10 11895 40
rect 11845 0 11895 10
rect 11930 40 11980 50
rect 11930 10 11940 40
rect 11970 10 11980 40
rect 11930 0 11980 10
rect 12015 40 12065 50
rect 12015 10 12025 40
rect 12055 10 12065 40
rect 12015 0 12065 10
rect 12100 40 12150 50
rect 12100 10 12110 40
rect 12140 10 12150 40
rect 12100 0 12150 10
rect 12185 40 12235 50
rect 12185 10 12195 40
rect 12225 10 12235 40
rect 12185 0 12235 10
rect 12270 40 12320 50
rect 12270 10 12280 40
rect 12310 10 12320 40
rect 12270 0 12320 10
rect 12355 40 12405 50
rect 12355 10 12365 40
rect 12395 10 12405 40
rect 12355 0 12405 10
rect 12440 40 12490 50
rect 12440 10 12450 40
rect 12480 10 12490 40
rect 12440 0 12490 10
rect 12525 40 12575 50
rect 12525 10 12535 40
rect 12565 10 12575 40
rect 12525 0 12575 10
rect 12610 40 12660 50
rect 12610 10 12620 40
rect 12650 10 12660 40
rect 12610 0 12660 10
rect 12695 40 12745 50
rect 12695 10 12705 40
rect 12735 10 12745 40
rect 12695 0 12745 10
rect 12780 40 12830 50
rect 12780 10 12790 40
rect 12820 10 12830 40
rect 12780 0 12830 10
rect 12865 40 12915 50
rect 12865 10 12875 40
rect 12905 10 12915 40
rect 12865 0 12915 10
rect 12950 40 13000 50
rect 12950 10 12960 40
rect 12990 10 13000 40
rect 12950 0 13000 10
rect 13035 40 13085 50
rect 13035 10 13045 40
rect 13075 10 13085 40
rect 13035 0 13085 10
rect 13120 40 13170 50
rect 13120 10 13130 40
rect 13160 10 13170 40
rect 13120 0 13170 10
rect 13205 40 13255 50
rect 13205 10 13215 40
rect 13245 10 13255 40
rect 13205 0 13255 10
rect 13290 40 13340 50
rect 13290 10 13300 40
rect 13330 10 13340 40
rect 13290 0 13340 10
rect 13375 40 13425 50
rect 13375 10 13385 40
rect 13415 10 13425 40
rect 13375 0 13425 10
rect 13460 40 13510 50
rect 13460 10 13470 40
rect 13500 10 13510 40
rect 13460 0 13510 10
rect 13545 40 13595 50
rect 13545 10 13555 40
rect 13585 10 13595 40
rect 13545 0 13595 10
rect 13630 40 13680 50
rect 13630 10 13640 40
rect 13670 10 13680 40
rect 13630 0 13680 10
rect 13715 40 13765 50
rect 13715 10 13725 40
rect 13755 10 13765 40
rect 13715 0 13765 10
rect 13800 40 13850 50
rect 13800 10 13810 40
rect 13840 10 13850 40
rect 13800 0 13850 10
rect 13885 40 13935 50
rect 13885 10 13895 40
rect 13925 10 13935 40
rect 13885 0 13935 10
rect 13970 40 14020 50
rect 13970 10 13980 40
rect 14010 10 14020 40
rect 13970 0 14020 10
rect 14055 40 14105 50
rect 14055 10 14065 40
rect 14095 10 14105 40
rect 14055 0 14105 10
rect 14140 40 14190 50
rect 14140 10 14150 40
rect 14180 10 14190 40
rect 14140 0 14190 10
rect 14225 40 14275 50
rect 14225 10 14235 40
rect 14265 10 14275 40
rect 14225 0 14275 10
rect 14310 40 14360 50
rect 14310 10 14320 40
rect 14350 10 14360 40
rect 14310 0 14360 10
rect 14395 40 14445 50
rect 14395 10 14405 40
rect 14435 10 14445 40
rect 14395 0 14445 10
rect 14480 40 14530 50
rect 14480 10 14490 40
rect 14520 10 14530 40
rect 14480 0 14530 10
rect 14565 40 14615 50
rect 14565 10 14575 40
rect 14605 10 14615 40
rect 14565 0 14615 10
rect 14650 40 14700 50
rect 14650 10 14660 40
rect 14690 10 14700 40
rect 14650 0 14700 10
rect 14735 40 14785 50
rect 14735 10 14745 40
rect 14775 10 14785 40
rect 14735 0 14785 10
rect 14820 40 14870 50
rect 14820 10 14830 40
rect 14860 10 14870 40
rect 14820 0 14870 10
rect 14905 40 14955 50
rect 14905 10 14915 40
rect 14945 10 14955 40
rect 14905 0 14955 10
rect 14990 40 15040 50
rect 14990 10 15000 40
rect 15030 10 15040 40
rect 14990 0 15040 10
rect 15075 40 15125 50
rect 15075 10 15085 40
rect 15115 10 15125 40
rect 15075 0 15125 10
rect 15160 40 15210 50
rect 15160 10 15170 40
rect 15200 10 15210 40
rect 15160 0 15210 10
rect 15245 40 15295 50
rect 15245 10 15255 40
rect 15285 10 15295 40
rect 15245 0 15295 10
rect 15330 40 15380 50
rect 15330 10 15340 40
rect 15370 10 15380 40
rect 15330 0 15380 10
rect 15415 40 15465 50
rect 15415 10 15425 40
rect 15455 10 15465 40
rect 15415 0 15465 10
rect 15500 40 15550 50
rect 15500 10 15510 40
rect 15540 10 15550 40
rect 15500 0 15550 10
rect 15585 40 15635 50
rect 15585 10 15595 40
rect 15625 10 15635 40
rect 15585 0 15635 10
rect 15670 40 15720 50
rect 15670 10 15680 40
rect 15710 10 15720 40
rect 15670 0 15720 10
rect 15755 40 15805 50
rect 15755 10 15765 40
rect 15795 10 15805 40
rect 15755 0 15805 10
rect 15840 40 15890 50
rect 15840 10 15850 40
rect 15880 10 15890 40
rect 15840 0 15890 10
rect 15925 40 15975 50
rect 15925 10 15935 40
rect 15965 10 15975 40
rect 15925 0 15975 10
rect 16010 40 16060 50
rect 16010 10 16020 40
rect 16050 10 16060 40
rect 16010 0 16060 10
rect 16095 40 16145 50
rect 16095 10 16105 40
rect 16135 10 16145 40
rect 16095 0 16145 10
rect 16180 40 16230 50
rect 16180 10 16190 40
rect 16220 10 16230 40
rect 16180 0 16230 10
rect 16265 40 16315 50
rect 16265 10 16275 40
rect 16305 10 16315 40
rect 16265 0 16315 10
rect 16350 40 16400 50
rect 16350 10 16360 40
rect 16390 10 16400 40
rect 16350 0 16400 10
rect 16435 40 16485 50
rect 16435 10 16445 40
rect 16475 10 16485 40
rect 16435 0 16485 10
rect 16520 40 16570 50
rect 16520 10 16530 40
rect 16560 10 16570 40
rect 16520 0 16570 10
rect 16605 40 16655 50
rect 16605 10 16615 40
rect 16645 10 16655 40
rect 16605 0 16655 10
rect 16690 40 16740 50
rect 16690 10 16700 40
rect 16730 10 16740 40
rect 16690 0 16740 10
rect 16775 40 16825 50
rect 16775 10 16785 40
rect 16815 10 16825 40
rect 16775 0 16825 10
rect 16860 40 16910 50
rect 16860 10 16870 40
rect 16900 10 16910 40
rect 16860 0 16910 10
rect 16945 40 16995 50
rect 16945 10 16955 40
rect 16985 10 16995 40
rect 16945 0 16995 10
rect 17030 40 17080 50
rect 17030 10 17040 40
rect 17070 10 17080 40
rect 17030 0 17080 10
rect 17115 40 17165 50
rect 17115 10 17125 40
rect 17155 10 17165 40
rect 17115 0 17165 10
rect 17200 40 17250 50
rect 17200 10 17210 40
rect 17240 10 17250 40
rect 17200 0 17250 10
rect 17285 40 17335 50
rect 17285 10 17295 40
rect 17325 10 17335 40
rect 17285 0 17335 10
rect 17370 40 17420 50
rect 17370 10 17380 40
rect 17410 10 17420 40
rect 17370 0 17420 10
rect 17455 40 17505 50
rect 17455 10 17465 40
rect 17495 10 17505 40
rect 17455 0 17505 10
rect 17540 40 17590 50
rect 17540 10 17550 40
rect 17580 10 17590 40
rect 17540 0 17590 10
rect 17625 40 17675 50
rect 17625 10 17635 40
rect 17665 10 17675 40
rect 17625 0 17675 10
rect 17710 40 17760 50
rect 17710 10 17720 40
rect 17750 10 17760 40
rect 17710 0 17760 10
rect 17795 40 17845 50
rect 17795 10 17805 40
rect 17835 10 17845 40
rect 17795 0 17845 10
rect 17880 40 17930 50
rect 17880 10 17890 40
rect 17920 10 17930 40
rect 17880 0 17930 10
rect 17965 40 18015 50
rect 17965 10 17975 40
rect 18005 10 18015 40
rect 17965 0 18015 10
rect 18050 40 18100 50
rect 18050 10 18060 40
rect 18090 10 18100 40
rect 18050 0 18100 10
rect 18135 40 18185 50
rect 18135 10 18145 40
rect 18175 10 18185 40
rect 18135 0 18185 10
rect 18220 40 18270 50
rect 18220 10 18230 40
rect 18260 10 18270 40
rect 18220 0 18270 10
rect 18305 40 18355 50
rect 18305 10 18315 40
rect 18345 10 18355 40
rect 18305 0 18355 10
rect 18390 40 18440 50
rect 18390 10 18400 40
rect 18430 10 18440 40
rect 18390 0 18440 10
rect 18475 40 18525 50
rect 18475 10 18485 40
rect 18515 10 18525 40
rect 18475 0 18525 10
rect 18560 40 18610 50
rect 18560 10 18570 40
rect 18600 10 18610 40
rect 18560 0 18610 10
rect 18645 40 18695 50
rect 18645 10 18655 40
rect 18685 10 18695 40
rect 18645 0 18695 10
rect 18730 40 18780 50
rect 18730 10 18740 40
rect 18770 10 18780 40
rect 18730 0 18780 10
rect 18815 40 18865 50
rect 18815 10 18825 40
rect 18855 10 18865 40
rect 18815 0 18865 10
rect 18900 40 18950 50
rect 18900 10 18910 40
rect 18940 10 18950 40
rect 18900 0 18950 10
rect 18985 40 19035 50
rect 18985 10 18995 40
rect 19025 10 19035 40
rect 18985 0 19035 10
rect 19070 40 19120 50
rect 19070 10 19080 40
rect 19110 10 19120 40
rect 19070 0 19120 10
rect 19155 40 19205 50
rect 19155 10 19165 40
rect 19195 10 19205 40
rect 19155 0 19205 10
rect 19240 40 19290 50
rect 19240 10 19250 40
rect 19280 10 19290 40
rect 19240 0 19290 10
rect 19325 40 19375 50
rect 19325 10 19335 40
rect 19365 10 19375 40
rect 19325 0 19375 10
rect 19410 40 19460 50
rect 19410 10 19420 40
rect 19450 10 19460 40
rect 19410 0 19460 10
rect 19495 40 19545 50
rect 19495 10 19505 40
rect 19535 10 19545 40
rect 19495 0 19545 10
rect 19580 40 19630 50
rect 19580 10 19590 40
rect 19620 10 19630 40
rect 19580 0 19630 10
rect 19665 40 19715 50
rect 19665 10 19675 40
rect 19705 10 19715 40
rect 19665 0 19715 10
rect 19750 40 19800 50
rect 19750 10 19760 40
rect 19790 10 19800 40
rect 19750 0 19800 10
rect 19835 40 19885 50
rect 19835 10 19845 40
rect 19875 10 19885 40
rect 19835 0 19885 10
rect 19920 40 19970 50
rect 19920 10 19930 40
rect 19960 10 19970 40
rect 19920 0 19970 10
rect 20005 40 20055 50
rect 20005 10 20015 40
rect 20045 10 20055 40
rect 20005 0 20055 10
rect 20090 40 20140 50
rect 20090 10 20100 40
rect 20130 10 20140 40
rect 20090 0 20140 10
rect 20175 40 20225 50
rect 20175 10 20185 40
rect 20215 10 20225 40
rect 20175 0 20225 10
rect 20260 40 20310 50
rect 20260 10 20270 40
rect 20300 10 20310 40
rect 20260 0 20310 10
rect 20345 40 20395 50
rect 20345 10 20355 40
rect 20385 10 20395 40
rect 20345 0 20395 10
rect 20430 40 20480 50
rect 20430 10 20440 40
rect 20470 10 20480 40
rect 20430 0 20480 10
rect 20515 40 20565 50
rect 20515 10 20525 40
rect 20555 10 20565 40
rect 20515 0 20565 10
rect 20600 40 20650 50
rect 20600 10 20610 40
rect 20640 10 20650 40
rect 20600 0 20650 10
rect 20685 40 20735 50
rect 20685 10 20695 40
rect 20725 10 20735 40
rect 20685 0 20735 10
rect 20770 40 20820 50
rect 20770 10 20780 40
rect 20810 10 20820 40
rect 20770 0 20820 10
rect 20855 40 20905 50
rect 20855 10 20865 40
rect 20895 10 20905 40
rect 20855 0 20905 10
rect 20940 40 20990 50
rect 20940 10 20950 40
rect 20980 10 20990 40
rect 20940 0 20990 10
rect 21025 40 21075 50
rect 21025 10 21035 40
rect 21065 10 21075 40
rect 21025 0 21075 10
rect 21110 40 21160 50
rect 21110 10 21120 40
rect 21150 10 21160 40
rect 21110 0 21160 10
rect 21195 40 21245 50
rect 21195 10 21205 40
rect 21235 10 21245 40
rect 21195 0 21245 10
rect 21280 40 21330 50
rect 21280 10 21290 40
rect 21320 10 21330 40
rect 21280 0 21330 10
rect 21365 40 21415 50
rect 21365 10 21375 40
rect 21405 10 21415 40
rect 21365 0 21415 10
rect 21450 40 21500 50
rect 21450 10 21460 40
rect 21490 10 21500 40
rect 21450 0 21500 10
rect 21535 40 21585 50
rect 21535 10 21545 40
rect 21575 10 21585 40
rect 21535 0 21585 10
rect 21620 40 21670 50
rect 21620 10 21630 40
rect 21660 10 21670 40
rect 21620 0 21670 10
rect 21705 40 21755 50
rect 21705 10 21715 40
rect 21745 10 21755 40
rect 21705 0 21755 10
rect 21790 40 21840 50
rect 21790 10 21800 40
rect 21830 10 21840 40
rect 21790 0 21840 10
rect 21875 40 21925 50
rect 21875 10 21885 40
rect 21915 10 21925 40
rect 21875 0 21925 10
rect 21960 40 22010 50
rect 21960 10 21970 40
rect 22000 10 22010 40
rect 21960 0 22010 10
rect 22045 40 22095 50
rect 22045 10 22055 40
rect 22085 10 22095 40
rect 22045 0 22095 10
rect 22130 40 22180 50
rect 22130 10 22140 40
rect 22170 10 22180 40
rect 22130 0 22180 10
rect 22215 40 22265 50
rect 22215 10 22225 40
rect 22255 10 22265 40
rect 22215 0 22265 10
rect 22300 40 22350 50
rect 22300 10 22310 40
rect 22340 10 22350 40
rect 22300 0 22350 10
rect 22385 40 22435 50
rect 22385 10 22395 40
rect 22425 10 22435 40
rect 22385 0 22435 10
rect 22470 40 22520 50
rect 22470 10 22480 40
rect 22510 10 22520 40
rect 22470 0 22520 10
rect 22555 40 22605 50
rect 22555 10 22565 40
rect 22595 10 22605 40
rect 22555 0 22605 10
rect 22640 40 22690 50
rect 22640 10 22650 40
rect 22680 10 22690 40
rect 22640 0 22690 10
rect 22725 40 22775 50
rect 22725 10 22735 40
rect 22765 10 22775 40
rect 22725 0 22775 10
rect 22810 40 22860 50
rect 22810 10 22820 40
rect 22850 10 22860 40
rect 22810 0 22860 10
rect 22895 40 22945 50
rect 22895 10 22905 40
rect 22935 10 22945 40
rect 22895 0 22945 10
rect 22980 40 23030 50
rect 22980 10 22990 40
rect 23020 10 23030 40
rect 22980 0 23030 10
rect 23065 40 23115 50
rect 23065 10 23075 40
rect 23105 10 23115 40
rect 23065 0 23115 10
rect 23150 40 23200 50
rect 23150 10 23160 40
rect 23190 10 23200 40
rect 23150 0 23200 10
rect 23235 40 23285 50
rect 23235 10 23245 40
rect 23275 10 23285 40
rect 23235 0 23285 10
rect 23320 40 23370 50
rect 23320 10 23330 40
rect 23360 10 23370 40
rect 23320 0 23370 10
rect 23405 40 23455 50
rect 23405 10 23415 40
rect 23445 10 23455 40
rect 23405 0 23455 10
rect 23490 40 23540 50
rect 23490 10 23500 40
rect 23530 10 23540 40
rect 23490 0 23540 10
rect 23575 40 23625 50
rect 23575 10 23585 40
rect 23615 10 23625 40
rect 23575 0 23625 10
rect 23660 40 23710 50
rect 23660 10 23670 40
rect 23700 10 23710 40
rect 23660 0 23710 10
rect 23745 40 23795 50
rect 23745 10 23755 40
rect 23785 10 23795 40
rect 23745 0 23795 10
rect 23830 40 23880 50
rect 23830 10 23840 40
rect 23870 10 23880 40
rect 23830 0 23880 10
rect 23915 40 23965 50
rect 23915 10 23925 40
rect 23955 10 23965 40
rect 23915 0 23965 10
rect 24000 40 24050 50
rect 24000 10 24010 40
rect 24040 10 24050 40
rect 24000 0 24050 10
rect 24085 40 24135 50
rect 24085 10 24095 40
rect 24125 10 24135 40
rect 24085 0 24135 10
rect 24170 40 24220 50
rect 24170 10 24180 40
rect 24210 10 24220 40
rect 24170 0 24220 10
rect 24255 40 24305 50
rect 24255 10 24265 40
rect 24295 10 24305 40
rect 24255 0 24305 10
rect 24340 40 24390 50
rect 24340 10 24350 40
rect 24380 10 24390 40
rect 24340 0 24390 10
rect 24425 40 24475 50
rect 24425 10 24435 40
rect 24465 10 24475 40
rect 24425 0 24475 10
rect 24510 40 24560 50
rect 24510 10 24520 40
rect 24550 10 24560 40
rect 24510 0 24560 10
rect 24595 40 24645 50
rect 24595 10 24605 40
rect 24635 10 24645 40
rect 24595 0 24645 10
rect 24680 40 24730 50
rect 24680 10 24690 40
rect 24720 10 24730 40
rect 24680 0 24730 10
rect 24765 40 24815 50
rect 24765 10 24775 40
rect 24805 10 24815 40
rect 24765 0 24815 10
rect 24850 40 24900 50
rect 24850 10 24860 40
rect 24890 10 24900 40
rect 24850 0 24900 10
rect 24935 40 24985 50
rect 24935 10 24945 40
rect 24975 10 24985 40
rect 24935 0 24985 10
rect 25020 40 25070 50
rect 25020 10 25030 40
rect 25060 10 25070 40
rect 25020 0 25070 10
rect 25105 40 25155 50
rect 25105 10 25115 40
rect 25145 10 25155 40
rect 25105 0 25155 10
rect 25190 40 25240 50
rect 25190 10 25200 40
rect 25230 10 25240 40
rect 25190 0 25240 10
rect 25275 40 25325 50
rect 25275 10 25285 40
rect 25315 10 25325 40
rect 25275 0 25325 10
rect 25360 40 25410 50
rect 25360 10 25370 40
rect 25400 10 25410 40
rect 25360 0 25410 10
rect 25445 40 25495 50
rect 25445 10 25455 40
rect 25485 10 25495 40
rect 25445 0 25495 10
rect 25530 40 25580 50
rect 25530 10 25540 40
rect 25570 10 25580 40
rect 25530 0 25580 10
rect 25615 40 25665 50
rect 25615 10 25625 40
rect 25655 10 25665 40
rect 25615 0 25665 10
rect 25700 40 25750 50
rect 25700 10 25710 40
rect 25740 10 25750 40
rect 25700 0 25750 10
rect 25785 40 25835 50
rect 25785 10 25795 40
rect 25825 10 25835 40
rect 25785 0 25835 10
rect 25870 40 25920 50
rect 25870 10 25880 40
rect 25910 10 25920 40
rect 25870 0 25920 10
rect 25955 40 26005 50
rect 25955 10 25965 40
rect 25995 10 26005 40
rect 25955 0 26005 10
rect 26040 40 26090 50
rect 26040 10 26050 40
rect 26080 10 26090 40
rect 26040 0 26090 10
rect 26125 40 26175 50
rect 26125 10 26135 40
rect 26165 10 26175 40
rect 26125 0 26175 10
rect 26210 40 26260 50
rect 26210 10 26220 40
rect 26250 10 26260 40
rect 26210 0 26260 10
rect 26295 40 26345 50
rect 26295 10 26305 40
rect 26335 10 26345 40
rect 26295 0 26345 10
rect 26380 40 26430 50
rect 26380 10 26390 40
rect 26420 10 26430 40
rect 26380 0 26430 10
rect 26465 40 26515 50
rect 26465 10 26475 40
rect 26505 10 26515 40
rect 26465 0 26515 10
rect 26550 40 26600 50
rect 26550 10 26560 40
rect 26590 10 26600 40
rect 26550 0 26600 10
rect 26635 40 26685 50
rect 26635 10 26645 40
rect 26675 10 26685 40
rect 26635 0 26685 10
rect 26720 40 26770 50
rect 26720 10 26730 40
rect 26760 10 26770 40
rect 26720 0 26770 10
rect 26805 40 26855 50
rect 26805 10 26815 40
rect 26845 10 26855 40
rect 26805 0 26855 10
rect 26890 40 26940 50
rect 26890 10 26900 40
rect 26930 10 26940 40
rect 26890 0 26940 10
rect 26975 40 27025 50
rect 26975 10 26985 40
rect 27015 10 27025 40
rect 26975 0 27025 10
rect 27060 40 27110 50
rect 27060 10 27070 40
rect 27100 10 27110 40
rect 27060 0 27110 10
rect 27145 40 27195 50
rect 27145 10 27155 40
rect 27185 10 27195 40
rect 27145 0 27195 10
rect 27230 40 27280 50
rect 27230 10 27240 40
rect 27270 10 27280 40
rect 27230 0 27280 10
rect 27315 40 27365 50
rect 27315 10 27325 40
rect 27355 10 27365 40
rect 27315 0 27365 10
rect 27400 40 27450 50
rect 27400 10 27410 40
rect 27440 10 27450 40
rect 27400 0 27450 10
rect 27485 40 27535 50
rect 27485 10 27495 40
rect 27525 10 27535 40
rect 27485 0 27535 10
rect 27570 40 27620 50
rect 27570 10 27580 40
rect 27610 10 27620 40
rect 27570 0 27620 10
rect 27655 40 27705 50
rect 27655 10 27665 40
rect 27695 10 27705 40
rect 27655 0 27705 10
rect 27740 40 27790 50
rect 27740 10 27750 40
rect 27780 10 27790 40
rect 27740 0 27790 10
rect 27825 40 27875 50
rect 27825 10 27835 40
rect 27865 10 27875 40
rect 27825 0 27875 10
rect 27910 40 27960 50
rect 27910 10 27920 40
rect 27950 10 27960 40
rect 27910 0 27960 10
rect 27995 40 28045 50
rect 27995 10 28005 40
rect 28035 10 28045 40
rect 27995 0 28045 10
rect 28080 40 28130 50
rect 28080 10 28090 40
rect 28120 10 28130 40
rect 28080 0 28130 10
rect 28165 40 28215 50
rect 28165 10 28175 40
rect 28205 10 28215 40
rect 28165 0 28215 10
rect 28250 40 28300 50
rect 28250 10 28260 40
rect 28290 10 28300 40
rect 28250 0 28300 10
rect 28335 40 28385 50
rect 28335 10 28345 40
rect 28375 10 28385 40
rect 28335 0 28385 10
rect 28420 40 28470 50
rect 28420 10 28430 40
rect 28460 10 28470 40
rect 28420 0 28470 10
rect 28505 40 28555 50
rect 28505 10 28515 40
rect 28545 10 28555 40
rect 28505 0 28555 10
rect 28590 40 28640 50
rect 28590 10 28600 40
rect 28630 10 28640 40
rect 28590 0 28640 10
rect 28675 40 28725 50
rect 28675 10 28685 40
rect 28715 10 28725 40
rect 28675 0 28725 10
rect 28760 40 28810 50
rect 28760 10 28770 40
rect 28800 10 28810 40
rect 28760 0 28810 10
rect 28845 40 28895 50
rect 28845 10 28855 40
rect 28885 10 28895 40
rect 28845 0 28895 10
rect 28930 40 28980 50
rect 28930 10 28940 40
rect 28970 10 28980 40
rect 28930 0 28980 10
rect 29015 40 29065 50
rect 29015 10 29025 40
rect 29055 10 29065 40
rect 29015 0 29065 10
rect 29100 40 29150 50
rect 29100 10 29110 40
rect 29140 10 29150 40
rect 29100 0 29150 10
rect 29185 40 29235 50
rect 29185 10 29195 40
rect 29225 10 29235 40
rect 29185 0 29235 10
rect 29270 40 29320 50
rect 29270 10 29280 40
rect 29310 10 29320 40
rect 29270 0 29320 10
rect 29355 40 29405 50
rect 29355 10 29365 40
rect 29395 10 29405 40
rect 29355 0 29405 10
rect 29440 40 29490 50
rect 29440 10 29450 40
rect 29480 10 29490 40
rect 29440 0 29490 10
rect 29525 40 29575 50
rect 29525 10 29535 40
rect 29565 10 29575 40
rect 29525 0 29575 10
rect 29610 40 29660 50
rect 29610 10 29620 40
rect 29650 10 29660 40
rect 29610 0 29660 10
rect 5 -30 55 -20
rect 5 -60 15 -30
rect 45 -60 55 -30
rect 5 -70 55 -60
rect 90 -30 140 -20
rect 90 -60 100 -30
rect 130 -60 140 -30
rect 90 -70 140 -60
rect 255 -30 310 -20
rect 255 -60 265 -30
rect 300 -60 310 -30
rect 255 -70 310 -60
rect 340 -30 395 -20
rect 340 -60 350 -30
rect 385 -60 395 -30
rect 340 -70 395 -60
rect 425 -30 480 -20
rect 425 -60 435 -30
rect 470 -60 480 -30
rect 425 -70 480 -60
rect 510 -30 565 -20
rect 510 -60 520 -30
rect 555 -60 565 -30
rect 510 -70 565 -60
rect 790 -30 845 -20
rect 790 -60 800 -30
rect 835 -60 845 -30
rect 790 -70 845 -60
rect 875 -30 930 -20
rect 875 -60 885 -30
rect 920 -60 930 -30
rect 875 -70 930 -60
rect 960 -30 1015 -20
rect 960 -60 970 -30
rect 1005 -60 1015 -30
rect 960 -70 1015 -60
rect 1045 -30 1100 -20
rect 1045 -60 1055 -30
rect 1090 -60 1100 -30
rect 1045 -70 1100 -60
rect 1130 -30 1185 -20
rect 1130 -60 1140 -30
rect 1175 -60 1185 -30
rect 1130 -70 1185 -60
rect 1215 -30 1270 -20
rect 1215 -60 1225 -30
rect 1260 -60 1270 -30
rect 1215 -70 1270 -60
rect 1300 -30 1355 -20
rect 1300 -60 1310 -30
rect 1345 -60 1355 -30
rect 1300 -70 1355 -60
rect 1385 -30 1440 -20
rect 1385 -60 1395 -30
rect 1430 -60 1440 -30
rect 1385 -70 1440 -60
rect 1470 -30 1525 -20
rect 1470 -60 1480 -30
rect 1515 -60 1525 -30
rect 1470 -70 1525 -60
rect 1555 -30 1610 -20
rect 1555 -60 1565 -30
rect 1600 -60 1610 -30
rect 1555 -70 1610 -60
rect 1640 -30 1695 -20
rect 1640 -60 1650 -30
rect 1685 -60 1695 -30
rect 1640 -70 1695 -60
rect 1725 -30 1780 -20
rect 1725 -60 1735 -30
rect 1770 -60 1780 -30
rect 1725 -70 1780 -60
rect 1810 -30 1865 -20
rect 1810 -60 1820 -30
rect 1855 -60 1865 -30
rect 1810 -70 1865 -60
rect 1895 -30 1950 -20
rect 1895 -60 1905 -30
rect 1940 -60 1950 -30
rect 1895 -70 1950 -60
rect 1980 -30 2035 -20
rect 1980 -60 1990 -30
rect 2025 -60 2035 -30
rect 1980 -70 2035 -60
rect 2065 -30 2120 -20
rect 2065 -60 2075 -30
rect 2110 -60 2120 -30
rect 2065 -70 2120 -60
rect 2300 -30 2355 -20
rect 2300 -60 2310 -30
rect 2345 -60 2355 -30
rect 2300 -70 2355 -60
rect 2385 -30 2440 -20
rect 2385 -60 2395 -30
rect 2430 -60 2440 -30
rect 2385 -70 2440 -60
rect 2470 -30 2525 -20
rect 2470 -60 2480 -30
rect 2515 -60 2525 -30
rect 2470 -70 2525 -60
rect 2555 -30 2610 -20
rect 2555 -60 2565 -30
rect 2600 -60 2610 -30
rect 2555 -70 2610 -60
rect 2640 -30 2695 -20
rect 2640 -60 2650 -30
rect 2685 -60 2695 -30
rect 2640 -70 2695 -60
rect 2725 -30 2780 -20
rect 2725 -60 2735 -30
rect 2770 -60 2780 -30
rect 2725 -70 2780 -60
rect 2810 -30 2865 -20
rect 2810 -60 2820 -30
rect 2855 -60 2865 -30
rect 2810 -70 2865 -60
rect 2895 -30 2950 -20
rect 2895 -60 2905 -30
rect 2940 -60 2950 -30
rect 2895 -70 2950 -60
rect 2980 -30 3035 -20
rect 2980 -60 2990 -30
rect 3025 -60 3035 -30
rect 2980 -70 3035 -60
rect 3065 -30 3120 -20
rect 3065 -60 3075 -30
rect 3110 -60 3120 -30
rect 3065 -70 3120 -60
rect 3150 -30 3205 -20
rect 3150 -60 3160 -30
rect 3195 -60 3205 -30
rect 3150 -70 3205 -60
rect 3235 -30 3290 -20
rect 3235 -60 3245 -30
rect 3280 -60 3290 -30
rect 3235 -70 3290 -60
rect 3320 -30 3375 -20
rect 3320 -60 3330 -30
rect 3365 -60 3375 -30
rect 3320 -70 3375 -60
rect 3405 -30 3460 -20
rect 3405 -60 3415 -30
rect 3450 -60 3460 -30
rect 3405 -70 3460 -60
rect 3490 -30 3545 -20
rect 3490 -60 3500 -30
rect 3535 -60 3545 -30
rect 3490 -70 3545 -60
rect 3575 -30 3630 -20
rect 3575 -60 3585 -30
rect 3620 -60 3630 -30
rect 3575 -70 3630 -60
rect 3660 -30 3715 -20
rect 3660 -60 3670 -30
rect 3705 -60 3715 -30
rect 3660 -70 3715 -60
rect 3745 -30 3800 -20
rect 3745 -60 3755 -30
rect 3790 -60 3800 -30
rect 3745 -70 3800 -60
rect 3830 -30 3885 -20
rect 3830 -60 3840 -30
rect 3875 -60 3885 -30
rect 3830 -70 3885 -60
rect 3915 -30 3970 -20
rect 3915 -60 3925 -30
rect 3960 -60 3970 -30
rect 3915 -70 3970 -60
rect 4000 -30 4055 -20
rect 4000 -60 4010 -30
rect 4045 -60 4055 -30
rect 4000 -70 4055 -60
rect 4085 -30 4140 -20
rect 4085 -60 4095 -30
rect 4130 -60 4140 -30
rect 4085 -70 4140 -60
rect 4170 -30 4225 -20
rect 4170 -60 4180 -30
rect 4215 -60 4225 -30
rect 4170 -70 4225 -60
rect 4255 -30 4310 -20
rect 4255 -60 4265 -30
rect 4300 -60 4310 -30
rect 4255 -70 4310 -60
rect 4340 -30 4395 -20
rect 4340 -60 4350 -30
rect 4385 -60 4395 -30
rect 4340 -70 4395 -60
rect 4425 -30 4480 -20
rect 4425 -60 4435 -30
rect 4470 -60 4480 -30
rect 4425 -70 4480 -60
rect 4510 -30 4565 -20
rect 4510 -60 4520 -30
rect 4555 -60 4565 -30
rect 4510 -70 4565 -60
rect 4595 -30 4650 -20
rect 4595 -60 4605 -30
rect 4640 -60 4650 -30
rect 4595 -70 4650 -60
rect 4680 -30 4735 -20
rect 4680 -60 4690 -30
rect 4725 -60 4735 -30
rect 4680 -70 4735 -60
rect 4765 -30 4820 -20
rect 4765 -60 4775 -30
rect 4810 -60 4820 -30
rect 4765 -70 4820 -60
rect 4850 -30 4905 -20
rect 4850 -60 4860 -30
rect 4895 -60 4905 -30
rect 4850 -70 4905 -60
rect 4935 -30 4990 -20
rect 4935 -60 4945 -30
rect 4980 -60 4990 -30
rect 4935 -70 4990 -60
rect 5020 -30 5075 -20
rect 5020 -60 5030 -30
rect 5065 -60 5075 -30
rect 5020 -70 5075 -60
rect 5105 -30 5160 -20
rect 5105 -60 5115 -30
rect 5150 -60 5160 -30
rect 5105 -70 5160 -60
rect 5190 -30 5245 -20
rect 5190 -60 5200 -30
rect 5235 -60 5245 -30
rect 5190 -70 5245 -60
rect 5275 -30 5330 -20
rect 5275 -60 5285 -30
rect 5320 -60 5330 -30
rect 5275 -70 5330 -60
rect 5360 -30 5415 -20
rect 5360 -60 5370 -30
rect 5405 -60 5415 -30
rect 5360 -70 5415 -60
rect 5445 -30 5500 -20
rect 5445 -60 5455 -30
rect 5490 -60 5500 -30
rect 5445 -70 5500 -60
rect 5530 -30 5585 -20
rect 5530 -60 5540 -30
rect 5575 -60 5585 -30
rect 5530 -70 5585 -60
rect 5615 -30 5670 -20
rect 5615 -60 5625 -30
rect 5660 -60 5670 -30
rect 5615 -70 5670 -60
rect 5700 -30 5755 -20
rect 5700 -60 5710 -30
rect 5745 -60 5755 -30
rect 5700 -70 5755 -60
rect 5785 -30 5840 -20
rect 5785 -60 5795 -30
rect 5830 -60 5840 -30
rect 5785 -70 5840 -60
rect 5870 -30 5925 -20
rect 5870 -60 5880 -30
rect 5915 -60 5925 -30
rect 5870 -70 5925 -60
rect 5955 -30 6010 -20
rect 5955 -60 5965 -30
rect 6000 -60 6010 -30
rect 5955 -70 6010 -60
rect 6040 -30 6095 -20
rect 6040 -60 6050 -30
rect 6085 -60 6095 -30
rect 6040 -70 6095 -60
rect 6125 -30 6180 -20
rect 6125 -60 6135 -30
rect 6170 -60 6180 -30
rect 6125 -70 6180 -60
rect 6210 -30 6265 -20
rect 6210 -60 6220 -30
rect 6255 -60 6265 -30
rect 6210 -70 6265 -60
rect 6295 -30 6350 -20
rect 6295 -60 6305 -30
rect 6340 -60 6350 -30
rect 6295 -70 6350 -60
rect 6380 -30 6435 -20
rect 6380 -60 6390 -30
rect 6425 -60 6435 -30
rect 6380 -70 6435 -60
rect 6465 -30 6520 -20
rect 6465 -60 6475 -30
rect 6510 -60 6520 -30
rect 6465 -70 6520 -60
rect 6550 -30 6605 -20
rect 6550 -60 6560 -30
rect 6595 -60 6605 -30
rect 6550 -70 6605 -60
rect 6635 -30 6690 -20
rect 6635 -60 6645 -30
rect 6680 -60 6690 -30
rect 6635 -70 6690 -60
rect 6720 -30 6775 -20
rect 6720 -60 6730 -30
rect 6765 -60 6775 -30
rect 6720 -70 6775 -60
rect 6805 -30 6860 -20
rect 6805 -60 6815 -30
rect 6850 -60 6860 -30
rect 6805 -70 6860 -60
rect 6890 -30 6945 -20
rect 6890 -60 6900 -30
rect 6935 -60 6945 -30
rect 6890 -70 6945 -60
rect 6975 -30 7030 -20
rect 6975 -60 6985 -30
rect 7020 -60 7030 -30
rect 6975 -70 7030 -60
rect 7060 -30 7115 -20
rect 7060 -60 7070 -30
rect 7105 -60 7115 -30
rect 7060 -70 7115 -60
rect 7145 -30 7200 -20
rect 7145 -60 7155 -30
rect 7190 -60 7200 -30
rect 7145 -70 7200 -60
rect 7230 -30 7285 -20
rect 7230 -60 7240 -30
rect 7275 -60 7285 -30
rect 7230 -70 7285 -60
rect 7315 -30 7370 -20
rect 7315 -60 7325 -30
rect 7360 -60 7370 -30
rect 7315 -70 7370 -60
rect 7400 -30 7455 -20
rect 7400 -60 7410 -30
rect 7445 -60 7455 -30
rect 7400 -70 7455 -60
rect 7485 -30 7540 -20
rect 7485 -60 7495 -30
rect 7530 -60 7540 -30
rect 7485 -70 7540 -60
rect 7570 -30 7625 -20
rect 7570 -60 7580 -30
rect 7615 -60 7625 -30
rect 7570 -70 7625 -60
rect 7655 -30 7710 -20
rect 7655 -60 7665 -30
rect 7700 -60 7710 -30
rect 7655 -70 7710 -60
rect 7890 -30 7945 -20
rect 7890 -60 7900 -30
rect 7935 -60 7945 -30
rect 7890 -70 7945 -60
rect 7975 -30 8030 -20
rect 7975 -60 7985 -30
rect 8020 -60 8030 -30
rect 7975 -70 8030 -60
rect 8060 -30 8115 -20
rect 8060 -60 8070 -30
rect 8105 -60 8115 -30
rect 8060 -70 8115 -60
rect 8145 -30 8200 -20
rect 8145 -60 8155 -30
rect 8190 -60 8200 -30
rect 8145 -70 8200 -60
rect 8230 -30 8285 -20
rect 8230 -60 8240 -30
rect 8275 -60 8285 -30
rect 8230 -70 8285 -60
rect 8315 -30 8370 -20
rect 8315 -60 8325 -30
rect 8360 -60 8370 -30
rect 8315 -70 8370 -60
rect 8400 -30 8455 -20
rect 8400 -60 8410 -30
rect 8445 -60 8455 -30
rect 8400 -70 8455 -60
rect 8485 -30 8540 -20
rect 8485 -60 8495 -30
rect 8530 -60 8540 -30
rect 8485 -70 8540 -60
rect 8570 -30 8625 -20
rect 8570 -60 8580 -30
rect 8615 -60 8625 -30
rect 8570 -70 8625 -60
rect 8655 -30 8710 -20
rect 8655 -60 8665 -30
rect 8700 -60 8710 -30
rect 8655 -70 8710 -60
rect 8740 -30 8795 -20
rect 8740 -60 8750 -30
rect 8785 -60 8795 -30
rect 8740 -70 8795 -60
rect 8825 -30 8880 -20
rect 8825 -60 8835 -30
rect 8870 -60 8880 -30
rect 8825 -70 8880 -60
rect 8910 -30 8965 -20
rect 8910 -60 8920 -30
rect 8955 -60 8965 -30
rect 8910 -70 8965 -60
rect 8995 -30 9050 -20
rect 8995 -60 9005 -30
rect 9040 -60 9050 -30
rect 8995 -70 9050 -60
rect 9080 -30 9135 -20
rect 9080 -60 9090 -30
rect 9125 -60 9135 -30
rect 9080 -70 9135 -60
rect 9165 -30 9220 -20
rect 9165 -60 9175 -30
rect 9210 -60 9220 -30
rect 9165 -70 9220 -60
rect 9250 -30 9305 -20
rect 9250 -60 9260 -30
rect 9295 -60 9305 -30
rect 9250 -70 9305 -60
rect 9335 -30 9390 -20
rect 9335 -60 9345 -30
rect 9380 -60 9390 -30
rect 9335 -70 9390 -60
rect 9420 -30 9475 -20
rect 9420 -60 9430 -30
rect 9465 -60 9475 -30
rect 9420 -70 9475 -60
rect 9505 -30 9560 -20
rect 9505 -60 9515 -30
rect 9550 -60 9560 -30
rect 9505 -70 9560 -60
rect 9590 -30 9645 -20
rect 9590 -60 9600 -30
rect 9635 -60 9645 -30
rect 9590 -70 9645 -60
rect 9675 -30 9730 -20
rect 9675 -60 9685 -30
rect 9720 -60 9730 -30
rect 9675 -70 9730 -60
rect 9760 -30 9815 -20
rect 9760 -60 9770 -30
rect 9805 -60 9815 -30
rect 9760 -70 9815 -60
rect 9845 -30 9900 -20
rect 9845 -60 9855 -30
rect 9890 -60 9900 -30
rect 9845 -70 9900 -60
rect 9930 -30 9985 -20
rect 9930 -60 9940 -30
rect 9975 -60 9985 -30
rect 9930 -70 9985 -60
rect 10015 -30 10070 -20
rect 10015 -60 10025 -30
rect 10060 -60 10070 -30
rect 10015 -70 10070 -60
rect 10100 -30 10155 -20
rect 10100 -60 10110 -30
rect 10145 -60 10155 -30
rect 10100 -70 10155 -60
rect 10185 -30 10240 -20
rect 10185 -60 10195 -30
rect 10230 -60 10240 -30
rect 10185 -70 10240 -60
rect 10270 -30 10325 -20
rect 10270 -60 10280 -30
rect 10315 -60 10325 -30
rect 10270 -70 10325 -60
rect 10355 -30 10410 -20
rect 10355 -60 10365 -30
rect 10400 -60 10410 -30
rect 10355 -70 10410 -60
rect 10440 -30 10495 -20
rect 10440 -60 10450 -30
rect 10485 -60 10495 -30
rect 10440 -70 10495 -60
rect 10525 -30 10580 -20
rect 10525 -60 10535 -30
rect 10570 -60 10580 -30
rect 10525 -70 10580 -60
rect 10610 -30 10665 -20
rect 10610 -60 10620 -30
rect 10655 -60 10665 -30
rect 10610 -70 10665 -60
rect 10695 -30 10750 -20
rect 10695 -60 10705 -30
rect 10740 -60 10750 -30
rect 10695 -70 10750 -60
rect 10780 -30 10835 -20
rect 10780 -60 10790 -30
rect 10825 -60 10835 -30
rect 10780 -70 10835 -60
rect 10865 -30 10920 -20
rect 10865 -60 10875 -30
rect 10910 -60 10920 -30
rect 10865 -70 10920 -60
rect 10950 -30 11005 -20
rect 10950 -60 10960 -30
rect 10995 -60 11005 -30
rect 10950 -70 11005 -60
rect 11035 -30 11090 -20
rect 11035 -60 11045 -30
rect 11080 -60 11090 -30
rect 11035 -70 11090 -60
rect 11120 -30 11175 -20
rect 11120 -60 11130 -30
rect 11165 -60 11175 -30
rect 11120 -70 11175 -60
rect 11205 -30 11260 -20
rect 11205 -60 11215 -30
rect 11250 -60 11260 -30
rect 11205 -70 11260 -60
rect 11290 -30 11345 -20
rect 11290 -60 11300 -30
rect 11335 -60 11345 -30
rect 11290 -70 11345 -60
rect 11375 -30 11430 -20
rect 11375 -60 11385 -30
rect 11420 -60 11430 -30
rect 11375 -70 11430 -60
rect 11460 -30 11515 -20
rect 11460 -60 11470 -30
rect 11505 -60 11515 -30
rect 11460 -70 11515 -60
rect 11545 -30 11600 -20
rect 11545 -60 11555 -30
rect 11590 -60 11600 -30
rect 11545 -70 11600 -60
rect 11630 -30 11685 -20
rect 11630 -60 11640 -30
rect 11675 -60 11685 -30
rect 11630 -70 11685 -60
rect 11715 -30 11770 -20
rect 11715 -60 11725 -30
rect 11760 -60 11770 -30
rect 11715 -70 11770 -60
rect 11800 -30 11855 -20
rect 11800 -60 11810 -30
rect 11845 -60 11855 -30
rect 11800 -70 11855 -60
rect 11885 -30 11940 -20
rect 11885 -60 11895 -30
rect 11930 -60 11940 -30
rect 11885 -70 11940 -60
rect 11970 -30 12025 -20
rect 11970 -60 11980 -30
rect 12015 -60 12025 -30
rect 11970 -70 12025 -60
rect 12055 -30 12110 -20
rect 12055 -60 12065 -30
rect 12100 -60 12110 -30
rect 12055 -70 12110 -60
rect 12140 -30 12195 -20
rect 12140 -60 12150 -30
rect 12185 -60 12195 -30
rect 12140 -70 12195 -60
rect 12225 -30 12280 -20
rect 12225 -60 12235 -30
rect 12270 -60 12280 -30
rect 12225 -70 12280 -60
rect 12310 -30 12365 -20
rect 12310 -60 12320 -30
rect 12355 -60 12365 -30
rect 12310 -70 12365 -60
rect 12395 -30 12450 -20
rect 12395 -60 12405 -30
rect 12440 -60 12450 -30
rect 12395 -70 12450 -60
rect 12480 -30 12535 -20
rect 12480 -60 12490 -30
rect 12525 -60 12535 -30
rect 12480 -70 12535 -60
rect 12565 -30 12620 -20
rect 12565 -60 12575 -30
rect 12610 -60 12620 -30
rect 12565 -70 12620 -60
rect 12650 -30 12705 -20
rect 12650 -60 12660 -30
rect 12695 -60 12705 -30
rect 12650 -70 12705 -60
rect 12735 -30 12790 -20
rect 12735 -60 12745 -30
rect 12780 -60 12790 -30
rect 12735 -70 12790 -60
rect 12820 -30 12875 -20
rect 12820 -60 12830 -30
rect 12865 -60 12875 -30
rect 12820 -70 12875 -60
rect 12905 -30 12960 -20
rect 12905 -60 12915 -30
rect 12950 -60 12960 -30
rect 12905 -70 12960 -60
rect 12990 -30 13045 -20
rect 12990 -60 13000 -30
rect 13035 -60 13045 -30
rect 12990 -70 13045 -60
rect 13075 -30 13130 -20
rect 13075 -60 13085 -30
rect 13120 -60 13130 -30
rect 13075 -70 13130 -60
rect 13160 -30 13215 -20
rect 13160 -60 13170 -30
rect 13205 -60 13215 -30
rect 13160 -70 13215 -60
rect 13245 -30 13300 -20
rect 13245 -60 13255 -30
rect 13290 -60 13300 -30
rect 13245 -70 13300 -60
rect 13330 -30 13385 -20
rect 13330 -60 13340 -30
rect 13375 -60 13385 -30
rect 13330 -70 13385 -60
rect 13415 -30 13470 -20
rect 13415 -60 13425 -30
rect 13460 -60 13470 -30
rect 13415 -70 13470 -60
rect 13500 -30 13555 -20
rect 13500 -60 13510 -30
rect 13545 -60 13555 -30
rect 13500 -70 13555 -60
rect 13585 -30 13640 -20
rect 13585 -60 13595 -30
rect 13630 -60 13640 -30
rect 13585 -70 13640 -60
rect 13670 -30 13725 -20
rect 13670 -60 13680 -30
rect 13715 -60 13725 -30
rect 13670 -70 13725 -60
rect 13755 -30 13810 -20
rect 13755 -60 13765 -30
rect 13800 -60 13810 -30
rect 13755 -70 13810 -60
rect 13840 -30 13895 -20
rect 13840 -60 13850 -30
rect 13885 -60 13895 -30
rect 13840 -70 13895 -60
rect 13925 -30 13980 -20
rect 13925 -60 13935 -30
rect 13970 -60 13980 -30
rect 13925 -70 13980 -60
rect 14010 -30 14065 -20
rect 14010 -60 14020 -30
rect 14055 -60 14065 -30
rect 14010 -70 14065 -60
rect 14095 -30 14150 -20
rect 14095 -60 14105 -30
rect 14140 -60 14150 -30
rect 14095 -70 14150 -60
rect 14180 -30 14235 -20
rect 14180 -60 14190 -30
rect 14225 -60 14235 -30
rect 14180 -70 14235 -60
rect 14265 -30 14320 -20
rect 14265 -60 14275 -30
rect 14310 -60 14320 -30
rect 14265 -70 14320 -60
rect 14350 -30 14405 -20
rect 14350 -60 14360 -30
rect 14395 -60 14405 -30
rect 14350 -70 14405 -60
rect 14435 -30 14490 -20
rect 14435 -60 14445 -30
rect 14480 -60 14490 -30
rect 14435 -70 14490 -60
rect 14520 -30 14575 -20
rect 14520 -60 14530 -30
rect 14565 -60 14575 -30
rect 14520 -70 14575 -60
rect 14605 -30 14660 -20
rect 14605 -60 14615 -30
rect 14650 -60 14660 -30
rect 14605 -70 14660 -60
rect 14690 -30 14745 -20
rect 14690 -60 14700 -30
rect 14735 -60 14745 -30
rect 14690 -70 14745 -60
rect 14775 -30 14830 -20
rect 14775 -60 14785 -30
rect 14820 -60 14830 -30
rect 14775 -70 14830 -60
rect 14860 -30 14915 -20
rect 14860 -60 14870 -30
rect 14905 -60 14915 -30
rect 14860 -70 14915 -60
rect 14945 -30 15000 -20
rect 14945 -60 14955 -30
rect 14990 -60 15000 -30
rect 14945 -70 15000 -60
rect 15030 -30 15085 -20
rect 15030 -60 15040 -30
rect 15075 -60 15085 -30
rect 15030 -70 15085 -60
rect 15115 -30 15170 -20
rect 15115 -60 15125 -30
rect 15160 -60 15170 -30
rect 15115 -70 15170 -60
rect 15200 -30 15255 -20
rect 15200 -60 15210 -30
rect 15245 -60 15255 -30
rect 15200 -70 15255 -60
rect 15285 -30 15340 -20
rect 15285 -60 15295 -30
rect 15330 -60 15340 -30
rect 15285 -70 15340 -60
rect 15370 -30 15425 -20
rect 15370 -60 15380 -30
rect 15415 -60 15425 -30
rect 15370 -70 15425 -60
rect 15455 -30 15510 -20
rect 15455 -60 15465 -30
rect 15500 -60 15510 -30
rect 15455 -70 15510 -60
rect 15540 -30 15595 -20
rect 15540 -60 15550 -30
rect 15585 -60 15595 -30
rect 15540 -70 15595 -60
rect 15625 -30 15680 -20
rect 15625 -60 15635 -30
rect 15670 -60 15680 -30
rect 15625 -70 15680 -60
rect 15710 -30 15765 -20
rect 15710 -60 15720 -30
rect 15755 -60 15765 -30
rect 15710 -70 15765 -60
rect 15795 -30 15850 -20
rect 15795 -60 15805 -30
rect 15840 -60 15850 -30
rect 15795 -70 15850 -60
rect 15880 -30 15935 -20
rect 15880 -60 15890 -30
rect 15925 -60 15935 -30
rect 15880 -70 15935 -60
rect 15965 -30 16020 -20
rect 15965 -60 15975 -30
rect 16010 -60 16020 -30
rect 15965 -70 16020 -60
rect 16050 -30 16105 -20
rect 16050 -60 16060 -30
rect 16095 -60 16105 -30
rect 16050 -70 16105 -60
rect 16135 -30 16190 -20
rect 16135 -60 16145 -30
rect 16180 -60 16190 -30
rect 16135 -70 16190 -60
rect 16220 -30 16275 -20
rect 16220 -60 16230 -30
rect 16265 -60 16275 -30
rect 16220 -70 16275 -60
rect 16305 -30 16360 -20
rect 16305 -60 16315 -30
rect 16350 -60 16360 -30
rect 16305 -70 16360 -60
rect 16390 -30 16445 -20
rect 16390 -60 16400 -30
rect 16435 -60 16445 -30
rect 16390 -70 16445 -60
rect 16475 -30 16530 -20
rect 16475 -60 16485 -30
rect 16520 -60 16530 -30
rect 16475 -70 16530 -60
rect 16560 -30 16615 -20
rect 16560 -60 16570 -30
rect 16605 -60 16615 -30
rect 16560 -70 16615 -60
rect 16645 -30 16700 -20
rect 16645 -60 16655 -30
rect 16690 -60 16700 -30
rect 16645 -70 16700 -60
rect 16730 -30 16785 -20
rect 16730 -60 16740 -30
rect 16775 -60 16785 -30
rect 16730 -70 16785 -60
rect 16815 -30 16870 -20
rect 16815 -60 16825 -30
rect 16860 -60 16870 -30
rect 16815 -70 16870 -60
rect 16900 -30 16955 -20
rect 16900 -60 16910 -30
rect 16945 -60 16955 -30
rect 16900 -70 16955 -60
rect 16985 -30 17040 -20
rect 16985 -60 16995 -30
rect 17030 -60 17040 -30
rect 16985 -70 17040 -60
rect 17070 -30 17125 -20
rect 17070 -60 17080 -30
rect 17115 -60 17125 -30
rect 17070 -70 17125 -60
rect 17155 -30 17210 -20
rect 17155 -60 17165 -30
rect 17200 -60 17210 -30
rect 17155 -70 17210 -60
rect 17240 -30 17295 -20
rect 17240 -60 17250 -30
rect 17285 -60 17295 -30
rect 17240 -70 17295 -60
rect 17325 -30 17380 -20
rect 17325 -60 17335 -30
rect 17370 -60 17380 -30
rect 17325 -70 17380 -60
rect 17410 -30 17465 -20
rect 17410 -60 17420 -30
rect 17455 -60 17465 -30
rect 17410 -70 17465 -60
rect 17495 -30 17550 -20
rect 17495 -60 17505 -30
rect 17540 -60 17550 -30
rect 17495 -70 17550 -60
rect 17580 -30 17635 -20
rect 17580 -60 17590 -30
rect 17625 -60 17635 -30
rect 17580 -70 17635 -60
rect 17665 -30 17720 -20
rect 17665 -60 17675 -30
rect 17710 -60 17720 -30
rect 17665 -70 17720 -60
rect 17750 -30 17805 -20
rect 17750 -60 17760 -30
rect 17795 -60 17805 -30
rect 17750 -70 17805 -60
rect 17835 -30 17890 -20
rect 17835 -60 17845 -30
rect 17880 -60 17890 -30
rect 17835 -70 17890 -60
rect 17920 -30 17975 -20
rect 17920 -60 17930 -30
rect 17965 -60 17975 -30
rect 17920 -70 17975 -60
rect 18005 -30 18060 -20
rect 18005 -60 18015 -30
rect 18050 -60 18060 -30
rect 18005 -70 18060 -60
rect 18090 -30 18145 -20
rect 18090 -60 18100 -30
rect 18135 -60 18145 -30
rect 18090 -70 18145 -60
rect 18175 -30 18230 -20
rect 18175 -60 18185 -30
rect 18220 -60 18230 -30
rect 18175 -70 18230 -60
rect 18260 -30 18315 -20
rect 18260 -60 18270 -30
rect 18305 -60 18315 -30
rect 18260 -70 18315 -60
rect 18345 -30 18400 -20
rect 18345 -60 18355 -30
rect 18390 -60 18400 -30
rect 18345 -70 18400 -60
rect 18430 -30 18485 -20
rect 18430 -60 18440 -30
rect 18475 -60 18485 -30
rect 18430 -70 18485 -60
rect 18515 -30 18570 -20
rect 18515 -60 18525 -30
rect 18560 -60 18570 -30
rect 18515 -70 18570 -60
rect 18600 -30 18655 -20
rect 18600 -60 18610 -30
rect 18645 -60 18655 -30
rect 18600 -70 18655 -60
rect 18685 -30 18740 -20
rect 18685 -60 18695 -30
rect 18730 -60 18740 -30
rect 18685 -70 18740 -60
rect 18770 -30 18825 -20
rect 18770 -60 18780 -30
rect 18815 -60 18825 -30
rect 18770 -70 18825 -60
rect 18855 -30 18910 -20
rect 18855 -60 18865 -30
rect 18900 -60 18910 -30
rect 18855 -70 18910 -60
rect 18940 -30 18995 -20
rect 18940 -60 18950 -30
rect 18985 -60 18995 -30
rect 18940 -70 18995 -60
rect 19025 -30 19080 -20
rect 19025 -60 19035 -30
rect 19070 -60 19080 -30
rect 19025 -70 19080 -60
rect 19110 -30 19165 -20
rect 19110 -60 19120 -30
rect 19155 -60 19165 -30
rect 19110 -70 19165 -60
rect 19195 -30 19250 -20
rect 19195 -60 19205 -30
rect 19240 -60 19250 -30
rect 19195 -70 19250 -60
rect 19280 -30 19335 -20
rect 19280 -60 19290 -30
rect 19325 -60 19335 -30
rect 19280 -70 19335 -60
rect 19365 -30 19420 -20
rect 19365 -60 19375 -30
rect 19410 -60 19420 -30
rect 19365 -70 19420 -60
rect 19450 -30 19505 -20
rect 19450 -60 19460 -30
rect 19495 -60 19505 -30
rect 19450 -70 19505 -60
rect 19535 -30 19590 -20
rect 19535 -60 19545 -30
rect 19580 -60 19590 -30
rect 19535 -70 19590 -60
rect 19620 -30 19675 -20
rect 19620 -60 19630 -30
rect 19665 -60 19675 -30
rect 19620 -70 19675 -60
rect 19705 -30 19760 -20
rect 19705 -60 19715 -30
rect 19750 -60 19760 -30
rect 19705 -70 19760 -60
rect 19790 -30 19845 -20
rect 19790 -60 19800 -30
rect 19835 -60 19845 -30
rect 19790 -70 19845 -60
rect 19875 -30 19930 -20
rect 19875 -60 19885 -30
rect 19920 -60 19930 -30
rect 19875 -70 19930 -60
rect 19960 -30 20015 -20
rect 19960 -60 19970 -30
rect 20005 -60 20015 -30
rect 19960 -70 20015 -60
rect 20045 -30 20100 -20
rect 20045 -60 20055 -30
rect 20090 -60 20100 -30
rect 20045 -70 20100 -60
rect 20130 -30 20185 -20
rect 20130 -60 20140 -30
rect 20175 -60 20185 -30
rect 20130 -70 20185 -60
rect 20215 -30 20270 -20
rect 20215 -60 20225 -30
rect 20260 -60 20270 -30
rect 20215 -70 20270 -60
rect 20300 -30 20355 -20
rect 20300 -60 20310 -30
rect 20345 -60 20355 -30
rect 20300 -70 20355 -60
rect 20385 -30 20440 -20
rect 20385 -60 20395 -30
rect 20430 -60 20440 -30
rect 20385 -70 20440 -60
rect 20470 -30 20525 -20
rect 20470 -60 20480 -30
rect 20515 -60 20525 -30
rect 20470 -70 20525 -60
rect 20555 -30 20610 -20
rect 20555 -60 20565 -30
rect 20600 -60 20610 -30
rect 20555 -70 20610 -60
rect 20640 -30 20695 -20
rect 20640 -60 20650 -30
rect 20685 -60 20695 -30
rect 20640 -70 20695 -60
rect 20725 -30 20780 -20
rect 20725 -60 20735 -30
rect 20770 -60 20780 -30
rect 20725 -70 20780 -60
rect 20810 -30 20865 -20
rect 20810 -60 20820 -30
rect 20855 -60 20865 -30
rect 20810 -70 20865 -60
rect 20895 -30 20950 -20
rect 20895 -60 20905 -30
rect 20940 -60 20950 -30
rect 20895 -70 20950 -60
rect 20980 -30 21035 -20
rect 20980 -60 20990 -30
rect 21025 -60 21035 -30
rect 20980 -70 21035 -60
rect 21065 -30 21120 -20
rect 21065 -60 21075 -30
rect 21110 -60 21120 -30
rect 21065 -70 21120 -60
rect 21150 -30 21205 -20
rect 21150 -60 21160 -30
rect 21195 -60 21205 -30
rect 21150 -70 21205 -60
rect 21235 -30 21290 -20
rect 21235 -60 21245 -30
rect 21280 -60 21290 -30
rect 21235 -70 21290 -60
rect 21320 -30 21375 -20
rect 21320 -60 21330 -30
rect 21365 -60 21375 -30
rect 21320 -70 21375 -60
rect 21405 -30 21460 -20
rect 21405 -60 21415 -30
rect 21450 -60 21460 -30
rect 21405 -70 21460 -60
rect 21490 -30 21545 -20
rect 21490 -60 21500 -30
rect 21535 -60 21545 -30
rect 21490 -70 21545 -60
rect 21575 -30 21630 -20
rect 21575 -60 21585 -30
rect 21620 -60 21630 -30
rect 21575 -70 21630 -60
rect 21660 -30 21715 -20
rect 21660 -60 21670 -30
rect 21705 -60 21715 -30
rect 21660 -70 21715 -60
rect 21745 -30 21800 -20
rect 21745 -60 21755 -30
rect 21790 -60 21800 -30
rect 21745 -70 21800 -60
rect 21830 -30 21885 -20
rect 21830 -60 21840 -30
rect 21875 -60 21885 -30
rect 21830 -70 21885 -60
rect 21915 -30 21970 -20
rect 21915 -60 21925 -30
rect 21960 -60 21970 -30
rect 21915 -70 21970 -60
rect 22000 -30 22055 -20
rect 22000 -60 22010 -30
rect 22045 -60 22055 -30
rect 22000 -70 22055 -60
rect 22085 -30 22140 -20
rect 22085 -60 22095 -30
rect 22130 -60 22140 -30
rect 22085 -70 22140 -60
rect 22170 -30 22225 -20
rect 22170 -60 22180 -30
rect 22215 -60 22225 -30
rect 22170 -70 22225 -60
rect 22255 -30 22310 -20
rect 22255 -60 22265 -30
rect 22300 -60 22310 -30
rect 22255 -70 22310 -60
rect 22340 -30 22395 -20
rect 22340 -60 22350 -30
rect 22385 -60 22395 -30
rect 22340 -70 22395 -60
rect 22425 -30 22480 -20
rect 22425 -60 22435 -30
rect 22470 -60 22480 -30
rect 22425 -70 22480 -60
rect 22510 -30 22565 -20
rect 22510 -60 22520 -30
rect 22555 -60 22565 -30
rect 22510 -70 22565 -60
rect 22595 -30 22650 -20
rect 22595 -60 22605 -30
rect 22640 -60 22650 -30
rect 22595 -70 22650 -60
rect 22680 -30 22735 -20
rect 22680 -60 22690 -30
rect 22725 -60 22735 -30
rect 22680 -70 22735 -60
rect 22765 -30 22820 -20
rect 22765 -60 22775 -30
rect 22810 -60 22820 -30
rect 22765 -70 22820 -60
rect 22850 -30 22905 -20
rect 22850 -60 22860 -30
rect 22895 -60 22905 -30
rect 22850 -70 22905 -60
rect 22935 -30 22990 -20
rect 22935 -60 22945 -30
rect 22980 -60 22990 -30
rect 22935 -70 22990 -60
rect 23020 -30 23075 -20
rect 23020 -60 23030 -30
rect 23065 -60 23075 -30
rect 23020 -70 23075 -60
rect 23105 -30 23160 -20
rect 23105 -60 23115 -30
rect 23150 -60 23160 -30
rect 23105 -70 23160 -60
rect 23190 -30 23245 -20
rect 23190 -60 23200 -30
rect 23235 -60 23245 -30
rect 23190 -70 23245 -60
rect 23275 -30 23330 -20
rect 23275 -60 23285 -30
rect 23320 -60 23330 -30
rect 23275 -70 23330 -60
rect 23360 -30 23415 -20
rect 23360 -60 23370 -30
rect 23405 -60 23415 -30
rect 23360 -70 23415 -60
rect 23445 -30 23500 -20
rect 23445 -60 23455 -30
rect 23490 -60 23500 -30
rect 23445 -70 23500 -60
rect 23530 -30 23585 -20
rect 23530 -60 23540 -30
rect 23575 -60 23585 -30
rect 23530 -70 23585 -60
rect 23615 -30 23670 -20
rect 23615 -60 23625 -30
rect 23660 -60 23670 -30
rect 23615 -70 23670 -60
rect 23700 -30 23755 -20
rect 23700 -60 23710 -30
rect 23745 -60 23755 -30
rect 23700 -70 23755 -60
rect 23785 -30 23840 -20
rect 23785 -60 23795 -30
rect 23830 -60 23840 -30
rect 23785 -70 23840 -60
rect 23870 -30 23925 -20
rect 23870 -60 23880 -30
rect 23915 -60 23925 -30
rect 23870 -70 23925 -60
rect 23955 -30 24010 -20
rect 23955 -60 23965 -30
rect 24000 -60 24010 -30
rect 23955 -70 24010 -60
rect 24040 -30 24095 -20
rect 24040 -60 24050 -30
rect 24085 -60 24095 -30
rect 24040 -70 24095 -60
rect 24125 -30 24180 -20
rect 24125 -60 24135 -30
rect 24170 -60 24180 -30
rect 24125 -70 24180 -60
rect 24210 -30 24265 -20
rect 24210 -60 24220 -30
rect 24255 -60 24265 -30
rect 24210 -70 24265 -60
rect 24295 -30 24350 -20
rect 24295 -60 24305 -30
rect 24340 -60 24350 -30
rect 24295 -70 24350 -60
rect 24380 -30 24435 -20
rect 24380 -60 24390 -30
rect 24425 -60 24435 -30
rect 24380 -70 24435 -60
rect 24465 -30 24520 -20
rect 24465 -60 24475 -30
rect 24510 -60 24520 -30
rect 24465 -70 24520 -60
rect 24550 -30 24605 -20
rect 24550 -60 24560 -30
rect 24595 -60 24605 -30
rect 24550 -70 24605 -60
rect 24635 -30 24690 -20
rect 24635 -60 24645 -30
rect 24680 -60 24690 -30
rect 24635 -70 24690 -60
rect 24720 -30 24775 -20
rect 24720 -60 24730 -30
rect 24765 -60 24775 -30
rect 24720 -70 24775 -60
rect 24805 -30 24860 -20
rect 24805 -60 24815 -30
rect 24850 -60 24860 -30
rect 24805 -70 24860 -60
rect 24890 -30 24945 -20
rect 24890 -60 24900 -30
rect 24935 -60 24945 -30
rect 24890 -70 24945 -60
rect 24975 -30 25030 -20
rect 24975 -60 24985 -30
rect 25020 -60 25030 -30
rect 24975 -70 25030 -60
rect 25060 -30 25115 -20
rect 25060 -60 25070 -30
rect 25105 -60 25115 -30
rect 25060 -70 25115 -60
rect 25145 -30 25200 -20
rect 25145 -60 25155 -30
rect 25190 -60 25200 -30
rect 25145 -70 25200 -60
rect 25230 -30 25285 -20
rect 25230 -60 25240 -30
rect 25275 -60 25285 -30
rect 25230 -70 25285 -60
rect 25315 -30 25370 -20
rect 25315 -60 25325 -30
rect 25360 -60 25370 -30
rect 25315 -70 25370 -60
rect 25400 -30 25455 -20
rect 25400 -60 25410 -30
rect 25445 -60 25455 -30
rect 25400 -70 25455 -60
rect 25485 -30 25540 -20
rect 25485 -60 25495 -30
rect 25530 -60 25540 -30
rect 25485 -70 25540 -60
rect 25570 -30 25625 -20
rect 25570 -60 25580 -30
rect 25615 -60 25625 -30
rect 25570 -70 25625 -60
rect 25655 -30 25710 -20
rect 25655 -60 25665 -30
rect 25700 -60 25710 -30
rect 25655 -70 25710 -60
rect 25740 -30 25795 -20
rect 25740 -60 25750 -30
rect 25785 -60 25795 -30
rect 25740 -70 25795 -60
rect 25825 -30 25880 -20
rect 25825 -60 25835 -30
rect 25870 -60 25880 -30
rect 25825 -70 25880 -60
rect 25910 -30 25965 -20
rect 25910 -60 25920 -30
rect 25955 -60 25965 -30
rect 25910 -70 25965 -60
rect 25995 -30 26050 -20
rect 25995 -60 26005 -30
rect 26040 -60 26050 -30
rect 25995 -70 26050 -60
rect 26080 -30 26135 -20
rect 26080 -60 26090 -30
rect 26125 -60 26135 -30
rect 26080 -70 26135 -60
rect 26165 -30 26220 -20
rect 26165 -60 26175 -30
rect 26210 -60 26220 -30
rect 26165 -70 26220 -60
rect 26250 -30 26305 -20
rect 26250 -60 26260 -30
rect 26295 -60 26305 -30
rect 26250 -70 26305 -60
rect 26335 -30 26390 -20
rect 26335 -60 26345 -30
rect 26380 -60 26390 -30
rect 26335 -70 26390 -60
rect 26420 -30 26475 -20
rect 26420 -60 26430 -30
rect 26465 -60 26475 -30
rect 26420 -70 26475 -60
rect 26505 -30 26560 -20
rect 26505 -60 26515 -30
rect 26550 -60 26560 -30
rect 26505 -70 26560 -60
rect 26590 -30 26645 -20
rect 26590 -60 26600 -30
rect 26635 -60 26645 -30
rect 26590 -70 26645 -60
rect 26675 -30 26730 -20
rect 26675 -60 26685 -30
rect 26720 -60 26730 -30
rect 26675 -70 26730 -60
rect 26760 -30 26815 -20
rect 26760 -60 26770 -30
rect 26805 -60 26815 -30
rect 26760 -70 26815 -60
rect 26845 -30 26900 -20
rect 26845 -60 26855 -30
rect 26890 -60 26900 -30
rect 26845 -70 26900 -60
rect 26930 -30 26985 -20
rect 26930 -60 26940 -30
rect 26975 -60 26985 -30
rect 26930 -70 26985 -60
rect 27015 -30 27070 -20
rect 27015 -60 27025 -30
rect 27060 -60 27070 -30
rect 27015 -70 27070 -60
rect 27100 -30 27155 -20
rect 27100 -60 27110 -30
rect 27145 -60 27155 -30
rect 27100 -70 27155 -60
rect 27185 -30 27240 -20
rect 27185 -60 27195 -30
rect 27230 -60 27240 -30
rect 27185 -70 27240 -60
rect 27270 -30 27325 -20
rect 27270 -60 27280 -30
rect 27315 -60 27325 -30
rect 27270 -70 27325 -60
rect 27355 -30 27410 -20
rect 27355 -60 27365 -30
rect 27400 -60 27410 -30
rect 27355 -70 27410 -60
rect 27440 -30 27495 -20
rect 27440 -60 27450 -30
rect 27485 -60 27495 -30
rect 27440 -70 27495 -60
rect 27525 -30 27580 -20
rect 27525 -60 27535 -30
rect 27570 -60 27580 -30
rect 27525 -70 27580 -60
rect 27610 -30 27665 -20
rect 27610 -60 27620 -30
rect 27655 -60 27665 -30
rect 27610 -70 27665 -60
rect 27695 -30 27750 -20
rect 27695 -60 27705 -30
rect 27740 -60 27750 -30
rect 27695 -70 27750 -60
rect 27780 -30 27835 -20
rect 27780 -60 27790 -30
rect 27825 -60 27835 -30
rect 27780 -70 27835 -60
rect 27865 -30 27920 -20
rect 27865 -60 27875 -30
rect 27910 -60 27920 -30
rect 27865 -70 27920 -60
rect 27950 -30 28005 -20
rect 27950 -60 27960 -30
rect 27995 -60 28005 -30
rect 27950 -70 28005 -60
rect 28035 -30 28090 -20
rect 28035 -60 28045 -30
rect 28080 -60 28090 -30
rect 28035 -70 28090 -60
rect 28120 -30 28175 -20
rect 28120 -60 28130 -30
rect 28165 -60 28175 -30
rect 28120 -70 28175 -60
rect 28205 -30 28260 -20
rect 28205 -60 28215 -30
rect 28250 -60 28260 -30
rect 28205 -70 28260 -60
rect 28290 -30 28345 -20
rect 28290 -60 28300 -30
rect 28335 -60 28345 -30
rect 28290 -70 28345 -60
rect 28375 -30 28430 -20
rect 28375 -60 28385 -30
rect 28420 -60 28430 -30
rect 28375 -70 28430 -60
rect 28460 -30 28515 -20
rect 28460 -60 28470 -30
rect 28505 -60 28515 -30
rect 28460 -70 28515 -60
rect 28545 -30 28600 -20
rect 28545 -60 28555 -30
rect 28590 -60 28600 -30
rect 28545 -70 28600 -60
rect 28630 -30 28685 -20
rect 28630 -60 28640 -30
rect 28675 -60 28685 -30
rect 28630 -70 28685 -60
rect 28715 -30 28770 -20
rect 28715 -60 28725 -30
rect 28760 -60 28770 -30
rect 28715 -70 28770 -60
rect 28800 -30 28855 -20
rect 28800 -60 28810 -30
rect 28845 -60 28855 -30
rect 28800 -70 28855 -60
rect 28885 -30 28940 -20
rect 28885 -60 28895 -30
rect 28930 -60 28940 -30
rect 28885 -70 28940 -60
rect 28970 -30 29025 -20
rect 28970 -60 28980 -30
rect 29015 -60 29025 -30
rect 28970 -70 29025 -60
rect 29055 -30 29110 -20
rect 29055 -60 29065 -30
rect 29100 -60 29110 -30
rect 29055 -70 29110 -60
rect 29140 -30 29195 -20
rect 29140 -60 29150 -30
rect 29185 -60 29195 -30
rect 29140 -70 29195 -60
rect 29225 -30 29280 -20
rect 29225 -60 29235 -30
rect 29270 -60 29280 -30
rect 29225 -70 29280 -60
rect 29310 -30 29365 -20
rect 29310 -60 29320 -30
rect 29355 -60 29365 -30
rect 29310 -70 29365 -60
rect 29395 -30 29450 -20
rect 29395 -60 29405 -30
rect 29440 -60 29450 -30
rect 29395 -70 29450 -60
rect 29480 -30 29535 -20
rect 29480 -60 29490 -30
rect 29525 -60 29535 -30
rect 29480 -70 29535 -60
rect 29565 -30 29620 -20
rect 29565 -60 29575 -30
rect 29610 -60 29620 -30
rect 29565 -70 29620 -60
rect 105 -265 160 -255
rect 105 -295 115 -265
rect 150 -295 160 -265
rect 105 -305 160 -295
rect 190 -265 245 -255
rect 190 -295 200 -265
rect 235 -295 245 -265
rect 190 -305 245 -295
rect 275 -265 330 -255
rect 275 -295 285 -265
rect 320 -295 330 -265
rect 275 -305 330 -295
rect 360 -265 415 -255
rect 360 -295 370 -265
rect 405 -295 415 -265
rect 360 -305 415 -295
rect 445 -265 500 -255
rect 445 -295 455 -265
rect 490 -295 500 -265
rect 445 -305 500 -295
rect 530 -265 585 -255
rect 530 -295 540 -265
rect 575 -295 585 -265
rect 530 -305 585 -295
rect 615 -265 670 -255
rect 615 -295 625 -265
rect 660 -295 670 -265
rect 615 -305 670 -295
rect 700 -265 755 -255
rect 700 -295 710 -265
rect 745 -295 755 -265
rect 700 -305 755 -295
rect 785 -265 840 -255
rect 785 -295 795 -265
rect 830 -295 840 -265
rect 785 -305 840 -295
rect 870 -265 925 -255
rect 870 -295 880 -265
rect 915 -295 925 -265
rect 870 -305 925 -295
rect 955 -265 1010 -255
rect 955 -295 965 -265
rect 1000 -295 1010 -265
rect 955 -305 1010 -295
rect 1040 -265 1095 -255
rect 1040 -295 1050 -265
rect 1085 -295 1095 -265
rect 1040 -305 1095 -295
rect 1125 -265 1180 -255
rect 1125 -295 1135 -265
rect 1170 -295 1180 -265
rect 1125 -305 1180 -295
rect 1210 -265 1265 -255
rect 1210 -295 1220 -265
rect 1255 -295 1265 -265
rect 1210 -305 1265 -295
rect 1295 -265 1350 -255
rect 1295 -295 1305 -265
rect 1340 -295 1350 -265
rect 1295 -305 1350 -295
rect 1380 -265 1435 -255
rect 1380 -295 1390 -265
rect 1425 -295 1435 -265
rect 1380 -305 1435 -295
rect 1465 -265 1520 -255
rect 1465 -295 1475 -265
rect 1510 -295 1520 -265
rect 1465 -305 1520 -295
rect 1550 -265 1605 -255
rect 1550 -295 1560 -265
rect 1595 -295 1605 -265
rect 1550 -305 1605 -295
rect 1635 -265 1690 -255
rect 1635 -295 1645 -265
rect 1680 -295 1690 -265
rect 1635 -305 1690 -295
rect 1720 -265 1775 -255
rect 1720 -295 1730 -265
rect 1765 -295 1775 -265
rect 1720 -305 1775 -295
rect 1805 -265 1860 -255
rect 1805 -295 1815 -265
rect 1850 -295 1860 -265
rect 1805 -305 1860 -295
rect 1890 -265 1945 -255
rect 1890 -295 1900 -265
rect 1935 -295 1945 -265
rect 1890 -305 1945 -295
rect 1975 -265 2030 -255
rect 1975 -295 1985 -265
rect 2020 -295 2030 -265
rect 1975 -305 2030 -295
rect 2060 -265 2115 -255
rect 2060 -295 2070 -265
rect 2105 -295 2115 -265
rect 2060 -305 2115 -295
rect 2145 -265 2200 -255
rect 2145 -295 2155 -265
rect 2190 -295 2200 -265
rect 2145 -305 2200 -295
rect 2230 -265 2285 -255
rect 2230 -295 2240 -265
rect 2275 -295 2285 -265
rect 2230 -305 2285 -295
rect 2315 -265 2370 -255
rect 2315 -295 2325 -265
rect 2360 -295 2370 -265
rect 2315 -305 2370 -295
rect 2400 -265 2455 -255
rect 2400 -295 2410 -265
rect 2445 -295 2455 -265
rect 2400 -305 2455 -295
rect 2485 -265 2540 -255
rect 2485 -295 2495 -265
rect 2530 -295 2540 -265
rect 2485 -305 2540 -295
rect 2570 -265 2625 -255
rect 2570 -295 2580 -265
rect 2615 -295 2625 -265
rect 2570 -305 2625 -295
rect 2655 -265 2710 -255
rect 2655 -295 2665 -265
rect 2700 -295 2710 -265
rect 2655 -305 2710 -295
rect 2740 -265 2795 -255
rect 2740 -295 2750 -265
rect 2785 -295 2795 -265
rect 2740 -305 2795 -295
rect 2825 -265 2880 -255
rect 2825 -295 2835 -265
rect 2870 -295 2880 -265
rect 2825 -305 2880 -295
rect 2910 -265 2965 -255
rect 2910 -295 2920 -265
rect 2955 -295 2965 -265
rect 2910 -305 2965 -295
rect 2995 -265 3050 -255
rect 2995 -295 3005 -265
rect 3040 -295 3050 -265
rect 2995 -305 3050 -295
rect 3080 -265 3135 -255
rect 3080 -295 3090 -265
rect 3125 -295 3135 -265
rect 3080 -305 3135 -295
rect 3165 -265 3220 -255
rect 3165 -295 3175 -265
rect 3210 -295 3220 -265
rect 3165 -305 3220 -295
rect 3250 -265 3305 -255
rect 3250 -295 3260 -265
rect 3295 -295 3305 -265
rect 3250 -305 3305 -295
rect 3335 -265 3390 -255
rect 3335 -295 3345 -265
rect 3380 -295 3390 -265
rect 3335 -305 3390 -295
rect 3420 -265 3475 -255
rect 3420 -295 3430 -265
rect 3465 -295 3475 -265
rect 3420 -305 3475 -295
rect 3505 -265 3560 -255
rect 3505 -295 3515 -265
rect 3550 -295 3560 -265
rect 3505 -305 3560 -295
rect 3590 -265 3645 -255
rect 3590 -295 3600 -265
rect 3635 -295 3645 -265
rect 3590 -305 3645 -295
rect 3675 -265 3730 -255
rect 3675 -295 3685 -265
rect 3720 -295 3730 -265
rect 3675 -305 3730 -295
rect 3760 -265 3815 -255
rect 3760 -295 3770 -265
rect 3805 -295 3815 -265
rect 3760 -305 3815 -295
rect 3845 -265 3900 -255
rect 3845 -295 3855 -265
rect 3890 -295 3900 -265
rect 3845 -305 3900 -295
rect 3930 -265 3985 -255
rect 3930 -295 3940 -265
rect 3975 -295 3985 -265
rect 3930 -305 3985 -295
rect 4015 -265 4070 -255
rect 4015 -295 4025 -265
rect 4060 -295 4070 -265
rect 4015 -305 4070 -295
rect 4100 -265 4155 -255
rect 4100 -295 4110 -265
rect 4145 -295 4155 -265
rect 4100 -305 4155 -295
rect 4185 -265 4240 -255
rect 4185 -295 4195 -265
rect 4230 -295 4240 -265
rect 4185 -305 4240 -295
rect 4270 -265 4325 -255
rect 4270 -295 4280 -265
rect 4315 -295 4325 -265
rect 4270 -305 4325 -295
rect 4355 -265 4410 -255
rect 4355 -295 4365 -265
rect 4400 -295 4410 -265
rect 4355 -305 4410 -295
rect 4440 -265 4495 -255
rect 4440 -295 4450 -265
rect 4485 -295 4495 -265
rect 4440 -305 4495 -295
rect 4525 -265 4580 -255
rect 4525 -295 4535 -265
rect 4570 -295 4580 -265
rect 4525 -305 4580 -295
rect 4610 -265 4665 -255
rect 4610 -295 4620 -265
rect 4655 -295 4665 -265
rect 4610 -305 4665 -295
rect 4695 -265 4750 -255
rect 4695 -295 4705 -265
rect 4740 -295 4750 -265
rect 4695 -305 4750 -295
rect 4780 -265 4835 -255
rect 4780 -295 4790 -265
rect 4825 -295 4835 -265
rect 4780 -305 4835 -295
rect 4865 -265 4920 -255
rect 4865 -295 4875 -265
rect 4910 -295 4920 -265
rect 4865 -305 4920 -295
rect 4950 -265 5005 -255
rect 4950 -295 4960 -265
rect 4995 -295 5005 -265
rect 4950 -305 5005 -295
rect 5035 -265 5090 -255
rect 5035 -295 5045 -265
rect 5080 -295 5090 -265
rect 5035 -305 5090 -295
rect 5120 -265 5175 -255
rect 5120 -295 5130 -265
rect 5165 -295 5175 -265
rect 5120 -305 5175 -295
rect 5205 -265 5260 -255
rect 5205 -295 5215 -265
rect 5250 -295 5260 -265
rect 5205 -305 5260 -295
rect 5290 -265 5345 -255
rect 5290 -295 5300 -265
rect 5335 -295 5345 -265
rect 5290 -305 5345 -295
rect 5375 -265 5430 -255
rect 5375 -295 5385 -265
rect 5420 -295 5430 -265
rect 5375 -305 5430 -295
rect 5460 -265 5515 -255
rect 5460 -295 5470 -265
rect 5505 -295 5515 -265
rect 5460 -305 5515 -295
rect 5545 -265 5600 -255
rect 5545 -295 5555 -265
rect 5590 -295 5600 -265
rect 5545 -305 5600 -295
rect 5630 -265 5685 -255
rect 5630 -295 5640 -265
rect 5675 -295 5685 -265
rect 5630 -305 5685 -295
rect 5715 -265 5770 -255
rect 5715 -295 5725 -265
rect 5760 -295 5770 -265
rect 5715 -305 5770 -295
rect 5800 -265 5855 -255
rect 5800 -295 5810 -265
rect 5845 -295 5855 -265
rect 5800 -305 5855 -295
rect 5885 -265 5940 -255
rect 5885 -295 5895 -265
rect 5930 -295 5940 -265
rect 5885 -305 5940 -295
rect 5970 -265 6025 -255
rect 5970 -295 5980 -265
rect 6015 -295 6025 -265
rect 5970 -305 6025 -295
rect 6055 -265 6110 -255
rect 6055 -295 6065 -265
rect 6100 -295 6110 -265
rect 6055 -305 6110 -295
rect 6140 -265 6195 -255
rect 6140 -295 6150 -265
rect 6185 -295 6195 -265
rect 6140 -305 6195 -295
rect 6225 -265 6280 -255
rect 6225 -295 6235 -265
rect 6270 -295 6280 -265
rect 6225 -305 6280 -295
rect 6310 -265 6365 -255
rect 6310 -295 6320 -265
rect 6355 -295 6365 -265
rect 6310 -305 6365 -295
rect 6395 -265 6450 -255
rect 6395 -295 6405 -265
rect 6440 -295 6450 -265
rect 6395 -305 6450 -295
rect 6480 -265 6535 -255
rect 6480 -295 6490 -265
rect 6525 -295 6535 -265
rect 6480 -305 6535 -295
rect 6565 -265 6620 -255
rect 6565 -295 6575 -265
rect 6610 -295 6620 -265
rect 6565 -305 6620 -295
rect 6650 -265 6705 -255
rect 6650 -295 6660 -265
rect 6695 -295 6705 -265
rect 6650 -305 6705 -295
rect 6735 -265 6790 -255
rect 6735 -295 6745 -265
rect 6780 -295 6790 -265
rect 6735 -305 6790 -295
rect 6820 -265 6875 -255
rect 6820 -295 6830 -265
rect 6865 -295 6875 -265
rect 6820 -305 6875 -295
rect 6905 -265 6960 -255
rect 6905 -295 6915 -265
rect 6950 -295 6960 -265
rect 6905 -305 6960 -295
rect 6990 -265 7045 -255
rect 6990 -295 7000 -265
rect 7035 -295 7045 -265
rect 6990 -305 7045 -295
rect 7075 -265 7130 -255
rect 7075 -295 7085 -265
rect 7120 -295 7130 -265
rect 7075 -305 7130 -295
rect 7160 -265 7215 -255
rect 7160 -295 7170 -265
rect 7205 -295 7215 -265
rect 7160 -305 7215 -295
rect 7245 -265 7300 -255
rect 7245 -295 7255 -265
rect 7290 -295 7300 -265
rect 7245 -305 7300 -295
rect 7330 -265 7385 -255
rect 7330 -295 7340 -265
rect 7375 -295 7385 -265
rect 7330 -305 7385 -295
rect 7415 -265 7470 -255
rect 7415 -295 7425 -265
rect 7460 -295 7470 -265
rect 7415 -305 7470 -295
rect 7500 -265 7555 -255
rect 7500 -295 7510 -265
rect 7545 -295 7555 -265
rect 7500 -305 7555 -295
rect 7585 -265 7640 -255
rect 7585 -295 7595 -265
rect 7630 -295 7640 -265
rect 7585 -305 7640 -295
rect 7670 -265 7725 -255
rect 7670 -295 7680 -265
rect 7715 -295 7725 -265
rect 7670 -305 7725 -295
rect 7755 -265 7810 -255
rect 7755 -295 7765 -265
rect 7800 -295 7810 -265
rect 7755 -305 7810 -295
rect 7840 -265 7895 -255
rect 7840 -295 7850 -265
rect 7885 -295 7895 -265
rect 7840 -305 7895 -295
rect 7925 -265 7980 -255
rect 7925 -295 7935 -265
rect 7970 -295 7980 -265
rect 7925 -305 7980 -295
rect 8010 -265 8065 -255
rect 8010 -295 8020 -265
rect 8055 -295 8065 -265
rect 8010 -305 8065 -295
rect 8095 -265 8150 -255
rect 8095 -295 8105 -265
rect 8140 -295 8150 -265
rect 8095 -305 8150 -295
rect 8180 -265 8235 -255
rect 8180 -295 8190 -265
rect 8225 -295 8235 -265
rect 8180 -305 8235 -295
rect 8265 -265 8320 -255
rect 8265 -295 8275 -265
rect 8310 -295 8320 -265
rect 8265 -305 8320 -295
rect 8350 -265 8405 -255
rect 8350 -295 8360 -265
rect 8395 -295 8405 -265
rect 8350 -305 8405 -295
rect 8435 -265 8490 -255
rect 8435 -295 8445 -265
rect 8480 -295 8490 -265
rect 8435 -305 8490 -295
rect 8520 -265 8575 -255
rect 8520 -295 8530 -265
rect 8565 -295 8575 -265
rect 8520 -305 8575 -295
rect 8605 -265 8660 -255
rect 8605 -295 8615 -265
rect 8650 -295 8660 -265
rect 8605 -305 8660 -295
rect 8690 -265 8745 -255
rect 8690 -295 8700 -265
rect 8735 -295 8745 -265
rect 8690 -305 8745 -295
rect 8775 -265 8830 -255
rect 8775 -295 8785 -265
rect 8820 -295 8830 -265
rect 8775 -305 8830 -295
rect 8860 -265 8915 -255
rect 8860 -295 8870 -265
rect 8905 -295 8915 -265
rect 8860 -305 8915 -295
rect 8945 -265 9000 -255
rect 8945 -295 8955 -265
rect 8990 -295 9000 -265
rect 8945 -305 9000 -295
rect 9030 -265 9085 -255
rect 9030 -295 9040 -265
rect 9075 -295 9085 -265
rect 9030 -305 9085 -295
rect 9115 -265 9170 -255
rect 9115 -295 9125 -265
rect 9160 -295 9170 -265
rect 9115 -305 9170 -295
rect 9200 -265 9255 -255
rect 9200 -295 9210 -265
rect 9245 -295 9255 -265
rect 9200 -305 9255 -295
rect 9285 -265 9340 -255
rect 9285 -295 9295 -265
rect 9330 -295 9340 -265
rect 9285 -305 9340 -295
rect 9370 -265 9425 -255
rect 9370 -295 9380 -265
rect 9415 -295 9425 -265
rect 9370 -305 9425 -295
rect 9455 -265 9510 -255
rect 9455 -295 9465 -265
rect 9500 -295 9510 -265
rect 9455 -305 9510 -295
rect 9540 -265 9595 -255
rect 9540 -295 9550 -265
rect 9585 -295 9595 -265
rect 9540 -305 9595 -295
rect 9625 -265 9680 -255
rect 9625 -295 9635 -265
rect 9670 -295 9680 -265
rect 9625 -305 9680 -295
rect 9710 -265 9765 -255
rect 9710 -295 9720 -265
rect 9755 -295 9765 -265
rect 9710 -305 9765 -295
rect 9795 -265 9850 -255
rect 9795 -295 9805 -265
rect 9840 -295 9850 -265
rect 9795 -305 9850 -295
rect 9880 -265 9935 -255
rect 9880 -295 9890 -265
rect 9925 -295 9935 -265
rect 9880 -305 9935 -295
rect 9965 -265 10020 -255
rect 9965 -295 9975 -265
rect 10010 -295 10020 -265
rect 9965 -305 10020 -295
rect 10050 -265 10105 -255
rect 10050 -295 10060 -265
rect 10095 -295 10105 -265
rect 10050 -305 10105 -295
rect 10135 -265 10190 -255
rect 10135 -295 10145 -265
rect 10180 -295 10190 -265
rect 10135 -305 10190 -295
rect 10220 -265 10275 -255
rect 10220 -295 10230 -265
rect 10265 -295 10275 -265
rect 10220 -305 10275 -295
rect 10305 -265 10360 -255
rect 10305 -295 10315 -265
rect 10350 -295 10360 -265
rect 10305 -305 10360 -295
rect 10390 -265 10445 -255
rect 10390 -295 10400 -265
rect 10435 -295 10445 -265
rect 10390 -305 10445 -295
rect 10475 -265 10530 -255
rect 10475 -295 10485 -265
rect 10520 -295 10530 -265
rect 10475 -305 10530 -295
rect 10560 -265 10615 -255
rect 10560 -295 10570 -265
rect 10605 -295 10615 -265
rect 10560 -305 10615 -295
rect 10645 -265 10700 -255
rect 10645 -295 10655 -265
rect 10690 -295 10700 -265
rect 10645 -305 10700 -295
rect 10730 -265 10785 -255
rect 10730 -295 10740 -265
rect 10775 -295 10785 -265
rect 10730 -305 10785 -295
rect 10815 -265 10870 -255
rect 10815 -295 10825 -265
rect 10860 -295 10870 -265
rect 10815 -305 10870 -295
rect 10900 -265 10955 -255
rect 10900 -295 10910 -265
rect 10945 -295 10955 -265
rect 10900 -305 10955 -295
rect 10985 -265 11040 -255
rect 10985 -295 10995 -265
rect 11030 -295 11040 -265
rect 10985 -305 11040 -295
rect 11070 -265 11125 -255
rect 11070 -295 11080 -265
rect 11115 -295 11125 -265
rect 11070 -305 11125 -295
rect 11155 -265 11210 -255
rect 11155 -295 11165 -265
rect 11200 -295 11210 -265
rect 11155 -305 11210 -295
rect 11240 -265 11295 -255
rect 11240 -295 11250 -265
rect 11285 -295 11295 -265
rect 11240 -305 11295 -295
rect 11325 -265 11380 -255
rect 11325 -295 11335 -265
rect 11370 -295 11380 -265
rect 11325 -305 11380 -295
rect 11410 -265 11465 -255
rect 11410 -295 11420 -265
rect 11455 -295 11465 -265
rect 11410 -305 11465 -295
rect 11495 -265 11550 -255
rect 11495 -295 11505 -265
rect 11540 -295 11550 -265
rect 11495 -305 11550 -295
rect 11580 -265 11635 -255
rect 11580 -295 11590 -265
rect 11625 -295 11635 -265
rect 11580 -305 11635 -295
rect 11665 -265 11720 -255
rect 11665 -295 11675 -265
rect 11710 -295 11720 -265
rect 11665 -305 11720 -295
rect 11750 -265 11805 -255
rect 11750 -295 11760 -265
rect 11795 -295 11805 -265
rect 11750 -305 11805 -295
rect 11835 -265 11890 -255
rect 11835 -295 11845 -265
rect 11880 -295 11890 -265
rect 11835 -305 11890 -295
rect 11920 -265 11975 -255
rect 11920 -295 11930 -265
rect 11965 -295 11975 -265
rect 11920 -305 11975 -295
rect 12005 -265 12060 -255
rect 12005 -295 12015 -265
rect 12050 -295 12060 -265
rect 12005 -305 12060 -295
rect 12090 -265 12145 -255
rect 12090 -295 12100 -265
rect 12135 -295 12145 -265
rect 12090 -305 12145 -295
rect 12175 -265 12230 -255
rect 12175 -295 12185 -265
rect 12220 -295 12230 -265
rect 12175 -305 12230 -295
rect 12260 -265 12315 -255
rect 12260 -295 12270 -265
rect 12305 -295 12315 -265
rect 12260 -305 12315 -295
rect 12345 -265 12400 -255
rect 12345 -295 12355 -265
rect 12390 -295 12400 -265
rect 12345 -305 12400 -295
rect 12430 -265 12485 -255
rect 12430 -295 12440 -265
rect 12475 -295 12485 -265
rect 12430 -305 12485 -295
rect 12515 -265 12570 -255
rect 12515 -295 12525 -265
rect 12560 -295 12570 -265
rect 12515 -305 12570 -295
rect 12600 -265 12655 -255
rect 12600 -295 12610 -265
rect 12645 -295 12655 -265
rect 12600 -305 12655 -295
rect 12685 -265 12740 -255
rect 12685 -295 12695 -265
rect 12730 -295 12740 -265
rect 12685 -305 12740 -295
rect 12770 -265 12825 -255
rect 12770 -295 12780 -265
rect 12815 -295 12825 -265
rect 12770 -305 12825 -295
rect 12855 -265 12910 -255
rect 12855 -295 12865 -265
rect 12900 -295 12910 -265
rect 12855 -305 12910 -295
rect 12940 -265 12995 -255
rect 12940 -295 12950 -265
rect 12985 -295 12995 -265
rect 12940 -305 12995 -295
rect 13025 -265 13080 -255
rect 13025 -295 13035 -265
rect 13070 -295 13080 -265
rect 13025 -305 13080 -295
rect 13110 -265 13165 -255
rect 13110 -295 13120 -265
rect 13155 -295 13165 -265
rect 13110 -305 13165 -295
rect 13195 -265 13250 -255
rect 13195 -295 13205 -265
rect 13240 -295 13250 -265
rect 13195 -305 13250 -295
rect 13280 -265 13335 -255
rect 13280 -295 13290 -265
rect 13325 -295 13335 -265
rect 13280 -305 13335 -295
rect 13365 -265 13420 -255
rect 13365 -295 13375 -265
rect 13410 -295 13420 -265
rect 13365 -305 13420 -295
rect 13450 -265 13505 -255
rect 13450 -295 13460 -265
rect 13495 -295 13505 -265
rect 13450 -305 13505 -295
rect 13535 -265 13590 -255
rect 13535 -295 13545 -265
rect 13580 -295 13590 -265
rect 13535 -305 13590 -295
rect 13620 -265 13675 -255
rect 13620 -295 13630 -265
rect 13665 -295 13675 -265
rect 13620 -305 13675 -295
rect 13705 -265 13760 -255
rect 13705 -295 13715 -265
rect 13750 -295 13760 -265
rect 13705 -305 13760 -295
rect 13790 -265 13845 -255
rect 13790 -295 13800 -265
rect 13835 -295 13845 -265
rect 13790 -305 13845 -295
rect 13875 -265 13930 -255
rect 13875 -295 13885 -265
rect 13920 -295 13930 -265
rect 13875 -305 13930 -295
rect 13960 -265 14015 -255
rect 13960 -295 13970 -265
rect 14005 -295 14015 -265
rect 13960 -305 14015 -295
rect 14045 -265 14100 -255
rect 14045 -295 14055 -265
rect 14090 -295 14100 -265
rect 14045 -305 14100 -295
rect 14130 -265 14185 -255
rect 14130 -295 14140 -265
rect 14175 -295 14185 -265
rect 14130 -305 14185 -295
rect 14215 -265 14270 -255
rect 14215 -295 14225 -265
rect 14260 -295 14270 -265
rect 14215 -305 14270 -295
rect 14300 -265 14355 -255
rect 14300 -295 14310 -265
rect 14345 -295 14355 -265
rect 14300 -305 14355 -295
rect 14385 -265 14440 -255
rect 14385 -295 14395 -265
rect 14430 -295 14440 -265
rect 14385 -305 14440 -295
rect 14470 -265 14525 -255
rect 14470 -295 14480 -265
rect 14515 -295 14525 -265
rect 14470 -305 14525 -295
rect 14555 -265 14610 -255
rect 14555 -295 14565 -265
rect 14600 -295 14610 -265
rect 14555 -305 14610 -295
rect 14640 -265 14695 -255
rect 14640 -295 14650 -265
rect 14685 -295 14695 -265
rect 14640 -305 14695 -295
rect 14725 -265 14780 -255
rect 14725 -295 14735 -265
rect 14770 -295 14780 -265
rect 14725 -305 14780 -295
rect 14810 -265 14865 -255
rect 14810 -295 14820 -265
rect 14855 -295 14865 -265
rect 14810 -305 14865 -295
rect 14895 -265 14950 -255
rect 14895 -295 14905 -265
rect 14940 -295 14950 -265
rect 14895 -305 14950 -295
rect 14980 -265 15035 -255
rect 14980 -295 14990 -265
rect 15025 -295 15035 -265
rect 14980 -305 15035 -295
rect 15065 -265 15120 -255
rect 15065 -295 15075 -265
rect 15110 -295 15120 -265
rect 15065 -305 15120 -295
rect 15150 -265 15205 -255
rect 15150 -295 15160 -265
rect 15195 -295 15205 -265
rect 15150 -305 15205 -295
rect 15235 -265 15290 -255
rect 15235 -295 15245 -265
rect 15280 -295 15290 -265
rect 15235 -305 15290 -295
rect 15320 -265 15375 -255
rect 15320 -295 15330 -265
rect 15365 -295 15375 -265
rect 15320 -305 15375 -295
rect 15405 -265 15460 -255
rect 15405 -295 15415 -265
rect 15450 -295 15460 -265
rect 15405 -305 15460 -295
rect 15490 -265 15545 -255
rect 15490 -295 15500 -265
rect 15535 -295 15545 -265
rect 15490 -305 15545 -295
rect 15575 -265 15630 -255
rect 15575 -295 15585 -265
rect 15620 -295 15630 -265
rect 15575 -305 15630 -295
rect 15660 -265 15715 -255
rect 15660 -295 15670 -265
rect 15705 -295 15715 -265
rect 15660 -305 15715 -295
rect 15745 -265 15800 -255
rect 15745 -295 15755 -265
rect 15790 -295 15800 -265
rect 15745 -305 15800 -295
rect 15830 -265 15885 -255
rect 15830 -295 15840 -265
rect 15875 -295 15885 -265
rect 15830 -305 15885 -295
rect 15915 -265 15970 -255
rect 15915 -295 15925 -265
rect 15960 -295 15970 -265
rect 15915 -305 15970 -295
rect 16000 -265 16055 -255
rect 16000 -295 16010 -265
rect 16045 -295 16055 -265
rect 16000 -305 16055 -295
rect 16085 -265 16140 -255
rect 16085 -295 16095 -265
rect 16130 -295 16140 -265
rect 16085 -305 16140 -295
rect 16170 -265 16225 -255
rect 16170 -295 16180 -265
rect 16215 -295 16225 -265
rect 16170 -305 16225 -295
rect 16255 -265 16310 -255
rect 16255 -295 16265 -265
rect 16300 -295 16310 -265
rect 16255 -305 16310 -295
rect 16340 -265 16395 -255
rect 16340 -295 16350 -265
rect 16385 -295 16395 -265
rect 16340 -305 16395 -295
rect 16425 -265 16480 -255
rect 16425 -295 16435 -265
rect 16470 -295 16480 -265
rect 16425 -305 16480 -295
rect 16510 -265 16565 -255
rect 16510 -295 16520 -265
rect 16555 -295 16565 -265
rect 16510 -305 16565 -295
rect 16595 -265 16650 -255
rect 16595 -295 16605 -265
rect 16640 -295 16650 -265
rect 16595 -305 16650 -295
rect 16680 -265 16735 -255
rect 16680 -295 16690 -265
rect 16725 -295 16735 -265
rect 16680 -305 16735 -295
rect 16765 -265 16820 -255
rect 16765 -295 16775 -265
rect 16810 -295 16820 -265
rect 16765 -305 16820 -295
rect 16850 -265 16905 -255
rect 16850 -295 16860 -265
rect 16895 -295 16905 -265
rect 16850 -305 16905 -295
rect 16935 -265 16990 -255
rect 16935 -295 16945 -265
rect 16980 -295 16990 -265
rect 16935 -305 16990 -295
rect 17020 -265 17075 -255
rect 17020 -295 17030 -265
rect 17065 -295 17075 -265
rect 17020 -305 17075 -295
rect 17105 -265 17160 -255
rect 17105 -295 17115 -265
rect 17150 -295 17160 -265
rect 17105 -305 17160 -295
rect 17190 -265 17245 -255
rect 17190 -295 17200 -265
rect 17235 -295 17245 -265
rect 17190 -305 17245 -295
rect 17275 -265 17330 -255
rect 17275 -295 17285 -265
rect 17320 -295 17330 -265
rect 17275 -305 17330 -295
rect 17360 -265 17415 -255
rect 17360 -295 17370 -265
rect 17405 -295 17415 -265
rect 17360 -305 17415 -295
rect 17445 -265 17500 -255
rect 17445 -295 17455 -265
rect 17490 -295 17500 -265
rect 17445 -305 17500 -295
rect 17530 -265 17585 -255
rect 17530 -295 17540 -265
rect 17575 -295 17585 -265
rect 17530 -305 17585 -295
rect 17615 -265 17670 -255
rect 17615 -295 17625 -265
rect 17660 -295 17670 -265
rect 17615 -305 17670 -295
rect 17700 -265 17755 -255
rect 17700 -295 17710 -265
rect 17745 -295 17755 -265
rect 17700 -305 17755 -295
rect 17785 -265 17840 -255
rect 17785 -295 17795 -265
rect 17830 -295 17840 -265
rect 17785 -305 17840 -295
rect 17870 -265 17925 -255
rect 17870 -295 17880 -265
rect 17915 -295 17925 -265
rect 17870 -305 17925 -295
rect 17955 -265 18010 -255
rect 17955 -295 17965 -265
rect 18000 -295 18010 -265
rect 17955 -305 18010 -295
rect 18040 -265 18095 -255
rect 18040 -295 18050 -265
rect 18085 -295 18095 -265
rect 18040 -305 18095 -295
rect 18125 -265 18180 -255
rect 18125 -295 18135 -265
rect 18170 -295 18180 -265
rect 18125 -305 18180 -295
rect 18210 -265 18265 -255
rect 18210 -295 18220 -265
rect 18255 -295 18265 -265
rect 18210 -305 18265 -295
rect 18295 -265 18350 -255
rect 18295 -295 18305 -265
rect 18340 -295 18350 -265
rect 18295 -305 18350 -295
rect 18380 -265 18435 -255
rect 18380 -295 18390 -265
rect 18425 -295 18435 -265
rect 18380 -305 18435 -295
rect 18465 -265 18520 -255
rect 18465 -295 18475 -265
rect 18510 -295 18520 -265
rect 18465 -305 18520 -295
rect 18550 -265 18605 -255
rect 18550 -295 18560 -265
rect 18595 -295 18605 -265
rect 18550 -305 18605 -295
rect 18635 -265 18690 -255
rect 18635 -295 18645 -265
rect 18680 -295 18690 -265
rect 18635 -305 18690 -295
rect 18720 -265 18775 -255
rect 18720 -295 18730 -265
rect 18765 -295 18775 -265
rect 18720 -305 18775 -295
rect 18805 -265 18860 -255
rect 18805 -295 18815 -265
rect 18850 -295 18860 -265
rect 18805 -305 18860 -295
rect 18890 -265 18945 -255
rect 18890 -295 18900 -265
rect 18935 -295 18945 -265
rect 18890 -305 18945 -295
rect 18975 -265 19030 -255
rect 18975 -295 18985 -265
rect 19020 -295 19030 -265
rect 18975 -305 19030 -295
rect 19060 -265 19115 -255
rect 19060 -295 19070 -265
rect 19105 -295 19115 -265
rect 19060 -305 19115 -295
rect 19145 -265 19200 -255
rect 19145 -295 19155 -265
rect 19190 -295 19200 -265
rect 19145 -305 19200 -295
rect 19230 -265 19285 -255
rect 19230 -295 19240 -265
rect 19275 -295 19285 -265
rect 19230 -305 19285 -295
rect 19315 -265 19370 -255
rect 19315 -295 19325 -265
rect 19360 -295 19370 -265
rect 19315 -305 19370 -295
rect 19400 -265 19455 -255
rect 19400 -295 19410 -265
rect 19445 -295 19455 -265
rect 19400 -305 19455 -295
rect 19485 -265 19540 -255
rect 19485 -295 19495 -265
rect 19530 -295 19540 -265
rect 19485 -305 19540 -295
rect 19570 -265 19625 -255
rect 19570 -295 19580 -265
rect 19615 -295 19625 -265
rect 19570 -305 19625 -295
rect 19655 -265 19710 -255
rect 19655 -295 19665 -265
rect 19700 -295 19710 -265
rect 19655 -305 19710 -295
rect 19740 -265 19795 -255
rect 19740 -295 19750 -265
rect 19785 -295 19795 -265
rect 19740 -305 19795 -295
rect 19825 -265 19880 -255
rect 19825 -295 19835 -265
rect 19870 -295 19880 -265
rect 19825 -305 19880 -295
rect 19910 -265 19965 -255
rect 19910 -295 19920 -265
rect 19955 -295 19965 -265
rect 19910 -305 19965 -295
rect 19995 -265 20050 -255
rect 19995 -295 20005 -265
rect 20040 -295 20050 -265
rect 19995 -305 20050 -295
rect 20080 -265 20135 -255
rect 20080 -295 20090 -265
rect 20125 -295 20135 -265
rect 20080 -305 20135 -295
rect 20165 -265 20220 -255
rect 20165 -295 20175 -265
rect 20210 -295 20220 -265
rect 20165 -305 20220 -295
rect 20250 -265 20305 -255
rect 20250 -295 20260 -265
rect 20295 -295 20305 -265
rect 20250 -305 20305 -295
rect 20335 -265 20390 -255
rect 20335 -295 20345 -265
rect 20380 -295 20390 -265
rect 20335 -305 20390 -295
rect 20420 -265 20475 -255
rect 20420 -295 20430 -265
rect 20465 -295 20475 -265
rect 20420 -305 20475 -295
rect 20505 -265 20560 -255
rect 20505 -295 20515 -265
rect 20550 -295 20560 -265
rect 20505 -305 20560 -295
rect 20590 -265 20645 -255
rect 20590 -295 20600 -265
rect 20635 -295 20645 -265
rect 20590 -305 20645 -295
rect 20675 -265 20730 -255
rect 20675 -295 20685 -265
rect 20720 -295 20730 -265
rect 20675 -305 20730 -295
rect 20760 -265 20815 -255
rect 20760 -295 20770 -265
rect 20805 -295 20815 -265
rect 20760 -305 20815 -295
rect 20845 -265 20900 -255
rect 20845 -295 20855 -265
rect 20890 -295 20900 -265
rect 20845 -305 20900 -295
rect 20930 -265 20985 -255
rect 20930 -295 20940 -265
rect 20975 -295 20985 -265
rect 20930 -305 20985 -295
rect 21015 -265 21070 -255
rect 21015 -295 21025 -265
rect 21060 -295 21070 -265
rect 21015 -305 21070 -295
rect 21100 -265 21155 -255
rect 21100 -295 21110 -265
rect 21145 -295 21155 -265
rect 21100 -305 21155 -295
rect 21185 -265 21240 -255
rect 21185 -295 21195 -265
rect 21230 -295 21240 -265
rect 21185 -305 21240 -295
rect 21270 -265 21325 -255
rect 21270 -295 21280 -265
rect 21315 -295 21325 -265
rect 21270 -305 21325 -295
rect 21355 -265 21410 -255
rect 21355 -295 21365 -265
rect 21400 -295 21410 -265
rect 21355 -305 21410 -295
rect 21440 -265 21495 -255
rect 21440 -295 21450 -265
rect 21485 -295 21495 -265
rect 21440 -305 21495 -295
rect 21525 -265 21580 -255
rect 21525 -295 21535 -265
rect 21570 -295 21580 -265
rect 21525 -305 21580 -295
rect 21610 -265 21665 -255
rect 21610 -295 21620 -265
rect 21655 -295 21665 -265
rect 21610 -305 21665 -295
rect 21695 -265 21750 -255
rect 21695 -295 21705 -265
rect 21740 -295 21750 -265
rect 21695 -305 21750 -295
rect 21780 -265 21835 -255
rect 21780 -295 21790 -265
rect 21825 -295 21835 -265
rect 21780 -305 21835 -295
rect 21865 -265 21920 -255
rect 21865 -295 21875 -265
rect 21910 -295 21920 -265
rect 21865 -305 21920 -295
rect 21950 -265 22005 -255
rect 21950 -295 21960 -265
rect 21995 -295 22005 -265
rect 21950 -305 22005 -295
rect 22035 -265 22090 -255
rect 22035 -295 22045 -265
rect 22080 -295 22090 -265
rect 22035 -305 22090 -295
rect 22120 -265 22175 -255
rect 22120 -295 22130 -265
rect 22165 -295 22175 -265
rect 22120 -305 22175 -295
rect 22205 -265 22260 -255
rect 22205 -295 22215 -265
rect 22250 -295 22260 -265
rect 22205 -305 22260 -295
rect 22290 -265 22345 -255
rect 22290 -295 22300 -265
rect 22335 -295 22345 -265
rect 22290 -305 22345 -295
rect 22375 -265 22430 -255
rect 22375 -295 22385 -265
rect 22420 -295 22430 -265
rect 22375 -305 22430 -295
rect 22460 -265 22515 -255
rect 22460 -295 22470 -265
rect 22505 -295 22515 -265
rect 22460 -305 22515 -295
rect 22545 -265 22600 -255
rect 22545 -295 22555 -265
rect 22590 -295 22600 -265
rect 22545 -305 22600 -295
rect 22630 -265 22685 -255
rect 22630 -295 22640 -265
rect 22675 -295 22685 -265
rect 22630 -305 22685 -295
rect 22715 -265 22770 -255
rect 22715 -295 22725 -265
rect 22760 -295 22770 -265
rect 22715 -305 22770 -295
rect 22800 -265 22855 -255
rect 22800 -295 22810 -265
rect 22845 -295 22855 -265
rect 22800 -305 22855 -295
rect 22885 -265 22940 -255
rect 22885 -295 22895 -265
rect 22930 -295 22940 -265
rect 22885 -305 22940 -295
rect 22970 -265 23025 -255
rect 22970 -295 22980 -265
rect 23015 -295 23025 -265
rect 22970 -305 23025 -295
rect 23055 -265 23110 -255
rect 23055 -295 23065 -265
rect 23100 -295 23110 -265
rect 23055 -305 23110 -295
rect 23140 -265 23195 -255
rect 23140 -295 23150 -265
rect 23185 -295 23195 -265
rect 23140 -305 23195 -295
rect 23225 -265 23280 -255
rect 23225 -295 23235 -265
rect 23270 -295 23280 -265
rect 23225 -305 23280 -295
rect 23310 -265 23365 -255
rect 23310 -295 23320 -265
rect 23355 -295 23365 -265
rect 23310 -305 23365 -295
rect 23395 -265 23450 -255
rect 23395 -295 23405 -265
rect 23440 -295 23450 -265
rect 23395 -305 23450 -295
rect 23480 -265 23535 -255
rect 23480 -295 23490 -265
rect 23525 -295 23535 -265
rect 23480 -305 23535 -295
rect 23565 -265 23620 -255
rect 23565 -295 23575 -265
rect 23610 -295 23620 -265
rect 23565 -305 23620 -295
rect 23650 -265 23705 -255
rect 23650 -295 23660 -265
rect 23695 -295 23705 -265
rect 23650 -305 23705 -295
rect 23735 -265 23790 -255
rect 23735 -295 23745 -265
rect 23780 -295 23790 -265
rect 23735 -305 23790 -295
rect 23820 -265 23875 -255
rect 23820 -295 23830 -265
rect 23865 -295 23875 -265
rect 23820 -305 23875 -295
rect 23905 -265 23960 -255
rect 23905 -295 23915 -265
rect 23950 -295 23960 -265
rect 23905 -305 23960 -295
rect 23990 -265 24045 -255
rect 23990 -295 24000 -265
rect 24035 -295 24045 -265
rect 23990 -305 24045 -295
rect 24075 -265 24130 -255
rect 24075 -295 24085 -265
rect 24120 -295 24130 -265
rect 24075 -305 24130 -295
rect 24160 -265 24215 -255
rect 24160 -295 24170 -265
rect 24205 -295 24215 -265
rect 24160 -305 24215 -295
rect 24245 -265 24300 -255
rect 24245 -295 24255 -265
rect 24290 -295 24300 -265
rect 24245 -305 24300 -295
rect 24330 -265 24385 -255
rect 24330 -295 24340 -265
rect 24375 -295 24385 -265
rect 24330 -305 24385 -295
rect 24415 -265 24470 -255
rect 24415 -295 24425 -265
rect 24460 -295 24470 -265
rect 24415 -305 24470 -295
rect 24500 -265 24555 -255
rect 24500 -295 24510 -265
rect 24545 -295 24555 -265
rect 24500 -305 24555 -295
rect 24585 -265 24640 -255
rect 24585 -295 24595 -265
rect 24630 -295 24640 -265
rect 24585 -305 24640 -295
rect 24670 -265 24725 -255
rect 24670 -295 24680 -265
rect 24715 -295 24725 -265
rect 24670 -305 24725 -295
rect 24755 -265 24810 -255
rect 24755 -295 24765 -265
rect 24800 -295 24810 -265
rect 24755 -305 24810 -295
rect 24840 -265 24895 -255
rect 24840 -295 24850 -265
rect 24885 -295 24895 -265
rect 24840 -305 24895 -295
rect 24925 -265 24980 -255
rect 24925 -295 24935 -265
rect 24970 -295 24980 -265
rect 24925 -305 24980 -295
rect 25010 -265 25065 -255
rect 25010 -295 25020 -265
rect 25055 -295 25065 -265
rect 25010 -305 25065 -295
rect 25095 -265 25150 -255
rect 25095 -295 25105 -265
rect 25140 -295 25150 -265
rect 25095 -305 25150 -295
rect 25180 -265 25235 -255
rect 25180 -295 25190 -265
rect 25225 -295 25235 -265
rect 25180 -305 25235 -295
rect 25265 -265 25320 -255
rect 25265 -295 25275 -265
rect 25310 -295 25320 -265
rect 25265 -305 25320 -295
rect 25350 -265 25405 -255
rect 25350 -295 25360 -265
rect 25395 -295 25405 -265
rect 25350 -305 25405 -295
rect 25435 -265 25490 -255
rect 25435 -295 25445 -265
rect 25480 -295 25490 -265
rect 25435 -305 25490 -295
rect 25520 -265 25575 -255
rect 25520 -295 25530 -265
rect 25565 -295 25575 -265
rect 25520 -305 25575 -295
rect 25605 -265 25660 -255
rect 25605 -295 25615 -265
rect 25650 -295 25660 -265
rect 25605 -305 25660 -295
rect 25690 -265 25745 -255
rect 25690 -295 25700 -265
rect 25735 -295 25745 -265
rect 25690 -305 25745 -295
rect 25775 -265 25830 -255
rect 25775 -295 25785 -265
rect 25820 -295 25830 -265
rect 25775 -305 25830 -295
rect 25860 -265 25915 -255
rect 25860 -295 25870 -265
rect 25905 -295 25915 -265
rect 25860 -305 25915 -295
rect 25945 -265 26000 -255
rect 25945 -295 25955 -265
rect 25990 -295 26000 -265
rect 25945 -305 26000 -295
rect 26030 -265 26085 -255
rect 26030 -295 26040 -265
rect 26075 -295 26085 -265
rect 26030 -305 26085 -295
rect 26115 -265 26170 -255
rect 26115 -295 26125 -265
rect 26160 -295 26170 -265
rect 26115 -305 26170 -295
rect 26200 -265 26255 -255
rect 26200 -295 26210 -265
rect 26245 -295 26255 -265
rect 26200 -305 26255 -295
rect 26285 -265 26340 -255
rect 26285 -295 26295 -265
rect 26330 -295 26340 -265
rect 26285 -305 26340 -295
rect 26370 -265 26425 -255
rect 26370 -295 26380 -265
rect 26415 -295 26425 -265
rect 26370 -305 26425 -295
rect 26455 -265 26510 -255
rect 26455 -295 26465 -265
rect 26500 -295 26510 -265
rect 26455 -305 26510 -295
rect 26540 -265 26595 -255
rect 26540 -295 26550 -265
rect 26585 -295 26595 -265
rect 26540 -305 26595 -295
rect 26625 -265 26680 -255
rect 26625 -295 26635 -265
rect 26670 -295 26680 -265
rect 26625 -305 26680 -295
rect 26710 -265 26765 -255
rect 26710 -295 26720 -265
rect 26755 -295 26765 -265
rect 26710 -305 26765 -295
rect 26795 -265 26850 -255
rect 26795 -295 26805 -265
rect 26840 -295 26850 -265
rect 26795 -305 26850 -295
rect 26880 -265 26935 -255
rect 26880 -295 26890 -265
rect 26925 -295 26935 -265
rect 26880 -305 26935 -295
rect 26965 -265 27020 -255
rect 26965 -295 26975 -265
rect 27010 -295 27020 -265
rect 26965 -305 27020 -295
rect 27050 -265 27105 -255
rect 27050 -295 27060 -265
rect 27095 -295 27105 -265
rect 27050 -305 27105 -295
rect 27135 -265 27190 -255
rect 27135 -295 27145 -265
rect 27180 -295 27190 -265
rect 27135 -305 27190 -295
rect 27220 -265 27275 -255
rect 27220 -295 27230 -265
rect 27265 -295 27275 -265
rect 27220 -305 27275 -295
rect 27305 -265 27360 -255
rect 27305 -295 27315 -265
rect 27350 -295 27360 -265
rect 27305 -305 27360 -295
rect 27390 -265 27445 -255
rect 27390 -295 27400 -265
rect 27435 -295 27445 -265
rect 27390 -305 27445 -295
rect 27475 -265 27530 -255
rect 27475 -295 27485 -265
rect 27520 -295 27530 -265
rect 27475 -305 27530 -295
rect 27560 -265 27615 -255
rect 27560 -295 27570 -265
rect 27605 -295 27615 -265
rect 27560 -305 27615 -295
rect 27645 -265 27700 -255
rect 27645 -295 27655 -265
rect 27690 -295 27700 -265
rect 27645 -305 27700 -295
rect 27730 -265 27785 -255
rect 27730 -295 27740 -265
rect 27775 -295 27785 -265
rect 27730 -305 27785 -295
rect 27815 -265 27870 -255
rect 27815 -295 27825 -265
rect 27860 -295 27870 -265
rect 27815 -305 27870 -295
rect 27900 -265 27955 -255
rect 27900 -295 27910 -265
rect 27945 -295 27955 -265
rect 27900 -305 27955 -295
rect 27985 -265 28040 -255
rect 27985 -295 27995 -265
rect 28030 -295 28040 -265
rect 27985 -305 28040 -295
rect 28070 -265 28125 -255
rect 28070 -295 28080 -265
rect 28115 -295 28125 -265
rect 28070 -305 28125 -295
rect 28155 -265 28210 -255
rect 28155 -295 28165 -265
rect 28200 -295 28210 -265
rect 28155 -305 28210 -295
rect 28240 -265 28295 -255
rect 28240 -295 28250 -265
rect 28285 -295 28295 -265
rect 28240 -305 28295 -295
rect 28325 -265 28380 -255
rect 28325 -295 28335 -265
rect 28370 -295 28380 -265
rect 28325 -305 28380 -295
rect 28410 -265 28465 -255
rect 28410 -295 28420 -265
rect 28455 -295 28465 -265
rect 28410 -305 28465 -295
rect 28495 -265 28550 -255
rect 28495 -295 28505 -265
rect 28540 -295 28550 -265
rect 28495 -305 28550 -295
rect 28580 -265 28635 -255
rect 28580 -295 28590 -265
rect 28625 -295 28635 -265
rect 28580 -305 28635 -295
rect 28665 -265 28720 -255
rect 28665 -295 28675 -265
rect 28710 -295 28720 -265
rect 28665 -305 28720 -295
rect 28750 -265 28805 -255
rect 28750 -295 28760 -265
rect 28795 -295 28805 -265
rect 28750 -305 28805 -295
rect 28835 -265 28890 -255
rect 28835 -295 28845 -265
rect 28880 -295 28890 -265
rect 28835 -305 28890 -295
rect 28920 -265 28975 -255
rect 28920 -295 28930 -265
rect 28965 -295 28975 -265
rect 28920 -305 28975 -295
rect 29005 -265 29060 -255
rect 29005 -295 29015 -265
rect 29050 -295 29060 -265
rect 29005 -305 29060 -295
rect 29090 -265 29145 -255
rect 29090 -295 29100 -265
rect 29135 -295 29145 -265
rect 29090 -305 29145 -295
rect 29175 -265 29230 -255
rect 29175 -295 29185 -265
rect 29220 -295 29230 -265
rect 29175 -305 29230 -295
rect 29260 -265 29315 -255
rect 29260 -295 29270 -265
rect 29305 -295 29315 -265
rect 29260 -305 29315 -295
rect 29345 -265 29400 -255
rect 29345 -295 29355 -265
rect 29390 -295 29400 -265
rect 29345 -305 29400 -295
rect 29430 -265 29485 -255
rect 29430 -295 29440 -265
rect 29475 -295 29485 -265
rect 29430 -305 29485 -295
rect 29515 -265 29570 -255
rect 29515 -295 29525 -265
rect 29560 -295 29570 -265
rect 29515 -305 29570 -295
rect 29600 -265 29655 -255
rect 29600 -295 29610 -265
rect 29645 -295 29655 -265
rect 29600 -305 29655 -295
rect 29685 -265 29740 -255
rect 29685 -295 29695 -265
rect 29730 -295 29740 -265
rect 29685 -305 29740 -295
rect 29770 -265 29825 -255
rect 29770 -295 29780 -265
rect 29815 -295 29825 -265
rect 29770 -305 29825 -295
rect 29855 -265 29910 -255
rect 29855 -295 29865 -265
rect 29900 -295 29910 -265
rect 29855 -305 29910 -295
rect 29940 -265 29995 -255
rect 29940 -295 29950 -265
rect 29985 -295 29995 -265
rect 29940 -305 29995 -295
rect 30025 -265 30080 -255
rect 30025 -295 30035 -265
rect 30070 -295 30080 -265
rect 30025 -305 30080 -295
rect 30110 -265 30165 -255
rect 30110 -295 30120 -265
rect 30155 -295 30165 -265
rect 30110 -305 30165 -295
rect 30195 -265 30250 -255
rect 30195 -295 30205 -265
rect 30240 -295 30250 -265
rect 30195 -305 30250 -295
rect 30280 -265 30335 -255
rect 30280 -295 30290 -265
rect 30325 -295 30335 -265
rect 30280 -305 30335 -295
rect 30365 -265 30420 -255
rect 30365 -295 30375 -265
rect 30410 -295 30420 -265
rect 30365 -305 30420 -295
rect 30450 -265 30505 -255
rect 30450 -295 30460 -265
rect 30495 -295 30505 -265
rect 30450 -305 30505 -295
rect 30535 -265 30590 -255
rect 30535 -295 30545 -265
rect 30580 -295 30590 -265
rect 30535 -305 30590 -295
rect 30620 -265 30675 -255
rect 30620 -295 30630 -265
rect 30665 -295 30675 -265
rect 30620 -305 30675 -295
rect 30705 -265 30760 -255
rect 30705 -295 30715 -265
rect 30750 -295 30760 -265
rect 30705 -305 30760 -295
rect 30790 -265 30845 -255
rect 30790 -295 30800 -265
rect 30835 -295 30845 -265
rect 30790 -305 30845 -295
rect 30875 -265 30930 -255
rect 30875 -295 30885 -265
rect 30920 -295 30930 -265
rect 30875 -305 30930 -295
rect 30960 -265 31015 -255
rect 30960 -295 30970 -265
rect 31005 -295 31015 -265
rect 30960 -305 31015 -295
rect 31045 -265 31100 -255
rect 31045 -295 31055 -265
rect 31090 -295 31100 -265
rect 31045 -305 31100 -295
rect 31130 -265 31185 -255
rect 31130 -295 31140 -265
rect 31175 -295 31185 -265
rect 31130 -305 31185 -295
rect 31215 -265 31270 -255
rect 31215 -295 31225 -265
rect 31260 -295 31270 -265
rect 31215 -305 31270 -295
rect 31300 -265 31355 -255
rect 31300 -295 31310 -265
rect 31345 -295 31355 -265
rect 31300 -305 31355 -295
rect 31385 -265 31440 -255
rect 31385 -295 31395 -265
rect 31430 -295 31440 -265
rect 31385 -305 31440 -295
rect 31470 -265 31525 -255
rect 31470 -295 31480 -265
rect 31515 -295 31525 -265
rect 31470 -305 31525 -295
rect 31555 -265 31610 -255
rect 31555 -295 31565 -265
rect 31600 -295 31610 -265
rect 31555 -305 31610 -295
rect 31640 -265 31695 -255
rect 31640 -295 31650 -265
rect 31685 -295 31695 -265
rect 31640 -305 31695 -295
rect 31725 -265 31780 -255
rect 31725 -295 31735 -265
rect 31770 -295 31780 -265
rect 31725 -305 31780 -295
rect 31810 -265 31865 -255
rect 31810 -295 31820 -265
rect 31855 -295 31865 -265
rect 31810 -305 31865 -295
rect 31895 -265 31950 -255
rect 31895 -295 31905 -265
rect 31940 -295 31950 -265
rect 31895 -305 31950 -295
rect 31980 -265 32035 -255
rect 31980 -295 31990 -265
rect 32025 -295 32035 -265
rect 31980 -305 32035 -295
rect 32065 -265 32120 -255
rect 32065 -295 32075 -265
rect 32110 -295 32120 -265
rect 32065 -305 32120 -295
rect 32150 -265 32205 -255
rect 32150 -295 32160 -265
rect 32195 -295 32205 -265
rect 32150 -305 32205 -295
rect 32235 -265 32290 -255
rect 32235 -295 32245 -265
rect 32280 -295 32290 -265
rect 32235 -305 32290 -295
rect 32320 -265 32375 -255
rect 32320 -295 32330 -265
rect 32365 -295 32375 -265
rect 32320 -305 32375 -295
rect 32405 -265 32460 -255
rect 32405 -295 32415 -265
rect 32450 -295 32460 -265
rect 32405 -305 32460 -295
rect 32490 -265 32545 -255
rect 32490 -295 32500 -265
rect 32535 -295 32545 -265
rect 32490 -305 32545 -295
rect 32575 -265 32630 -255
rect 32575 -295 32585 -265
rect 32620 -295 32630 -265
rect 32575 -305 32630 -295
rect 32660 -265 32715 -255
rect 32660 -295 32670 -265
rect 32705 -295 32715 -265
rect 32660 -305 32715 -295
rect 32745 -265 32800 -255
rect 32745 -295 32755 -265
rect 32790 -295 32800 -265
rect 32745 -305 32800 -295
rect 32830 -265 32885 -255
rect 32830 -295 32840 -265
rect 32875 -295 32885 -265
rect 32830 -305 32885 -295
rect 32915 -265 32970 -255
rect 32915 -295 32925 -265
rect 32960 -295 32970 -265
rect 32915 -305 32970 -295
rect 33000 -265 33055 -255
rect 33000 -295 33010 -265
rect 33045 -295 33055 -265
rect 33000 -305 33055 -295
rect 33085 -265 33140 -255
rect 33085 -295 33095 -265
rect 33130 -295 33140 -265
rect 33085 -305 33140 -295
rect 33170 -265 33225 -255
rect 33170 -295 33180 -265
rect 33215 -295 33225 -265
rect 33170 -305 33225 -295
rect 33255 -265 33310 -255
rect 33255 -295 33265 -265
rect 33300 -295 33310 -265
rect 33255 -305 33310 -295
rect 33340 -265 33395 -255
rect 33340 -295 33350 -265
rect 33385 -295 33395 -265
rect 33340 -305 33395 -295
rect 33425 -265 33480 -255
rect 33425 -295 33435 -265
rect 33470 -295 33480 -265
rect 33425 -305 33480 -295
rect 33510 -265 33565 -255
rect 33510 -295 33520 -265
rect 33555 -295 33565 -265
rect 33510 -305 33565 -295
rect 33595 -265 33650 -255
rect 33595 -295 33605 -265
rect 33640 -295 33650 -265
rect 33595 -305 33650 -295
rect 33680 -265 33735 -255
rect 33680 -295 33690 -265
rect 33725 -295 33735 -265
rect 33680 -305 33735 -295
rect 33765 -265 33820 -255
rect 33765 -295 33775 -265
rect 33810 -295 33820 -265
rect 33765 -305 33820 -295
rect 33850 -265 33905 -255
rect 33850 -295 33860 -265
rect 33895 -295 33905 -265
rect 33850 -305 33905 -295
rect 33935 -265 33990 -255
rect 33935 -295 33945 -265
rect 33980 -295 33990 -265
rect 33935 -305 33990 -295
rect 34020 -265 34075 -255
rect 34020 -295 34030 -265
rect 34065 -295 34075 -265
rect 34020 -305 34075 -295
rect 34105 -265 34160 -255
rect 34105 -295 34115 -265
rect 34150 -295 34160 -265
rect 34105 -305 34160 -295
rect 34190 -265 34245 -255
rect 34190 -295 34200 -265
rect 34235 -295 34245 -265
rect 34190 -305 34245 -295
rect 34275 -265 34330 -255
rect 34275 -295 34285 -265
rect 34320 -295 34330 -265
rect 34275 -305 34330 -295
rect 34360 -265 34415 -255
rect 34360 -295 34370 -265
rect 34405 -295 34415 -265
rect 34360 -305 34415 -295
rect 34445 -265 34500 -255
rect 34445 -295 34455 -265
rect 34490 -295 34500 -265
rect 34445 -305 34500 -295
rect 34530 -265 34585 -255
rect 34530 -295 34540 -265
rect 34575 -295 34585 -265
rect 34530 -305 34585 -295
rect 34615 -265 34670 -255
rect 34615 -295 34625 -265
rect 34660 -295 34670 -265
rect 34615 -305 34670 -295
rect 34700 -265 34755 -255
rect 34700 -295 34710 -265
rect 34745 -295 34755 -265
rect 34700 -305 34755 -295
rect 34785 -265 34840 -255
rect 34785 -295 34795 -265
rect 34830 -295 34840 -265
rect 34785 -305 34840 -295
rect 34870 -265 34925 -255
rect 34870 -295 34880 -265
rect 34915 -295 34925 -265
rect 34870 -305 34925 -295
rect 34955 -265 35010 -255
rect 34955 -295 34965 -265
rect 35000 -295 35010 -265
rect 34955 -305 35010 -295
rect 35040 -265 35095 -255
rect 35040 -295 35050 -265
rect 35085 -295 35095 -265
rect 35040 -305 35095 -295
rect 35125 -265 35180 -255
rect 35125 -295 35135 -265
rect 35170 -295 35180 -265
rect 35125 -305 35180 -295
rect 35210 -265 35265 -255
rect 35210 -295 35220 -265
rect 35255 -295 35265 -265
rect 35210 -305 35265 -295
rect 35295 -265 35350 -255
rect 35295 -295 35305 -265
rect 35340 -295 35350 -265
rect 35295 -305 35350 -295
rect 35380 -265 35435 -255
rect 35380 -295 35390 -265
rect 35425 -295 35435 -265
rect 35380 -305 35435 -295
rect 35465 -265 35520 -255
rect 35465 -295 35475 -265
rect 35510 -295 35520 -265
rect 35465 -305 35520 -295
rect 35550 -265 35605 -255
rect 35550 -295 35560 -265
rect 35595 -295 35605 -265
rect 35550 -305 35605 -295
rect 35635 -265 35690 -255
rect 35635 -295 35645 -265
rect 35680 -295 35690 -265
rect 35635 -305 35690 -295
rect 35720 -265 35775 -255
rect 35720 -295 35730 -265
rect 35765 -295 35775 -265
rect 35720 -305 35775 -295
rect 35805 -265 35860 -255
rect 35805 -295 35815 -265
rect 35850 -295 35860 -265
rect 35805 -305 35860 -295
rect 35890 -265 35945 -255
rect 35890 -295 35900 -265
rect 35935 -295 35945 -265
rect 35890 -305 35945 -295
rect 35975 -265 36030 -255
rect 35975 -295 35985 -265
rect 36020 -295 36030 -265
rect 35975 -305 36030 -295
rect 36060 -265 36115 -255
rect 36060 -295 36070 -265
rect 36105 -295 36115 -265
rect 36060 -305 36115 -295
rect 36145 -265 36200 -255
rect 36145 -295 36155 -265
rect 36190 -295 36200 -265
rect 36145 -305 36200 -295
rect 36230 -265 36285 -255
rect 36230 -295 36240 -265
rect 36275 -295 36285 -265
rect 36230 -305 36285 -295
rect 36315 -265 36370 -255
rect 36315 -295 36325 -265
rect 36360 -295 36370 -265
rect 36315 -305 36370 -295
rect 36400 -265 36455 -255
rect 36400 -295 36410 -265
rect 36445 -295 36455 -265
rect 36400 -305 36455 -295
rect 36485 -265 36540 -255
rect 36485 -295 36495 -265
rect 36530 -295 36540 -265
rect 36485 -305 36540 -295
rect 36570 -265 36625 -255
rect 36570 -295 36580 -265
rect 36615 -295 36625 -265
rect 36570 -305 36625 -295
rect 36655 -265 36710 -255
rect 36655 -295 36665 -265
rect 36700 -295 36710 -265
rect 36655 -305 36710 -295
rect 36740 -265 36795 -255
rect 36740 -295 36750 -265
rect 36785 -295 36795 -265
rect 36740 -305 36795 -295
rect 36825 -265 36880 -255
rect 36825 -295 36835 -265
rect 36870 -295 36880 -265
rect 36825 -305 36880 -295
rect 36910 -265 36965 -255
rect 36910 -295 36920 -265
rect 36955 -295 36965 -265
rect 36910 -305 36965 -295
rect 36995 -265 37050 -255
rect 36995 -295 37005 -265
rect 37040 -295 37050 -265
rect 36995 -305 37050 -295
rect 37080 -265 37135 -255
rect 37080 -295 37090 -265
rect 37125 -295 37135 -265
rect 37080 -305 37135 -295
rect 37165 -265 37220 -255
rect 37165 -295 37175 -265
rect 37210 -295 37220 -265
rect 37165 -305 37220 -295
rect 37250 -265 37305 -255
rect 37250 -295 37260 -265
rect 37295 -295 37305 -265
rect 37250 -305 37305 -295
rect 37335 -265 37390 -255
rect 37335 -295 37345 -265
rect 37380 -295 37390 -265
rect 37335 -305 37390 -295
rect 37420 -265 37475 -255
rect 37420 -295 37430 -265
rect 37465 -295 37475 -265
rect 37420 -305 37475 -295
rect 37505 -265 37560 -255
rect 37505 -295 37515 -265
rect 37550 -295 37560 -265
rect 37505 -305 37560 -295
rect 37590 -265 37645 -255
rect 37590 -295 37600 -265
rect 37635 -295 37645 -265
rect 37590 -305 37645 -295
rect 37675 -265 37730 -255
rect 37675 -295 37685 -265
rect 37720 -295 37730 -265
rect 37675 -305 37730 -295
rect 37760 -265 37815 -255
rect 37760 -295 37770 -265
rect 37805 -295 37815 -265
rect 37760 -305 37815 -295
rect 37845 -265 37900 -255
rect 37845 -295 37855 -265
rect 37890 -295 37900 -265
rect 37845 -305 37900 -295
rect 37930 -265 37985 -255
rect 37930 -295 37940 -265
rect 37975 -295 37985 -265
rect 37930 -305 37985 -295
rect 38015 -265 38070 -255
rect 38015 -295 38025 -265
rect 38060 -295 38070 -265
rect 38015 -305 38070 -295
rect 38100 -265 38155 -255
rect 38100 -295 38110 -265
rect 38145 -295 38155 -265
rect 38100 -305 38155 -295
rect 38185 -265 38240 -255
rect 38185 -295 38195 -265
rect 38230 -295 38240 -265
rect 38185 -305 38240 -295
rect 38270 -265 38325 -255
rect 38270 -295 38280 -265
rect 38315 -295 38325 -265
rect 38270 -305 38325 -295
rect 38355 -265 38410 -255
rect 38355 -295 38365 -265
rect 38400 -295 38410 -265
rect 38355 -305 38410 -295
rect 38440 -265 38495 -255
rect 38440 -295 38450 -265
rect 38485 -295 38495 -265
rect 38440 -305 38495 -295
rect 38525 -265 38580 -255
rect 38525 -295 38535 -265
rect 38570 -295 38580 -265
rect 38525 -305 38580 -295
rect 38610 -265 38665 -255
rect 38610 -295 38620 -265
rect 38655 -295 38665 -265
rect 38610 -305 38665 -295
rect 38695 -265 38750 -255
rect 38695 -295 38705 -265
rect 38740 -295 38750 -265
rect 38695 -305 38750 -295
rect 38780 -265 38835 -255
rect 38780 -295 38790 -265
rect 38825 -295 38835 -265
rect 38780 -305 38835 -295
rect 38865 -265 38920 -255
rect 38865 -295 38875 -265
rect 38910 -295 38920 -265
rect 38865 -305 38920 -295
rect 38950 -265 39005 -255
rect 38950 -295 38960 -265
rect 38995 -295 39005 -265
rect 38950 -305 39005 -295
rect 39035 -265 39090 -255
rect 39035 -295 39045 -265
rect 39080 -295 39090 -265
rect 39035 -305 39090 -295
rect 39120 -265 39175 -255
rect 39120 -295 39130 -265
rect 39165 -295 39175 -265
rect 39120 -305 39175 -295
rect 39205 -265 39260 -255
rect 39205 -295 39215 -265
rect 39250 -295 39260 -265
rect 39205 -305 39260 -295
rect 39290 -265 39345 -255
rect 39290 -295 39300 -265
rect 39335 -295 39345 -265
rect 39290 -305 39345 -295
rect 39375 -265 39430 -255
rect 39375 -295 39385 -265
rect 39420 -295 39430 -265
rect 39375 -305 39430 -295
rect 39460 -265 39515 -255
rect 39460 -295 39470 -265
rect 39505 -295 39515 -265
rect 39460 -305 39515 -295
rect 39545 -265 39600 -255
rect 39545 -295 39555 -265
rect 39590 -295 39600 -265
rect 39545 -305 39600 -295
rect 39630 -265 39685 -255
rect 39630 -295 39640 -265
rect 39675 -295 39685 -265
rect 39630 -305 39685 -295
rect 39715 -265 39770 -255
rect 39715 -295 39725 -265
rect 39760 -295 39770 -265
rect 39715 -305 39770 -295
rect 39800 -265 39855 -255
rect 39800 -295 39810 -265
rect 39845 -295 39855 -265
rect 39800 -305 39855 -295
rect 39885 -265 39940 -255
rect 39885 -295 39895 -265
rect 39930 -295 39940 -265
rect 39885 -305 39940 -295
rect 39970 -265 40025 -255
rect 39970 -295 39980 -265
rect 40015 -295 40025 -265
rect 39970 -305 40025 -295
rect 40055 -265 40110 -255
rect 40055 -295 40065 -265
rect 40100 -295 40110 -265
rect 40055 -305 40110 -295
rect 40140 -265 40195 -255
rect 40140 -295 40150 -265
rect 40185 -295 40195 -265
rect 40140 -305 40195 -295
rect 40225 -265 40280 -255
rect 40225 -295 40235 -265
rect 40270 -295 40280 -265
rect 40225 -305 40280 -295
rect 40310 -265 40365 -255
rect 40310 -295 40320 -265
rect 40355 -295 40365 -265
rect 40310 -305 40365 -295
rect 40395 -265 40450 -255
rect 40395 -295 40405 -265
rect 40440 -295 40450 -265
rect 40395 -305 40450 -295
rect 40480 -265 40535 -255
rect 40480 -295 40490 -265
rect 40525 -295 40535 -265
rect 40480 -305 40535 -295
rect 40565 -265 40620 -255
rect 40565 -295 40575 -265
rect 40610 -295 40620 -265
rect 40565 -305 40620 -295
rect 40650 -265 40705 -255
rect 40650 -295 40660 -265
rect 40695 -295 40705 -265
rect 40650 -305 40705 -295
rect 40735 -265 40790 -255
rect 40735 -295 40745 -265
rect 40780 -295 40790 -265
rect 40735 -305 40790 -295
rect 40820 -265 40875 -255
rect 40820 -295 40830 -265
rect 40865 -295 40875 -265
rect 40820 -305 40875 -295
rect 40905 -265 40960 -255
rect 40905 -295 40915 -265
rect 40950 -295 40960 -265
rect 40905 -305 40960 -295
rect 40990 -265 41045 -255
rect 40990 -295 41000 -265
rect 41035 -295 41045 -265
rect 40990 -305 41045 -295
rect 41075 -265 41130 -255
rect 41075 -295 41085 -265
rect 41120 -295 41130 -265
rect 41075 -305 41130 -295
rect 41160 -265 41215 -255
rect 41160 -295 41170 -265
rect 41205 -295 41215 -265
rect 41160 -305 41215 -295
rect 41245 -265 41300 -255
rect 41245 -295 41255 -265
rect 41290 -295 41300 -265
rect 41245 -305 41300 -295
rect 41330 -265 41385 -255
rect 41330 -295 41340 -265
rect 41375 -295 41385 -265
rect 41330 -305 41385 -295
rect 41415 -265 41470 -255
rect 41415 -295 41425 -265
rect 41460 -295 41470 -265
rect 41415 -305 41470 -295
rect 41500 -265 41555 -255
rect 41500 -295 41510 -265
rect 41545 -295 41555 -265
rect 41500 -305 41555 -295
rect 41585 -265 41640 -255
rect 41585 -295 41595 -265
rect 41630 -295 41640 -265
rect 41585 -305 41640 -295
rect 41670 -265 41725 -255
rect 41670 -295 41680 -265
rect 41715 -295 41725 -265
rect 41670 -305 41725 -295
rect 41755 -265 41810 -255
rect 41755 -295 41765 -265
rect 41800 -295 41810 -265
rect 41755 -305 41810 -295
rect 41840 -265 41895 -255
rect 41840 -295 41850 -265
rect 41885 -295 41895 -265
rect 41840 -305 41895 -295
rect 41925 -265 41980 -255
rect 41925 -295 41935 -265
rect 41970 -295 41980 -265
rect 41925 -305 41980 -295
rect 42010 -265 42065 -255
rect 42010 -295 42020 -265
rect 42055 -295 42065 -265
rect 42010 -305 42065 -295
rect 42095 -265 42150 -255
rect 42095 -295 42105 -265
rect 42140 -295 42150 -265
rect 42095 -305 42150 -295
rect 42180 -265 42235 -255
rect 42180 -295 42190 -265
rect 42225 -295 42235 -265
rect 42180 -305 42235 -295
rect 42265 -265 42320 -255
rect 42265 -295 42275 -265
rect 42310 -295 42320 -265
rect 42265 -305 42320 -295
rect 42350 -265 42405 -255
rect 42350 -295 42360 -265
rect 42395 -295 42405 -265
rect 42350 -305 42405 -295
rect 42435 -265 42490 -255
rect 42435 -295 42445 -265
rect 42480 -295 42490 -265
rect 42435 -305 42490 -295
rect 42520 -265 42575 -255
rect 42520 -295 42530 -265
rect 42565 -295 42575 -265
rect 42520 -305 42575 -295
rect 42605 -265 42660 -255
rect 42605 -295 42615 -265
rect 42650 -295 42660 -265
rect 42605 -305 42660 -295
rect 42690 -265 42745 -255
rect 42690 -295 42700 -265
rect 42735 -295 42745 -265
rect 42690 -305 42745 -295
rect 42775 -265 42830 -255
rect 42775 -295 42785 -265
rect 42820 -295 42830 -265
rect 42775 -305 42830 -295
rect 42860 -265 42915 -255
rect 42860 -295 42870 -265
rect 42905 -295 42915 -265
rect 42860 -305 42915 -295
rect 42945 -265 43000 -255
rect 42945 -295 42955 -265
rect 42990 -295 43000 -265
rect 42945 -305 43000 -295
rect 43030 -265 43085 -255
rect 43030 -295 43040 -265
rect 43075 -295 43085 -265
rect 43030 -305 43085 -295
rect 43115 -265 43170 -255
rect 43115 -295 43125 -265
rect 43160 -295 43170 -265
rect 43115 -305 43170 -295
rect 43200 -265 43255 -255
rect 43200 -295 43210 -265
rect 43245 -295 43255 -265
rect 43200 -305 43255 -295
rect 43285 -265 43340 -255
rect 43285 -295 43295 -265
rect 43330 -295 43340 -265
rect 43285 -305 43340 -295
rect 43370 -265 43425 -255
rect 43370 -295 43380 -265
rect 43415 -295 43425 -265
rect 43370 -305 43425 -295
rect 43455 -265 43510 -255
rect 43455 -295 43465 -265
rect 43500 -295 43510 -265
rect 43455 -305 43510 -295
rect 43540 -265 43595 -255
rect 43540 -295 43550 -265
rect 43585 -295 43595 -265
rect 43540 -305 43595 -295
rect 65 -335 115 -325
rect 65 -365 75 -335
rect 105 -365 115 -335
rect 65 -385 115 -365
rect 65 -415 75 -385
rect 105 -415 115 -385
rect 65 -425 115 -415
rect 150 -335 200 -325
rect 150 -365 160 -335
rect 190 -365 200 -335
rect 150 -385 200 -365
rect 150 -415 160 -385
rect 190 -415 200 -385
rect 150 -425 200 -415
rect 235 -335 285 -325
rect 235 -365 245 -335
rect 275 -365 285 -335
rect 235 -385 285 -365
rect 235 -415 245 -385
rect 275 -415 285 -385
rect 235 -425 285 -415
rect 320 -335 370 -325
rect 320 -365 330 -335
rect 360 -365 370 -335
rect 320 -385 370 -365
rect 320 -415 330 -385
rect 360 -415 370 -385
rect 320 -425 370 -415
rect 405 -335 455 -325
rect 405 -365 415 -335
rect 445 -365 455 -335
rect 405 -385 455 -365
rect 405 -415 415 -385
rect 445 -415 455 -385
rect 405 -425 455 -415
rect 490 -335 540 -325
rect 490 -365 500 -335
rect 530 -365 540 -335
rect 490 -385 540 -365
rect 490 -415 500 -385
rect 530 -415 540 -385
rect 490 -425 540 -415
rect 575 -335 625 -325
rect 575 -365 585 -335
rect 615 -365 625 -335
rect 575 -385 625 -365
rect 575 -415 585 -385
rect 615 -415 625 -385
rect 575 -425 625 -415
rect 660 -335 710 -325
rect 660 -365 670 -335
rect 700 -365 710 -335
rect 660 -385 710 -365
rect 660 -415 670 -385
rect 700 -415 710 -385
rect 660 -425 710 -415
rect 745 -335 795 -325
rect 745 -365 755 -335
rect 785 -365 795 -335
rect 745 -385 795 -365
rect 745 -415 755 -385
rect 785 -415 795 -385
rect 745 -425 795 -415
rect 830 -335 880 -325
rect 830 -365 840 -335
rect 870 -365 880 -335
rect 830 -385 880 -365
rect 830 -415 840 -385
rect 870 -415 880 -385
rect 830 -425 880 -415
rect 915 -335 965 -325
rect 915 -365 925 -335
rect 955 -365 965 -335
rect 915 -385 965 -365
rect 915 -415 925 -385
rect 955 -415 965 -385
rect 915 -425 965 -415
rect 1000 -335 1050 -325
rect 1000 -365 1010 -335
rect 1040 -365 1050 -335
rect 1000 -385 1050 -365
rect 1000 -415 1010 -385
rect 1040 -415 1050 -385
rect 1000 -425 1050 -415
rect 1085 -335 1135 -325
rect 1085 -365 1095 -335
rect 1125 -365 1135 -335
rect 1085 -385 1135 -365
rect 1085 -415 1095 -385
rect 1125 -415 1135 -385
rect 1085 -425 1135 -415
rect 1170 -335 1220 -325
rect 1170 -365 1180 -335
rect 1210 -365 1220 -335
rect 1170 -385 1220 -365
rect 1170 -415 1180 -385
rect 1210 -415 1220 -385
rect 1170 -425 1220 -415
rect 1255 -335 1305 -325
rect 1255 -365 1265 -335
rect 1295 -365 1305 -335
rect 1255 -385 1305 -365
rect 1255 -415 1265 -385
rect 1295 -415 1305 -385
rect 1255 -425 1305 -415
rect 1340 -335 1390 -325
rect 1340 -365 1350 -335
rect 1380 -365 1390 -335
rect 1340 -385 1390 -365
rect 1340 -415 1350 -385
rect 1380 -415 1390 -385
rect 1340 -425 1390 -415
rect 1425 -335 1475 -325
rect 1425 -365 1435 -335
rect 1465 -365 1475 -335
rect 1425 -385 1475 -365
rect 1425 -415 1435 -385
rect 1465 -415 1475 -385
rect 1425 -425 1475 -415
rect 1510 -335 1560 -325
rect 1510 -365 1520 -335
rect 1550 -365 1560 -335
rect 1510 -385 1560 -365
rect 1510 -415 1520 -385
rect 1550 -415 1560 -385
rect 1510 -425 1560 -415
rect 1595 -335 1645 -325
rect 1595 -365 1605 -335
rect 1635 -365 1645 -335
rect 1595 -385 1645 -365
rect 1595 -415 1605 -385
rect 1635 -415 1645 -385
rect 1595 -425 1645 -415
rect 1680 -335 1730 -325
rect 1680 -365 1690 -335
rect 1720 -365 1730 -335
rect 1680 -385 1730 -365
rect 1680 -415 1690 -385
rect 1720 -415 1730 -385
rect 1680 -425 1730 -415
rect 1765 -335 1815 -325
rect 1765 -365 1775 -335
rect 1805 -365 1815 -335
rect 1765 -385 1815 -365
rect 1765 -415 1775 -385
rect 1805 -415 1815 -385
rect 1765 -425 1815 -415
rect 1850 -335 1900 -325
rect 1850 -365 1860 -335
rect 1890 -365 1900 -335
rect 1850 -385 1900 -365
rect 1850 -415 1860 -385
rect 1890 -415 1900 -385
rect 1850 -425 1900 -415
rect 1935 -335 1985 -325
rect 1935 -365 1945 -335
rect 1975 -365 1985 -335
rect 1935 -385 1985 -365
rect 1935 -415 1945 -385
rect 1975 -415 1985 -385
rect 1935 -425 1985 -415
rect 2020 -335 2070 -325
rect 2020 -365 2030 -335
rect 2060 -365 2070 -335
rect 2020 -385 2070 -365
rect 2020 -415 2030 -385
rect 2060 -415 2070 -385
rect 2020 -425 2070 -415
rect 2105 -335 2155 -325
rect 2105 -365 2115 -335
rect 2145 -365 2155 -335
rect 2105 -385 2155 -365
rect 2105 -415 2115 -385
rect 2145 -415 2155 -385
rect 2105 -425 2155 -415
rect 2190 -335 2240 -325
rect 2190 -365 2200 -335
rect 2230 -365 2240 -335
rect 2190 -385 2240 -365
rect 2190 -415 2200 -385
rect 2230 -415 2240 -385
rect 2190 -425 2240 -415
rect 2275 -335 2325 -325
rect 2275 -365 2285 -335
rect 2315 -365 2325 -335
rect 2275 -385 2325 -365
rect 2275 -415 2285 -385
rect 2315 -415 2325 -385
rect 2275 -425 2325 -415
rect 2360 -335 2410 -325
rect 2360 -365 2370 -335
rect 2400 -365 2410 -335
rect 2360 -385 2410 -365
rect 2360 -415 2370 -385
rect 2400 -415 2410 -385
rect 2360 -425 2410 -415
rect 2445 -335 2495 -325
rect 2445 -365 2455 -335
rect 2485 -365 2495 -335
rect 2445 -385 2495 -365
rect 2445 -415 2455 -385
rect 2485 -415 2495 -385
rect 2445 -425 2495 -415
rect 2530 -335 2580 -325
rect 2530 -365 2540 -335
rect 2570 -365 2580 -335
rect 2530 -385 2580 -365
rect 2530 -415 2540 -385
rect 2570 -415 2580 -385
rect 2530 -425 2580 -415
rect 2615 -335 2665 -325
rect 2615 -365 2625 -335
rect 2655 -365 2665 -335
rect 2615 -385 2665 -365
rect 2615 -415 2625 -385
rect 2655 -415 2665 -385
rect 2615 -425 2665 -415
rect 2700 -335 2750 -325
rect 2700 -365 2710 -335
rect 2740 -365 2750 -335
rect 2700 -385 2750 -365
rect 2700 -415 2710 -385
rect 2740 -415 2750 -385
rect 2700 -425 2750 -415
rect 2785 -335 2835 -325
rect 2785 -365 2795 -335
rect 2825 -365 2835 -335
rect 2785 -385 2835 -365
rect 2785 -415 2795 -385
rect 2825 -415 2835 -385
rect 2785 -425 2835 -415
rect 2870 -335 2920 -325
rect 2870 -365 2880 -335
rect 2910 -365 2920 -335
rect 2870 -385 2920 -365
rect 2870 -415 2880 -385
rect 2910 -415 2920 -385
rect 2870 -425 2920 -415
rect 2955 -335 3005 -325
rect 2955 -365 2965 -335
rect 2995 -365 3005 -335
rect 2955 -385 3005 -365
rect 2955 -415 2965 -385
rect 2995 -415 3005 -385
rect 2955 -425 3005 -415
rect 3040 -335 3090 -325
rect 3040 -365 3050 -335
rect 3080 -365 3090 -335
rect 3040 -385 3090 -365
rect 3040 -415 3050 -385
rect 3080 -415 3090 -385
rect 3040 -425 3090 -415
rect 3125 -335 3175 -325
rect 3125 -365 3135 -335
rect 3165 -365 3175 -335
rect 3125 -385 3175 -365
rect 3125 -415 3135 -385
rect 3165 -415 3175 -385
rect 3125 -425 3175 -415
rect 3210 -335 3260 -325
rect 3210 -365 3220 -335
rect 3250 -365 3260 -335
rect 3210 -385 3260 -365
rect 3210 -415 3220 -385
rect 3250 -415 3260 -385
rect 3210 -425 3260 -415
rect 3295 -335 3345 -325
rect 3295 -365 3305 -335
rect 3335 -365 3345 -335
rect 3295 -385 3345 -365
rect 3295 -415 3305 -385
rect 3335 -415 3345 -385
rect 3295 -425 3345 -415
rect 3380 -335 3430 -325
rect 3380 -365 3390 -335
rect 3420 -365 3430 -335
rect 3380 -385 3430 -365
rect 3380 -415 3390 -385
rect 3420 -415 3430 -385
rect 3380 -425 3430 -415
rect 3465 -335 3515 -325
rect 3465 -365 3475 -335
rect 3505 -365 3515 -335
rect 3465 -385 3515 -365
rect 3465 -415 3475 -385
rect 3505 -415 3515 -385
rect 3465 -425 3515 -415
rect 3550 -335 3600 -325
rect 3550 -365 3560 -335
rect 3590 -365 3600 -335
rect 3550 -385 3600 -365
rect 3550 -415 3560 -385
rect 3590 -415 3600 -385
rect 3550 -425 3600 -415
rect 3635 -335 3685 -325
rect 3635 -365 3645 -335
rect 3675 -365 3685 -335
rect 3635 -385 3685 -365
rect 3635 -415 3645 -385
rect 3675 -415 3685 -385
rect 3635 -425 3685 -415
rect 3720 -335 3770 -325
rect 3720 -365 3730 -335
rect 3760 -365 3770 -335
rect 3720 -385 3770 -365
rect 3720 -415 3730 -385
rect 3760 -415 3770 -385
rect 3720 -425 3770 -415
rect 3805 -335 3855 -325
rect 3805 -365 3815 -335
rect 3845 -365 3855 -335
rect 3805 -385 3855 -365
rect 3805 -415 3815 -385
rect 3845 -415 3855 -385
rect 3805 -425 3855 -415
rect 3890 -335 3940 -325
rect 3890 -365 3900 -335
rect 3930 -365 3940 -335
rect 3890 -385 3940 -365
rect 3890 -415 3900 -385
rect 3930 -415 3940 -385
rect 3890 -425 3940 -415
rect 3975 -335 4025 -325
rect 3975 -365 3985 -335
rect 4015 -365 4025 -335
rect 3975 -385 4025 -365
rect 3975 -415 3985 -385
rect 4015 -415 4025 -385
rect 3975 -425 4025 -415
rect 4060 -335 4110 -325
rect 4060 -365 4070 -335
rect 4100 -365 4110 -335
rect 4060 -385 4110 -365
rect 4060 -415 4070 -385
rect 4100 -415 4110 -385
rect 4060 -425 4110 -415
rect 4145 -335 4195 -325
rect 4145 -365 4155 -335
rect 4185 -365 4195 -335
rect 4145 -385 4195 -365
rect 4145 -415 4155 -385
rect 4185 -415 4195 -385
rect 4145 -425 4195 -415
rect 4230 -335 4280 -325
rect 4230 -365 4240 -335
rect 4270 -365 4280 -335
rect 4230 -385 4280 -365
rect 4230 -415 4240 -385
rect 4270 -415 4280 -385
rect 4230 -425 4280 -415
rect 4315 -335 4365 -325
rect 4315 -365 4325 -335
rect 4355 -365 4365 -335
rect 4315 -385 4365 -365
rect 4315 -415 4325 -385
rect 4355 -415 4365 -385
rect 4315 -425 4365 -415
rect 4400 -335 4450 -325
rect 4400 -365 4410 -335
rect 4440 -365 4450 -335
rect 4400 -385 4450 -365
rect 4400 -415 4410 -385
rect 4440 -415 4450 -385
rect 4400 -425 4450 -415
rect 4485 -335 4535 -325
rect 4485 -365 4495 -335
rect 4525 -365 4535 -335
rect 4485 -385 4535 -365
rect 4485 -415 4495 -385
rect 4525 -415 4535 -385
rect 4485 -425 4535 -415
rect 4570 -335 4620 -325
rect 4570 -365 4580 -335
rect 4610 -365 4620 -335
rect 4570 -385 4620 -365
rect 4570 -415 4580 -385
rect 4610 -415 4620 -385
rect 4570 -425 4620 -415
rect 4655 -335 4705 -325
rect 4655 -365 4665 -335
rect 4695 -365 4705 -335
rect 4655 -385 4705 -365
rect 4655 -415 4665 -385
rect 4695 -415 4705 -385
rect 4655 -425 4705 -415
rect 4740 -335 4790 -325
rect 4740 -365 4750 -335
rect 4780 -365 4790 -335
rect 4740 -385 4790 -365
rect 4740 -415 4750 -385
rect 4780 -415 4790 -385
rect 4740 -425 4790 -415
rect 4825 -335 4875 -325
rect 4825 -365 4835 -335
rect 4865 -365 4875 -335
rect 4825 -385 4875 -365
rect 4825 -415 4835 -385
rect 4865 -415 4875 -385
rect 4825 -425 4875 -415
rect 4910 -335 4960 -325
rect 4910 -365 4920 -335
rect 4950 -365 4960 -335
rect 4910 -385 4960 -365
rect 4910 -415 4920 -385
rect 4950 -415 4960 -385
rect 4910 -425 4960 -415
rect 4995 -335 5045 -325
rect 4995 -365 5005 -335
rect 5035 -365 5045 -335
rect 4995 -385 5045 -365
rect 4995 -415 5005 -385
rect 5035 -415 5045 -385
rect 4995 -425 5045 -415
rect 5080 -335 5130 -325
rect 5080 -365 5090 -335
rect 5120 -365 5130 -335
rect 5080 -385 5130 -365
rect 5080 -415 5090 -385
rect 5120 -415 5130 -385
rect 5080 -425 5130 -415
rect 5165 -335 5215 -325
rect 5165 -365 5175 -335
rect 5205 -365 5215 -335
rect 5165 -385 5215 -365
rect 5165 -415 5175 -385
rect 5205 -415 5215 -385
rect 5165 -425 5215 -415
rect 5250 -335 5300 -325
rect 5250 -365 5260 -335
rect 5290 -365 5300 -335
rect 5250 -385 5300 -365
rect 5250 -415 5260 -385
rect 5290 -415 5300 -385
rect 5250 -425 5300 -415
rect 5335 -335 5385 -325
rect 5335 -365 5345 -335
rect 5375 -365 5385 -335
rect 5335 -385 5385 -365
rect 5335 -415 5345 -385
rect 5375 -415 5385 -385
rect 5335 -425 5385 -415
rect 5420 -335 5470 -325
rect 5420 -365 5430 -335
rect 5460 -365 5470 -335
rect 5420 -385 5470 -365
rect 5420 -415 5430 -385
rect 5460 -415 5470 -385
rect 5420 -425 5470 -415
rect 5505 -335 5555 -325
rect 5505 -365 5515 -335
rect 5545 -365 5555 -335
rect 5505 -385 5555 -365
rect 5505 -415 5515 -385
rect 5545 -415 5555 -385
rect 5505 -425 5555 -415
rect 5590 -335 5640 -325
rect 5590 -365 5600 -335
rect 5630 -365 5640 -335
rect 5590 -385 5640 -365
rect 5590 -415 5600 -385
rect 5630 -415 5640 -385
rect 5590 -425 5640 -415
rect 5675 -335 5725 -325
rect 5675 -365 5685 -335
rect 5715 -365 5725 -335
rect 5675 -385 5725 -365
rect 5675 -415 5685 -385
rect 5715 -415 5725 -385
rect 5675 -425 5725 -415
rect 5760 -335 5810 -325
rect 5760 -365 5770 -335
rect 5800 -365 5810 -335
rect 5760 -385 5810 -365
rect 5760 -415 5770 -385
rect 5800 -415 5810 -385
rect 5760 -425 5810 -415
rect 5845 -335 5895 -325
rect 5845 -365 5855 -335
rect 5885 -365 5895 -335
rect 5845 -385 5895 -365
rect 5845 -415 5855 -385
rect 5885 -415 5895 -385
rect 5845 -425 5895 -415
rect 5930 -335 5980 -325
rect 5930 -365 5940 -335
rect 5970 -365 5980 -335
rect 5930 -385 5980 -365
rect 5930 -415 5940 -385
rect 5970 -415 5980 -385
rect 5930 -425 5980 -415
rect 6015 -335 6065 -325
rect 6015 -365 6025 -335
rect 6055 -365 6065 -335
rect 6015 -385 6065 -365
rect 6015 -415 6025 -385
rect 6055 -415 6065 -385
rect 6015 -425 6065 -415
rect 6100 -335 6150 -325
rect 6100 -365 6110 -335
rect 6140 -365 6150 -335
rect 6100 -385 6150 -365
rect 6100 -415 6110 -385
rect 6140 -415 6150 -385
rect 6100 -425 6150 -415
rect 6185 -335 6235 -325
rect 6185 -365 6195 -335
rect 6225 -365 6235 -335
rect 6185 -385 6235 -365
rect 6185 -415 6195 -385
rect 6225 -415 6235 -385
rect 6185 -425 6235 -415
rect 6270 -335 6320 -325
rect 6270 -365 6280 -335
rect 6310 -365 6320 -335
rect 6270 -385 6320 -365
rect 6270 -415 6280 -385
rect 6310 -415 6320 -385
rect 6270 -425 6320 -415
rect 6355 -335 6405 -325
rect 6355 -365 6365 -335
rect 6395 -365 6405 -335
rect 6355 -385 6405 -365
rect 6355 -415 6365 -385
rect 6395 -415 6405 -385
rect 6355 -425 6405 -415
rect 6440 -335 6490 -325
rect 6440 -365 6450 -335
rect 6480 -365 6490 -335
rect 6440 -385 6490 -365
rect 6440 -415 6450 -385
rect 6480 -415 6490 -385
rect 6440 -425 6490 -415
rect 6525 -335 6575 -325
rect 6525 -365 6535 -335
rect 6565 -365 6575 -335
rect 6525 -385 6575 -365
rect 6525 -415 6535 -385
rect 6565 -415 6575 -385
rect 6525 -425 6575 -415
rect 6610 -335 6660 -325
rect 6610 -365 6620 -335
rect 6650 -365 6660 -335
rect 6610 -385 6660 -365
rect 6610 -415 6620 -385
rect 6650 -415 6660 -385
rect 6610 -425 6660 -415
rect 6695 -335 6745 -325
rect 6695 -365 6705 -335
rect 6735 -365 6745 -335
rect 6695 -385 6745 -365
rect 6695 -415 6705 -385
rect 6735 -415 6745 -385
rect 6695 -425 6745 -415
rect 6780 -335 6830 -325
rect 6780 -365 6790 -335
rect 6820 -365 6830 -335
rect 6780 -385 6830 -365
rect 6780 -415 6790 -385
rect 6820 -415 6830 -385
rect 6780 -425 6830 -415
rect 6865 -335 6915 -325
rect 6865 -365 6875 -335
rect 6905 -365 6915 -335
rect 6865 -385 6915 -365
rect 6865 -415 6875 -385
rect 6905 -415 6915 -385
rect 6865 -425 6915 -415
rect 6950 -335 7000 -325
rect 6950 -365 6960 -335
rect 6990 -365 7000 -335
rect 6950 -385 7000 -365
rect 6950 -415 6960 -385
rect 6990 -415 7000 -385
rect 6950 -425 7000 -415
rect 7035 -335 7085 -325
rect 7035 -365 7045 -335
rect 7075 -365 7085 -335
rect 7035 -385 7085 -365
rect 7035 -415 7045 -385
rect 7075 -415 7085 -385
rect 7035 -425 7085 -415
rect 7120 -335 7170 -325
rect 7120 -365 7130 -335
rect 7160 -365 7170 -335
rect 7120 -385 7170 -365
rect 7120 -415 7130 -385
rect 7160 -415 7170 -385
rect 7120 -425 7170 -415
rect 7205 -335 7255 -325
rect 7205 -365 7215 -335
rect 7245 -365 7255 -335
rect 7205 -385 7255 -365
rect 7205 -415 7215 -385
rect 7245 -415 7255 -385
rect 7205 -425 7255 -415
rect 7290 -335 7340 -325
rect 7290 -365 7300 -335
rect 7330 -365 7340 -335
rect 7290 -385 7340 -365
rect 7290 -415 7300 -385
rect 7330 -415 7340 -385
rect 7290 -425 7340 -415
rect 7375 -335 7425 -325
rect 7375 -365 7385 -335
rect 7415 -365 7425 -335
rect 7375 -385 7425 -365
rect 7375 -415 7385 -385
rect 7415 -415 7425 -385
rect 7375 -425 7425 -415
rect 7460 -335 7510 -325
rect 7460 -365 7470 -335
rect 7500 -365 7510 -335
rect 7460 -385 7510 -365
rect 7460 -415 7470 -385
rect 7500 -415 7510 -385
rect 7460 -425 7510 -415
rect 7545 -335 7595 -325
rect 7545 -365 7555 -335
rect 7585 -365 7595 -335
rect 7545 -385 7595 -365
rect 7545 -415 7555 -385
rect 7585 -415 7595 -385
rect 7545 -425 7595 -415
rect 7630 -335 7680 -325
rect 7630 -365 7640 -335
rect 7670 -365 7680 -335
rect 7630 -385 7680 -365
rect 7630 -415 7640 -385
rect 7670 -415 7680 -385
rect 7630 -425 7680 -415
rect 7715 -335 7765 -325
rect 7715 -365 7725 -335
rect 7755 -365 7765 -335
rect 7715 -385 7765 -365
rect 7715 -415 7725 -385
rect 7755 -415 7765 -385
rect 7715 -425 7765 -415
rect 7800 -335 7850 -325
rect 7800 -365 7810 -335
rect 7840 -365 7850 -335
rect 7800 -385 7850 -365
rect 7800 -415 7810 -385
rect 7840 -415 7850 -385
rect 7800 -425 7850 -415
rect 7885 -335 7935 -325
rect 7885 -365 7895 -335
rect 7925 -365 7935 -335
rect 7885 -385 7935 -365
rect 7885 -415 7895 -385
rect 7925 -415 7935 -385
rect 7885 -425 7935 -415
rect 7970 -335 8020 -325
rect 7970 -365 7980 -335
rect 8010 -365 8020 -335
rect 7970 -385 8020 -365
rect 7970 -415 7980 -385
rect 8010 -415 8020 -385
rect 7970 -425 8020 -415
rect 8055 -335 8105 -325
rect 8055 -365 8065 -335
rect 8095 -365 8105 -335
rect 8055 -385 8105 -365
rect 8055 -415 8065 -385
rect 8095 -415 8105 -385
rect 8055 -425 8105 -415
rect 8140 -335 8190 -325
rect 8140 -365 8150 -335
rect 8180 -365 8190 -335
rect 8140 -385 8190 -365
rect 8140 -415 8150 -385
rect 8180 -415 8190 -385
rect 8140 -425 8190 -415
rect 8225 -335 8275 -325
rect 8225 -365 8235 -335
rect 8265 -365 8275 -335
rect 8225 -385 8275 -365
rect 8225 -415 8235 -385
rect 8265 -415 8275 -385
rect 8225 -425 8275 -415
rect 8310 -335 8360 -325
rect 8310 -365 8320 -335
rect 8350 -365 8360 -335
rect 8310 -385 8360 -365
rect 8310 -415 8320 -385
rect 8350 -415 8360 -385
rect 8310 -425 8360 -415
rect 8395 -335 8445 -325
rect 8395 -365 8405 -335
rect 8435 -365 8445 -335
rect 8395 -385 8445 -365
rect 8395 -415 8405 -385
rect 8435 -415 8445 -385
rect 8395 -425 8445 -415
rect 8480 -335 8530 -325
rect 8480 -365 8490 -335
rect 8520 -365 8530 -335
rect 8480 -385 8530 -365
rect 8480 -415 8490 -385
rect 8520 -415 8530 -385
rect 8480 -425 8530 -415
rect 8565 -335 8615 -325
rect 8565 -365 8575 -335
rect 8605 -365 8615 -335
rect 8565 -385 8615 -365
rect 8565 -415 8575 -385
rect 8605 -415 8615 -385
rect 8565 -425 8615 -415
rect 8650 -335 8700 -325
rect 8650 -365 8660 -335
rect 8690 -365 8700 -335
rect 8650 -385 8700 -365
rect 8650 -415 8660 -385
rect 8690 -415 8700 -385
rect 8650 -425 8700 -415
rect 8735 -335 8785 -325
rect 8735 -365 8745 -335
rect 8775 -365 8785 -335
rect 8735 -385 8785 -365
rect 8735 -415 8745 -385
rect 8775 -415 8785 -385
rect 8735 -425 8785 -415
rect 8820 -335 8870 -325
rect 8820 -365 8830 -335
rect 8860 -365 8870 -335
rect 8820 -385 8870 -365
rect 8820 -415 8830 -385
rect 8860 -415 8870 -385
rect 8820 -425 8870 -415
rect 8905 -335 8955 -325
rect 8905 -365 8915 -335
rect 8945 -365 8955 -335
rect 8905 -385 8955 -365
rect 8905 -415 8915 -385
rect 8945 -415 8955 -385
rect 8905 -425 8955 -415
rect 8990 -335 9040 -325
rect 8990 -365 9000 -335
rect 9030 -365 9040 -335
rect 8990 -385 9040 -365
rect 8990 -415 9000 -385
rect 9030 -415 9040 -385
rect 8990 -425 9040 -415
rect 9075 -335 9125 -325
rect 9075 -365 9085 -335
rect 9115 -365 9125 -335
rect 9075 -385 9125 -365
rect 9075 -415 9085 -385
rect 9115 -415 9125 -385
rect 9075 -425 9125 -415
rect 9160 -335 9210 -325
rect 9160 -365 9170 -335
rect 9200 -365 9210 -335
rect 9160 -385 9210 -365
rect 9160 -415 9170 -385
rect 9200 -415 9210 -385
rect 9160 -425 9210 -415
rect 9245 -335 9295 -325
rect 9245 -365 9255 -335
rect 9285 -365 9295 -335
rect 9245 -385 9295 -365
rect 9245 -415 9255 -385
rect 9285 -415 9295 -385
rect 9245 -425 9295 -415
rect 9330 -335 9380 -325
rect 9330 -365 9340 -335
rect 9370 -365 9380 -335
rect 9330 -385 9380 -365
rect 9330 -415 9340 -385
rect 9370 -415 9380 -385
rect 9330 -425 9380 -415
rect 9415 -335 9465 -325
rect 9415 -365 9425 -335
rect 9455 -365 9465 -335
rect 9415 -385 9465 -365
rect 9415 -415 9425 -385
rect 9455 -415 9465 -385
rect 9415 -425 9465 -415
rect 9500 -335 9550 -325
rect 9500 -365 9510 -335
rect 9540 -365 9550 -335
rect 9500 -385 9550 -365
rect 9500 -415 9510 -385
rect 9540 -415 9550 -385
rect 9500 -425 9550 -415
rect 9585 -335 9635 -325
rect 9585 -365 9595 -335
rect 9625 -365 9635 -335
rect 9585 -385 9635 -365
rect 9585 -415 9595 -385
rect 9625 -415 9635 -385
rect 9585 -425 9635 -415
rect 9670 -335 9720 -325
rect 9670 -365 9680 -335
rect 9710 -365 9720 -335
rect 9670 -385 9720 -365
rect 9670 -415 9680 -385
rect 9710 -415 9720 -385
rect 9670 -425 9720 -415
rect 9755 -335 9805 -325
rect 9755 -365 9765 -335
rect 9795 -365 9805 -335
rect 9755 -385 9805 -365
rect 9755 -415 9765 -385
rect 9795 -415 9805 -385
rect 9755 -425 9805 -415
rect 9840 -335 9890 -325
rect 9840 -365 9850 -335
rect 9880 -365 9890 -335
rect 9840 -385 9890 -365
rect 9840 -415 9850 -385
rect 9880 -415 9890 -385
rect 9840 -425 9890 -415
rect 9925 -335 9975 -325
rect 9925 -365 9935 -335
rect 9965 -365 9975 -335
rect 9925 -385 9975 -365
rect 9925 -415 9935 -385
rect 9965 -415 9975 -385
rect 9925 -425 9975 -415
rect 10010 -335 10060 -325
rect 10010 -365 10020 -335
rect 10050 -365 10060 -335
rect 10010 -385 10060 -365
rect 10010 -415 10020 -385
rect 10050 -415 10060 -385
rect 10010 -425 10060 -415
rect 10095 -335 10145 -325
rect 10095 -365 10105 -335
rect 10135 -365 10145 -335
rect 10095 -385 10145 -365
rect 10095 -415 10105 -385
rect 10135 -415 10145 -385
rect 10095 -425 10145 -415
rect 10180 -335 10230 -325
rect 10180 -365 10190 -335
rect 10220 -365 10230 -335
rect 10180 -385 10230 -365
rect 10180 -415 10190 -385
rect 10220 -415 10230 -385
rect 10180 -425 10230 -415
rect 10265 -335 10315 -325
rect 10265 -365 10275 -335
rect 10305 -365 10315 -335
rect 10265 -385 10315 -365
rect 10265 -415 10275 -385
rect 10305 -415 10315 -385
rect 10265 -425 10315 -415
rect 10350 -335 10400 -325
rect 10350 -365 10360 -335
rect 10390 -365 10400 -335
rect 10350 -385 10400 -365
rect 10350 -415 10360 -385
rect 10390 -415 10400 -385
rect 10350 -425 10400 -415
rect 10435 -335 10485 -325
rect 10435 -365 10445 -335
rect 10475 -365 10485 -335
rect 10435 -385 10485 -365
rect 10435 -415 10445 -385
rect 10475 -415 10485 -385
rect 10435 -425 10485 -415
rect 10520 -335 10570 -325
rect 10520 -365 10530 -335
rect 10560 -365 10570 -335
rect 10520 -385 10570 -365
rect 10520 -415 10530 -385
rect 10560 -415 10570 -385
rect 10520 -425 10570 -415
rect 10605 -335 10655 -325
rect 10605 -365 10615 -335
rect 10645 -365 10655 -335
rect 10605 -385 10655 -365
rect 10605 -415 10615 -385
rect 10645 -415 10655 -385
rect 10605 -425 10655 -415
rect 10690 -335 10740 -325
rect 10690 -365 10700 -335
rect 10730 -365 10740 -335
rect 10690 -385 10740 -365
rect 10690 -415 10700 -385
rect 10730 -415 10740 -385
rect 10690 -425 10740 -415
rect 10775 -335 10825 -325
rect 10775 -365 10785 -335
rect 10815 -365 10825 -335
rect 10775 -385 10825 -365
rect 10775 -415 10785 -385
rect 10815 -415 10825 -385
rect 10775 -425 10825 -415
rect 10860 -335 10910 -325
rect 10860 -365 10870 -335
rect 10900 -365 10910 -335
rect 10860 -385 10910 -365
rect 10860 -415 10870 -385
rect 10900 -415 10910 -385
rect 10860 -425 10910 -415
rect 10945 -335 10995 -325
rect 10945 -365 10955 -335
rect 10985 -365 10995 -335
rect 10945 -385 10995 -365
rect 10945 -415 10955 -385
rect 10985 -415 10995 -385
rect 10945 -425 10995 -415
rect 11030 -335 11080 -325
rect 11030 -365 11040 -335
rect 11070 -365 11080 -335
rect 11030 -385 11080 -365
rect 11030 -415 11040 -385
rect 11070 -415 11080 -385
rect 11030 -425 11080 -415
rect 11115 -335 11165 -325
rect 11115 -365 11125 -335
rect 11155 -365 11165 -335
rect 11115 -385 11165 -365
rect 11115 -415 11125 -385
rect 11155 -415 11165 -385
rect 11115 -425 11165 -415
rect 11200 -335 11250 -325
rect 11200 -365 11210 -335
rect 11240 -365 11250 -335
rect 11200 -385 11250 -365
rect 11200 -415 11210 -385
rect 11240 -415 11250 -385
rect 11200 -425 11250 -415
rect 11285 -335 11335 -325
rect 11285 -365 11295 -335
rect 11325 -365 11335 -335
rect 11285 -385 11335 -365
rect 11285 -415 11295 -385
rect 11325 -415 11335 -385
rect 11285 -425 11335 -415
rect 11370 -335 11420 -325
rect 11370 -365 11380 -335
rect 11410 -365 11420 -335
rect 11370 -385 11420 -365
rect 11370 -415 11380 -385
rect 11410 -415 11420 -385
rect 11370 -425 11420 -415
rect 11455 -335 11505 -325
rect 11455 -365 11465 -335
rect 11495 -365 11505 -335
rect 11455 -385 11505 -365
rect 11455 -415 11465 -385
rect 11495 -415 11505 -385
rect 11455 -425 11505 -415
rect 11540 -335 11590 -325
rect 11540 -365 11550 -335
rect 11580 -365 11590 -335
rect 11540 -385 11590 -365
rect 11540 -415 11550 -385
rect 11580 -415 11590 -385
rect 11540 -425 11590 -415
rect 11625 -335 11675 -325
rect 11625 -365 11635 -335
rect 11665 -365 11675 -335
rect 11625 -385 11675 -365
rect 11625 -415 11635 -385
rect 11665 -415 11675 -385
rect 11625 -425 11675 -415
rect 11710 -335 11760 -325
rect 11710 -365 11720 -335
rect 11750 -365 11760 -335
rect 11710 -385 11760 -365
rect 11710 -415 11720 -385
rect 11750 -415 11760 -385
rect 11710 -425 11760 -415
rect 11795 -335 11845 -325
rect 11795 -365 11805 -335
rect 11835 -365 11845 -335
rect 11795 -385 11845 -365
rect 11795 -415 11805 -385
rect 11835 -415 11845 -385
rect 11795 -425 11845 -415
rect 11880 -335 11930 -325
rect 11880 -365 11890 -335
rect 11920 -365 11930 -335
rect 11880 -385 11930 -365
rect 11880 -415 11890 -385
rect 11920 -415 11930 -385
rect 11880 -425 11930 -415
rect 11965 -335 12015 -325
rect 11965 -365 11975 -335
rect 12005 -365 12015 -335
rect 11965 -385 12015 -365
rect 11965 -415 11975 -385
rect 12005 -415 12015 -385
rect 11965 -425 12015 -415
rect 12050 -335 12100 -325
rect 12050 -365 12060 -335
rect 12090 -365 12100 -335
rect 12050 -385 12100 -365
rect 12050 -415 12060 -385
rect 12090 -415 12100 -385
rect 12050 -425 12100 -415
rect 12135 -335 12185 -325
rect 12135 -365 12145 -335
rect 12175 -365 12185 -335
rect 12135 -385 12185 -365
rect 12135 -415 12145 -385
rect 12175 -415 12185 -385
rect 12135 -425 12185 -415
rect 12220 -335 12270 -325
rect 12220 -365 12230 -335
rect 12260 -365 12270 -335
rect 12220 -385 12270 -365
rect 12220 -415 12230 -385
rect 12260 -415 12270 -385
rect 12220 -425 12270 -415
rect 12305 -335 12355 -325
rect 12305 -365 12315 -335
rect 12345 -365 12355 -335
rect 12305 -385 12355 -365
rect 12305 -415 12315 -385
rect 12345 -415 12355 -385
rect 12305 -425 12355 -415
rect 12390 -335 12440 -325
rect 12390 -365 12400 -335
rect 12430 -365 12440 -335
rect 12390 -385 12440 -365
rect 12390 -415 12400 -385
rect 12430 -415 12440 -385
rect 12390 -425 12440 -415
rect 12475 -335 12525 -325
rect 12475 -365 12485 -335
rect 12515 -365 12525 -335
rect 12475 -385 12525 -365
rect 12475 -415 12485 -385
rect 12515 -415 12525 -385
rect 12475 -425 12525 -415
rect 12560 -335 12610 -325
rect 12560 -365 12570 -335
rect 12600 -365 12610 -335
rect 12560 -385 12610 -365
rect 12560 -415 12570 -385
rect 12600 -415 12610 -385
rect 12560 -425 12610 -415
rect 12645 -335 12695 -325
rect 12645 -365 12655 -335
rect 12685 -365 12695 -335
rect 12645 -385 12695 -365
rect 12645 -415 12655 -385
rect 12685 -415 12695 -385
rect 12645 -425 12695 -415
rect 12730 -335 12780 -325
rect 12730 -365 12740 -335
rect 12770 -365 12780 -335
rect 12730 -385 12780 -365
rect 12730 -415 12740 -385
rect 12770 -415 12780 -385
rect 12730 -425 12780 -415
rect 12815 -335 12865 -325
rect 12815 -365 12825 -335
rect 12855 -365 12865 -335
rect 12815 -385 12865 -365
rect 12815 -415 12825 -385
rect 12855 -415 12865 -385
rect 12815 -425 12865 -415
rect 12900 -335 12950 -325
rect 12900 -365 12910 -335
rect 12940 -365 12950 -335
rect 12900 -385 12950 -365
rect 12900 -415 12910 -385
rect 12940 -415 12950 -385
rect 12900 -425 12950 -415
rect 12985 -335 13035 -325
rect 12985 -365 12995 -335
rect 13025 -365 13035 -335
rect 12985 -385 13035 -365
rect 12985 -415 12995 -385
rect 13025 -415 13035 -385
rect 12985 -425 13035 -415
rect 13070 -335 13120 -325
rect 13070 -365 13080 -335
rect 13110 -365 13120 -335
rect 13070 -385 13120 -365
rect 13070 -415 13080 -385
rect 13110 -415 13120 -385
rect 13070 -425 13120 -415
rect 13155 -335 13205 -325
rect 13155 -365 13165 -335
rect 13195 -365 13205 -335
rect 13155 -385 13205 -365
rect 13155 -415 13165 -385
rect 13195 -415 13205 -385
rect 13155 -425 13205 -415
rect 13240 -335 13290 -325
rect 13240 -365 13250 -335
rect 13280 -365 13290 -335
rect 13240 -385 13290 -365
rect 13240 -415 13250 -385
rect 13280 -415 13290 -385
rect 13240 -425 13290 -415
rect 13325 -335 13375 -325
rect 13325 -365 13335 -335
rect 13365 -365 13375 -335
rect 13325 -385 13375 -365
rect 13325 -415 13335 -385
rect 13365 -415 13375 -385
rect 13325 -425 13375 -415
rect 13410 -335 13460 -325
rect 13410 -365 13420 -335
rect 13450 -365 13460 -335
rect 13410 -385 13460 -365
rect 13410 -415 13420 -385
rect 13450 -415 13460 -385
rect 13410 -425 13460 -415
rect 13495 -335 13545 -325
rect 13495 -365 13505 -335
rect 13535 -365 13545 -335
rect 13495 -385 13545 -365
rect 13495 -415 13505 -385
rect 13535 -415 13545 -385
rect 13495 -425 13545 -415
rect 13580 -335 13630 -325
rect 13580 -365 13590 -335
rect 13620 -365 13630 -335
rect 13580 -385 13630 -365
rect 13580 -415 13590 -385
rect 13620 -415 13630 -385
rect 13580 -425 13630 -415
rect 13665 -335 13715 -325
rect 13665 -365 13675 -335
rect 13705 -365 13715 -335
rect 13665 -385 13715 -365
rect 13665 -415 13675 -385
rect 13705 -415 13715 -385
rect 13665 -425 13715 -415
rect 13750 -335 13800 -325
rect 13750 -365 13760 -335
rect 13790 -365 13800 -335
rect 13750 -385 13800 -365
rect 13750 -415 13760 -385
rect 13790 -415 13800 -385
rect 13750 -425 13800 -415
rect 13835 -335 13885 -325
rect 13835 -365 13845 -335
rect 13875 -365 13885 -335
rect 13835 -385 13885 -365
rect 13835 -415 13845 -385
rect 13875 -415 13885 -385
rect 13835 -425 13885 -415
rect 13920 -335 13970 -325
rect 13920 -365 13930 -335
rect 13960 -365 13970 -335
rect 13920 -385 13970 -365
rect 13920 -415 13930 -385
rect 13960 -415 13970 -385
rect 13920 -425 13970 -415
rect 14005 -335 14055 -325
rect 14005 -365 14015 -335
rect 14045 -365 14055 -335
rect 14005 -385 14055 -365
rect 14005 -415 14015 -385
rect 14045 -415 14055 -385
rect 14005 -425 14055 -415
rect 14090 -335 14140 -325
rect 14090 -365 14100 -335
rect 14130 -365 14140 -335
rect 14090 -385 14140 -365
rect 14090 -415 14100 -385
rect 14130 -415 14140 -385
rect 14090 -425 14140 -415
rect 14175 -335 14225 -325
rect 14175 -365 14185 -335
rect 14215 -365 14225 -335
rect 14175 -385 14225 -365
rect 14175 -415 14185 -385
rect 14215 -415 14225 -385
rect 14175 -425 14225 -415
rect 14260 -335 14310 -325
rect 14260 -365 14270 -335
rect 14300 -365 14310 -335
rect 14260 -385 14310 -365
rect 14260 -415 14270 -385
rect 14300 -415 14310 -385
rect 14260 -425 14310 -415
rect 14345 -335 14395 -325
rect 14345 -365 14355 -335
rect 14385 -365 14395 -335
rect 14345 -385 14395 -365
rect 14345 -415 14355 -385
rect 14385 -415 14395 -385
rect 14345 -425 14395 -415
rect 14430 -335 14480 -325
rect 14430 -365 14440 -335
rect 14470 -365 14480 -335
rect 14430 -385 14480 -365
rect 14430 -415 14440 -385
rect 14470 -415 14480 -385
rect 14430 -425 14480 -415
rect 14515 -335 14565 -325
rect 14515 -365 14525 -335
rect 14555 -365 14565 -335
rect 14515 -385 14565 -365
rect 14515 -415 14525 -385
rect 14555 -415 14565 -385
rect 14515 -425 14565 -415
rect 14600 -335 14650 -325
rect 14600 -365 14610 -335
rect 14640 -365 14650 -335
rect 14600 -385 14650 -365
rect 14600 -415 14610 -385
rect 14640 -415 14650 -385
rect 14600 -425 14650 -415
rect 14685 -335 14735 -325
rect 14685 -365 14695 -335
rect 14725 -365 14735 -335
rect 14685 -385 14735 -365
rect 14685 -415 14695 -385
rect 14725 -415 14735 -385
rect 14685 -425 14735 -415
rect 14770 -335 14820 -325
rect 14770 -365 14780 -335
rect 14810 -365 14820 -335
rect 14770 -385 14820 -365
rect 14770 -415 14780 -385
rect 14810 -415 14820 -385
rect 14770 -425 14820 -415
rect 14855 -335 14905 -325
rect 14855 -365 14865 -335
rect 14895 -365 14905 -335
rect 14855 -385 14905 -365
rect 14855 -415 14865 -385
rect 14895 -415 14905 -385
rect 14855 -425 14905 -415
rect 14940 -335 14990 -325
rect 14940 -365 14950 -335
rect 14980 -365 14990 -335
rect 14940 -385 14990 -365
rect 14940 -415 14950 -385
rect 14980 -415 14990 -385
rect 14940 -425 14990 -415
rect 15025 -335 15075 -325
rect 15025 -365 15035 -335
rect 15065 -365 15075 -335
rect 15025 -385 15075 -365
rect 15025 -415 15035 -385
rect 15065 -415 15075 -385
rect 15025 -425 15075 -415
rect 15110 -335 15160 -325
rect 15110 -365 15120 -335
rect 15150 -365 15160 -335
rect 15110 -385 15160 -365
rect 15110 -415 15120 -385
rect 15150 -415 15160 -385
rect 15110 -425 15160 -415
rect 15195 -335 15245 -325
rect 15195 -365 15205 -335
rect 15235 -365 15245 -335
rect 15195 -385 15245 -365
rect 15195 -415 15205 -385
rect 15235 -415 15245 -385
rect 15195 -425 15245 -415
rect 15280 -335 15330 -325
rect 15280 -365 15290 -335
rect 15320 -365 15330 -335
rect 15280 -385 15330 -365
rect 15280 -415 15290 -385
rect 15320 -415 15330 -385
rect 15280 -425 15330 -415
rect 15365 -335 15415 -325
rect 15365 -365 15375 -335
rect 15405 -365 15415 -335
rect 15365 -385 15415 -365
rect 15365 -415 15375 -385
rect 15405 -415 15415 -385
rect 15365 -425 15415 -415
rect 15450 -335 15500 -325
rect 15450 -365 15460 -335
rect 15490 -365 15500 -335
rect 15450 -385 15500 -365
rect 15450 -415 15460 -385
rect 15490 -415 15500 -385
rect 15450 -425 15500 -415
rect 15535 -335 15585 -325
rect 15535 -365 15545 -335
rect 15575 -365 15585 -335
rect 15535 -385 15585 -365
rect 15535 -415 15545 -385
rect 15575 -415 15585 -385
rect 15535 -425 15585 -415
rect 15620 -335 15670 -325
rect 15620 -365 15630 -335
rect 15660 -365 15670 -335
rect 15620 -385 15670 -365
rect 15620 -415 15630 -385
rect 15660 -415 15670 -385
rect 15620 -425 15670 -415
rect 15705 -335 15755 -325
rect 15705 -365 15715 -335
rect 15745 -365 15755 -335
rect 15705 -385 15755 -365
rect 15705 -415 15715 -385
rect 15745 -415 15755 -385
rect 15705 -425 15755 -415
rect 15790 -335 15840 -325
rect 15790 -365 15800 -335
rect 15830 -365 15840 -335
rect 15790 -385 15840 -365
rect 15790 -415 15800 -385
rect 15830 -415 15840 -385
rect 15790 -425 15840 -415
rect 15875 -335 15925 -325
rect 15875 -365 15885 -335
rect 15915 -365 15925 -335
rect 15875 -385 15925 -365
rect 15875 -415 15885 -385
rect 15915 -415 15925 -385
rect 15875 -425 15925 -415
rect 15960 -335 16010 -325
rect 15960 -365 15970 -335
rect 16000 -365 16010 -335
rect 15960 -385 16010 -365
rect 15960 -415 15970 -385
rect 16000 -415 16010 -385
rect 15960 -425 16010 -415
rect 16045 -335 16095 -325
rect 16045 -365 16055 -335
rect 16085 -365 16095 -335
rect 16045 -385 16095 -365
rect 16045 -415 16055 -385
rect 16085 -415 16095 -385
rect 16045 -425 16095 -415
rect 16130 -335 16180 -325
rect 16130 -365 16140 -335
rect 16170 -365 16180 -335
rect 16130 -385 16180 -365
rect 16130 -415 16140 -385
rect 16170 -415 16180 -385
rect 16130 -425 16180 -415
rect 16215 -335 16265 -325
rect 16215 -365 16225 -335
rect 16255 -365 16265 -335
rect 16215 -385 16265 -365
rect 16215 -415 16225 -385
rect 16255 -415 16265 -385
rect 16215 -425 16265 -415
rect 16300 -335 16350 -325
rect 16300 -365 16310 -335
rect 16340 -365 16350 -335
rect 16300 -385 16350 -365
rect 16300 -415 16310 -385
rect 16340 -415 16350 -385
rect 16300 -425 16350 -415
rect 16385 -335 16435 -325
rect 16385 -365 16395 -335
rect 16425 -365 16435 -335
rect 16385 -385 16435 -365
rect 16385 -415 16395 -385
rect 16425 -415 16435 -385
rect 16385 -425 16435 -415
rect 16470 -335 16520 -325
rect 16470 -365 16480 -335
rect 16510 -365 16520 -335
rect 16470 -385 16520 -365
rect 16470 -415 16480 -385
rect 16510 -415 16520 -385
rect 16470 -425 16520 -415
rect 16555 -335 16605 -325
rect 16555 -365 16565 -335
rect 16595 -365 16605 -335
rect 16555 -385 16605 -365
rect 16555 -415 16565 -385
rect 16595 -415 16605 -385
rect 16555 -425 16605 -415
rect 16640 -335 16690 -325
rect 16640 -365 16650 -335
rect 16680 -365 16690 -335
rect 16640 -385 16690 -365
rect 16640 -415 16650 -385
rect 16680 -415 16690 -385
rect 16640 -425 16690 -415
rect 16725 -335 16775 -325
rect 16725 -365 16735 -335
rect 16765 -365 16775 -335
rect 16725 -385 16775 -365
rect 16725 -415 16735 -385
rect 16765 -415 16775 -385
rect 16725 -425 16775 -415
rect 16810 -335 16860 -325
rect 16810 -365 16820 -335
rect 16850 -365 16860 -335
rect 16810 -385 16860 -365
rect 16810 -415 16820 -385
rect 16850 -415 16860 -385
rect 16810 -425 16860 -415
rect 16895 -335 16945 -325
rect 16895 -365 16905 -335
rect 16935 -365 16945 -335
rect 16895 -385 16945 -365
rect 16895 -415 16905 -385
rect 16935 -415 16945 -385
rect 16895 -425 16945 -415
rect 16980 -335 17030 -325
rect 16980 -365 16990 -335
rect 17020 -365 17030 -335
rect 16980 -385 17030 -365
rect 16980 -415 16990 -385
rect 17020 -415 17030 -385
rect 16980 -425 17030 -415
rect 17065 -335 17115 -325
rect 17065 -365 17075 -335
rect 17105 -365 17115 -335
rect 17065 -385 17115 -365
rect 17065 -415 17075 -385
rect 17105 -415 17115 -385
rect 17065 -425 17115 -415
rect 17150 -335 17200 -325
rect 17150 -365 17160 -335
rect 17190 -365 17200 -335
rect 17150 -385 17200 -365
rect 17150 -415 17160 -385
rect 17190 -415 17200 -385
rect 17150 -425 17200 -415
rect 17235 -335 17285 -325
rect 17235 -365 17245 -335
rect 17275 -365 17285 -335
rect 17235 -385 17285 -365
rect 17235 -415 17245 -385
rect 17275 -415 17285 -385
rect 17235 -425 17285 -415
rect 17320 -335 17370 -325
rect 17320 -365 17330 -335
rect 17360 -365 17370 -335
rect 17320 -385 17370 -365
rect 17320 -415 17330 -385
rect 17360 -415 17370 -385
rect 17320 -425 17370 -415
rect 17405 -335 17455 -325
rect 17405 -365 17415 -335
rect 17445 -365 17455 -335
rect 17405 -385 17455 -365
rect 17405 -415 17415 -385
rect 17445 -415 17455 -385
rect 17405 -425 17455 -415
rect 17490 -335 17540 -325
rect 17490 -365 17500 -335
rect 17530 -365 17540 -335
rect 17490 -385 17540 -365
rect 17490 -415 17500 -385
rect 17530 -415 17540 -385
rect 17490 -425 17540 -415
rect 17575 -335 17625 -325
rect 17575 -365 17585 -335
rect 17615 -365 17625 -335
rect 17575 -385 17625 -365
rect 17575 -415 17585 -385
rect 17615 -415 17625 -385
rect 17575 -425 17625 -415
rect 17660 -335 17710 -325
rect 17660 -365 17670 -335
rect 17700 -365 17710 -335
rect 17660 -385 17710 -365
rect 17660 -415 17670 -385
rect 17700 -415 17710 -385
rect 17660 -425 17710 -415
rect 17745 -335 17795 -325
rect 17745 -365 17755 -335
rect 17785 -365 17795 -335
rect 17745 -385 17795 -365
rect 17745 -415 17755 -385
rect 17785 -415 17795 -385
rect 17745 -425 17795 -415
rect 17830 -335 17880 -325
rect 17830 -365 17840 -335
rect 17870 -365 17880 -335
rect 17830 -385 17880 -365
rect 17830 -415 17840 -385
rect 17870 -415 17880 -385
rect 17830 -425 17880 -415
rect 17915 -335 17965 -325
rect 17915 -365 17925 -335
rect 17955 -365 17965 -335
rect 17915 -385 17965 -365
rect 17915 -415 17925 -385
rect 17955 -415 17965 -385
rect 17915 -425 17965 -415
rect 18000 -335 18050 -325
rect 18000 -365 18010 -335
rect 18040 -365 18050 -335
rect 18000 -385 18050 -365
rect 18000 -415 18010 -385
rect 18040 -415 18050 -385
rect 18000 -425 18050 -415
rect 18085 -335 18135 -325
rect 18085 -365 18095 -335
rect 18125 -365 18135 -335
rect 18085 -385 18135 -365
rect 18085 -415 18095 -385
rect 18125 -415 18135 -385
rect 18085 -425 18135 -415
rect 18170 -335 18220 -325
rect 18170 -365 18180 -335
rect 18210 -365 18220 -335
rect 18170 -385 18220 -365
rect 18170 -415 18180 -385
rect 18210 -415 18220 -385
rect 18170 -425 18220 -415
rect 18255 -335 18305 -325
rect 18255 -365 18265 -335
rect 18295 -365 18305 -335
rect 18255 -385 18305 -365
rect 18255 -415 18265 -385
rect 18295 -415 18305 -385
rect 18255 -425 18305 -415
rect 18340 -335 18390 -325
rect 18340 -365 18350 -335
rect 18380 -365 18390 -335
rect 18340 -385 18390 -365
rect 18340 -415 18350 -385
rect 18380 -415 18390 -385
rect 18340 -425 18390 -415
rect 18425 -335 18475 -325
rect 18425 -365 18435 -335
rect 18465 -365 18475 -335
rect 18425 -385 18475 -365
rect 18425 -415 18435 -385
rect 18465 -415 18475 -385
rect 18425 -425 18475 -415
rect 18510 -335 18560 -325
rect 18510 -365 18520 -335
rect 18550 -365 18560 -335
rect 18510 -385 18560 -365
rect 18510 -415 18520 -385
rect 18550 -415 18560 -385
rect 18510 -425 18560 -415
rect 18595 -335 18645 -325
rect 18595 -365 18605 -335
rect 18635 -365 18645 -335
rect 18595 -385 18645 -365
rect 18595 -415 18605 -385
rect 18635 -415 18645 -385
rect 18595 -425 18645 -415
rect 18680 -335 18730 -325
rect 18680 -365 18690 -335
rect 18720 -365 18730 -335
rect 18680 -385 18730 -365
rect 18680 -415 18690 -385
rect 18720 -415 18730 -385
rect 18680 -425 18730 -415
rect 18765 -335 18815 -325
rect 18765 -365 18775 -335
rect 18805 -365 18815 -335
rect 18765 -385 18815 -365
rect 18765 -415 18775 -385
rect 18805 -415 18815 -385
rect 18765 -425 18815 -415
rect 18850 -335 18900 -325
rect 18850 -365 18860 -335
rect 18890 -365 18900 -335
rect 18850 -385 18900 -365
rect 18850 -415 18860 -385
rect 18890 -415 18900 -385
rect 18850 -425 18900 -415
rect 18935 -335 18985 -325
rect 18935 -365 18945 -335
rect 18975 -365 18985 -335
rect 18935 -385 18985 -365
rect 18935 -415 18945 -385
rect 18975 -415 18985 -385
rect 18935 -425 18985 -415
rect 19020 -335 19070 -325
rect 19020 -365 19030 -335
rect 19060 -365 19070 -335
rect 19020 -385 19070 -365
rect 19020 -415 19030 -385
rect 19060 -415 19070 -385
rect 19020 -425 19070 -415
rect 19105 -335 19155 -325
rect 19105 -365 19115 -335
rect 19145 -365 19155 -335
rect 19105 -385 19155 -365
rect 19105 -415 19115 -385
rect 19145 -415 19155 -385
rect 19105 -425 19155 -415
rect 19190 -335 19240 -325
rect 19190 -365 19200 -335
rect 19230 -365 19240 -335
rect 19190 -385 19240 -365
rect 19190 -415 19200 -385
rect 19230 -415 19240 -385
rect 19190 -425 19240 -415
rect 19275 -335 19325 -325
rect 19275 -365 19285 -335
rect 19315 -365 19325 -335
rect 19275 -385 19325 -365
rect 19275 -415 19285 -385
rect 19315 -415 19325 -385
rect 19275 -425 19325 -415
rect 19360 -335 19410 -325
rect 19360 -365 19370 -335
rect 19400 -365 19410 -335
rect 19360 -385 19410 -365
rect 19360 -415 19370 -385
rect 19400 -415 19410 -385
rect 19360 -425 19410 -415
rect 19445 -335 19495 -325
rect 19445 -365 19455 -335
rect 19485 -365 19495 -335
rect 19445 -385 19495 -365
rect 19445 -415 19455 -385
rect 19485 -415 19495 -385
rect 19445 -425 19495 -415
rect 19530 -335 19580 -325
rect 19530 -365 19540 -335
rect 19570 -365 19580 -335
rect 19530 -385 19580 -365
rect 19530 -415 19540 -385
rect 19570 -415 19580 -385
rect 19530 -425 19580 -415
rect 19615 -335 19665 -325
rect 19615 -365 19625 -335
rect 19655 -365 19665 -335
rect 19615 -385 19665 -365
rect 19615 -415 19625 -385
rect 19655 -415 19665 -385
rect 19615 -425 19665 -415
rect 19700 -335 19750 -325
rect 19700 -365 19710 -335
rect 19740 -365 19750 -335
rect 19700 -385 19750 -365
rect 19700 -415 19710 -385
rect 19740 -415 19750 -385
rect 19700 -425 19750 -415
rect 19785 -335 19835 -325
rect 19785 -365 19795 -335
rect 19825 -365 19835 -335
rect 19785 -385 19835 -365
rect 19785 -415 19795 -385
rect 19825 -415 19835 -385
rect 19785 -425 19835 -415
rect 19870 -335 19920 -325
rect 19870 -365 19880 -335
rect 19910 -365 19920 -335
rect 19870 -385 19920 -365
rect 19870 -415 19880 -385
rect 19910 -415 19920 -385
rect 19870 -425 19920 -415
rect 19955 -335 20005 -325
rect 19955 -365 19965 -335
rect 19995 -365 20005 -335
rect 19955 -385 20005 -365
rect 19955 -415 19965 -385
rect 19995 -415 20005 -385
rect 19955 -425 20005 -415
rect 20040 -335 20090 -325
rect 20040 -365 20050 -335
rect 20080 -365 20090 -335
rect 20040 -385 20090 -365
rect 20040 -415 20050 -385
rect 20080 -415 20090 -385
rect 20040 -425 20090 -415
rect 20125 -335 20175 -325
rect 20125 -365 20135 -335
rect 20165 -365 20175 -335
rect 20125 -385 20175 -365
rect 20125 -415 20135 -385
rect 20165 -415 20175 -385
rect 20125 -425 20175 -415
rect 20210 -335 20260 -325
rect 20210 -365 20220 -335
rect 20250 -365 20260 -335
rect 20210 -385 20260 -365
rect 20210 -415 20220 -385
rect 20250 -415 20260 -385
rect 20210 -425 20260 -415
rect 20295 -335 20345 -325
rect 20295 -365 20305 -335
rect 20335 -365 20345 -335
rect 20295 -385 20345 -365
rect 20295 -415 20305 -385
rect 20335 -415 20345 -385
rect 20295 -425 20345 -415
rect 20380 -335 20430 -325
rect 20380 -365 20390 -335
rect 20420 -365 20430 -335
rect 20380 -385 20430 -365
rect 20380 -415 20390 -385
rect 20420 -415 20430 -385
rect 20380 -425 20430 -415
rect 20465 -335 20515 -325
rect 20465 -365 20475 -335
rect 20505 -365 20515 -335
rect 20465 -385 20515 -365
rect 20465 -415 20475 -385
rect 20505 -415 20515 -385
rect 20465 -425 20515 -415
rect 20550 -335 20600 -325
rect 20550 -365 20560 -335
rect 20590 -365 20600 -335
rect 20550 -385 20600 -365
rect 20550 -415 20560 -385
rect 20590 -415 20600 -385
rect 20550 -425 20600 -415
rect 20635 -335 20685 -325
rect 20635 -365 20645 -335
rect 20675 -365 20685 -335
rect 20635 -385 20685 -365
rect 20635 -415 20645 -385
rect 20675 -415 20685 -385
rect 20635 -425 20685 -415
rect 20720 -335 20770 -325
rect 20720 -365 20730 -335
rect 20760 -365 20770 -335
rect 20720 -385 20770 -365
rect 20720 -415 20730 -385
rect 20760 -415 20770 -385
rect 20720 -425 20770 -415
rect 20805 -335 20855 -325
rect 20805 -365 20815 -335
rect 20845 -365 20855 -335
rect 20805 -385 20855 -365
rect 20805 -415 20815 -385
rect 20845 -415 20855 -385
rect 20805 -425 20855 -415
rect 20890 -335 20940 -325
rect 20890 -365 20900 -335
rect 20930 -365 20940 -335
rect 20890 -385 20940 -365
rect 20890 -415 20900 -385
rect 20930 -415 20940 -385
rect 20890 -425 20940 -415
rect 20975 -335 21025 -325
rect 20975 -365 20985 -335
rect 21015 -365 21025 -335
rect 20975 -385 21025 -365
rect 20975 -415 20985 -385
rect 21015 -415 21025 -385
rect 20975 -425 21025 -415
rect 21060 -335 21110 -325
rect 21060 -365 21070 -335
rect 21100 -365 21110 -335
rect 21060 -385 21110 -365
rect 21060 -415 21070 -385
rect 21100 -415 21110 -385
rect 21060 -425 21110 -415
rect 21145 -335 21195 -325
rect 21145 -365 21155 -335
rect 21185 -365 21195 -335
rect 21145 -385 21195 -365
rect 21145 -415 21155 -385
rect 21185 -415 21195 -385
rect 21145 -425 21195 -415
rect 21230 -335 21280 -325
rect 21230 -365 21240 -335
rect 21270 -365 21280 -335
rect 21230 -385 21280 -365
rect 21230 -415 21240 -385
rect 21270 -415 21280 -385
rect 21230 -425 21280 -415
rect 21315 -335 21365 -325
rect 21315 -365 21325 -335
rect 21355 -365 21365 -335
rect 21315 -385 21365 -365
rect 21315 -415 21325 -385
rect 21355 -415 21365 -385
rect 21315 -425 21365 -415
rect 21400 -335 21450 -325
rect 21400 -365 21410 -335
rect 21440 -365 21450 -335
rect 21400 -385 21450 -365
rect 21400 -415 21410 -385
rect 21440 -415 21450 -385
rect 21400 -425 21450 -415
rect 21485 -335 21535 -325
rect 21485 -365 21495 -335
rect 21525 -365 21535 -335
rect 21485 -385 21535 -365
rect 21485 -415 21495 -385
rect 21525 -415 21535 -385
rect 21485 -425 21535 -415
rect 21570 -335 21620 -325
rect 21570 -365 21580 -335
rect 21610 -365 21620 -335
rect 21570 -385 21620 -365
rect 21570 -415 21580 -385
rect 21610 -415 21620 -385
rect 21570 -425 21620 -415
rect 21655 -335 21705 -325
rect 21655 -365 21665 -335
rect 21695 -365 21705 -335
rect 21655 -385 21705 -365
rect 21655 -415 21665 -385
rect 21695 -415 21705 -385
rect 21655 -425 21705 -415
rect 21740 -335 21790 -325
rect 21740 -365 21750 -335
rect 21780 -365 21790 -335
rect 21740 -385 21790 -365
rect 21740 -415 21750 -385
rect 21780 -415 21790 -385
rect 21740 -425 21790 -415
rect 21825 -335 21875 -325
rect 21825 -365 21835 -335
rect 21865 -365 21875 -335
rect 21825 -385 21875 -365
rect 21825 -415 21835 -385
rect 21865 -415 21875 -385
rect 21825 -425 21875 -415
rect 21910 -335 21960 -325
rect 21910 -365 21920 -335
rect 21950 -365 21960 -335
rect 21910 -385 21960 -365
rect 21910 -415 21920 -385
rect 21950 -415 21960 -385
rect 21910 -425 21960 -415
rect 21995 -335 22045 -325
rect 21995 -365 22005 -335
rect 22035 -365 22045 -335
rect 21995 -385 22045 -365
rect 21995 -415 22005 -385
rect 22035 -415 22045 -385
rect 21995 -425 22045 -415
rect 22080 -335 22130 -325
rect 22080 -365 22090 -335
rect 22120 -365 22130 -335
rect 22080 -385 22130 -365
rect 22080 -415 22090 -385
rect 22120 -415 22130 -385
rect 22080 -425 22130 -415
rect 22165 -335 22215 -325
rect 22165 -365 22175 -335
rect 22205 -365 22215 -335
rect 22165 -385 22215 -365
rect 22165 -415 22175 -385
rect 22205 -415 22215 -385
rect 22165 -425 22215 -415
rect 22250 -335 22300 -325
rect 22250 -365 22260 -335
rect 22290 -365 22300 -335
rect 22250 -385 22300 -365
rect 22250 -415 22260 -385
rect 22290 -415 22300 -385
rect 22250 -425 22300 -415
rect 22335 -335 22385 -325
rect 22335 -365 22345 -335
rect 22375 -365 22385 -335
rect 22335 -385 22385 -365
rect 22335 -415 22345 -385
rect 22375 -415 22385 -385
rect 22335 -425 22385 -415
rect 22420 -335 22470 -325
rect 22420 -365 22430 -335
rect 22460 -365 22470 -335
rect 22420 -385 22470 -365
rect 22420 -415 22430 -385
rect 22460 -415 22470 -385
rect 22420 -425 22470 -415
rect 22505 -335 22555 -325
rect 22505 -365 22515 -335
rect 22545 -365 22555 -335
rect 22505 -385 22555 -365
rect 22505 -415 22515 -385
rect 22545 -415 22555 -385
rect 22505 -425 22555 -415
rect 22590 -335 22640 -325
rect 22590 -365 22600 -335
rect 22630 -365 22640 -335
rect 22590 -385 22640 -365
rect 22590 -415 22600 -385
rect 22630 -415 22640 -385
rect 22590 -425 22640 -415
rect 22675 -335 22725 -325
rect 22675 -365 22685 -335
rect 22715 -365 22725 -335
rect 22675 -385 22725 -365
rect 22675 -415 22685 -385
rect 22715 -415 22725 -385
rect 22675 -425 22725 -415
rect 22760 -335 22810 -325
rect 22760 -365 22770 -335
rect 22800 -365 22810 -335
rect 22760 -385 22810 -365
rect 22760 -415 22770 -385
rect 22800 -415 22810 -385
rect 22760 -425 22810 -415
rect 22845 -335 22895 -325
rect 22845 -365 22855 -335
rect 22885 -365 22895 -335
rect 22845 -385 22895 -365
rect 22845 -415 22855 -385
rect 22885 -415 22895 -385
rect 22845 -425 22895 -415
rect 22930 -335 22980 -325
rect 22930 -365 22940 -335
rect 22970 -365 22980 -335
rect 22930 -385 22980 -365
rect 22930 -415 22940 -385
rect 22970 -415 22980 -385
rect 22930 -425 22980 -415
rect 23015 -335 23065 -325
rect 23015 -365 23025 -335
rect 23055 -365 23065 -335
rect 23015 -385 23065 -365
rect 23015 -415 23025 -385
rect 23055 -415 23065 -385
rect 23015 -425 23065 -415
rect 23100 -335 23150 -325
rect 23100 -365 23110 -335
rect 23140 -365 23150 -335
rect 23100 -385 23150 -365
rect 23100 -415 23110 -385
rect 23140 -415 23150 -385
rect 23100 -425 23150 -415
rect 23185 -335 23235 -325
rect 23185 -365 23195 -335
rect 23225 -365 23235 -335
rect 23185 -385 23235 -365
rect 23185 -415 23195 -385
rect 23225 -415 23235 -385
rect 23185 -425 23235 -415
rect 23270 -335 23320 -325
rect 23270 -365 23280 -335
rect 23310 -365 23320 -335
rect 23270 -385 23320 -365
rect 23270 -415 23280 -385
rect 23310 -415 23320 -385
rect 23270 -425 23320 -415
rect 23355 -335 23405 -325
rect 23355 -365 23365 -335
rect 23395 -365 23405 -335
rect 23355 -385 23405 -365
rect 23355 -415 23365 -385
rect 23395 -415 23405 -385
rect 23355 -425 23405 -415
rect 23440 -335 23490 -325
rect 23440 -365 23450 -335
rect 23480 -365 23490 -335
rect 23440 -385 23490 -365
rect 23440 -415 23450 -385
rect 23480 -415 23490 -385
rect 23440 -425 23490 -415
rect 23525 -335 23575 -325
rect 23525 -365 23535 -335
rect 23565 -365 23575 -335
rect 23525 -385 23575 -365
rect 23525 -415 23535 -385
rect 23565 -415 23575 -385
rect 23525 -425 23575 -415
rect 23610 -335 23660 -325
rect 23610 -365 23620 -335
rect 23650 -365 23660 -335
rect 23610 -385 23660 -365
rect 23610 -415 23620 -385
rect 23650 -415 23660 -385
rect 23610 -425 23660 -415
rect 23695 -335 23745 -325
rect 23695 -365 23705 -335
rect 23735 -365 23745 -335
rect 23695 -385 23745 -365
rect 23695 -415 23705 -385
rect 23735 -415 23745 -385
rect 23695 -425 23745 -415
rect 23780 -335 23830 -325
rect 23780 -365 23790 -335
rect 23820 -365 23830 -335
rect 23780 -385 23830 -365
rect 23780 -415 23790 -385
rect 23820 -415 23830 -385
rect 23780 -425 23830 -415
rect 23865 -335 23915 -325
rect 23865 -365 23875 -335
rect 23905 -365 23915 -335
rect 23865 -385 23915 -365
rect 23865 -415 23875 -385
rect 23905 -415 23915 -385
rect 23865 -425 23915 -415
rect 23950 -335 24000 -325
rect 23950 -365 23960 -335
rect 23990 -365 24000 -335
rect 23950 -385 24000 -365
rect 23950 -415 23960 -385
rect 23990 -415 24000 -385
rect 23950 -425 24000 -415
rect 24035 -335 24085 -325
rect 24035 -365 24045 -335
rect 24075 -365 24085 -335
rect 24035 -385 24085 -365
rect 24035 -415 24045 -385
rect 24075 -415 24085 -385
rect 24035 -425 24085 -415
rect 24120 -335 24170 -325
rect 24120 -365 24130 -335
rect 24160 -365 24170 -335
rect 24120 -385 24170 -365
rect 24120 -415 24130 -385
rect 24160 -415 24170 -385
rect 24120 -425 24170 -415
rect 24205 -335 24255 -325
rect 24205 -365 24215 -335
rect 24245 -365 24255 -335
rect 24205 -385 24255 -365
rect 24205 -415 24215 -385
rect 24245 -415 24255 -385
rect 24205 -425 24255 -415
rect 24290 -335 24340 -325
rect 24290 -365 24300 -335
rect 24330 -365 24340 -335
rect 24290 -385 24340 -365
rect 24290 -415 24300 -385
rect 24330 -415 24340 -385
rect 24290 -425 24340 -415
rect 24375 -335 24425 -325
rect 24375 -365 24385 -335
rect 24415 -365 24425 -335
rect 24375 -385 24425 -365
rect 24375 -415 24385 -385
rect 24415 -415 24425 -385
rect 24375 -425 24425 -415
rect 24460 -335 24510 -325
rect 24460 -365 24470 -335
rect 24500 -365 24510 -335
rect 24460 -385 24510 -365
rect 24460 -415 24470 -385
rect 24500 -415 24510 -385
rect 24460 -425 24510 -415
rect 24545 -335 24595 -325
rect 24545 -365 24555 -335
rect 24585 -365 24595 -335
rect 24545 -385 24595 -365
rect 24545 -415 24555 -385
rect 24585 -415 24595 -385
rect 24545 -425 24595 -415
rect 24630 -335 24680 -325
rect 24630 -365 24640 -335
rect 24670 -365 24680 -335
rect 24630 -385 24680 -365
rect 24630 -415 24640 -385
rect 24670 -415 24680 -385
rect 24630 -425 24680 -415
rect 24715 -335 24765 -325
rect 24715 -365 24725 -335
rect 24755 -365 24765 -335
rect 24715 -385 24765 -365
rect 24715 -415 24725 -385
rect 24755 -415 24765 -385
rect 24715 -425 24765 -415
rect 24800 -335 24850 -325
rect 24800 -365 24810 -335
rect 24840 -365 24850 -335
rect 24800 -385 24850 -365
rect 24800 -415 24810 -385
rect 24840 -415 24850 -385
rect 24800 -425 24850 -415
rect 24885 -335 24935 -325
rect 24885 -365 24895 -335
rect 24925 -365 24935 -335
rect 24885 -385 24935 -365
rect 24885 -415 24895 -385
rect 24925 -415 24935 -385
rect 24885 -425 24935 -415
rect 24970 -335 25020 -325
rect 24970 -365 24980 -335
rect 25010 -365 25020 -335
rect 24970 -385 25020 -365
rect 24970 -415 24980 -385
rect 25010 -415 25020 -385
rect 24970 -425 25020 -415
rect 25055 -335 25105 -325
rect 25055 -365 25065 -335
rect 25095 -365 25105 -335
rect 25055 -385 25105 -365
rect 25055 -415 25065 -385
rect 25095 -415 25105 -385
rect 25055 -425 25105 -415
rect 25140 -335 25190 -325
rect 25140 -365 25150 -335
rect 25180 -365 25190 -335
rect 25140 -385 25190 -365
rect 25140 -415 25150 -385
rect 25180 -415 25190 -385
rect 25140 -425 25190 -415
rect 25225 -335 25275 -325
rect 25225 -365 25235 -335
rect 25265 -365 25275 -335
rect 25225 -385 25275 -365
rect 25225 -415 25235 -385
rect 25265 -415 25275 -385
rect 25225 -425 25275 -415
rect 25310 -335 25360 -325
rect 25310 -365 25320 -335
rect 25350 -365 25360 -335
rect 25310 -385 25360 -365
rect 25310 -415 25320 -385
rect 25350 -415 25360 -385
rect 25310 -425 25360 -415
rect 25395 -335 25445 -325
rect 25395 -365 25405 -335
rect 25435 -365 25445 -335
rect 25395 -385 25445 -365
rect 25395 -415 25405 -385
rect 25435 -415 25445 -385
rect 25395 -425 25445 -415
rect 25480 -335 25530 -325
rect 25480 -365 25490 -335
rect 25520 -365 25530 -335
rect 25480 -385 25530 -365
rect 25480 -415 25490 -385
rect 25520 -415 25530 -385
rect 25480 -425 25530 -415
rect 25565 -335 25615 -325
rect 25565 -365 25575 -335
rect 25605 -365 25615 -335
rect 25565 -385 25615 -365
rect 25565 -415 25575 -385
rect 25605 -415 25615 -385
rect 25565 -425 25615 -415
rect 25650 -335 25700 -325
rect 25650 -365 25660 -335
rect 25690 -365 25700 -335
rect 25650 -385 25700 -365
rect 25650 -415 25660 -385
rect 25690 -415 25700 -385
rect 25650 -425 25700 -415
rect 25735 -335 25785 -325
rect 25735 -365 25745 -335
rect 25775 -365 25785 -335
rect 25735 -385 25785 -365
rect 25735 -415 25745 -385
rect 25775 -415 25785 -385
rect 25735 -425 25785 -415
rect 25820 -335 25870 -325
rect 25820 -365 25830 -335
rect 25860 -365 25870 -335
rect 25820 -385 25870 -365
rect 25820 -415 25830 -385
rect 25860 -415 25870 -385
rect 25820 -425 25870 -415
rect 25905 -335 25955 -325
rect 25905 -365 25915 -335
rect 25945 -365 25955 -335
rect 25905 -385 25955 -365
rect 25905 -415 25915 -385
rect 25945 -415 25955 -385
rect 25905 -425 25955 -415
rect 25990 -335 26040 -325
rect 25990 -365 26000 -335
rect 26030 -365 26040 -335
rect 25990 -385 26040 -365
rect 25990 -415 26000 -385
rect 26030 -415 26040 -385
rect 25990 -425 26040 -415
rect 26075 -335 26125 -325
rect 26075 -365 26085 -335
rect 26115 -365 26125 -335
rect 26075 -385 26125 -365
rect 26075 -415 26085 -385
rect 26115 -415 26125 -385
rect 26075 -425 26125 -415
rect 26160 -335 26210 -325
rect 26160 -365 26170 -335
rect 26200 -365 26210 -335
rect 26160 -385 26210 -365
rect 26160 -415 26170 -385
rect 26200 -415 26210 -385
rect 26160 -425 26210 -415
rect 26245 -335 26295 -325
rect 26245 -365 26255 -335
rect 26285 -365 26295 -335
rect 26245 -385 26295 -365
rect 26245 -415 26255 -385
rect 26285 -415 26295 -385
rect 26245 -425 26295 -415
rect 26330 -335 26380 -325
rect 26330 -365 26340 -335
rect 26370 -365 26380 -335
rect 26330 -385 26380 -365
rect 26330 -415 26340 -385
rect 26370 -415 26380 -385
rect 26330 -425 26380 -415
rect 26415 -335 26465 -325
rect 26415 -365 26425 -335
rect 26455 -365 26465 -335
rect 26415 -385 26465 -365
rect 26415 -415 26425 -385
rect 26455 -415 26465 -385
rect 26415 -425 26465 -415
rect 26500 -335 26550 -325
rect 26500 -365 26510 -335
rect 26540 -365 26550 -335
rect 26500 -385 26550 -365
rect 26500 -415 26510 -385
rect 26540 -415 26550 -385
rect 26500 -425 26550 -415
rect 26585 -335 26635 -325
rect 26585 -365 26595 -335
rect 26625 -365 26635 -335
rect 26585 -385 26635 -365
rect 26585 -415 26595 -385
rect 26625 -415 26635 -385
rect 26585 -425 26635 -415
rect 26670 -335 26720 -325
rect 26670 -365 26680 -335
rect 26710 -365 26720 -335
rect 26670 -385 26720 -365
rect 26670 -415 26680 -385
rect 26710 -415 26720 -385
rect 26670 -425 26720 -415
rect 26755 -335 26805 -325
rect 26755 -365 26765 -335
rect 26795 -365 26805 -335
rect 26755 -385 26805 -365
rect 26755 -415 26765 -385
rect 26795 -415 26805 -385
rect 26755 -425 26805 -415
rect 26840 -335 26890 -325
rect 26840 -365 26850 -335
rect 26880 -365 26890 -335
rect 26840 -385 26890 -365
rect 26840 -415 26850 -385
rect 26880 -415 26890 -385
rect 26840 -425 26890 -415
rect 26925 -335 26975 -325
rect 26925 -365 26935 -335
rect 26965 -365 26975 -335
rect 26925 -385 26975 -365
rect 26925 -415 26935 -385
rect 26965 -415 26975 -385
rect 26925 -425 26975 -415
rect 27010 -335 27060 -325
rect 27010 -365 27020 -335
rect 27050 -365 27060 -335
rect 27010 -385 27060 -365
rect 27010 -415 27020 -385
rect 27050 -415 27060 -385
rect 27010 -425 27060 -415
rect 27095 -335 27145 -325
rect 27095 -365 27105 -335
rect 27135 -365 27145 -335
rect 27095 -385 27145 -365
rect 27095 -415 27105 -385
rect 27135 -415 27145 -385
rect 27095 -425 27145 -415
rect 27180 -335 27230 -325
rect 27180 -365 27190 -335
rect 27220 -365 27230 -335
rect 27180 -385 27230 -365
rect 27180 -415 27190 -385
rect 27220 -415 27230 -385
rect 27180 -425 27230 -415
rect 27265 -335 27315 -325
rect 27265 -365 27275 -335
rect 27305 -365 27315 -335
rect 27265 -385 27315 -365
rect 27265 -415 27275 -385
rect 27305 -415 27315 -385
rect 27265 -425 27315 -415
rect 27350 -335 27400 -325
rect 27350 -365 27360 -335
rect 27390 -365 27400 -335
rect 27350 -385 27400 -365
rect 27350 -415 27360 -385
rect 27390 -415 27400 -385
rect 27350 -425 27400 -415
rect 27435 -335 27485 -325
rect 27435 -365 27445 -335
rect 27475 -365 27485 -335
rect 27435 -385 27485 -365
rect 27435 -415 27445 -385
rect 27475 -415 27485 -385
rect 27435 -425 27485 -415
rect 27520 -335 27570 -325
rect 27520 -365 27530 -335
rect 27560 -365 27570 -335
rect 27520 -385 27570 -365
rect 27520 -415 27530 -385
rect 27560 -415 27570 -385
rect 27520 -425 27570 -415
rect 27605 -335 27655 -325
rect 27605 -365 27615 -335
rect 27645 -365 27655 -335
rect 27605 -385 27655 -365
rect 27605 -415 27615 -385
rect 27645 -415 27655 -385
rect 27605 -425 27655 -415
rect 27690 -335 27740 -325
rect 27690 -365 27700 -335
rect 27730 -365 27740 -335
rect 27690 -385 27740 -365
rect 27690 -415 27700 -385
rect 27730 -415 27740 -385
rect 27690 -425 27740 -415
rect 27775 -335 27825 -325
rect 27775 -365 27785 -335
rect 27815 -365 27825 -335
rect 27775 -385 27825 -365
rect 27775 -415 27785 -385
rect 27815 -415 27825 -385
rect 27775 -425 27825 -415
rect 27860 -335 27910 -325
rect 27860 -365 27870 -335
rect 27900 -365 27910 -335
rect 27860 -385 27910 -365
rect 27860 -415 27870 -385
rect 27900 -415 27910 -385
rect 27860 -425 27910 -415
rect 27945 -335 27995 -325
rect 27945 -365 27955 -335
rect 27985 -365 27995 -335
rect 27945 -385 27995 -365
rect 27945 -415 27955 -385
rect 27985 -415 27995 -385
rect 27945 -425 27995 -415
rect 28030 -335 28080 -325
rect 28030 -365 28040 -335
rect 28070 -365 28080 -335
rect 28030 -385 28080 -365
rect 28030 -415 28040 -385
rect 28070 -415 28080 -385
rect 28030 -425 28080 -415
rect 28115 -335 28165 -325
rect 28115 -365 28125 -335
rect 28155 -365 28165 -335
rect 28115 -385 28165 -365
rect 28115 -415 28125 -385
rect 28155 -415 28165 -385
rect 28115 -425 28165 -415
rect 28200 -335 28250 -325
rect 28200 -365 28210 -335
rect 28240 -365 28250 -335
rect 28200 -385 28250 -365
rect 28200 -415 28210 -385
rect 28240 -415 28250 -385
rect 28200 -425 28250 -415
rect 28285 -335 28335 -325
rect 28285 -365 28295 -335
rect 28325 -365 28335 -335
rect 28285 -385 28335 -365
rect 28285 -415 28295 -385
rect 28325 -415 28335 -385
rect 28285 -425 28335 -415
rect 28370 -335 28420 -325
rect 28370 -365 28380 -335
rect 28410 -365 28420 -335
rect 28370 -385 28420 -365
rect 28370 -415 28380 -385
rect 28410 -415 28420 -385
rect 28370 -425 28420 -415
rect 28455 -335 28505 -325
rect 28455 -365 28465 -335
rect 28495 -365 28505 -335
rect 28455 -385 28505 -365
rect 28455 -415 28465 -385
rect 28495 -415 28505 -385
rect 28455 -425 28505 -415
rect 28540 -335 28590 -325
rect 28540 -365 28550 -335
rect 28580 -365 28590 -335
rect 28540 -385 28590 -365
rect 28540 -415 28550 -385
rect 28580 -415 28590 -385
rect 28540 -425 28590 -415
rect 28625 -335 28675 -325
rect 28625 -365 28635 -335
rect 28665 -365 28675 -335
rect 28625 -385 28675 -365
rect 28625 -415 28635 -385
rect 28665 -415 28675 -385
rect 28625 -425 28675 -415
rect 28710 -335 28760 -325
rect 28710 -365 28720 -335
rect 28750 -365 28760 -335
rect 28710 -385 28760 -365
rect 28710 -415 28720 -385
rect 28750 -415 28760 -385
rect 28710 -425 28760 -415
rect 28795 -335 28845 -325
rect 28795 -365 28805 -335
rect 28835 -365 28845 -335
rect 28795 -385 28845 -365
rect 28795 -415 28805 -385
rect 28835 -415 28845 -385
rect 28795 -425 28845 -415
rect 28880 -335 28930 -325
rect 28880 -365 28890 -335
rect 28920 -365 28930 -335
rect 28880 -385 28930 -365
rect 28880 -415 28890 -385
rect 28920 -415 28930 -385
rect 28880 -425 28930 -415
rect 28965 -335 29015 -325
rect 28965 -365 28975 -335
rect 29005 -365 29015 -335
rect 28965 -385 29015 -365
rect 28965 -415 28975 -385
rect 29005 -415 29015 -385
rect 28965 -425 29015 -415
rect 29050 -335 29100 -325
rect 29050 -365 29060 -335
rect 29090 -365 29100 -335
rect 29050 -385 29100 -365
rect 29050 -415 29060 -385
rect 29090 -415 29100 -385
rect 29050 -425 29100 -415
rect 29135 -335 29185 -325
rect 29135 -365 29145 -335
rect 29175 -365 29185 -335
rect 29135 -385 29185 -365
rect 29135 -415 29145 -385
rect 29175 -415 29185 -385
rect 29135 -425 29185 -415
rect 29220 -335 29270 -325
rect 29220 -365 29230 -335
rect 29260 -365 29270 -335
rect 29220 -385 29270 -365
rect 29220 -415 29230 -385
rect 29260 -415 29270 -385
rect 29220 -425 29270 -415
rect 29305 -335 29355 -325
rect 29305 -365 29315 -335
rect 29345 -365 29355 -335
rect 29305 -385 29355 -365
rect 29305 -415 29315 -385
rect 29345 -415 29355 -385
rect 29305 -425 29355 -415
rect 29390 -335 29440 -325
rect 29390 -365 29400 -335
rect 29430 -365 29440 -335
rect 29390 -385 29440 -365
rect 29390 -415 29400 -385
rect 29430 -415 29440 -385
rect 29390 -425 29440 -415
rect 29475 -335 29525 -325
rect 29475 -365 29485 -335
rect 29515 -365 29525 -335
rect 29475 -385 29525 -365
rect 29475 -415 29485 -385
rect 29515 -415 29525 -385
rect 29475 -425 29525 -415
rect 29560 -335 29610 -325
rect 29560 -365 29570 -335
rect 29600 -365 29610 -335
rect 29560 -385 29610 -365
rect 29560 -415 29570 -385
rect 29600 -415 29610 -385
rect 29560 -425 29610 -415
rect 29645 -335 29695 -325
rect 29645 -365 29655 -335
rect 29685 -365 29695 -335
rect 29645 -385 29695 -365
rect 29645 -415 29655 -385
rect 29685 -415 29695 -385
rect 29645 -425 29695 -415
rect 29730 -335 29780 -325
rect 29730 -365 29740 -335
rect 29770 -365 29780 -335
rect 29730 -385 29780 -365
rect 29730 -415 29740 -385
rect 29770 -415 29780 -385
rect 29730 -425 29780 -415
rect 29815 -335 29865 -325
rect 29815 -365 29825 -335
rect 29855 -365 29865 -335
rect 29815 -385 29865 -365
rect 29815 -415 29825 -385
rect 29855 -415 29865 -385
rect 29815 -425 29865 -415
rect 29900 -335 29950 -325
rect 29900 -365 29910 -335
rect 29940 -365 29950 -335
rect 29900 -385 29950 -365
rect 29900 -415 29910 -385
rect 29940 -415 29950 -385
rect 29900 -425 29950 -415
rect 29985 -335 30035 -325
rect 29985 -365 29995 -335
rect 30025 -365 30035 -335
rect 29985 -385 30035 -365
rect 29985 -415 29995 -385
rect 30025 -415 30035 -385
rect 29985 -425 30035 -415
rect 30070 -335 30120 -325
rect 30070 -365 30080 -335
rect 30110 -365 30120 -335
rect 30070 -385 30120 -365
rect 30070 -415 30080 -385
rect 30110 -415 30120 -385
rect 30070 -425 30120 -415
rect 30155 -335 30205 -325
rect 30155 -365 30165 -335
rect 30195 -365 30205 -335
rect 30155 -385 30205 -365
rect 30155 -415 30165 -385
rect 30195 -415 30205 -385
rect 30155 -425 30205 -415
rect 30240 -335 30290 -325
rect 30240 -365 30250 -335
rect 30280 -365 30290 -335
rect 30240 -385 30290 -365
rect 30240 -415 30250 -385
rect 30280 -415 30290 -385
rect 30240 -425 30290 -415
rect 30325 -335 30375 -325
rect 30325 -365 30335 -335
rect 30365 -365 30375 -335
rect 30325 -385 30375 -365
rect 30325 -415 30335 -385
rect 30365 -415 30375 -385
rect 30325 -425 30375 -415
rect 30410 -335 30460 -325
rect 30410 -365 30420 -335
rect 30450 -365 30460 -335
rect 30410 -385 30460 -365
rect 30410 -415 30420 -385
rect 30450 -415 30460 -385
rect 30410 -425 30460 -415
rect 30495 -335 30545 -325
rect 30495 -365 30505 -335
rect 30535 -365 30545 -335
rect 30495 -385 30545 -365
rect 30495 -415 30505 -385
rect 30535 -415 30545 -385
rect 30495 -425 30545 -415
rect 30580 -335 30630 -325
rect 30580 -365 30590 -335
rect 30620 -365 30630 -335
rect 30580 -385 30630 -365
rect 30580 -415 30590 -385
rect 30620 -415 30630 -385
rect 30580 -425 30630 -415
rect 30665 -335 30715 -325
rect 30665 -365 30675 -335
rect 30705 -365 30715 -335
rect 30665 -385 30715 -365
rect 30665 -415 30675 -385
rect 30705 -415 30715 -385
rect 30665 -425 30715 -415
rect 30750 -335 30800 -325
rect 30750 -365 30760 -335
rect 30790 -365 30800 -335
rect 30750 -385 30800 -365
rect 30750 -415 30760 -385
rect 30790 -415 30800 -385
rect 30750 -425 30800 -415
rect 30835 -335 30885 -325
rect 30835 -365 30845 -335
rect 30875 -365 30885 -335
rect 30835 -385 30885 -365
rect 30835 -415 30845 -385
rect 30875 -415 30885 -385
rect 30835 -425 30885 -415
rect 30920 -335 30970 -325
rect 30920 -365 30930 -335
rect 30960 -365 30970 -335
rect 30920 -385 30970 -365
rect 30920 -415 30930 -385
rect 30960 -415 30970 -385
rect 30920 -425 30970 -415
rect 31005 -335 31055 -325
rect 31005 -365 31015 -335
rect 31045 -365 31055 -335
rect 31005 -385 31055 -365
rect 31005 -415 31015 -385
rect 31045 -415 31055 -385
rect 31005 -425 31055 -415
rect 31090 -335 31140 -325
rect 31090 -365 31100 -335
rect 31130 -365 31140 -335
rect 31090 -385 31140 -365
rect 31090 -415 31100 -385
rect 31130 -415 31140 -385
rect 31090 -425 31140 -415
rect 31175 -335 31225 -325
rect 31175 -365 31185 -335
rect 31215 -365 31225 -335
rect 31175 -385 31225 -365
rect 31175 -415 31185 -385
rect 31215 -415 31225 -385
rect 31175 -425 31225 -415
rect 31260 -335 31310 -325
rect 31260 -365 31270 -335
rect 31300 -365 31310 -335
rect 31260 -385 31310 -365
rect 31260 -415 31270 -385
rect 31300 -415 31310 -385
rect 31260 -425 31310 -415
rect 31345 -335 31395 -325
rect 31345 -365 31355 -335
rect 31385 -365 31395 -335
rect 31345 -385 31395 -365
rect 31345 -415 31355 -385
rect 31385 -415 31395 -385
rect 31345 -425 31395 -415
rect 31430 -335 31480 -325
rect 31430 -365 31440 -335
rect 31470 -365 31480 -335
rect 31430 -385 31480 -365
rect 31430 -415 31440 -385
rect 31470 -415 31480 -385
rect 31430 -425 31480 -415
rect 31515 -335 31565 -325
rect 31515 -365 31525 -335
rect 31555 -365 31565 -335
rect 31515 -385 31565 -365
rect 31515 -415 31525 -385
rect 31555 -415 31565 -385
rect 31515 -425 31565 -415
rect 31600 -335 31650 -325
rect 31600 -365 31610 -335
rect 31640 -365 31650 -335
rect 31600 -385 31650 -365
rect 31600 -415 31610 -385
rect 31640 -415 31650 -385
rect 31600 -425 31650 -415
rect 31685 -335 31735 -325
rect 31685 -365 31695 -335
rect 31725 -365 31735 -335
rect 31685 -385 31735 -365
rect 31685 -415 31695 -385
rect 31725 -415 31735 -385
rect 31685 -425 31735 -415
rect 31770 -335 31820 -325
rect 31770 -365 31780 -335
rect 31810 -365 31820 -335
rect 31770 -385 31820 -365
rect 31770 -415 31780 -385
rect 31810 -415 31820 -385
rect 31770 -425 31820 -415
rect 31855 -335 31905 -325
rect 31855 -365 31865 -335
rect 31895 -365 31905 -335
rect 31855 -385 31905 -365
rect 31855 -415 31865 -385
rect 31895 -415 31905 -385
rect 31855 -425 31905 -415
rect 31940 -335 31990 -325
rect 31940 -365 31950 -335
rect 31980 -365 31990 -335
rect 31940 -385 31990 -365
rect 31940 -415 31950 -385
rect 31980 -415 31990 -385
rect 31940 -425 31990 -415
rect 32025 -335 32075 -325
rect 32025 -365 32035 -335
rect 32065 -365 32075 -335
rect 32025 -385 32075 -365
rect 32025 -415 32035 -385
rect 32065 -415 32075 -385
rect 32025 -425 32075 -415
rect 32110 -335 32160 -325
rect 32110 -365 32120 -335
rect 32150 -365 32160 -335
rect 32110 -385 32160 -365
rect 32110 -415 32120 -385
rect 32150 -415 32160 -385
rect 32110 -425 32160 -415
rect 32195 -335 32245 -325
rect 32195 -365 32205 -335
rect 32235 -365 32245 -335
rect 32195 -385 32245 -365
rect 32195 -415 32205 -385
rect 32235 -415 32245 -385
rect 32195 -425 32245 -415
rect 32280 -335 32330 -325
rect 32280 -365 32290 -335
rect 32320 -365 32330 -335
rect 32280 -385 32330 -365
rect 32280 -415 32290 -385
rect 32320 -415 32330 -385
rect 32280 -425 32330 -415
rect 32365 -335 32415 -325
rect 32365 -365 32375 -335
rect 32405 -365 32415 -335
rect 32365 -385 32415 -365
rect 32365 -415 32375 -385
rect 32405 -415 32415 -385
rect 32365 -425 32415 -415
rect 32450 -335 32500 -325
rect 32450 -365 32460 -335
rect 32490 -365 32500 -335
rect 32450 -385 32500 -365
rect 32450 -415 32460 -385
rect 32490 -415 32500 -385
rect 32450 -425 32500 -415
rect 32535 -335 32585 -325
rect 32535 -365 32545 -335
rect 32575 -365 32585 -335
rect 32535 -385 32585 -365
rect 32535 -415 32545 -385
rect 32575 -415 32585 -385
rect 32535 -425 32585 -415
rect 32620 -335 32670 -325
rect 32620 -365 32630 -335
rect 32660 -365 32670 -335
rect 32620 -385 32670 -365
rect 32620 -415 32630 -385
rect 32660 -415 32670 -385
rect 32620 -425 32670 -415
rect 32705 -335 32755 -325
rect 32705 -365 32715 -335
rect 32745 -365 32755 -335
rect 32705 -385 32755 -365
rect 32705 -415 32715 -385
rect 32745 -415 32755 -385
rect 32705 -425 32755 -415
rect 32790 -335 32840 -325
rect 32790 -365 32800 -335
rect 32830 -365 32840 -335
rect 32790 -385 32840 -365
rect 32790 -415 32800 -385
rect 32830 -415 32840 -385
rect 32790 -425 32840 -415
rect 32875 -335 32925 -325
rect 32875 -365 32885 -335
rect 32915 -365 32925 -335
rect 32875 -385 32925 -365
rect 32875 -415 32885 -385
rect 32915 -415 32925 -385
rect 32875 -425 32925 -415
rect 32960 -335 33010 -325
rect 32960 -365 32970 -335
rect 33000 -365 33010 -335
rect 32960 -385 33010 -365
rect 32960 -415 32970 -385
rect 33000 -415 33010 -385
rect 32960 -425 33010 -415
rect 33045 -335 33095 -325
rect 33045 -365 33055 -335
rect 33085 -365 33095 -335
rect 33045 -385 33095 -365
rect 33045 -415 33055 -385
rect 33085 -415 33095 -385
rect 33045 -425 33095 -415
rect 33130 -335 33180 -325
rect 33130 -365 33140 -335
rect 33170 -365 33180 -335
rect 33130 -385 33180 -365
rect 33130 -415 33140 -385
rect 33170 -415 33180 -385
rect 33130 -425 33180 -415
rect 33215 -335 33265 -325
rect 33215 -365 33225 -335
rect 33255 -365 33265 -335
rect 33215 -385 33265 -365
rect 33215 -415 33225 -385
rect 33255 -415 33265 -385
rect 33215 -425 33265 -415
rect 33300 -335 33350 -325
rect 33300 -365 33310 -335
rect 33340 -365 33350 -335
rect 33300 -385 33350 -365
rect 33300 -415 33310 -385
rect 33340 -415 33350 -385
rect 33300 -425 33350 -415
rect 33385 -335 33435 -325
rect 33385 -365 33395 -335
rect 33425 -365 33435 -335
rect 33385 -385 33435 -365
rect 33385 -415 33395 -385
rect 33425 -415 33435 -385
rect 33385 -425 33435 -415
rect 33470 -335 33520 -325
rect 33470 -365 33480 -335
rect 33510 -365 33520 -335
rect 33470 -385 33520 -365
rect 33470 -415 33480 -385
rect 33510 -415 33520 -385
rect 33470 -425 33520 -415
rect 33555 -335 33605 -325
rect 33555 -365 33565 -335
rect 33595 -365 33605 -335
rect 33555 -385 33605 -365
rect 33555 -415 33565 -385
rect 33595 -415 33605 -385
rect 33555 -425 33605 -415
rect 33640 -335 33690 -325
rect 33640 -365 33650 -335
rect 33680 -365 33690 -335
rect 33640 -385 33690 -365
rect 33640 -415 33650 -385
rect 33680 -415 33690 -385
rect 33640 -425 33690 -415
rect 33725 -335 33775 -325
rect 33725 -365 33735 -335
rect 33765 -365 33775 -335
rect 33725 -385 33775 -365
rect 33725 -415 33735 -385
rect 33765 -415 33775 -385
rect 33725 -425 33775 -415
rect 33810 -335 33860 -325
rect 33810 -365 33820 -335
rect 33850 -365 33860 -335
rect 33810 -385 33860 -365
rect 33810 -415 33820 -385
rect 33850 -415 33860 -385
rect 33810 -425 33860 -415
rect 33895 -335 33945 -325
rect 33895 -365 33905 -335
rect 33935 -365 33945 -335
rect 33895 -385 33945 -365
rect 33895 -415 33905 -385
rect 33935 -415 33945 -385
rect 33895 -425 33945 -415
rect 33980 -335 34030 -325
rect 33980 -365 33990 -335
rect 34020 -365 34030 -335
rect 33980 -385 34030 -365
rect 33980 -415 33990 -385
rect 34020 -415 34030 -385
rect 33980 -425 34030 -415
rect 34065 -335 34115 -325
rect 34065 -365 34075 -335
rect 34105 -365 34115 -335
rect 34065 -385 34115 -365
rect 34065 -415 34075 -385
rect 34105 -415 34115 -385
rect 34065 -425 34115 -415
rect 34150 -335 34200 -325
rect 34150 -365 34160 -335
rect 34190 -365 34200 -335
rect 34150 -385 34200 -365
rect 34150 -415 34160 -385
rect 34190 -415 34200 -385
rect 34150 -425 34200 -415
rect 34235 -335 34285 -325
rect 34235 -365 34245 -335
rect 34275 -365 34285 -335
rect 34235 -385 34285 -365
rect 34235 -415 34245 -385
rect 34275 -415 34285 -385
rect 34235 -425 34285 -415
rect 34320 -335 34370 -325
rect 34320 -365 34330 -335
rect 34360 -365 34370 -335
rect 34320 -385 34370 -365
rect 34320 -415 34330 -385
rect 34360 -415 34370 -385
rect 34320 -425 34370 -415
rect 34405 -335 34455 -325
rect 34405 -365 34415 -335
rect 34445 -365 34455 -335
rect 34405 -385 34455 -365
rect 34405 -415 34415 -385
rect 34445 -415 34455 -385
rect 34405 -425 34455 -415
rect 34490 -335 34540 -325
rect 34490 -365 34500 -335
rect 34530 -365 34540 -335
rect 34490 -385 34540 -365
rect 34490 -415 34500 -385
rect 34530 -415 34540 -385
rect 34490 -425 34540 -415
rect 34575 -335 34625 -325
rect 34575 -365 34585 -335
rect 34615 -365 34625 -335
rect 34575 -385 34625 -365
rect 34575 -415 34585 -385
rect 34615 -415 34625 -385
rect 34575 -425 34625 -415
rect 34660 -335 34710 -325
rect 34660 -365 34670 -335
rect 34700 -365 34710 -335
rect 34660 -385 34710 -365
rect 34660 -415 34670 -385
rect 34700 -415 34710 -385
rect 34660 -425 34710 -415
rect 34745 -335 34795 -325
rect 34745 -365 34755 -335
rect 34785 -365 34795 -335
rect 34745 -385 34795 -365
rect 34745 -415 34755 -385
rect 34785 -415 34795 -385
rect 34745 -425 34795 -415
rect 34830 -335 34880 -325
rect 34830 -365 34840 -335
rect 34870 -365 34880 -335
rect 34830 -385 34880 -365
rect 34830 -415 34840 -385
rect 34870 -415 34880 -385
rect 34830 -425 34880 -415
rect 34915 -335 34965 -325
rect 34915 -365 34925 -335
rect 34955 -365 34965 -335
rect 34915 -385 34965 -365
rect 34915 -415 34925 -385
rect 34955 -415 34965 -385
rect 34915 -425 34965 -415
rect 35000 -335 35050 -325
rect 35000 -365 35010 -335
rect 35040 -365 35050 -335
rect 35000 -385 35050 -365
rect 35000 -415 35010 -385
rect 35040 -415 35050 -385
rect 35000 -425 35050 -415
rect 35085 -335 35135 -325
rect 35085 -365 35095 -335
rect 35125 -365 35135 -335
rect 35085 -385 35135 -365
rect 35085 -415 35095 -385
rect 35125 -415 35135 -385
rect 35085 -425 35135 -415
rect 35170 -335 35220 -325
rect 35170 -365 35180 -335
rect 35210 -365 35220 -335
rect 35170 -385 35220 -365
rect 35170 -415 35180 -385
rect 35210 -415 35220 -385
rect 35170 -425 35220 -415
rect 35255 -335 35305 -325
rect 35255 -365 35265 -335
rect 35295 -365 35305 -335
rect 35255 -385 35305 -365
rect 35255 -415 35265 -385
rect 35295 -415 35305 -385
rect 35255 -425 35305 -415
rect 35340 -335 35390 -325
rect 35340 -365 35350 -335
rect 35380 -365 35390 -335
rect 35340 -385 35390 -365
rect 35340 -415 35350 -385
rect 35380 -415 35390 -385
rect 35340 -425 35390 -415
rect 35425 -335 35475 -325
rect 35425 -365 35435 -335
rect 35465 -365 35475 -335
rect 35425 -385 35475 -365
rect 35425 -415 35435 -385
rect 35465 -415 35475 -385
rect 35425 -425 35475 -415
rect 35510 -335 35560 -325
rect 35510 -365 35520 -335
rect 35550 -365 35560 -335
rect 35510 -385 35560 -365
rect 35510 -415 35520 -385
rect 35550 -415 35560 -385
rect 35510 -425 35560 -415
rect 35595 -335 35645 -325
rect 35595 -365 35605 -335
rect 35635 -365 35645 -335
rect 35595 -385 35645 -365
rect 35595 -415 35605 -385
rect 35635 -415 35645 -385
rect 35595 -425 35645 -415
rect 35680 -335 35730 -325
rect 35680 -365 35690 -335
rect 35720 -365 35730 -335
rect 35680 -385 35730 -365
rect 35680 -415 35690 -385
rect 35720 -415 35730 -385
rect 35680 -425 35730 -415
rect 35765 -335 35815 -325
rect 35765 -365 35775 -335
rect 35805 -365 35815 -335
rect 35765 -385 35815 -365
rect 35765 -415 35775 -385
rect 35805 -415 35815 -385
rect 35765 -425 35815 -415
rect 35850 -335 35900 -325
rect 35850 -365 35860 -335
rect 35890 -365 35900 -335
rect 35850 -385 35900 -365
rect 35850 -415 35860 -385
rect 35890 -415 35900 -385
rect 35850 -425 35900 -415
rect 35935 -335 35985 -325
rect 35935 -365 35945 -335
rect 35975 -365 35985 -335
rect 35935 -385 35985 -365
rect 35935 -415 35945 -385
rect 35975 -415 35985 -385
rect 35935 -425 35985 -415
rect 36020 -335 36070 -325
rect 36020 -365 36030 -335
rect 36060 -365 36070 -335
rect 36020 -385 36070 -365
rect 36020 -415 36030 -385
rect 36060 -415 36070 -385
rect 36020 -425 36070 -415
rect 36105 -335 36155 -325
rect 36105 -365 36115 -335
rect 36145 -365 36155 -335
rect 36105 -385 36155 -365
rect 36105 -415 36115 -385
rect 36145 -415 36155 -385
rect 36105 -425 36155 -415
rect 36190 -335 36240 -325
rect 36190 -365 36200 -335
rect 36230 -365 36240 -335
rect 36190 -385 36240 -365
rect 36190 -415 36200 -385
rect 36230 -415 36240 -385
rect 36190 -425 36240 -415
rect 36275 -335 36325 -325
rect 36275 -365 36285 -335
rect 36315 -365 36325 -335
rect 36275 -385 36325 -365
rect 36275 -415 36285 -385
rect 36315 -415 36325 -385
rect 36275 -425 36325 -415
rect 36360 -335 36410 -325
rect 36360 -365 36370 -335
rect 36400 -365 36410 -335
rect 36360 -385 36410 -365
rect 36360 -415 36370 -385
rect 36400 -415 36410 -385
rect 36360 -425 36410 -415
rect 36445 -335 36495 -325
rect 36445 -365 36455 -335
rect 36485 -365 36495 -335
rect 36445 -385 36495 -365
rect 36445 -415 36455 -385
rect 36485 -415 36495 -385
rect 36445 -425 36495 -415
rect 36530 -335 36580 -325
rect 36530 -365 36540 -335
rect 36570 -365 36580 -335
rect 36530 -385 36580 -365
rect 36530 -415 36540 -385
rect 36570 -415 36580 -385
rect 36530 -425 36580 -415
rect 36615 -335 36665 -325
rect 36615 -365 36625 -335
rect 36655 -365 36665 -335
rect 36615 -385 36665 -365
rect 36615 -415 36625 -385
rect 36655 -415 36665 -385
rect 36615 -425 36665 -415
rect 36700 -335 36750 -325
rect 36700 -365 36710 -335
rect 36740 -365 36750 -335
rect 36700 -385 36750 -365
rect 36700 -415 36710 -385
rect 36740 -415 36750 -385
rect 36700 -425 36750 -415
rect 36785 -335 36835 -325
rect 36785 -365 36795 -335
rect 36825 -365 36835 -335
rect 36785 -385 36835 -365
rect 36785 -415 36795 -385
rect 36825 -415 36835 -385
rect 36785 -425 36835 -415
rect 36870 -335 36920 -325
rect 36870 -365 36880 -335
rect 36910 -365 36920 -335
rect 36870 -385 36920 -365
rect 36870 -415 36880 -385
rect 36910 -415 36920 -385
rect 36870 -425 36920 -415
rect 36955 -335 37005 -325
rect 36955 -365 36965 -335
rect 36995 -365 37005 -335
rect 36955 -385 37005 -365
rect 36955 -415 36965 -385
rect 36995 -415 37005 -385
rect 36955 -425 37005 -415
rect 37040 -335 37090 -325
rect 37040 -365 37050 -335
rect 37080 -365 37090 -335
rect 37040 -385 37090 -365
rect 37040 -415 37050 -385
rect 37080 -415 37090 -385
rect 37040 -425 37090 -415
rect 37125 -335 37175 -325
rect 37125 -365 37135 -335
rect 37165 -365 37175 -335
rect 37125 -385 37175 -365
rect 37125 -415 37135 -385
rect 37165 -415 37175 -385
rect 37125 -425 37175 -415
rect 37210 -335 37260 -325
rect 37210 -365 37220 -335
rect 37250 -365 37260 -335
rect 37210 -385 37260 -365
rect 37210 -415 37220 -385
rect 37250 -415 37260 -385
rect 37210 -425 37260 -415
rect 37295 -335 37345 -325
rect 37295 -365 37305 -335
rect 37335 -365 37345 -335
rect 37295 -385 37345 -365
rect 37295 -415 37305 -385
rect 37335 -415 37345 -385
rect 37295 -425 37345 -415
rect 37380 -335 37430 -325
rect 37380 -365 37390 -335
rect 37420 -365 37430 -335
rect 37380 -385 37430 -365
rect 37380 -415 37390 -385
rect 37420 -415 37430 -385
rect 37380 -425 37430 -415
rect 37465 -335 37515 -325
rect 37465 -365 37475 -335
rect 37505 -365 37515 -335
rect 37465 -385 37515 -365
rect 37465 -415 37475 -385
rect 37505 -415 37515 -385
rect 37465 -425 37515 -415
rect 37550 -335 37600 -325
rect 37550 -365 37560 -335
rect 37590 -365 37600 -335
rect 37550 -385 37600 -365
rect 37550 -415 37560 -385
rect 37590 -415 37600 -385
rect 37550 -425 37600 -415
rect 37635 -335 37685 -325
rect 37635 -365 37645 -335
rect 37675 -365 37685 -335
rect 37635 -385 37685 -365
rect 37635 -415 37645 -385
rect 37675 -415 37685 -385
rect 37635 -425 37685 -415
rect 37720 -335 37770 -325
rect 37720 -365 37730 -335
rect 37760 -365 37770 -335
rect 37720 -385 37770 -365
rect 37720 -415 37730 -385
rect 37760 -415 37770 -385
rect 37720 -425 37770 -415
rect 37805 -335 37855 -325
rect 37805 -365 37815 -335
rect 37845 -365 37855 -335
rect 37805 -385 37855 -365
rect 37805 -415 37815 -385
rect 37845 -415 37855 -385
rect 37805 -425 37855 -415
rect 37890 -335 37940 -325
rect 37890 -365 37900 -335
rect 37930 -365 37940 -335
rect 37890 -385 37940 -365
rect 37890 -415 37900 -385
rect 37930 -415 37940 -385
rect 37890 -425 37940 -415
rect 37975 -335 38025 -325
rect 37975 -365 37985 -335
rect 38015 -365 38025 -335
rect 37975 -385 38025 -365
rect 37975 -415 37985 -385
rect 38015 -415 38025 -385
rect 37975 -425 38025 -415
rect 38060 -335 38110 -325
rect 38060 -365 38070 -335
rect 38100 -365 38110 -335
rect 38060 -385 38110 -365
rect 38060 -415 38070 -385
rect 38100 -415 38110 -385
rect 38060 -425 38110 -415
rect 38145 -335 38195 -325
rect 38145 -365 38155 -335
rect 38185 -365 38195 -335
rect 38145 -385 38195 -365
rect 38145 -415 38155 -385
rect 38185 -415 38195 -385
rect 38145 -425 38195 -415
rect 38230 -335 38280 -325
rect 38230 -365 38240 -335
rect 38270 -365 38280 -335
rect 38230 -385 38280 -365
rect 38230 -415 38240 -385
rect 38270 -415 38280 -385
rect 38230 -425 38280 -415
rect 38315 -335 38365 -325
rect 38315 -365 38325 -335
rect 38355 -365 38365 -335
rect 38315 -385 38365 -365
rect 38315 -415 38325 -385
rect 38355 -415 38365 -385
rect 38315 -425 38365 -415
rect 38400 -335 38450 -325
rect 38400 -365 38410 -335
rect 38440 -365 38450 -335
rect 38400 -385 38450 -365
rect 38400 -415 38410 -385
rect 38440 -415 38450 -385
rect 38400 -425 38450 -415
rect 38485 -335 38535 -325
rect 38485 -365 38495 -335
rect 38525 -365 38535 -335
rect 38485 -385 38535 -365
rect 38485 -415 38495 -385
rect 38525 -415 38535 -385
rect 38485 -425 38535 -415
rect 38570 -335 38620 -325
rect 38570 -365 38580 -335
rect 38610 -365 38620 -335
rect 38570 -385 38620 -365
rect 38570 -415 38580 -385
rect 38610 -415 38620 -385
rect 38570 -425 38620 -415
rect 38655 -335 38705 -325
rect 38655 -365 38665 -335
rect 38695 -365 38705 -335
rect 38655 -385 38705 -365
rect 38655 -415 38665 -385
rect 38695 -415 38705 -385
rect 38655 -425 38705 -415
rect 38740 -335 38790 -325
rect 38740 -365 38750 -335
rect 38780 -365 38790 -335
rect 38740 -385 38790 -365
rect 38740 -415 38750 -385
rect 38780 -415 38790 -385
rect 38740 -425 38790 -415
rect 38825 -335 38875 -325
rect 38825 -365 38835 -335
rect 38865 -365 38875 -335
rect 38825 -385 38875 -365
rect 38825 -415 38835 -385
rect 38865 -415 38875 -385
rect 38825 -425 38875 -415
rect 38910 -335 38960 -325
rect 38910 -365 38920 -335
rect 38950 -365 38960 -335
rect 38910 -385 38960 -365
rect 38910 -415 38920 -385
rect 38950 -415 38960 -385
rect 38910 -425 38960 -415
rect 38995 -335 39045 -325
rect 38995 -365 39005 -335
rect 39035 -365 39045 -335
rect 38995 -385 39045 -365
rect 38995 -415 39005 -385
rect 39035 -415 39045 -385
rect 38995 -425 39045 -415
rect 39080 -335 39130 -325
rect 39080 -365 39090 -335
rect 39120 -365 39130 -335
rect 39080 -385 39130 -365
rect 39080 -415 39090 -385
rect 39120 -415 39130 -385
rect 39080 -425 39130 -415
rect 39165 -335 39215 -325
rect 39165 -365 39175 -335
rect 39205 -365 39215 -335
rect 39165 -385 39215 -365
rect 39165 -415 39175 -385
rect 39205 -415 39215 -385
rect 39165 -425 39215 -415
rect 39250 -335 39300 -325
rect 39250 -365 39260 -335
rect 39290 -365 39300 -335
rect 39250 -385 39300 -365
rect 39250 -415 39260 -385
rect 39290 -415 39300 -385
rect 39250 -425 39300 -415
rect 39335 -335 39385 -325
rect 39335 -365 39345 -335
rect 39375 -365 39385 -335
rect 39335 -385 39385 -365
rect 39335 -415 39345 -385
rect 39375 -415 39385 -385
rect 39335 -425 39385 -415
rect 39420 -335 39470 -325
rect 39420 -365 39430 -335
rect 39460 -365 39470 -335
rect 39420 -385 39470 -365
rect 39420 -415 39430 -385
rect 39460 -415 39470 -385
rect 39420 -425 39470 -415
rect 39505 -335 39555 -325
rect 39505 -365 39515 -335
rect 39545 -365 39555 -335
rect 39505 -385 39555 -365
rect 39505 -415 39515 -385
rect 39545 -415 39555 -385
rect 39505 -425 39555 -415
rect 39590 -335 39640 -325
rect 39590 -365 39600 -335
rect 39630 -365 39640 -335
rect 39590 -385 39640 -365
rect 39590 -415 39600 -385
rect 39630 -415 39640 -385
rect 39590 -425 39640 -415
rect 39675 -335 39725 -325
rect 39675 -365 39685 -335
rect 39715 -365 39725 -335
rect 39675 -385 39725 -365
rect 39675 -415 39685 -385
rect 39715 -415 39725 -385
rect 39675 -425 39725 -415
rect 39760 -335 39810 -325
rect 39760 -365 39770 -335
rect 39800 -365 39810 -335
rect 39760 -385 39810 -365
rect 39760 -415 39770 -385
rect 39800 -415 39810 -385
rect 39760 -425 39810 -415
rect 39845 -335 39895 -325
rect 39845 -365 39855 -335
rect 39885 -365 39895 -335
rect 39845 -385 39895 -365
rect 39845 -415 39855 -385
rect 39885 -415 39895 -385
rect 39845 -425 39895 -415
rect 39930 -335 39980 -325
rect 39930 -365 39940 -335
rect 39970 -365 39980 -335
rect 39930 -385 39980 -365
rect 39930 -415 39940 -385
rect 39970 -415 39980 -385
rect 39930 -425 39980 -415
rect 40015 -335 40065 -325
rect 40015 -365 40025 -335
rect 40055 -365 40065 -335
rect 40015 -385 40065 -365
rect 40015 -415 40025 -385
rect 40055 -415 40065 -385
rect 40015 -425 40065 -415
rect 40100 -335 40150 -325
rect 40100 -365 40110 -335
rect 40140 -365 40150 -335
rect 40100 -385 40150 -365
rect 40100 -415 40110 -385
rect 40140 -415 40150 -385
rect 40100 -425 40150 -415
rect 40185 -335 40235 -325
rect 40185 -365 40195 -335
rect 40225 -365 40235 -335
rect 40185 -385 40235 -365
rect 40185 -415 40195 -385
rect 40225 -415 40235 -385
rect 40185 -425 40235 -415
rect 40270 -335 40320 -325
rect 40270 -365 40280 -335
rect 40310 -365 40320 -335
rect 40270 -385 40320 -365
rect 40270 -415 40280 -385
rect 40310 -415 40320 -385
rect 40270 -425 40320 -415
rect 40355 -335 40405 -325
rect 40355 -365 40365 -335
rect 40395 -365 40405 -335
rect 40355 -385 40405 -365
rect 40355 -415 40365 -385
rect 40395 -415 40405 -385
rect 40355 -425 40405 -415
rect 40440 -335 40490 -325
rect 40440 -365 40450 -335
rect 40480 -365 40490 -335
rect 40440 -385 40490 -365
rect 40440 -415 40450 -385
rect 40480 -415 40490 -385
rect 40440 -425 40490 -415
rect 40525 -335 40575 -325
rect 40525 -365 40535 -335
rect 40565 -365 40575 -335
rect 40525 -385 40575 -365
rect 40525 -415 40535 -385
rect 40565 -415 40575 -385
rect 40525 -425 40575 -415
rect 40610 -335 40660 -325
rect 40610 -365 40620 -335
rect 40650 -365 40660 -335
rect 40610 -385 40660 -365
rect 40610 -415 40620 -385
rect 40650 -415 40660 -385
rect 40610 -425 40660 -415
rect 40695 -335 40745 -325
rect 40695 -365 40705 -335
rect 40735 -365 40745 -335
rect 40695 -385 40745 -365
rect 40695 -415 40705 -385
rect 40735 -415 40745 -385
rect 40695 -425 40745 -415
rect 40780 -335 40830 -325
rect 40780 -365 40790 -335
rect 40820 -365 40830 -335
rect 40780 -385 40830 -365
rect 40780 -415 40790 -385
rect 40820 -415 40830 -385
rect 40780 -425 40830 -415
rect 40865 -335 40915 -325
rect 40865 -365 40875 -335
rect 40905 -365 40915 -335
rect 40865 -385 40915 -365
rect 40865 -415 40875 -385
rect 40905 -415 40915 -385
rect 40865 -425 40915 -415
rect 40950 -335 41000 -325
rect 40950 -365 40960 -335
rect 40990 -365 41000 -335
rect 40950 -385 41000 -365
rect 40950 -415 40960 -385
rect 40990 -415 41000 -385
rect 40950 -425 41000 -415
rect 41035 -335 41085 -325
rect 41035 -365 41045 -335
rect 41075 -365 41085 -335
rect 41035 -385 41085 -365
rect 41035 -415 41045 -385
rect 41075 -415 41085 -385
rect 41035 -425 41085 -415
rect 41120 -335 41170 -325
rect 41120 -365 41130 -335
rect 41160 -365 41170 -335
rect 41120 -385 41170 -365
rect 41120 -415 41130 -385
rect 41160 -415 41170 -385
rect 41120 -425 41170 -415
rect 41205 -335 41255 -325
rect 41205 -365 41215 -335
rect 41245 -365 41255 -335
rect 41205 -385 41255 -365
rect 41205 -415 41215 -385
rect 41245 -415 41255 -385
rect 41205 -425 41255 -415
rect 41290 -335 41340 -325
rect 41290 -365 41300 -335
rect 41330 -365 41340 -335
rect 41290 -385 41340 -365
rect 41290 -415 41300 -385
rect 41330 -415 41340 -385
rect 41290 -425 41340 -415
rect 41375 -335 41425 -325
rect 41375 -365 41385 -335
rect 41415 -365 41425 -335
rect 41375 -385 41425 -365
rect 41375 -415 41385 -385
rect 41415 -415 41425 -385
rect 41375 -425 41425 -415
rect 41460 -335 41510 -325
rect 41460 -365 41470 -335
rect 41500 -365 41510 -335
rect 41460 -385 41510 -365
rect 41460 -415 41470 -385
rect 41500 -415 41510 -385
rect 41460 -425 41510 -415
rect 41545 -335 41595 -325
rect 41545 -365 41555 -335
rect 41585 -365 41595 -335
rect 41545 -385 41595 -365
rect 41545 -415 41555 -385
rect 41585 -415 41595 -385
rect 41545 -425 41595 -415
rect 41630 -335 41680 -325
rect 41630 -365 41640 -335
rect 41670 -365 41680 -335
rect 41630 -385 41680 -365
rect 41630 -415 41640 -385
rect 41670 -415 41680 -385
rect 41630 -425 41680 -415
rect 41715 -335 41765 -325
rect 41715 -365 41725 -335
rect 41755 -365 41765 -335
rect 41715 -385 41765 -365
rect 41715 -415 41725 -385
rect 41755 -415 41765 -385
rect 41715 -425 41765 -415
rect 41800 -335 41850 -325
rect 41800 -365 41810 -335
rect 41840 -365 41850 -335
rect 41800 -385 41850 -365
rect 41800 -415 41810 -385
rect 41840 -415 41850 -385
rect 41800 -425 41850 -415
rect 41885 -335 41935 -325
rect 41885 -365 41895 -335
rect 41925 -365 41935 -335
rect 41885 -385 41935 -365
rect 41885 -415 41895 -385
rect 41925 -415 41935 -385
rect 41885 -425 41935 -415
rect 41970 -335 42020 -325
rect 41970 -365 41980 -335
rect 42010 -365 42020 -335
rect 41970 -385 42020 -365
rect 41970 -415 41980 -385
rect 42010 -415 42020 -385
rect 41970 -425 42020 -415
rect 42055 -335 42105 -325
rect 42055 -365 42065 -335
rect 42095 -365 42105 -335
rect 42055 -385 42105 -365
rect 42055 -415 42065 -385
rect 42095 -415 42105 -385
rect 42055 -425 42105 -415
rect 42140 -335 42190 -325
rect 42140 -365 42150 -335
rect 42180 -365 42190 -335
rect 42140 -385 42190 -365
rect 42140 -415 42150 -385
rect 42180 -415 42190 -385
rect 42140 -425 42190 -415
rect 42225 -335 42275 -325
rect 42225 -365 42235 -335
rect 42265 -365 42275 -335
rect 42225 -385 42275 -365
rect 42225 -415 42235 -385
rect 42265 -415 42275 -385
rect 42225 -425 42275 -415
rect 42310 -335 42360 -325
rect 42310 -365 42320 -335
rect 42350 -365 42360 -335
rect 42310 -385 42360 -365
rect 42310 -415 42320 -385
rect 42350 -415 42360 -385
rect 42310 -425 42360 -415
rect 42395 -335 42445 -325
rect 42395 -365 42405 -335
rect 42435 -365 42445 -335
rect 42395 -385 42445 -365
rect 42395 -415 42405 -385
rect 42435 -415 42445 -385
rect 42395 -425 42445 -415
rect 42480 -335 42530 -325
rect 42480 -365 42490 -335
rect 42520 -365 42530 -335
rect 42480 -385 42530 -365
rect 42480 -415 42490 -385
rect 42520 -415 42530 -385
rect 42480 -425 42530 -415
rect 42565 -335 42615 -325
rect 42565 -365 42575 -335
rect 42605 -365 42615 -335
rect 42565 -385 42615 -365
rect 42565 -415 42575 -385
rect 42605 -415 42615 -385
rect 42565 -425 42615 -415
rect 42650 -335 42700 -325
rect 42650 -365 42660 -335
rect 42690 -365 42700 -335
rect 42650 -385 42700 -365
rect 42650 -415 42660 -385
rect 42690 -415 42700 -385
rect 42650 -425 42700 -415
rect 42735 -335 42785 -325
rect 42735 -365 42745 -335
rect 42775 -365 42785 -335
rect 42735 -385 42785 -365
rect 42735 -415 42745 -385
rect 42775 -415 42785 -385
rect 42735 -425 42785 -415
rect 42820 -335 42870 -325
rect 42820 -365 42830 -335
rect 42860 -365 42870 -335
rect 42820 -385 42870 -365
rect 42820 -415 42830 -385
rect 42860 -415 42870 -385
rect 42820 -425 42870 -415
rect 42905 -335 42955 -325
rect 42905 -365 42915 -335
rect 42945 -365 42955 -335
rect 42905 -385 42955 -365
rect 42905 -415 42915 -385
rect 42945 -415 42955 -385
rect 42905 -425 42955 -415
rect 42990 -335 43040 -325
rect 42990 -365 43000 -335
rect 43030 -365 43040 -335
rect 42990 -385 43040 -365
rect 42990 -415 43000 -385
rect 43030 -415 43040 -385
rect 42990 -425 43040 -415
rect 43075 -335 43125 -325
rect 43075 -365 43085 -335
rect 43115 -365 43125 -335
rect 43075 -385 43125 -365
rect 43075 -415 43085 -385
rect 43115 -415 43125 -385
rect 43075 -425 43125 -415
rect 43160 -335 43210 -325
rect 43160 -365 43170 -335
rect 43200 -365 43210 -335
rect 43160 -385 43210 -365
rect 43160 -415 43170 -385
rect 43200 -415 43210 -385
rect 43160 -425 43210 -415
rect 43245 -335 43295 -325
rect 43245 -365 43255 -335
rect 43285 -365 43295 -335
rect 43245 -385 43295 -365
rect 43245 -415 43255 -385
rect 43285 -415 43295 -385
rect 43245 -425 43295 -415
rect 43330 -335 43380 -325
rect 43330 -365 43340 -335
rect 43370 -365 43380 -335
rect 43330 -385 43380 -365
rect 43330 -415 43340 -385
rect 43370 -415 43380 -385
rect 43330 -425 43380 -415
rect 43415 -335 43465 -325
rect 43415 -365 43425 -335
rect 43455 -365 43465 -335
rect 43415 -385 43465 -365
rect 43415 -415 43425 -385
rect 43455 -415 43465 -385
rect 43415 -425 43465 -415
rect 43500 -335 43550 -325
rect 43500 -365 43510 -335
rect 43540 -365 43550 -335
rect 43500 -385 43550 -365
rect 43500 -415 43510 -385
rect 43540 -415 43550 -385
rect 43500 -425 43550 -415
rect 43585 -335 43635 -325
rect 43585 -365 43595 -335
rect 43625 -365 43635 -335
rect 43585 -385 43635 -365
rect 43585 -415 43595 -385
rect 43625 -415 43635 -385
rect 43585 -425 43635 -415
rect 65 -500 115 -490
rect 65 -530 75 -500
rect 105 -530 115 -500
rect 65 -550 115 -530
rect 65 -580 75 -550
rect 105 -580 115 -550
rect 65 -600 115 -580
rect 65 -630 75 -600
rect 105 -630 115 -600
rect 65 -650 115 -630
rect 65 -680 75 -650
rect 105 -680 115 -650
rect 65 -690 115 -680
rect 150 -500 200 -490
rect 150 -530 160 -500
rect 190 -530 200 -500
rect 150 -550 200 -530
rect 150 -580 160 -550
rect 190 -580 200 -550
rect 150 -600 200 -580
rect 150 -630 160 -600
rect 190 -630 200 -600
rect 150 -650 200 -630
rect 150 -680 160 -650
rect 190 -680 200 -650
rect 150 -690 200 -680
rect 235 -500 285 -490
rect 235 -530 245 -500
rect 275 -530 285 -500
rect 235 -550 285 -530
rect 235 -580 245 -550
rect 275 -580 285 -550
rect 235 -600 285 -580
rect 235 -630 245 -600
rect 275 -630 285 -600
rect 235 -650 285 -630
rect 235 -680 245 -650
rect 275 -680 285 -650
rect 235 -690 285 -680
rect 320 -500 370 -490
rect 320 -530 330 -500
rect 360 -530 370 -500
rect 320 -550 370 -530
rect 320 -580 330 -550
rect 360 -580 370 -550
rect 320 -600 370 -580
rect 320 -630 330 -600
rect 360 -630 370 -600
rect 320 -650 370 -630
rect 320 -680 330 -650
rect 360 -680 370 -650
rect 320 -690 370 -680
rect 405 -500 455 -490
rect 405 -530 415 -500
rect 445 -530 455 -500
rect 405 -550 455 -530
rect 405 -580 415 -550
rect 445 -580 455 -550
rect 405 -600 455 -580
rect 405 -630 415 -600
rect 445 -630 455 -600
rect 405 -650 455 -630
rect 405 -680 415 -650
rect 445 -680 455 -650
rect 405 -690 455 -680
rect 490 -500 540 -490
rect 490 -530 500 -500
rect 530 -530 540 -500
rect 490 -550 540 -530
rect 490 -580 500 -550
rect 530 -580 540 -550
rect 490 -600 540 -580
rect 490 -630 500 -600
rect 530 -630 540 -600
rect 490 -650 540 -630
rect 490 -680 500 -650
rect 530 -680 540 -650
rect 490 -690 540 -680
rect 575 -500 625 -490
rect 575 -530 585 -500
rect 615 -530 625 -500
rect 575 -550 625 -530
rect 575 -580 585 -550
rect 615 -580 625 -550
rect 575 -600 625 -580
rect 575 -630 585 -600
rect 615 -630 625 -600
rect 575 -650 625 -630
rect 575 -680 585 -650
rect 615 -680 625 -650
rect 575 -690 625 -680
rect 660 -500 710 -490
rect 660 -530 670 -500
rect 700 -530 710 -500
rect 660 -550 710 -530
rect 660 -580 670 -550
rect 700 -580 710 -550
rect 660 -600 710 -580
rect 660 -630 670 -600
rect 700 -630 710 -600
rect 660 -650 710 -630
rect 660 -680 670 -650
rect 700 -680 710 -650
rect 660 -690 710 -680
rect 745 -500 795 -490
rect 745 -530 755 -500
rect 785 -530 795 -500
rect 745 -550 795 -530
rect 745 -580 755 -550
rect 785 -580 795 -550
rect 745 -600 795 -580
rect 745 -630 755 -600
rect 785 -630 795 -600
rect 745 -650 795 -630
rect 745 -680 755 -650
rect 785 -680 795 -650
rect 745 -690 795 -680
rect 830 -500 880 -490
rect 830 -530 840 -500
rect 870 -530 880 -500
rect 830 -550 880 -530
rect 830 -580 840 -550
rect 870 -580 880 -550
rect 830 -600 880 -580
rect 830 -630 840 -600
rect 870 -630 880 -600
rect 830 -650 880 -630
rect 830 -680 840 -650
rect 870 -680 880 -650
rect 830 -690 880 -680
rect 915 -500 965 -490
rect 915 -530 925 -500
rect 955 -530 965 -500
rect 915 -550 965 -530
rect 915 -580 925 -550
rect 955 -580 965 -550
rect 915 -600 965 -580
rect 915 -630 925 -600
rect 955 -630 965 -600
rect 915 -650 965 -630
rect 915 -680 925 -650
rect 955 -680 965 -650
rect 915 -690 965 -680
rect 1000 -500 1050 -490
rect 1000 -530 1010 -500
rect 1040 -530 1050 -500
rect 1000 -550 1050 -530
rect 1000 -580 1010 -550
rect 1040 -580 1050 -550
rect 1000 -600 1050 -580
rect 1000 -630 1010 -600
rect 1040 -630 1050 -600
rect 1000 -650 1050 -630
rect 1000 -680 1010 -650
rect 1040 -680 1050 -650
rect 1000 -690 1050 -680
rect 1085 -500 1135 -490
rect 1085 -530 1095 -500
rect 1125 -530 1135 -500
rect 1085 -550 1135 -530
rect 1085 -580 1095 -550
rect 1125 -580 1135 -550
rect 1085 -600 1135 -580
rect 1085 -630 1095 -600
rect 1125 -630 1135 -600
rect 1085 -650 1135 -630
rect 1085 -680 1095 -650
rect 1125 -680 1135 -650
rect 1085 -690 1135 -680
rect 1170 -500 1220 -490
rect 1170 -530 1180 -500
rect 1210 -530 1220 -500
rect 1170 -550 1220 -530
rect 1170 -580 1180 -550
rect 1210 -580 1220 -550
rect 1170 -600 1220 -580
rect 1170 -630 1180 -600
rect 1210 -630 1220 -600
rect 1170 -650 1220 -630
rect 1170 -680 1180 -650
rect 1210 -680 1220 -650
rect 1170 -690 1220 -680
rect 1255 -500 1305 -490
rect 1255 -530 1265 -500
rect 1295 -530 1305 -500
rect 1255 -550 1305 -530
rect 1255 -580 1265 -550
rect 1295 -580 1305 -550
rect 1255 -600 1305 -580
rect 1255 -630 1265 -600
rect 1295 -630 1305 -600
rect 1255 -650 1305 -630
rect 1255 -680 1265 -650
rect 1295 -680 1305 -650
rect 1255 -690 1305 -680
rect 1340 -500 1390 -490
rect 1340 -530 1350 -500
rect 1380 -530 1390 -500
rect 1340 -550 1390 -530
rect 1340 -580 1350 -550
rect 1380 -580 1390 -550
rect 1340 -600 1390 -580
rect 1340 -630 1350 -600
rect 1380 -630 1390 -600
rect 1340 -650 1390 -630
rect 1340 -680 1350 -650
rect 1380 -680 1390 -650
rect 1340 -690 1390 -680
rect 1425 -500 1475 -490
rect 1425 -530 1435 -500
rect 1465 -530 1475 -500
rect 1425 -550 1475 -530
rect 1425 -580 1435 -550
rect 1465 -580 1475 -550
rect 1425 -600 1475 -580
rect 1425 -630 1435 -600
rect 1465 -630 1475 -600
rect 1425 -650 1475 -630
rect 1425 -680 1435 -650
rect 1465 -680 1475 -650
rect 1425 -690 1475 -680
rect 1510 -500 1560 -490
rect 1510 -530 1520 -500
rect 1550 -530 1560 -500
rect 1510 -550 1560 -530
rect 1510 -580 1520 -550
rect 1550 -580 1560 -550
rect 1510 -600 1560 -580
rect 1510 -630 1520 -600
rect 1550 -630 1560 -600
rect 1510 -650 1560 -630
rect 1510 -680 1520 -650
rect 1550 -680 1560 -650
rect 1510 -690 1560 -680
rect 1595 -500 1645 -490
rect 1595 -530 1605 -500
rect 1635 -530 1645 -500
rect 1595 -550 1645 -530
rect 1595 -580 1605 -550
rect 1635 -580 1645 -550
rect 1595 -600 1645 -580
rect 1595 -630 1605 -600
rect 1635 -630 1645 -600
rect 1595 -650 1645 -630
rect 1595 -680 1605 -650
rect 1635 -680 1645 -650
rect 1595 -690 1645 -680
rect 1680 -500 1730 -490
rect 1680 -530 1690 -500
rect 1720 -530 1730 -500
rect 1680 -550 1730 -530
rect 1680 -580 1690 -550
rect 1720 -580 1730 -550
rect 1680 -600 1730 -580
rect 1680 -630 1690 -600
rect 1720 -630 1730 -600
rect 1680 -650 1730 -630
rect 1680 -680 1690 -650
rect 1720 -680 1730 -650
rect 1680 -690 1730 -680
rect 1765 -500 1815 -490
rect 1765 -530 1775 -500
rect 1805 -530 1815 -500
rect 1765 -550 1815 -530
rect 1765 -580 1775 -550
rect 1805 -580 1815 -550
rect 1765 -600 1815 -580
rect 1765 -630 1775 -600
rect 1805 -630 1815 -600
rect 1765 -650 1815 -630
rect 1765 -680 1775 -650
rect 1805 -680 1815 -650
rect 1765 -690 1815 -680
rect 1850 -500 1900 -490
rect 1850 -530 1860 -500
rect 1890 -530 1900 -500
rect 1850 -550 1900 -530
rect 1850 -580 1860 -550
rect 1890 -580 1900 -550
rect 1850 -600 1900 -580
rect 1850 -630 1860 -600
rect 1890 -630 1900 -600
rect 1850 -650 1900 -630
rect 1850 -680 1860 -650
rect 1890 -680 1900 -650
rect 1850 -690 1900 -680
rect 1935 -500 1985 -490
rect 1935 -530 1945 -500
rect 1975 -530 1985 -500
rect 1935 -550 1985 -530
rect 1935 -580 1945 -550
rect 1975 -580 1985 -550
rect 1935 -600 1985 -580
rect 1935 -630 1945 -600
rect 1975 -630 1985 -600
rect 1935 -650 1985 -630
rect 1935 -680 1945 -650
rect 1975 -680 1985 -650
rect 1935 -690 1985 -680
rect 2020 -500 2070 -490
rect 2020 -530 2030 -500
rect 2060 -530 2070 -500
rect 2020 -550 2070 -530
rect 2020 -580 2030 -550
rect 2060 -580 2070 -550
rect 2020 -600 2070 -580
rect 2020 -630 2030 -600
rect 2060 -630 2070 -600
rect 2020 -650 2070 -630
rect 2020 -680 2030 -650
rect 2060 -680 2070 -650
rect 2020 -690 2070 -680
rect 2105 -500 2155 -490
rect 2105 -530 2115 -500
rect 2145 -530 2155 -500
rect 2105 -550 2155 -530
rect 2105 -580 2115 -550
rect 2145 -580 2155 -550
rect 2105 -600 2155 -580
rect 2105 -630 2115 -600
rect 2145 -630 2155 -600
rect 2105 -650 2155 -630
rect 2105 -680 2115 -650
rect 2145 -680 2155 -650
rect 2105 -690 2155 -680
rect 2190 -500 2240 -490
rect 2190 -530 2200 -500
rect 2230 -530 2240 -500
rect 2190 -550 2240 -530
rect 2190 -580 2200 -550
rect 2230 -580 2240 -550
rect 2190 -600 2240 -580
rect 2190 -630 2200 -600
rect 2230 -630 2240 -600
rect 2190 -650 2240 -630
rect 2190 -680 2200 -650
rect 2230 -680 2240 -650
rect 2190 -690 2240 -680
rect 2275 -500 2325 -490
rect 2275 -530 2285 -500
rect 2315 -530 2325 -500
rect 2275 -550 2325 -530
rect 2275 -580 2285 -550
rect 2315 -580 2325 -550
rect 2275 -600 2325 -580
rect 2275 -630 2285 -600
rect 2315 -630 2325 -600
rect 2275 -650 2325 -630
rect 2275 -680 2285 -650
rect 2315 -680 2325 -650
rect 2275 -690 2325 -680
rect 2360 -500 2410 -490
rect 2360 -530 2370 -500
rect 2400 -530 2410 -500
rect 2360 -550 2410 -530
rect 2360 -580 2370 -550
rect 2400 -580 2410 -550
rect 2360 -600 2410 -580
rect 2360 -630 2370 -600
rect 2400 -630 2410 -600
rect 2360 -650 2410 -630
rect 2360 -680 2370 -650
rect 2400 -680 2410 -650
rect 2360 -690 2410 -680
rect 2445 -500 2495 -490
rect 2445 -530 2455 -500
rect 2485 -530 2495 -500
rect 2445 -550 2495 -530
rect 2445 -580 2455 -550
rect 2485 -580 2495 -550
rect 2445 -600 2495 -580
rect 2445 -630 2455 -600
rect 2485 -630 2495 -600
rect 2445 -650 2495 -630
rect 2445 -680 2455 -650
rect 2485 -680 2495 -650
rect 2445 -690 2495 -680
rect 2530 -500 2580 -490
rect 2530 -530 2540 -500
rect 2570 -530 2580 -500
rect 2530 -550 2580 -530
rect 2530 -580 2540 -550
rect 2570 -580 2580 -550
rect 2530 -600 2580 -580
rect 2530 -630 2540 -600
rect 2570 -630 2580 -600
rect 2530 -650 2580 -630
rect 2530 -680 2540 -650
rect 2570 -680 2580 -650
rect 2530 -690 2580 -680
rect 2615 -500 2665 -490
rect 2615 -530 2625 -500
rect 2655 -530 2665 -500
rect 2615 -550 2665 -530
rect 2615 -580 2625 -550
rect 2655 -580 2665 -550
rect 2615 -600 2665 -580
rect 2615 -630 2625 -600
rect 2655 -630 2665 -600
rect 2615 -650 2665 -630
rect 2615 -680 2625 -650
rect 2655 -680 2665 -650
rect 2615 -690 2665 -680
rect 2700 -500 2750 -490
rect 2700 -530 2710 -500
rect 2740 -530 2750 -500
rect 2700 -550 2750 -530
rect 2700 -580 2710 -550
rect 2740 -580 2750 -550
rect 2700 -600 2750 -580
rect 2700 -630 2710 -600
rect 2740 -630 2750 -600
rect 2700 -650 2750 -630
rect 2700 -680 2710 -650
rect 2740 -680 2750 -650
rect 2700 -690 2750 -680
rect 2785 -500 2835 -490
rect 2785 -530 2795 -500
rect 2825 -530 2835 -500
rect 2785 -550 2835 -530
rect 2785 -580 2795 -550
rect 2825 -580 2835 -550
rect 2785 -600 2835 -580
rect 2785 -630 2795 -600
rect 2825 -630 2835 -600
rect 2785 -650 2835 -630
rect 2785 -680 2795 -650
rect 2825 -680 2835 -650
rect 2785 -690 2835 -680
rect 2870 -500 2920 -490
rect 2870 -530 2880 -500
rect 2910 -530 2920 -500
rect 2870 -550 2920 -530
rect 2870 -580 2880 -550
rect 2910 -580 2920 -550
rect 2870 -600 2920 -580
rect 2870 -630 2880 -600
rect 2910 -630 2920 -600
rect 2870 -650 2920 -630
rect 2870 -680 2880 -650
rect 2910 -680 2920 -650
rect 2870 -690 2920 -680
rect 2955 -500 3005 -490
rect 2955 -530 2965 -500
rect 2995 -530 3005 -500
rect 2955 -550 3005 -530
rect 2955 -580 2965 -550
rect 2995 -580 3005 -550
rect 2955 -600 3005 -580
rect 2955 -630 2965 -600
rect 2995 -630 3005 -600
rect 2955 -650 3005 -630
rect 2955 -680 2965 -650
rect 2995 -680 3005 -650
rect 2955 -690 3005 -680
rect 3040 -500 3090 -490
rect 3040 -530 3050 -500
rect 3080 -530 3090 -500
rect 3040 -550 3090 -530
rect 3040 -580 3050 -550
rect 3080 -580 3090 -550
rect 3040 -600 3090 -580
rect 3040 -630 3050 -600
rect 3080 -630 3090 -600
rect 3040 -650 3090 -630
rect 3040 -680 3050 -650
rect 3080 -680 3090 -650
rect 3040 -690 3090 -680
rect 3125 -500 3175 -490
rect 3125 -530 3135 -500
rect 3165 -530 3175 -500
rect 3125 -550 3175 -530
rect 3125 -580 3135 -550
rect 3165 -580 3175 -550
rect 3125 -600 3175 -580
rect 3125 -630 3135 -600
rect 3165 -630 3175 -600
rect 3125 -650 3175 -630
rect 3125 -680 3135 -650
rect 3165 -680 3175 -650
rect 3125 -690 3175 -680
rect 3210 -500 3260 -490
rect 3210 -530 3220 -500
rect 3250 -530 3260 -500
rect 3210 -550 3260 -530
rect 3210 -580 3220 -550
rect 3250 -580 3260 -550
rect 3210 -600 3260 -580
rect 3210 -630 3220 -600
rect 3250 -630 3260 -600
rect 3210 -650 3260 -630
rect 3210 -680 3220 -650
rect 3250 -680 3260 -650
rect 3210 -690 3260 -680
rect 3295 -500 3345 -490
rect 3295 -530 3305 -500
rect 3335 -530 3345 -500
rect 3295 -550 3345 -530
rect 3295 -580 3305 -550
rect 3335 -580 3345 -550
rect 3295 -600 3345 -580
rect 3295 -630 3305 -600
rect 3335 -630 3345 -600
rect 3295 -650 3345 -630
rect 3295 -680 3305 -650
rect 3335 -680 3345 -650
rect 3295 -690 3345 -680
rect 3380 -500 3430 -490
rect 3380 -530 3390 -500
rect 3420 -530 3430 -500
rect 3380 -550 3430 -530
rect 3380 -580 3390 -550
rect 3420 -580 3430 -550
rect 3380 -600 3430 -580
rect 3380 -630 3390 -600
rect 3420 -630 3430 -600
rect 3380 -650 3430 -630
rect 3380 -680 3390 -650
rect 3420 -680 3430 -650
rect 3380 -690 3430 -680
rect 3465 -500 3515 -490
rect 3465 -530 3475 -500
rect 3505 -530 3515 -500
rect 3465 -550 3515 -530
rect 3465 -580 3475 -550
rect 3505 -580 3515 -550
rect 3465 -600 3515 -580
rect 3465 -630 3475 -600
rect 3505 -630 3515 -600
rect 3465 -650 3515 -630
rect 3465 -680 3475 -650
rect 3505 -680 3515 -650
rect 3465 -690 3515 -680
rect 3550 -500 3600 -490
rect 3550 -530 3560 -500
rect 3590 -530 3600 -500
rect 3550 -550 3600 -530
rect 3550 -580 3560 -550
rect 3590 -580 3600 -550
rect 3550 -600 3600 -580
rect 3550 -630 3560 -600
rect 3590 -630 3600 -600
rect 3550 -650 3600 -630
rect 3550 -680 3560 -650
rect 3590 -680 3600 -650
rect 3550 -690 3600 -680
rect 3635 -500 3685 -490
rect 3635 -530 3645 -500
rect 3675 -530 3685 -500
rect 3635 -550 3685 -530
rect 3635 -580 3645 -550
rect 3675 -580 3685 -550
rect 3635 -600 3685 -580
rect 3635 -630 3645 -600
rect 3675 -630 3685 -600
rect 3635 -650 3685 -630
rect 3635 -680 3645 -650
rect 3675 -680 3685 -650
rect 3635 -690 3685 -680
rect 3720 -500 3770 -490
rect 3720 -530 3730 -500
rect 3760 -530 3770 -500
rect 3720 -550 3770 -530
rect 3720 -580 3730 -550
rect 3760 -580 3770 -550
rect 3720 -600 3770 -580
rect 3720 -630 3730 -600
rect 3760 -630 3770 -600
rect 3720 -650 3770 -630
rect 3720 -680 3730 -650
rect 3760 -680 3770 -650
rect 3720 -690 3770 -680
rect 3805 -500 3855 -490
rect 3805 -530 3815 -500
rect 3845 -530 3855 -500
rect 3805 -550 3855 -530
rect 3805 -580 3815 -550
rect 3845 -580 3855 -550
rect 3805 -600 3855 -580
rect 3805 -630 3815 -600
rect 3845 -630 3855 -600
rect 3805 -650 3855 -630
rect 3805 -680 3815 -650
rect 3845 -680 3855 -650
rect 3805 -690 3855 -680
rect 3890 -500 3940 -490
rect 3890 -530 3900 -500
rect 3930 -530 3940 -500
rect 3890 -550 3940 -530
rect 3890 -580 3900 -550
rect 3930 -580 3940 -550
rect 3890 -600 3940 -580
rect 3890 -630 3900 -600
rect 3930 -630 3940 -600
rect 3890 -650 3940 -630
rect 3890 -680 3900 -650
rect 3930 -680 3940 -650
rect 3890 -690 3940 -680
rect 3975 -500 4025 -490
rect 3975 -530 3985 -500
rect 4015 -530 4025 -500
rect 3975 -550 4025 -530
rect 3975 -580 3985 -550
rect 4015 -580 4025 -550
rect 3975 -600 4025 -580
rect 3975 -630 3985 -600
rect 4015 -630 4025 -600
rect 3975 -650 4025 -630
rect 3975 -680 3985 -650
rect 4015 -680 4025 -650
rect 3975 -690 4025 -680
rect 4060 -500 4110 -490
rect 4060 -530 4070 -500
rect 4100 -530 4110 -500
rect 4060 -550 4110 -530
rect 4060 -580 4070 -550
rect 4100 -580 4110 -550
rect 4060 -600 4110 -580
rect 4060 -630 4070 -600
rect 4100 -630 4110 -600
rect 4060 -650 4110 -630
rect 4060 -680 4070 -650
rect 4100 -680 4110 -650
rect 4060 -690 4110 -680
rect 4145 -500 4195 -490
rect 4145 -530 4155 -500
rect 4185 -530 4195 -500
rect 4145 -550 4195 -530
rect 4145 -580 4155 -550
rect 4185 -580 4195 -550
rect 4145 -600 4195 -580
rect 4145 -630 4155 -600
rect 4185 -630 4195 -600
rect 4145 -650 4195 -630
rect 4145 -680 4155 -650
rect 4185 -680 4195 -650
rect 4145 -690 4195 -680
rect 4230 -500 4280 -490
rect 4230 -530 4240 -500
rect 4270 -530 4280 -500
rect 4230 -550 4280 -530
rect 4230 -580 4240 -550
rect 4270 -580 4280 -550
rect 4230 -600 4280 -580
rect 4230 -630 4240 -600
rect 4270 -630 4280 -600
rect 4230 -650 4280 -630
rect 4230 -680 4240 -650
rect 4270 -680 4280 -650
rect 4230 -690 4280 -680
rect 4315 -500 4365 -490
rect 4315 -530 4325 -500
rect 4355 -530 4365 -500
rect 4315 -550 4365 -530
rect 4315 -580 4325 -550
rect 4355 -580 4365 -550
rect 4315 -600 4365 -580
rect 4315 -630 4325 -600
rect 4355 -630 4365 -600
rect 4315 -650 4365 -630
rect 4315 -680 4325 -650
rect 4355 -680 4365 -650
rect 4315 -690 4365 -680
rect 4400 -500 4450 -490
rect 4400 -530 4410 -500
rect 4440 -530 4450 -500
rect 4400 -550 4450 -530
rect 4400 -580 4410 -550
rect 4440 -580 4450 -550
rect 4400 -600 4450 -580
rect 4400 -630 4410 -600
rect 4440 -630 4450 -600
rect 4400 -650 4450 -630
rect 4400 -680 4410 -650
rect 4440 -680 4450 -650
rect 4400 -690 4450 -680
rect 4485 -500 4535 -490
rect 4485 -530 4495 -500
rect 4525 -530 4535 -500
rect 4485 -550 4535 -530
rect 4485 -580 4495 -550
rect 4525 -580 4535 -550
rect 4485 -600 4535 -580
rect 4485 -630 4495 -600
rect 4525 -630 4535 -600
rect 4485 -650 4535 -630
rect 4485 -680 4495 -650
rect 4525 -680 4535 -650
rect 4485 -690 4535 -680
rect 4570 -500 4620 -490
rect 4570 -530 4580 -500
rect 4610 -530 4620 -500
rect 4570 -550 4620 -530
rect 4570 -580 4580 -550
rect 4610 -580 4620 -550
rect 4570 -600 4620 -580
rect 4570 -630 4580 -600
rect 4610 -630 4620 -600
rect 4570 -650 4620 -630
rect 4570 -680 4580 -650
rect 4610 -680 4620 -650
rect 4570 -690 4620 -680
rect 4655 -500 4705 -490
rect 4655 -530 4665 -500
rect 4695 -530 4705 -500
rect 4655 -550 4705 -530
rect 4655 -580 4665 -550
rect 4695 -580 4705 -550
rect 4655 -600 4705 -580
rect 4655 -630 4665 -600
rect 4695 -630 4705 -600
rect 4655 -650 4705 -630
rect 4655 -680 4665 -650
rect 4695 -680 4705 -650
rect 4655 -690 4705 -680
rect 4740 -500 4790 -490
rect 4740 -530 4750 -500
rect 4780 -530 4790 -500
rect 4740 -550 4790 -530
rect 4740 -580 4750 -550
rect 4780 -580 4790 -550
rect 4740 -600 4790 -580
rect 4740 -630 4750 -600
rect 4780 -630 4790 -600
rect 4740 -650 4790 -630
rect 4740 -680 4750 -650
rect 4780 -680 4790 -650
rect 4740 -690 4790 -680
rect 4825 -500 4875 -490
rect 4825 -530 4835 -500
rect 4865 -530 4875 -500
rect 4825 -550 4875 -530
rect 4825 -580 4835 -550
rect 4865 -580 4875 -550
rect 4825 -600 4875 -580
rect 4825 -630 4835 -600
rect 4865 -630 4875 -600
rect 4825 -650 4875 -630
rect 4825 -680 4835 -650
rect 4865 -680 4875 -650
rect 4825 -690 4875 -680
rect 4910 -500 4960 -490
rect 4910 -530 4920 -500
rect 4950 -530 4960 -500
rect 4910 -550 4960 -530
rect 4910 -580 4920 -550
rect 4950 -580 4960 -550
rect 4910 -600 4960 -580
rect 4910 -630 4920 -600
rect 4950 -630 4960 -600
rect 4910 -650 4960 -630
rect 4910 -680 4920 -650
rect 4950 -680 4960 -650
rect 4910 -690 4960 -680
rect 4995 -500 5045 -490
rect 4995 -530 5005 -500
rect 5035 -530 5045 -500
rect 4995 -550 5045 -530
rect 4995 -580 5005 -550
rect 5035 -580 5045 -550
rect 4995 -600 5045 -580
rect 4995 -630 5005 -600
rect 5035 -630 5045 -600
rect 4995 -650 5045 -630
rect 4995 -680 5005 -650
rect 5035 -680 5045 -650
rect 4995 -690 5045 -680
rect 5080 -500 5130 -490
rect 5080 -530 5090 -500
rect 5120 -530 5130 -500
rect 5080 -550 5130 -530
rect 5080 -580 5090 -550
rect 5120 -580 5130 -550
rect 5080 -600 5130 -580
rect 5080 -630 5090 -600
rect 5120 -630 5130 -600
rect 5080 -650 5130 -630
rect 5080 -680 5090 -650
rect 5120 -680 5130 -650
rect 5080 -690 5130 -680
rect 5165 -500 5215 -490
rect 5165 -530 5175 -500
rect 5205 -530 5215 -500
rect 5165 -550 5215 -530
rect 5165 -580 5175 -550
rect 5205 -580 5215 -550
rect 5165 -600 5215 -580
rect 5165 -630 5175 -600
rect 5205 -630 5215 -600
rect 5165 -650 5215 -630
rect 5165 -680 5175 -650
rect 5205 -680 5215 -650
rect 5165 -690 5215 -680
rect 5250 -500 5300 -490
rect 5250 -530 5260 -500
rect 5290 -530 5300 -500
rect 5250 -550 5300 -530
rect 5250 -580 5260 -550
rect 5290 -580 5300 -550
rect 5250 -600 5300 -580
rect 5250 -630 5260 -600
rect 5290 -630 5300 -600
rect 5250 -650 5300 -630
rect 5250 -680 5260 -650
rect 5290 -680 5300 -650
rect 5250 -690 5300 -680
rect 5335 -500 5385 -490
rect 5335 -530 5345 -500
rect 5375 -530 5385 -500
rect 5335 -550 5385 -530
rect 5335 -580 5345 -550
rect 5375 -580 5385 -550
rect 5335 -600 5385 -580
rect 5335 -630 5345 -600
rect 5375 -630 5385 -600
rect 5335 -650 5385 -630
rect 5335 -680 5345 -650
rect 5375 -680 5385 -650
rect 5335 -690 5385 -680
rect 5420 -500 5470 -490
rect 5420 -530 5430 -500
rect 5460 -530 5470 -500
rect 5420 -550 5470 -530
rect 5420 -580 5430 -550
rect 5460 -580 5470 -550
rect 5420 -600 5470 -580
rect 5420 -630 5430 -600
rect 5460 -630 5470 -600
rect 5420 -650 5470 -630
rect 5420 -680 5430 -650
rect 5460 -680 5470 -650
rect 5420 -690 5470 -680
rect 5505 -500 5555 -490
rect 5505 -530 5515 -500
rect 5545 -530 5555 -500
rect 5505 -550 5555 -530
rect 5505 -580 5515 -550
rect 5545 -580 5555 -550
rect 5505 -600 5555 -580
rect 5505 -630 5515 -600
rect 5545 -630 5555 -600
rect 5505 -650 5555 -630
rect 5505 -680 5515 -650
rect 5545 -680 5555 -650
rect 5505 -690 5555 -680
rect 5590 -500 5640 -490
rect 5590 -530 5600 -500
rect 5630 -530 5640 -500
rect 5590 -550 5640 -530
rect 5590 -580 5600 -550
rect 5630 -580 5640 -550
rect 5590 -600 5640 -580
rect 5590 -630 5600 -600
rect 5630 -630 5640 -600
rect 5590 -650 5640 -630
rect 5590 -680 5600 -650
rect 5630 -680 5640 -650
rect 5590 -690 5640 -680
rect 5675 -500 5725 -490
rect 5675 -530 5685 -500
rect 5715 -530 5725 -500
rect 5675 -550 5725 -530
rect 5675 -580 5685 -550
rect 5715 -580 5725 -550
rect 5675 -600 5725 -580
rect 5675 -630 5685 -600
rect 5715 -630 5725 -600
rect 5675 -650 5725 -630
rect 5675 -680 5685 -650
rect 5715 -680 5725 -650
rect 5675 -690 5725 -680
rect 5760 -500 5810 -490
rect 5760 -530 5770 -500
rect 5800 -530 5810 -500
rect 5760 -550 5810 -530
rect 5760 -580 5770 -550
rect 5800 -580 5810 -550
rect 5760 -600 5810 -580
rect 5760 -630 5770 -600
rect 5800 -630 5810 -600
rect 5760 -650 5810 -630
rect 5760 -680 5770 -650
rect 5800 -680 5810 -650
rect 5760 -690 5810 -680
rect 5845 -500 5895 -490
rect 5845 -530 5855 -500
rect 5885 -530 5895 -500
rect 5845 -550 5895 -530
rect 5845 -580 5855 -550
rect 5885 -580 5895 -550
rect 5845 -600 5895 -580
rect 5845 -630 5855 -600
rect 5885 -630 5895 -600
rect 5845 -650 5895 -630
rect 5845 -680 5855 -650
rect 5885 -680 5895 -650
rect 5845 -690 5895 -680
rect 5930 -500 5980 -490
rect 5930 -530 5940 -500
rect 5970 -530 5980 -500
rect 5930 -550 5980 -530
rect 5930 -580 5940 -550
rect 5970 -580 5980 -550
rect 5930 -600 5980 -580
rect 5930 -630 5940 -600
rect 5970 -630 5980 -600
rect 5930 -650 5980 -630
rect 5930 -680 5940 -650
rect 5970 -680 5980 -650
rect 5930 -690 5980 -680
rect 6015 -500 6065 -490
rect 6015 -530 6025 -500
rect 6055 -530 6065 -500
rect 6015 -550 6065 -530
rect 6015 -580 6025 -550
rect 6055 -580 6065 -550
rect 6015 -600 6065 -580
rect 6015 -630 6025 -600
rect 6055 -630 6065 -600
rect 6015 -650 6065 -630
rect 6015 -680 6025 -650
rect 6055 -680 6065 -650
rect 6015 -690 6065 -680
rect 6100 -500 6150 -490
rect 6100 -530 6110 -500
rect 6140 -530 6150 -500
rect 6100 -550 6150 -530
rect 6100 -580 6110 -550
rect 6140 -580 6150 -550
rect 6100 -600 6150 -580
rect 6100 -630 6110 -600
rect 6140 -630 6150 -600
rect 6100 -650 6150 -630
rect 6100 -680 6110 -650
rect 6140 -680 6150 -650
rect 6100 -690 6150 -680
rect 6185 -500 6235 -490
rect 6185 -530 6195 -500
rect 6225 -530 6235 -500
rect 6185 -550 6235 -530
rect 6185 -580 6195 -550
rect 6225 -580 6235 -550
rect 6185 -600 6235 -580
rect 6185 -630 6195 -600
rect 6225 -630 6235 -600
rect 6185 -650 6235 -630
rect 6185 -680 6195 -650
rect 6225 -680 6235 -650
rect 6185 -690 6235 -680
rect 6270 -500 6320 -490
rect 6270 -530 6280 -500
rect 6310 -530 6320 -500
rect 6270 -550 6320 -530
rect 6270 -580 6280 -550
rect 6310 -580 6320 -550
rect 6270 -600 6320 -580
rect 6270 -630 6280 -600
rect 6310 -630 6320 -600
rect 6270 -650 6320 -630
rect 6270 -680 6280 -650
rect 6310 -680 6320 -650
rect 6270 -690 6320 -680
rect 6355 -500 6405 -490
rect 6355 -530 6365 -500
rect 6395 -530 6405 -500
rect 6355 -550 6405 -530
rect 6355 -580 6365 -550
rect 6395 -580 6405 -550
rect 6355 -600 6405 -580
rect 6355 -630 6365 -600
rect 6395 -630 6405 -600
rect 6355 -650 6405 -630
rect 6355 -680 6365 -650
rect 6395 -680 6405 -650
rect 6355 -690 6405 -680
rect 6440 -500 6490 -490
rect 6440 -530 6450 -500
rect 6480 -530 6490 -500
rect 6440 -550 6490 -530
rect 6440 -580 6450 -550
rect 6480 -580 6490 -550
rect 6440 -600 6490 -580
rect 6440 -630 6450 -600
rect 6480 -630 6490 -600
rect 6440 -650 6490 -630
rect 6440 -680 6450 -650
rect 6480 -680 6490 -650
rect 6440 -690 6490 -680
rect 6525 -500 6575 -490
rect 6525 -530 6535 -500
rect 6565 -530 6575 -500
rect 6525 -550 6575 -530
rect 6525 -580 6535 -550
rect 6565 -580 6575 -550
rect 6525 -600 6575 -580
rect 6525 -630 6535 -600
rect 6565 -630 6575 -600
rect 6525 -650 6575 -630
rect 6525 -680 6535 -650
rect 6565 -680 6575 -650
rect 6525 -690 6575 -680
rect 6610 -500 6660 -490
rect 6610 -530 6620 -500
rect 6650 -530 6660 -500
rect 6610 -550 6660 -530
rect 6610 -580 6620 -550
rect 6650 -580 6660 -550
rect 6610 -600 6660 -580
rect 6610 -630 6620 -600
rect 6650 -630 6660 -600
rect 6610 -650 6660 -630
rect 6610 -680 6620 -650
rect 6650 -680 6660 -650
rect 6610 -690 6660 -680
rect 6695 -500 6745 -490
rect 6695 -530 6705 -500
rect 6735 -530 6745 -500
rect 6695 -550 6745 -530
rect 6695 -580 6705 -550
rect 6735 -580 6745 -550
rect 6695 -600 6745 -580
rect 6695 -630 6705 -600
rect 6735 -630 6745 -600
rect 6695 -650 6745 -630
rect 6695 -680 6705 -650
rect 6735 -680 6745 -650
rect 6695 -690 6745 -680
rect 6780 -500 6830 -490
rect 6780 -530 6790 -500
rect 6820 -530 6830 -500
rect 6780 -550 6830 -530
rect 6780 -580 6790 -550
rect 6820 -580 6830 -550
rect 6780 -600 6830 -580
rect 6780 -630 6790 -600
rect 6820 -630 6830 -600
rect 6780 -650 6830 -630
rect 6780 -680 6790 -650
rect 6820 -680 6830 -650
rect 6780 -690 6830 -680
rect 6865 -500 6915 -490
rect 6865 -530 6875 -500
rect 6905 -530 6915 -500
rect 6865 -550 6915 -530
rect 6865 -580 6875 -550
rect 6905 -580 6915 -550
rect 6865 -600 6915 -580
rect 6865 -630 6875 -600
rect 6905 -630 6915 -600
rect 6865 -650 6915 -630
rect 6865 -680 6875 -650
rect 6905 -680 6915 -650
rect 6865 -690 6915 -680
rect 6950 -500 7000 -490
rect 6950 -530 6960 -500
rect 6990 -530 7000 -500
rect 6950 -550 7000 -530
rect 6950 -580 6960 -550
rect 6990 -580 7000 -550
rect 6950 -600 7000 -580
rect 6950 -630 6960 -600
rect 6990 -630 7000 -600
rect 6950 -650 7000 -630
rect 6950 -680 6960 -650
rect 6990 -680 7000 -650
rect 6950 -690 7000 -680
rect 7035 -500 7085 -490
rect 7035 -530 7045 -500
rect 7075 -530 7085 -500
rect 7035 -550 7085 -530
rect 7035 -580 7045 -550
rect 7075 -580 7085 -550
rect 7035 -600 7085 -580
rect 7035 -630 7045 -600
rect 7075 -630 7085 -600
rect 7035 -650 7085 -630
rect 7035 -680 7045 -650
rect 7075 -680 7085 -650
rect 7035 -690 7085 -680
rect 7120 -500 7170 -490
rect 7120 -530 7130 -500
rect 7160 -530 7170 -500
rect 7120 -550 7170 -530
rect 7120 -580 7130 -550
rect 7160 -580 7170 -550
rect 7120 -600 7170 -580
rect 7120 -630 7130 -600
rect 7160 -630 7170 -600
rect 7120 -650 7170 -630
rect 7120 -680 7130 -650
rect 7160 -680 7170 -650
rect 7120 -690 7170 -680
rect 7205 -500 7255 -490
rect 7205 -530 7215 -500
rect 7245 -530 7255 -500
rect 7205 -550 7255 -530
rect 7205 -580 7215 -550
rect 7245 -580 7255 -550
rect 7205 -600 7255 -580
rect 7205 -630 7215 -600
rect 7245 -630 7255 -600
rect 7205 -650 7255 -630
rect 7205 -680 7215 -650
rect 7245 -680 7255 -650
rect 7205 -690 7255 -680
rect 7290 -500 7340 -490
rect 7290 -530 7300 -500
rect 7330 -530 7340 -500
rect 7290 -550 7340 -530
rect 7290 -580 7300 -550
rect 7330 -580 7340 -550
rect 7290 -600 7340 -580
rect 7290 -630 7300 -600
rect 7330 -630 7340 -600
rect 7290 -650 7340 -630
rect 7290 -680 7300 -650
rect 7330 -680 7340 -650
rect 7290 -690 7340 -680
rect 7375 -500 7425 -490
rect 7375 -530 7385 -500
rect 7415 -530 7425 -500
rect 7375 -550 7425 -530
rect 7375 -580 7385 -550
rect 7415 -580 7425 -550
rect 7375 -600 7425 -580
rect 7375 -630 7385 -600
rect 7415 -630 7425 -600
rect 7375 -650 7425 -630
rect 7375 -680 7385 -650
rect 7415 -680 7425 -650
rect 7375 -690 7425 -680
rect 7460 -500 7510 -490
rect 7460 -530 7470 -500
rect 7500 -530 7510 -500
rect 7460 -550 7510 -530
rect 7460 -580 7470 -550
rect 7500 -580 7510 -550
rect 7460 -600 7510 -580
rect 7460 -630 7470 -600
rect 7500 -630 7510 -600
rect 7460 -650 7510 -630
rect 7460 -680 7470 -650
rect 7500 -680 7510 -650
rect 7460 -690 7510 -680
rect 7545 -500 7595 -490
rect 7545 -530 7555 -500
rect 7585 -530 7595 -500
rect 7545 -550 7595 -530
rect 7545 -580 7555 -550
rect 7585 -580 7595 -550
rect 7545 -600 7595 -580
rect 7545 -630 7555 -600
rect 7585 -630 7595 -600
rect 7545 -650 7595 -630
rect 7545 -680 7555 -650
rect 7585 -680 7595 -650
rect 7545 -690 7595 -680
rect 7630 -500 7680 -490
rect 7630 -530 7640 -500
rect 7670 -530 7680 -500
rect 7630 -550 7680 -530
rect 7630 -580 7640 -550
rect 7670 -580 7680 -550
rect 7630 -600 7680 -580
rect 7630 -630 7640 -600
rect 7670 -630 7680 -600
rect 7630 -650 7680 -630
rect 7630 -680 7640 -650
rect 7670 -680 7680 -650
rect 7630 -690 7680 -680
rect 7715 -500 7765 -490
rect 7715 -530 7725 -500
rect 7755 -530 7765 -500
rect 7715 -550 7765 -530
rect 7715 -580 7725 -550
rect 7755 -580 7765 -550
rect 7715 -600 7765 -580
rect 7715 -630 7725 -600
rect 7755 -630 7765 -600
rect 7715 -650 7765 -630
rect 7715 -680 7725 -650
rect 7755 -680 7765 -650
rect 7715 -690 7765 -680
rect 7800 -500 7850 -490
rect 7800 -530 7810 -500
rect 7840 -530 7850 -500
rect 7800 -550 7850 -530
rect 7800 -580 7810 -550
rect 7840 -580 7850 -550
rect 7800 -600 7850 -580
rect 7800 -630 7810 -600
rect 7840 -630 7850 -600
rect 7800 -650 7850 -630
rect 7800 -680 7810 -650
rect 7840 -680 7850 -650
rect 7800 -690 7850 -680
rect 7885 -500 7935 -490
rect 7885 -530 7895 -500
rect 7925 -530 7935 -500
rect 7885 -550 7935 -530
rect 7885 -580 7895 -550
rect 7925 -580 7935 -550
rect 7885 -600 7935 -580
rect 7885 -630 7895 -600
rect 7925 -630 7935 -600
rect 7885 -650 7935 -630
rect 7885 -680 7895 -650
rect 7925 -680 7935 -650
rect 7885 -690 7935 -680
rect 7970 -500 8020 -490
rect 7970 -530 7980 -500
rect 8010 -530 8020 -500
rect 7970 -550 8020 -530
rect 7970 -580 7980 -550
rect 8010 -580 8020 -550
rect 7970 -600 8020 -580
rect 7970 -630 7980 -600
rect 8010 -630 8020 -600
rect 7970 -650 8020 -630
rect 7970 -680 7980 -650
rect 8010 -680 8020 -650
rect 7970 -690 8020 -680
rect 8055 -500 8105 -490
rect 8055 -530 8065 -500
rect 8095 -530 8105 -500
rect 8055 -550 8105 -530
rect 8055 -580 8065 -550
rect 8095 -580 8105 -550
rect 8055 -600 8105 -580
rect 8055 -630 8065 -600
rect 8095 -630 8105 -600
rect 8055 -650 8105 -630
rect 8055 -680 8065 -650
rect 8095 -680 8105 -650
rect 8055 -690 8105 -680
rect 8140 -500 8190 -490
rect 8140 -530 8150 -500
rect 8180 -530 8190 -500
rect 8140 -550 8190 -530
rect 8140 -580 8150 -550
rect 8180 -580 8190 -550
rect 8140 -600 8190 -580
rect 8140 -630 8150 -600
rect 8180 -630 8190 -600
rect 8140 -650 8190 -630
rect 8140 -680 8150 -650
rect 8180 -680 8190 -650
rect 8140 -690 8190 -680
rect 8225 -500 8275 -490
rect 8225 -530 8235 -500
rect 8265 -530 8275 -500
rect 8225 -550 8275 -530
rect 8225 -580 8235 -550
rect 8265 -580 8275 -550
rect 8225 -600 8275 -580
rect 8225 -630 8235 -600
rect 8265 -630 8275 -600
rect 8225 -650 8275 -630
rect 8225 -680 8235 -650
rect 8265 -680 8275 -650
rect 8225 -690 8275 -680
rect 8310 -500 8360 -490
rect 8310 -530 8320 -500
rect 8350 -530 8360 -500
rect 8310 -550 8360 -530
rect 8310 -580 8320 -550
rect 8350 -580 8360 -550
rect 8310 -600 8360 -580
rect 8310 -630 8320 -600
rect 8350 -630 8360 -600
rect 8310 -650 8360 -630
rect 8310 -680 8320 -650
rect 8350 -680 8360 -650
rect 8310 -690 8360 -680
rect 8395 -500 8445 -490
rect 8395 -530 8405 -500
rect 8435 -530 8445 -500
rect 8395 -550 8445 -530
rect 8395 -580 8405 -550
rect 8435 -580 8445 -550
rect 8395 -600 8445 -580
rect 8395 -630 8405 -600
rect 8435 -630 8445 -600
rect 8395 -650 8445 -630
rect 8395 -680 8405 -650
rect 8435 -680 8445 -650
rect 8395 -690 8445 -680
rect 8480 -500 8530 -490
rect 8480 -530 8490 -500
rect 8520 -530 8530 -500
rect 8480 -550 8530 -530
rect 8480 -580 8490 -550
rect 8520 -580 8530 -550
rect 8480 -600 8530 -580
rect 8480 -630 8490 -600
rect 8520 -630 8530 -600
rect 8480 -650 8530 -630
rect 8480 -680 8490 -650
rect 8520 -680 8530 -650
rect 8480 -690 8530 -680
rect 8565 -500 8615 -490
rect 8565 -530 8575 -500
rect 8605 -530 8615 -500
rect 8565 -550 8615 -530
rect 8565 -580 8575 -550
rect 8605 -580 8615 -550
rect 8565 -600 8615 -580
rect 8565 -630 8575 -600
rect 8605 -630 8615 -600
rect 8565 -650 8615 -630
rect 8565 -680 8575 -650
rect 8605 -680 8615 -650
rect 8565 -690 8615 -680
rect 8650 -500 8700 -490
rect 8650 -530 8660 -500
rect 8690 -530 8700 -500
rect 8650 -550 8700 -530
rect 8650 -580 8660 -550
rect 8690 -580 8700 -550
rect 8650 -600 8700 -580
rect 8650 -630 8660 -600
rect 8690 -630 8700 -600
rect 8650 -650 8700 -630
rect 8650 -680 8660 -650
rect 8690 -680 8700 -650
rect 8650 -690 8700 -680
rect 8735 -500 8785 -490
rect 8735 -530 8745 -500
rect 8775 -530 8785 -500
rect 8735 -550 8785 -530
rect 8735 -580 8745 -550
rect 8775 -580 8785 -550
rect 8735 -600 8785 -580
rect 8735 -630 8745 -600
rect 8775 -630 8785 -600
rect 8735 -650 8785 -630
rect 8735 -680 8745 -650
rect 8775 -680 8785 -650
rect 8735 -690 8785 -680
rect 8820 -500 8870 -490
rect 8820 -530 8830 -500
rect 8860 -530 8870 -500
rect 8820 -550 8870 -530
rect 8820 -580 8830 -550
rect 8860 -580 8870 -550
rect 8820 -600 8870 -580
rect 8820 -630 8830 -600
rect 8860 -630 8870 -600
rect 8820 -650 8870 -630
rect 8820 -680 8830 -650
rect 8860 -680 8870 -650
rect 8820 -690 8870 -680
rect 8905 -500 8955 -490
rect 8905 -530 8915 -500
rect 8945 -530 8955 -500
rect 8905 -550 8955 -530
rect 8905 -580 8915 -550
rect 8945 -580 8955 -550
rect 8905 -600 8955 -580
rect 8905 -630 8915 -600
rect 8945 -630 8955 -600
rect 8905 -650 8955 -630
rect 8905 -680 8915 -650
rect 8945 -680 8955 -650
rect 8905 -690 8955 -680
rect 8990 -500 9040 -490
rect 8990 -530 9000 -500
rect 9030 -530 9040 -500
rect 8990 -550 9040 -530
rect 8990 -580 9000 -550
rect 9030 -580 9040 -550
rect 8990 -600 9040 -580
rect 8990 -630 9000 -600
rect 9030 -630 9040 -600
rect 8990 -650 9040 -630
rect 8990 -680 9000 -650
rect 9030 -680 9040 -650
rect 8990 -690 9040 -680
rect 9075 -500 9125 -490
rect 9075 -530 9085 -500
rect 9115 -530 9125 -500
rect 9075 -550 9125 -530
rect 9075 -580 9085 -550
rect 9115 -580 9125 -550
rect 9075 -600 9125 -580
rect 9075 -630 9085 -600
rect 9115 -630 9125 -600
rect 9075 -650 9125 -630
rect 9075 -680 9085 -650
rect 9115 -680 9125 -650
rect 9075 -690 9125 -680
rect 9160 -500 9210 -490
rect 9160 -530 9170 -500
rect 9200 -530 9210 -500
rect 9160 -550 9210 -530
rect 9160 -580 9170 -550
rect 9200 -580 9210 -550
rect 9160 -600 9210 -580
rect 9160 -630 9170 -600
rect 9200 -630 9210 -600
rect 9160 -650 9210 -630
rect 9160 -680 9170 -650
rect 9200 -680 9210 -650
rect 9160 -690 9210 -680
rect 9245 -500 9295 -490
rect 9245 -530 9255 -500
rect 9285 -530 9295 -500
rect 9245 -550 9295 -530
rect 9245 -580 9255 -550
rect 9285 -580 9295 -550
rect 9245 -600 9295 -580
rect 9245 -630 9255 -600
rect 9285 -630 9295 -600
rect 9245 -650 9295 -630
rect 9245 -680 9255 -650
rect 9285 -680 9295 -650
rect 9245 -690 9295 -680
rect 9330 -500 9380 -490
rect 9330 -530 9340 -500
rect 9370 -530 9380 -500
rect 9330 -550 9380 -530
rect 9330 -580 9340 -550
rect 9370 -580 9380 -550
rect 9330 -600 9380 -580
rect 9330 -630 9340 -600
rect 9370 -630 9380 -600
rect 9330 -650 9380 -630
rect 9330 -680 9340 -650
rect 9370 -680 9380 -650
rect 9330 -690 9380 -680
rect 9415 -500 9465 -490
rect 9415 -530 9425 -500
rect 9455 -530 9465 -500
rect 9415 -550 9465 -530
rect 9415 -580 9425 -550
rect 9455 -580 9465 -550
rect 9415 -600 9465 -580
rect 9415 -630 9425 -600
rect 9455 -630 9465 -600
rect 9415 -650 9465 -630
rect 9415 -680 9425 -650
rect 9455 -680 9465 -650
rect 9415 -690 9465 -680
rect 9500 -500 9550 -490
rect 9500 -530 9510 -500
rect 9540 -530 9550 -500
rect 9500 -550 9550 -530
rect 9500 -580 9510 -550
rect 9540 -580 9550 -550
rect 9500 -600 9550 -580
rect 9500 -630 9510 -600
rect 9540 -630 9550 -600
rect 9500 -650 9550 -630
rect 9500 -680 9510 -650
rect 9540 -680 9550 -650
rect 9500 -690 9550 -680
rect 9585 -500 9635 -490
rect 9585 -530 9595 -500
rect 9625 -530 9635 -500
rect 9585 -550 9635 -530
rect 9585 -580 9595 -550
rect 9625 -580 9635 -550
rect 9585 -600 9635 -580
rect 9585 -630 9595 -600
rect 9625 -630 9635 -600
rect 9585 -650 9635 -630
rect 9585 -680 9595 -650
rect 9625 -680 9635 -650
rect 9585 -690 9635 -680
rect 9670 -500 9720 -490
rect 9670 -530 9680 -500
rect 9710 -530 9720 -500
rect 9670 -550 9720 -530
rect 9670 -580 9680 -550
rect 9710 -580 9720 -550
rect 9670 -600 9720 -580
rect 9670 -630 9680 -600
rect 9710 -630 9720 -600
rect 9670 -650 9720 -630
rect 9670 -680 9680 -650
rect 9710 -680 9720 -650
rect 9670 -690 9720 -680
rect 9755 -500 9805 -490
rect 9755 -530 9765 -500
rect 9795 -530 9805 -500
rect 9755 -550 9805 -530
rect 9755 -580 9765 -550
rect 9795 -580 9805 -550
rect 9755 -600 9805 -580
rect 9755 -630 9765 -600
rect 9795 -630 9805 -600
rect 9755 -650 9805 -630
rect 9755 -680 9765 -650
rect 9795 -680 9805 -650
rect 9755 -690 9805 -680
rect 9840 -500 9890 -490
rect 9840 -530 9850 -500
rect 9880 -530 9890 -500
rect 9840 -550 9890 -530
rect 9840 -580 9850 -550
rect 9880 -580 9890 -550
rect 9840 -600 9890 -580
rect 9840 -630 9850 -600
rect 9880 -630 9890 -600
rect 9840 -650 9890 -630
rect 9840 -680 9850 -650
rect 9880 -680 9890 -650
rect 9840 -690 9890 -680
rect 9925 -500 9975 -490
rect 9925 -530 9935 -500
rect 9965 -530 9975 -500
rect 9925 -550 9975 -530
rect 9925 -580 9935 -550
rect 9965 -580 9975 -550
rect 9925 -600 9975 -580
rect 9925 -630 9935 -600
rect 9965 -630 9975 -600
rect 9925 -650 9975 -630
rect 9925 -680 9935 -650
rect 9965 -680 9975 -650
rect 9925 -690 9975 -680
rect 10010 -500 10060 -490
rect 10010 -530 10020 -500
rect 10050 -530 10060 -500
rect 10010 -550 10060 -530
rect 10010 -580 10020 -550
rect 10050 -580 10060 -550
rect 10010 -600 10060 -580
rect 10010 -630 10020 -600
rect 10050 -630 10060 -600
rect 10010 -650 10060 -630
rect 10010 -680 10020 -650
rect 10050 -680 10060 -650
rect 10010 -690 10060 -680
rect 10095 -500 10145 -490
rect 10095 -530 10105 -500
rect 10135 -530 10145 -500
rect 10095 -550 10145 -530
rect 10095 -580 10105 -550
rect 10135 -580 10145 -550
rect 10095 -600 10145 -580
rect 10095 -630 10105 -600
rect 10135 -630 10145 -600
rect 10095 -650 10145 -630
rect 10095 -680 10105 -650
rect 10135 -680 10145 -650
rect 10095 -690 10145 -680
rect 10180 -500 10230 -490
rect 10180 -530 10190 -500
rect 10220 -530 10230 -500
rect 10180 -550 10230 -530
rect 10180 -580 10190 -550
rect 10220 -580 10230 -550
rect 10180 -600 10230 -580
rect 10180 -630 10190 -600
rect 10220 -630 10230 -600
rect 10180 -650 10230 -630
rect 10180 -680 10190 -650
rect 10220 -680 10230 -650
rect 10180 -690 10230 -680
rect 10265 -500 10315 -490
rect 10265 -530 10275 -500
rect 10305 -530 10315 -500
rect 10265 -550 10315 -530
rect 10265 -580 10275 -550
rect 10305 -580 10315 -550
rect 10265 -600 10315 -580
rect 10265 -630 10275 -600
rect 10305 -630 10315 -600
rect 10265 -650 10315 -630
rect 10265 -680 10275 -650
rect 10305 -680 10315 -650
rect 10265 -690 10315 -680
rect 10350 -500 10400 -490
rect 10350 -530 10360 -500
rect 10390 -530 10400 -500
rect 10350 -550 10400 -530
rect 10350 -580 10360 -550
rect 10390 -580 10400 -550
rect 10350 -600 10400 -580
rect 10350 -630 10360 -600
rect 10390 -630 10400 -600
rect 10350 -650 10400 -630
rect 10350 -680 10360 -650
rect 10390 -680 10400 -650
rect 10350 -690 10400 -680
rect 10435 -500 10485 -490
rect 10435 -530 10445 -500
rect 10475 -530 10485 -500
rect 10435 -550 10485 -530
rect 10435 -580 10445 -550
rect 10475 -580 10485 -550
rect 10435 -600 10485 -580
rect 10435 -630 10445 -600
rect 10475 -630 10485 -600
rect 10435 -650 10485 -630
rect 10435 -680 10445 -650
rect 10475 -680 10485 -650
rect 10435 -690 10485 -680
rect 10520 -500 10570 -490
rect 10520 -530 10530 -500
rect 10560 -530 10570 -500
rect 10520 -550 10570 -530
rect 10520 -580 10530 -550
rect 10560 -580 10570 -550
rect 10520 -600 10570 -580
rect 10520 -630 10530 -600
rect 10560 -630 10570 -600
rect 10520 -650 10570 -630
rect 10520 -680 10530 -650
rect 10560 -680 10570 -650
rect 10520 -690 10570 -680
rect 10605 -500 10655 -490
rect 10605 -530 10615 -500
rect 10645 -530 10655 -500
rect 10605 -550 10655 -530
rect 10605 -580 10615 -550
rect 10645 -580 10655 -550
rect 10605 -600 10655 -580
rect 10605 -630 10615 -600
rect 10645 -630 10655 -600
rect 10605 -650 10655 -630
rect 10605 -680 10615 -650
rect 10645 -680 10655 -650
rect 10605 -690 10655 -680
rect 10690 -500 10740 -490
rect 10690 -530 10700 -500
rect 10730 -530 10740 -500
rect 10690 -550 10740 -530
rect 10690 -580 10700 -550
rect 10730 -580 10740 -550
rect 10690 -600 10740 -580
rect 10690 -630 10700 -600
rect 10730 -630 10740 -600
rect 10690 -650 10740 -630
rect 10690 -680 10700 -650
rect 10730 -680 10740 -650
rect 10690 -690 10740 -680
rect 10775 -500 10825 -490
rect 10775 -530 10785 -500
rect 10815 -530 10825 -500
rect 10775 -550 10825 -530
rect 10775 -580 10785 -550
rect 10815 -580 10825 -550
rect 10775 -600 10825 -580
rect 10775 -630 10785 -600
rect 10815 -630 10825 -600
rect 10775 -650 10825 -630
rect 10775 -680 10785 -650
rect 10815 -680 10825 -650
rect 10775 -690 10825 -680
rect 10860 -500 10910 -490
rect 10860 -530 10870 -500
rect 10900 -530 10910 -500
rect 10860 -550 10910 -530
rect 10860 -580 10870 -550
rect 10900 -580 10910 -550
rect 10860 -600 10910 -580
rect 10860 -630 10870 -600
rect 10900 -630 10910 -600
rect 10860 -650 10910 -630
rect 10860 -680 10870 -650
rect 10900 -680 10910 -650
rect 10860 -690 10910 -680
rect 10945 -500 10995 -490
rect 10945 -530 10955 -500
rect 10985 -530 10995 -500
rect 10945 -550 10995 -530
rect 10945 -580 10955 -550
rect 10985 -580 10995 -550
rect 10945 -600 10995 -580
rect 10945 -630 10955 -600
rect 10985 -630 10995 -600
rect 10945 -650 10995 -630
rect 10945 -680 10955 -650
rect 10985 -680 10995 -650
rect 10945 -690 10995 -680
rect 11030 -500 11080 -490
rect 11030 -530 11040 -500
rect 11070 -530 11080 -500
rect 11030 -550 11080 -530
rect 11030 -580 11040 -550
rect 11070 -580 11080 -550
rect 11030 -600 11080 -580
rect 11030 -630 11040 -600
rect 11070 -630 11080 -600
rect 11030 -650 11080 -630
rect 11030 -680 11040 -650
rect 11070 -680 11080 -650
rect 11030 -690 11080 -680
rect 11115 -500 11165 -490
rect 11115 -530 11125 -500
rect 11155 -530 11165 -500
rect 11115 -550 11165 -530
rect 11115 -580 11125 -550
rect 11155 -580 11165 -550
rect 11115 -600 11165 -580
rect 11115 -630 11125 -600
rect 11155 -630 11165 -600
rect 11115 -650 11165 -630
rect 11115 -680 11125 -650
rect 11155 -680 11165 -650
rect 11115 -690 11165 -680
rect 11200 -500 11250 -490
rect 11200 -530 11210 -500
rect 11240 -530 11250 -500
rect 11200 -550 11250 -530
rect 11200 -580 11210 -550
rect 11240 -580 11250 -550
rect 11200 -600 11250 -580
rect 11200 -630 11210 -600
rect 11240 -630 11250 -600
rect 11200 -650 11250 -630
rect 11200 -680 11210 -650
rect 11240 -680 11250 -650
rect 11200 -690 11250 -680
rect 11285 -500 11335 -490
rect 11285 -530 11295 -500
rect 11325 -530 11335 -500
rect 11285 -550 11335 -530
rect 11285 -580 11295 -550
rect 11325 -580 11335 -550
rect 11285 -600 11335 -580
rect 11285 -630 11295 -600
rect 11325 -630 11335 -600
rect 11285 -650 11335 -630
rect 11285 -680 11295 -650
rect 11325 -680 11335 -650
rect 11285 -690 11335 -680
rect 11370 -500 11420 -490
rect 11370 -530 11380 -500
rect 11410 -530 11420 -500
rect 11370 -550 11420 -530
rect 11370 -580 11380 -550
rect 11410 -580 11420 -550
rect 11370 -600 11420 -580
rect 11370 -630 11380 -600
rect 11410 -630 11420 -600
rect 11370 -650 11420 -630
rect 11370 -680 11380 -650
rect 11410 -680 11420 -650
rect 11370 -690 11420 -680
rect 11455 -500 11505 -490
rect 11455 -530 11465 -500
rect 11495 -530 11505 -500
rect 11455 -550 11505 -530
rect 11455 -580 11465 -550
rect 11495 -580 11505 -550
rect 11455 -600 11505 -580
rect 11455 -630 11465 -600
rect 11495 -630 11505 -600
rect 11455 -650 11505 -630
rect 11455 -680 11465 -650
rect 11495 -680 11505 -650
rect 11455 -690 11505 -680
rect 11540 -500 11590 -490
rect 11540 -530 11550 -500
rect 11580 -530 11590 -500
rect 11540 -550 11590 -530
rect 11540 -580 11550 -550
rect 11580 -580 11590 -550
rect 11540 -600 11590 -580
rect 11540 -630 11550 -600
rect 11580 -630 11590 -600
rect 11540 -650 11590 -630
rect 11540 -680 11550 -650
rect 11580 -680 11590 -650
rect 11540 -690 11590 -680
rect 11625 -500 11675 -490
rect 11625 -530 11635 -500
rect 11665 -530 11675 -500
rect 11625 -550 11675 -530
rect 11625 -580 11635 -550
rect 11665 -580 11675 -550
rect 11625 -600 11675 -580
rect 11625 -630 11635 -600
rect 11665 -630 11675 -600
rect 11625 -650 11675 -630
rect 11625 -680 11635 -650
rect 11665 -680 11675 -650
rect 11625 -690 11675 -680
rect 11710 -500 11760 -490
rect 11710 -530 11720 -500
rect 11750 -530 11760 -500
rect 11710 -550 11760 -530
rect 11710 -580 11720 -550
rect 11750 -580 11760 -550
rect 11710 -600 11760 -580
rect 11710 -630 11720 -600
rect 11750 -630 11760 -600
rect 11710 -650 11760 -630
rect 11710 -680 11720 -650
rect 11750 -680 11760 -650
rect 11710 -690 11760 -680
rect 11795 -500 11845 -490
rect 11795 -530 11805 -500
rect 11835 -530 11845 -500
rect 11795 -550 11845 -530
rect 11795 -580 11805 -550
rect 11835 -580 11845 -550
rect 11795 -600 11845 -580
rect 11795 -630 11805 -600
rect 11835 -630 11845 -600
rect 11795 -650 11845 -630
rect 11795 -680 11805 -650
rect 11835 -680 11845 -650
rect 11795 -690 11845 -680
rect 11880 -500 11930 -490
rect 11880 -530 11890 -500
rect 11920 -530 11930 -500
rect 11880 -550 11930 -530
rect 11880 -580 11890 -550
rect 11920 -580 11930 -550
rect 11880 -600 11930 -580
rect 11880 -630 11890 -600
rect 11920 -630 11930 -600
rect 11880 -650 11930 -630
rect 11880 -680 11890 -650
rect 11920 -680 11930 -650
rect 11880 -690 11930 -680
rect 11965 -500 12015 -490
rect 11965 -530 11975 -500
rect 12005 -530 12015 -500
rect 11965 -550 12015 -530
rect 11965 -580 11975 -550
rect 12005 -580 12015 -550
rect 11965 -600 12015 -580
rect 11965 -630 11975 -600
rect 12005 -630 12015 -600
rect 11965 -650 12015 -630
rect 11965 -680 11975 -650
rect 12005 -680 12015 -650
rect 11965 -690 12015 -680
rect 12050 -500 12100 -490
rect 12050 -530 12060 -500
rect 12090 -530 12100 -500
rect 12050 -550 12100 -530
rect 12050 -580 12060 -550
rect 12090 -580 12100 -550
rect 12050 -600 12100 -580
rect 12050 -630 12060 -600
rect 12090 -630 12100 -600
rect 12050 -650 12100 -630
rect 12050 -680 12060 -650
rect 12090 -680 12100 -650
rect 12050 -690 12100 -680
rect 12135 -500 12185 -490
rect 12135 -530 12145 -500
rect 12175 -530 12185 -500
rect 12135 -550 12185 -530
rect 12135 -580 12145 -550
rect 12175 -580 12185 -550
rect 12135 -600 12185 -580
rect 12135 -630 12145 -600
rect 12175 -630 12185 -600
rect 12135 -650 12185 -630
rect 12135 -680 12145 -650
rect 12175 -680 12185 -650
rect 12135 -690 12185 -680
rect 12220 -500 12270 -490
rect 12220 -530 12230 -500
rect 12260 -530 12270 -500
rect 12220 -550 12270 -530
rect 12220 -580 12230 -550
rect 12260 -580 12270 -550
rect 12220 -600 12270 -580
rect 12220 -630 12230 -600
rect 12260 -630 12270 -600
rect 12220 -650 12270 -630
rect 12220 -680 12230 -650
rect 12260 -680 12270 -650
rect 12220 -690 12270 -680
rect 12305 -500 12355 -490
rect 12305 -530 12315 -500
rect 12345 -530 12355 -500
rect 12305 -550 12355 -530
rect 12305 -580 12315 -550
rect 12345 -580 12355 -550
rect 12305 -600 12355 -580
rect 12305 -630 12315 -600
rect 12345 -630 12355 -600
rect 12305 -650 12355 -630
rect 12305 -680 12315 -650
rect 12345 -680 12355 -650
rect 12305 -690 12355 -680
rect 12390 -500 12440 -490
rect 12390 -530 12400 -500
rect 12430 -530 12440 -500
rect 12390 -550 12440 -530
rect 12390 -580 12400 -550
rect 12430 -580 12440 -550
rect 12390 -600 12440 -580
rect 12390 -630 12400 -600
rect 12430 -630 12440 -600
rect 12390 -650 12440 -630
rect 12390 -680 12400 -650
rect 12430 -680 12440 -650
rect 12390 -690 12440 -680
rect 12475 -500 12525 -490
rect 12475 -530 12485 -500
rect 12515 -530 12525 -500
rect 12475 -550 12525 -530
rect 12475 -580 12485 -550
rect 12515 -580 12525 -550
rect 12475 -600 12525 -580
rect 12475 -630 12485 -600
rect 12515 -630 12525 -600
rect 12475 -650 12525 -630
rect 12475 -680 12485 -650
rect 12515 -680 12525 -650
rect 12475 -690 12525 -680
rect 12560 -500 12610 -490
rect 12560 -530 12570 -500
rect 12600 -530 12610 -500
rect 12560 -550 12610 -530
rect 12560 -580 12570 -550
rect 12600 -580 12610 -550
rect 12560 -600 12610 -580
rect 12560 -630 12570 -600
rect 12600 -630 12610 -600
rect 12560 -650 12610 -630
rect 12560 -680 12570 -650
rect 12600 -680 12610 -650
rect 12560 -690 12610 -680
rect 12645 -500 12695 -490
rect 12645 -530 12655 -500
rect 12685 -530 12695 -500
rect 12645 -550 12695 -530
rect 12645 -580 12655 -550
rect 12685 -580 12695 -550
rect 12645 -600 12695 -580
rect 12645 -630 12655 -600
rect 12685 -630 12695 -600
rect 12645 -650 12695 -630
rect 12645 -680 12655 -650
rect 12685 -680 12695 -650
rect 12645 -690 12695 -680
rect 12730 -500 12780 -490
rect 12730 -530 12740 -500
rect 12770 -530 12780 -500
rect 12730 -550 12780 -530
rect 12730 -580 12740 -550
rect 12770 -580 12780 -550
rect 12730 -600 12780 -580
rect 12730 -630 12740 -600
rect 12770 -630 12780 -600
rect 12730 -650 12780 -630
rect 12730 -680 12740 -650
rect 12770 -680 12780 -650
rect 12730 -690 12780 -680
rect 12815 -500 12865 -490
rect 12815 -530 12825 -500
rect 12855 -530 12865 -500
rect 12815 -550 12865 -530
rect 12815 -580 12825 -550
rect 12855 -580 12865 -550
rect 12815 -600 12865 -580
rect 12815 -630 12825 -600
rect 12855 -630 12865 -600
rect 12815 -650 12865 -630
rect 12815 -680 12825 -650
rect 12855 -680 12865 -650
rect 12815 -690 12865 -680
rect 12900 -500 12950 -490
rect 12900 -530 12910 -500
rect 12940 -530 12950 -500
rect 12900 -550 12950 -530
rect 12900 -580 12910 -550
rect 12940 -580 12950 -550
rect 12900 -600 12950 -580
rect 12900 -630 12910 -600
rect 12940 -630 12950 -600
rect 12900 -650 12950 -630
rect 12900 -680 12910 -650
rect 12940 -680 12950 -650
rect 12900 -690 12950 -680
rect 12985 -500 13035 -490
rect 12985 -530 12995 -500
rect 13025 -530 13035 -500
rect 12985 -550 13035 -530
rect 12985 -580 12995 -550
rect 13025 -580 13035 -550
rect 12985 -600 13035 -580
rect 12985 -630 12995 -600
rect 13025 -630 13035 -600
rect 12985 -650 13035 -630
rect 12985 -680 12995 -650
rect 13025 -680 13035 -650
rect 12985 -690 13035 -680
rect 13070 -500 13120 -490
rect 13070 -530 13080 -500
rect 13110 -530 13120 -500
rect 13070 -550 13120 -530
rect 13070 -580 13080 -550
rect 13110 -580 13120 -550
rect 13070 -600 13120 -580
rect 13070 -630 13080 -600
rect 13110 -630 13120 -600
rect 13070 -650 13120 -630
rect 13070 -680 13080 -650
rect 13110 -680 13120 -650
rect 13070 -690 13120 -680
rect 13155 -500 13205 -490
rect 13155 -530 13165 -500
rect 13195 -530 13205 -500
rect 13155 -550 13205 -530
rect 13155 -580 13165 -550
rect 13195 -580 13205 -550
rect 13155 -600 13205 -580
rect 13155 -630 13165 -600
rect 13195 -630 13205 -600
rect 13155 -650 13205 -630
rect 13155 -680 13165 -650
rect 13195 -680 13205 -650
rect 13155 -690 13205 -680
rect 13240 -500 13290 -490
rect 13240 -530 13250 -500
rect 13280 -530 13290 -500
rect 13240 -550 13290 -530
rect 13240 -580 13250 -550
rect 13280 -580 13290 -550
rect 13240 -600 13290 -580
rect 13240 -630 13250 -600
rect 13280 -630 13290 -600
rect 13240 -650 13290 -630
rect 13240 -680 13250 -650
rect 13280 -680 13290 -650
rect 13240 -690 13290 -680
rect 13325 -500 13375 -490
rect 13325 -530 13335 -500
rect 13365 -530 13375 -500
rect 13325 -550 13375 -530
rect 13325 -580 13335 -550
rect 13365 -580 13375 -550
rect 13325 -600 13375 -580
rect 13325 -630 13335 -600
rect 13365 -630 13375 -600
rect 13325 -650 13375 -630
rect 13325 -680 13335 -650
rect 13365 -680 13375 -650
rect 13325 -690 13375 -680
rect 13410 -500 13460 -490
rect 13410 -530 13420 -500
rect 13450 -530 13460 -500
rect 13410 -550 13460 -530
rect 13410 -580 13420 -550
rect 13450 -580 13460 -550
rect 13410 -600 13460 -580
rect 13410 -630 13420 -600
rect 13450 -630 13460 -600
rect 13410 -650 13460 -630
rect 13410 -680 13420 -650
rect 13450 -680 13460 -650
rect 13410 -690 13460 -680
rect 13495 -500 13545 -490
rect 13495 -530 13505 -500
rect 13535 -530 13545 -500
rect 13495 -550 13545 -530
rect 13495 -580 13505 -550
rect 13535 -580 13545 -550
rect 13495 -600 13545 -580
rect 13495 -630 13505 -600
rect 13535 -630 13545 -600
rect 13495 -650 13545 -630
rect 13495 -680 13505 -650
rect 13535 -680 13545 -650
rect 13495 -690 13545 -680
rect 13580 -500 13630 -490
rect 13580 -530 13590 -500
rect 13620 -530 13630 -500
rect 13580 -550 13630 -530
rect 13580 -580 13590 -550
rect 13620 -580 13630 -550
rect 13580 -600 13630 -580
rect 13580 -630 13590 -600
rect 13620 -630 13630 -600
rect 13580 -650 13630 -630
rect 13580 -680 13590 -650
rect 13620 -680 13630 -650
rect 13580 -690 13630 -680
rect 13665 -500 13715 -490
rect 13665 -530 13675 -500
rect 13705 -530 13715 -500
rect 13665 -550 13715 -530
rect 13665 -580 13675 -550
rect 13705 -580 13715 -550
rect 13665 -600 13715 -580
rect 13665 -630 13675 -600
rect 13705 -630 13715 -600
rect 13665 -650 13715 -630
rect 13665 -680 13675 -650
rect 13705 -680 13715 -650
rect 13665 -690 13715 -680
rect 13750 -500 13800 -490
rect 13750 -530 13760 -500
rect 13790 -530 13800 -500
rect 13750 -550 13800 -530
rect 13750 -580 13760 -550
rect 13790 -580 13800 -550
rect 13750 -600 13800 -580
rect 13750 -630 13760 -600
rect 13790 -630 13800 -600
rect 13750 -650 13800 -630
rect 13750 -680 13760 -650
rect 13790 -680 13800 -650
rect 13750 -690 13800 -680
rect 13835 -500 13885 -490
rect 13835 -530 13845 -500
rect 13875 -530 13885 -500
rect 13835 -550 13885 -530
rect 13835 -580 13845 -550
rect 13875 -580 13885 -550
rect 13835 -600 13885 -580
rect 13835 -630 13845 -600
rect 13875 -630 13885 -600
rect 13835 -650 13885 -630
rect 13835 -680 13845 -650
rect 13875 -680 13885 -650
rect 13835 -690 13885 -680
rect 13920 -500 13970 -490
rect 13920 -530 13930 -500
rect 13960 -530 13970 -500
rect 13920 -550 13970 -530
rect 13920 -580 13930 -550
rect 13960 -580 13970 -550
rect 13920 -600 13970 -580
rect 13920 -630 13930 -600
rect 13960 -630 13970 -600
rect 13920 -650 13970 -630
rect 13920 -680 13930 -650
rect 13960 -680 13970 -650
rect 13920 -690 13970 -680
rect 14005 -500 14055 -490
rect 14005 -530 14015 -500
rect 14045 -530 14055 -500
rect 14005 -550 14055 -530
rect 14005 -580 14015 -550
rect 14045 -580 14055 -550
rect 14005 -600 14055 -580
rect 14005 -630 14015 -600
rect 14045 -630 14055 -600
rect 14005 -650 14055 -630
rect 14005 -680 14015 -650
rect 14045 -680 14055 -650
rect 14005 -690 14055 -680
rect 14090 -500 14140 -490
rect 14090 -530 14100 -500
rect 14130 -530 14140 -500
rect 14090 -550 14140 -530
rect 14090 -580 14100 -550
rect 14130 -580 14140 -550
rect 14090 -600 14140 -580
rect 14090 -630 14100 -600
rect 14130 -630 14140 -600
rect 14090 -650 14140 -630
rect 14090 -680 14100 -650
rect 14130 -680 14140 -650
rect 14090 -690 14140 -680
rect 14175 -500 14225 -490
rect 14175 -530 14185 -500
rect 14215 -530 14225 -500
rect 14175 -550 14225 -530
rect 14175 -580 14185 -550
rect 14215 -580 14225 -550
rect 14175 -600 14225 -580
rect 14175 -630 14185 -600
rect 14215 -630 14225 -600
rect 14175 -650 14225 -630
rect 14175 -680 14185 -650
rect 14215 -680 14225 -650
rect 14175 -690 14225 -680
rect 14260 -500 14310 -490
rect 14260 -530 14270 -500
rect 14300 -530 14310 -500
rect 14260 -550 14310 -530
rect 14260 -580 14270 -550
rect 14300 -580 14310 -550
rect 14260 -600 14310 -580
rect 14260 -630 14270 -600
rect 14300 -630 14310 -600
rect 14260 -650 14310 -630
rect 14260 -680 14270 -650
rect 14300 -680 14310 -650
rect 14260 -690 14310 -680
rect 14345 -500 14395 -490
rect 14345 -530 14355 -500
rect 14385 -530 14395 -500
rect 14345 -550 14395 -530
rect 14345 -580 14355 -550
rect 14385 -580 14395 -550
rect 14345 -600 14395 -580
rect 14345 -630 14355 -600
rect 14385 -630 14395 -600
rect 14345 -650 14395 -630
rect 14345 -680 14355 -650
rect 14385 -680 14395 -650
rect 14345 -690 14395 -680
rect 14430 -500 14480 -490
rect 14430 -530 14440 -500
rect 14470 -530 14480 -500
rect 14430 -550 14480 -530
rect 14430 -580 14440 -550
rect 14470 -580 14480 -550
rect 14430 -600 14480 -580
rect 14430 -630 14440 -600
rect 14470 -630 14480 -600
rect 14430 -650 14480 -630
rect 14430 -680 14440 -650
rect 14470 -680 14480 -650
rect 14430 -690 14480 -680
rect 14515 -500 14565 -490
rect 14515 -530 14525 -500
rect 14555 -530 14565 -500
rect 14515 -550 14565 -530
rect 14515 -580 14525 -550
rect 14555 -580 14565 -550
rect 14515 -600 14565 -580
rect 14515 -630 14525 -600
rect 14555 -630 14565 -600
rect 14515 -650 14565 -630
rect 14515 -680 14525 -650
rect 14555 -680 14565 -650
rect 14515 -690 14565 -680
rect 14600 -500 14650 -490
rect 14600 -530 14610 -500
rect 14640 -530 14650 -500
rect 14600 -550 14650 -530
rect 14600 -580 14610 -550
rect 14640 -580 14650 -550
rect 14600 -600 14650 -580
rect 14600 -630 14610 -600
rect 14640 -630 14650 -600
rect 14600 -650 14650 -630
rect 14600 -680 14610 -650
rect 14640 -680 14650 -650
rect 14600 -690 14650 -680
rect 14685 -500 14735 -490
rect 14685 -530 14695 -500
rect 14725 -530 14735 -500
rect 14685 -550 14735 -530
rect 14685 -580 14695 -550
rect 14725 -580 14735 -550
rect 14685 -600 14735 -580
rect 14685 -630 14695 -600
rect 14725 -630 14735 -600
rect 14685 -650 14735 -630
rect 14685 -680 14695 -650
rect 14725 -680 14735 -650
rect 14685 -690 14735 -680
rect 14770 -500 14820 -490
rect 14770 -530 14780 -500
rect 14810 -530 14820 -500
rect 14770 -550 14820 -530
rect 14770 -580 14780 -550
rect 14810 -580 14820 -550
rect 14770 -600 14820 -580
rect 14770 -630 14780 -600
rect 14810 -630 14820 -600
rect 14770 -650 14820 -630
rect 14770 -680 14780 -650
rect 14810 -680 14820 -650
rect 14770 -690 14820 -680
rect 14855 -500 14905 -490
rect 14855 -530 14865 -500
rect 14895 -530 14905 -500
rect 14855 -550 14905 -530
rect 14855 -580 14865 -550
rect 14895 -580 14905 -550
rect 14855 -600 14905 -580
rect 14855 -630 14865 -600
rect 14895 -630 14905 -600
rect 14855 -650 14905 -630
rect 14855 -680 14865 -650
rect 14895 -680 14905 -650
rect 14855 -690 14905 -680
rect 14940 -500 14990 -490
rect 14940 -530 14950 -500
rect 14980 -530 14990 -500
rect 14940 -550 14990 -530
rect 14940 -580 14950 -550
rect 14980 -580 14990 -550
rect 14940 -600 14990 -580
rect 14940 -630 14950 -600
rect 14980 -630 14990 -600
rect 14940 -650 14990 -630
rect 14940 -680 14950 -650
rect 14980 -680 14990 -650
rect 14940 -690 14990 -680
rect 15025 -500 15075 -490
rect 15025 -530 15035 -500
rect 15065 -530 15075 -500
rect 15025 -550 15075 -530
rect 15025 -580 15035 -550
rect 15065 -580 15075 -550
rect 15025 -600 15075 -580
rect 15025 -630 15035 -600
rect 15065 -630 15075 -600
rect 15025 -650 15075 -630
rect 15025 -680 15035 -650
rect 15065 -680 15075 -650
rect 15025 -690 15075 -680
rect 15110 -500 15160 -490
rect 15110 -530 15120 -500
rect 15150 -530 15160 -500
rect 15110 -550 15160 -530
rect 15110 -580 15120 -550
rect 15150 -580 15160 -550
rect 15110 -600 15160 -580
rect 15110 -630 15120 -600
rect 15150 -630 15160 -600
rect 15110 -650 15160 -630
rect 15110 -680 15120 -650
rect 15150 -680 15160 -650
rect 15110 -690 15160 -680
rect 15195 -500 15245 -490
rect 15195 -530 15205 -500
rect 15235 -530 15245 -500
rect 15195 -550 15245 -530
rect 15195 -580 15205 -550
rect 15235 -580 15245 -550
rect 15195 -600 15245 -580
rect 15195 -630 15205 -600
rect 15235 -630 15245 -600
rect 15195 -650 15245 -630
rect 15195 -680 15205 -650
rect 15235 -680 15245 -650
rect 15195 -690 15245 -680
rect 15280 -500 15330 -490
rect 15280 -530 15290 -500
rect 15320 -530 15330 -500
rect 15280 -550 15330 -530
rect 15280 -580 15290 -550
rect 15320 -580 15330 -550
rect 15280 -600 15330 -580
rect 15280 -630 15290 -600
rect 15320 -630 15330 -600
rect 15280 -650 15330 -630
rect 15280 -680 15290 -650
rect 15320 -680 15330 -650
rect 15280 -690 15330 -680
rect 15365 -500 15415 -490
rect 15365 -530 15375 -500
rect 15405 -530 15415 -500
rect 15365 -550 15415 -530
rect 15365 -580 15375 -550
rect 15405 -580 15415 -550
rect 15365 -600 15415 -580
rect 15365 -630 15375 -600
rect 15405 -630 15415 -600
rect 15365 -650 15415 -630
rect 15365 -680 15375 -650
rect 15405 -680 15415 -650
rect 15365 -690 15415 -680
rect 15450 -500 15500 -490
rect 15450 -530 15460 -500
rect 15490 -530 15500 -500
rect 15450 -550 15500 -530
rect 15450 -580 15460 -550
rect 15490 -580 15500 -550
rect 15450 -600 15500 -580
rect 15450 -630 15460 -600
rect 15490 -630 15500 -600
rect 15450 -650 15500 -630
rect 15450 -680 15460 -650
rect 15490 -680 15500 -650
rect 15450 -690 15500 -680
rect 15535 -500 15585 -490
rect 15535 -530 15545 -500
rect 15575 -530 15585 -500
rect 15535 -550 15585 -530
rect 15535 -580 15545 -550
rect 15575 -580 15585 -550
rect 15535 -600 15585 -580
rect 15535 -630 15545 -600
rect 15575 -630 15585 -600
rect 15535 -650 15585 -630
rect 15535 -680 15545 -650
rect 15575 -680 15585 -650
rect 15535 -690 15585 -680
rect 15620 -500 15670 -490
rect 15620 -530 15630 -500
rect 15660 -530 15670 -500
rect 15620 -550 15670 -530
rect 15620 -580 15630 -550
rect 15660 -580 15670 -550
rect 15620 -600 15670 -580
rect 15620 -630 15630 -600
rect 15660 -630 15670 -600
rect 15620 -650 15670 -630
rect 15620 -680 15630 -650
rect 15660 -680 15670 -650
rect 15620 -690 15670 -680
rect 15705 -500 15755 -490
rect 15705 -530 15715 -500
rect 15745 -530 15755 -500
rect 15705 -550 15755 -530
rect 15705 -580 15715 -550
rect 15745 -580 15755 -550
rect 15705 -600 15755 -580
rect 15705 -630 15715 -600
rect 15745 -630 15755 -600
rect 15705 -650 15755 -630
rect 15705 -680 15715 -650
rect 15745 -680 15755 -650
rect 15705 -690 15755 -680
rect 15790 -500 15840 -490
rect 15790 -530 15800 -500
rect 15830 -530 15840 -500
rect 15790 -550 15840 -530
rect 15790 -580 15800 -550
rect 15830 -580 15840 -550
rect 15790 -600 15840 -580
rect 15790 -630 15800 -600
rect 15830 -630 15840 -600
rect 15790 -650 15840 -630
rect 15790 -680 15800 -650
rect 15830 -680 15840 -650
rect 15790 -690 15840 -680
rect 15875 -500 15925 -490
rect 15875 -530 15885 -500
rect 15915 -530 15925 -500
rect 15875 -550 15925 -530
rect 15875 -580 15885 -550
rect 15915 -580 15925 -550
rect 15875 -600 15925 -580
rect 15875 -630 15885 -600
rect 15915 -630 15925 -600
rect 15875 -650 15925 -630
rect 15875 -680 15885 -650
rect 15915 -680 15925 -650
rect 15875 -690 15925 -680
rect 15960 -500 16010 -490
rect 15960 -530 15970 -500
rect 16000 -530 16010 -500
rect 15960 -550 16010 -530
rect 15960 -580 15970 -550
rect 16000 -580 16010 -550
rect 15960 -600 16010 -580
rect 15960 -630 15970 -600
rect 16000 -630 16010 -600
rect 15960 -650 16010 -630
rect 15960 -680 15970 -650
rect 16000 -680 16010 -650
rect 15960 -690 16010 -680
rect 16045 -500 16095 -490
rect 16045 -530 16055 -500
rect 16085 -530 16095 -500
rect 16045 -550 16095 -530
rect 16045 -580 16055 -550
rect 16085 -580 16095 -550
rect 16045 -600 16095 -580
rect 16045 -630 16055 -600
rect 16085 -630 16095 -600
rect 16045 -650 16095 -630
rect 16045 -680 16055 -650
rect 16085 -680 16095 -650
rect 16045 -690 16095 -680
rect 16130 -500 16180 -490
rect 16130 -530 16140 -500
rect 16170 -530 16180 -500
rect 16130 -550 16180 -530
rect 16130 -580 16140 -550
rect 16170 -580 16180 -550
rect 16130 -600 16180 -580
rect 16130 -630 16140 -600
rect 16170 -630 16180 -600
rect 16130 -650 16180 -630
rect 16130 -680 16140 -650
rect 16170 -680 16180 -650
rect 16130 -690 16180 -680
rect 16215 -500 16265 -490
rect 16215 -530 16225 -500
rect 16255 -530 16265 -500
rect 16215 -550 16265 -530
rect 16215 -580 16225 -550
rect 16255 -580 16265 -550
rect 16215 -600 16265 -580
rect 16215 -630 16225 -600
rect 16255 -630 16265 -600
rect 16215 -650 16265 -630
rect 16215 -680 16225 -650
rect 16255 -680 16265 -650
rect 16215 -690 16265 -680
rect 16300 -500 16350 -490
rect 16300 -530 16310 -500
rect 16340 -530 16350 -500
rect 16300 -550 16350 -530
rect 16300 -580 16310 -550
rect 16340 -580 16350 -550
rect 16300 -600 16350 -580
rect 16300 -630 16310 -600
rect 16340 -630 16350 -600
rect 16300 -650 16350 -630
rect 16300 -680 16310 -650
rect 16340 -680 16350 -650
rect 16300 -690 16350 -680
rect 16385 -500 16435 -490
rect 16385 -530 16395 -500
rect 16425 -530 16435 -500
rect 16385 -550 16435 -530
rect 16385 -580 16395 -550
rect 16425 -580 16435 -550
rect 16385 -600 16435 -580
rect 16385 -630 16395 -600
rect 16425 -630 16435 -600
rect 16385 -650 16435 -630
rect 16385 -680 16395 -650
rect 16425 -680 16435 -650
rect 16385 -690 16435 -680
rect 16470 -500 16520 -490
rect 16470 -530 16480 -500
rect 16510 -530 16520 -500
rect 16470 -550 16520 -530
rect 16470 -580 16480 -550
rect 16510 -580 16520 -550
rect 16470 -600 16520 -580
rect 16470 -630 16480 -600
rect 16510 -630 16520 -600
rect 16470 -650 16520 -630
rect 16470 -680 16480 -650
rect 16510 -680 16520 -650
rect 16470 -690 16520 -680
rect 16555 -500 16605 -490
rect 16555 -530 16565 -500
rect 16595 -530 16605 -500
rect 16555 -550 16605 -530
rect 16555 -580 16565 -550
rect 16595 -580 16605 -550
rect 16555 -600 16605 -580
rect 16555 -630 16565 -600
rect 16595 -630 16605 -600
rect 16555 -650 16605 -630
rect 16555 -680 16565 -650
rect 16595 -680 16605 -650
rect 16555 -690 16605 -680
rect 16640 -500 16690 -490
rect 16640 -530 16650 -500
rect 16680 -530 16690 -500
rect 16640 -550 16690 -530
rect 16640 -580 16650 -550
rect 16680 -580 16690 -550
rect 16640 -600 16690 -580
rect 16640 -630 16650 -600
rect 16680 -630 16690 -600
rect 16640 -650 16690 -630
rect 16640 -680 16650 -650
rect 16680 -680 16690 -650
rect 16640 -690 16690 -680
rect 16725 -500 16775 -490
rect 16725 -530 16735 -500
rect 16765 -530 16775 -500
rect 16725 -550 16775 -530
rect 16725 -580 16735 -550
rect 16765 -580 16775 -550
rect 16725 -600 16775 -580
rect 16725 -630 16735 -600
rect 16765 -630 16775 -600
rect 16725 -650 16775 -630
rect 16725 -680 16735 -650
rect 16765 -680 16775 -650
rect 16725 -690 16775 -680
rect 16810 -500 16860 -490
rect 16810 -530 16820 -500
rect 16850 -530 16860 -500
rect 16810 -550 16860 -530
rect 16810 -580 16820 -550
rect 16850 -580 16860 -550
rect 16810 -600 16860 -580
rect 16810 -630 16820 -600
rect 16850 -630 16860 -600
rect 16810 -650 16860 -630
rect 16810 -680 16820 -650
rect 16850 -680 16860 -650
rect 16810 -690 16860 -680
rect 16895 -500 16945 -490
rect 16895 -530 16905 -500
rect 16935 -530 16945 -500
rect 16895 -550 16945 -530
rect 16895 -580 16905 -550
rect 16935 -580 16945 -550
rect 16895 -600 16945 -580
rect 16895 -630 16905 -600
rect 16935 -630 16945 -600
rect 16895 -650 16945 -630
rect 16895 -680 16905 -650
rect 16935 -680 16945 -650
rect 16895 -690 16945 -680
rect 16980 -500 17030 -490
rect 16980 -530 16990 -500
rect 17020 -530 17030 -500
rect 16980 -550 17030 -530
rect 16980 -580 16990 -550
rect 17020 -580 17030 -550
rect 16980 -600 17030 -580
rect 16980 -630 16990 -600
rect 17020 -630 17030 -600
rect 16980 -650 17030 -630
rect 16980 -680 16990 -650
rect 17020 -680 17030 -650
rect 16980 -690 17030 -680
rect 17065 -500 17115 -490
rect 17065 -530 17075 -500
rect 17105 -530 17115 -500
rect 17065 -550 17115 -530
rect 17065 -580 17075 -550
rect 17105 -580 17115 -550
rect 17065 -600 17115 -580
rect 17065 -630 17075 -600
rect 17105 -630 17115 -600
rect 17065 -650 17115 -630
rect 17065 -680 17075 -650
rect 17105 -680 17115 -650
rect 17065 -690 17115 -680
rect 17150 -500 17200 -490
rect 17150 -530 17160 -500
rect 17190 -530 17200 -500
rect 17150 -550 17200 -530
rect 17150 -580 17160 -550
rect 17190 -580 17200 -550
rect 17150 -600 17200 -580
rect 17150 -630 17160 -600
rect 17190 -630 17200 -600
rect 17150 -650 17200 -630
rect 17150 -680 17160 -650
rect 17190 -680 17200 -650
rect 17150 -690 17200 -680
rect 17235 -500 17285 -490
rect 17235 -530 17245 -500
rect 17275 -530 17285 -500
rect 17235 -550 17285 -530
rect 17235 -580 17245 -550
rect 17275 -580 17285 -550
rect 17235 -600 17285 -580
rect 17235 -630 17245 -600
rect 17275 -630 17285 -600
rect 17235 -650 17285 -630
rect 17235 -680 17245 -650
rect 17275 -680 17285 -650
rect 17235 -690 17285 -680
rect 17320 -500 17370 -490
rect 17320 -530 17330 -500
rect 17360 -530 17370 -500
rect 17320 -550 17370 -530
rect 17320 -580 17330 -550
rect 17360 -580 17370 -550
rect 17320 -600 17370 -580
rect 17320 -630 17330 -600
rect 17360 -630 17370 -600
rect 17320 -650 17370 -630
rect 17320 -680 17330 -650
rect 17360 -680 17370 -650
rect 17320 -690 17370 -680
rect 17405 -500 17455 -490
rect 17405 -530 17415 -500
rect 17445 -530 17455 -500
rect 17405 -550 17455 -530
rect 17405 -580 17415 -550
rect 17445 -580 17455 -550
rect 17405 -600 17455 -580
rect 17405 -630 17415 -600
rect 17445 -630 17455 -600
rect 17405 -650 17455 -630
rect 17405 -680 17415 -650
rect 17445 -680 17455 -650
rect 17405 -690 17455 -680
rect 17490 -500 17540 -490
rect 17490 -530 17500 -500
rect 17530 -530 17540 -500
rect 17490 -550 17540 -530
rect 17490 -580 17500 -550
rect 17530 -580 17540 -550
rect 17490 -600 17540 -580
rect 17490 -630 17500 -600
rect 17530 -630 17540 -600
rect 17490 -650 17540 -630
rect 17490 -680 17500 -650
rect 17530 -680 17540 -650
rect 17490 -690 17540 -680
rect 17575 -500 17625 -490
rect 17575 -530 17585 -500
rect 17615 -530 17625 -500
rect 17575 -550 17625 -530
rect 17575 -580 17585 -550
rect 17615 -580 17625 -550
rect 17575 -600 17625 -580
rect 17575 -630 17585 -600
rect 17615 -630 17625 -600
rect 17575 -650 17625 -630
rect 17575 -680 17585 -650
rect 17615 -680 17625 -650
rect 17575 -690 17625 -680
rect 17660 -500 17710 -490
rect 17660 -530 17670 -500
rect 17700 -530 17710 -500
rect 17660 -550 17710 -530
rect 17660 -580 17670 -550
rect 17700 -580 17710 -550
rect 17660 -600 17710 -580
rect 17660 -630 17670 -600
rect 17700 -630 17710 -600
rect 17660 -650 17710 -630
rect 17660 -680 17670 -650
rect 17700 -680 17710 -650
rect 17660 -690 17710 -680
rect 17745 -500 17795 -490
rect 17745 -530 17755 -500
rect 17785 -530 17795 -500
rect 17745 -550 17795 -530
rect 17745 -580 17755 -550
rect 17785 -580 17795 -550
rect 17745 -600 17795 -580
rect 17745 -630 17755 -600
rect 17785 -630 17795 -600
rect 17745 -650 17795 -630
rect 17745 -680 17755 -650
rect 17785 -680 17795 -650
rect 17745 -690 17795 -680
rect 17830 -500 17880 -490
rect 17830 -530 17840 -500
rect 17870 -530 17880 -500
rect 17830 -550 17880 -530
rect 17830 -580 17840 -550
rect 17870 -580 17880 -550
rect 17830 -600 17880 -580
rect 17830 -630 17840 -600
rect 17870 -630 17880 -600
rect 17830 -650 17880 -630
rect 17830 -680 17840 -650
rect 17870 -680 17880 -650
rect 17830 -690 17880 -680
rect 17915 -500 17965 -490
rect 17915 -530 17925 -500
rect 17955 -530 17965 -500
rect 17915 -550 17965 -530
rect 17915 -580 17925 -550
rect 17955 -580 17965 -550
rect 17915 -600 17965 -580
rect 17915 -630 17925 -600
rect 17955 -630 17965 -600
rect 17915 -650 17965 -630
rect 17915 -680 17925 -650
rect 17955 -680 17965 -650
rect 17915 -690 17965 -680
rect 18000 -500 18050 -490
rect 18000 -530 18010 -500
rect 18040 -530 18050 -500
rect 18000 -550 18050 -530
rect 18000 -580 18010 -550
rect 18040 -580 18050 -550
rect 18000 -600 18050 -580
rect 18000 -630 18010 -600
rect 18040 -630 18050 -600
rect 18000 -650 18050 -630
rect 18000 -680 18010 -650
rect 18040 -680 18050 -650
rect 18000 -690 18050 -680
rect 18085 -500 18135 -490
rect 18085 -530 18095 -500
rect 18125 -530 18135 -500
rect 18085 -550 18135 -530
rect 18085 -580 18095 -550
rect 18125 -580 18135 -550
rect 18085 -600 18135 -580
rect 18085 -630 18095 -600
rect 18125 -630 18135 -600
rect 18085 -650 18135 -630
rect 18085 -680 18095 -650
rect 18125 -680 18135 -650
rect 18085 -690 18135 -680
rect 18170 -500 18220 -490
rect 18170 -530 18180 -500
rect 18210 -530 18220 -500
rect 18170 -550 18220 -530
rect 18170 -580 18180 -550
rect 18210 -580 18220 -550
rect 18170 -600 18220 -580
rect 18170 -630 18180 -600
rect 18210 -630 18220 -600
rect 18170 -650 18220 -630
rect 18170 -680 18180 -650
rect 18210 -680 18220 -650
rect 18170 -690 18220 -680
rect 18255 -500 18305 -490
rect 18255 -530 18265 -500
rect 18295 -530 18305 -500
rect 18255 -550 18305 -530
rect 18255 -580 18265 -550
rect 18295 -580 18305 -550
rect 18255 -600 18305 -580
rect 18255 -630 18265 -600
rect 18295 -630 18305 -600
rect 18255 -650 18305 -630
rect 18255 -680 18265 -650
rect 18295 -680 18305 -650
rect 18255 -690 18305 -680
rect 18340 -500 18390 -490
rect 18340 -530 18350 -500
rect 18380 -530 18390 -500
rect 18340 -550 18390 -530
rect 18340 -580 18350 -550
rect 18380 -580 18390 -550
rect 18340 -600 18390 -580
rect 18340 -630 18350 -600
rect 18380 -630 18390 -600
rect 18340 -650 18390 -630
rect 18340 -680 18350 -650
rect 18380 -680 18390 -650
rect 18340 -690 18390 -680
rect 18425 -500 18475 -490
rect 18425 -530 18435 -500
rect 18465 -530 18475 -500
rect 18425 -550 18475 -530
rect 18425 -580 18435 -550
rect 18465 -580 18475 -550
rect 18425 -600 18475 -580
rect 18425 -630 18435 -600
rect 18465 -630 18475 -600
rect 18425 -650 18475 -630
rect 18425 -680 18435 -650
rect 18465 -680 18475 -650
rect 18425 -690 18475 -680
rect 18510 -500 18560 -490
rect 18510 -530 18520 -500
rect 18550 -530 18560 -500
rect 18510 -550 18560 -530
rect 18510 -580 18520 -550
rect 18550 -580 18560 -550
rect 18510 -600 18560 -580
rect 18510 -630 18520 -600
rect 18550 -630 18560 -600
rect 18510 -650 18560 -630
rect 18510 -680 18520 -650
rect 18550 -680 18560 -650
rect 18510 -690 18560 -680
rect 18595 -500 18645 -490
rect 18595 -530 18605 -500
rect 18635 -530 18645 -500
rect 18595 -550 18645 -530
rect 18595 -580 18605 -550
rect 18635 -580 18645 -550
rect 18595 -600 18645 -580
rect 18595 -630 18605 -600
rect 18635 -630 18645 -600
rect 18595 -650 18645 -630
rect 18595 -680 18605 -650
rect 18635 -680 18645 -650
rect 18595 -690 18645 -680
rect 18680 -500 18730 -490
rect 18680 -530 18690 -500
rect 18720 -530 18730 -500
rect 18680 -550 18730 -530
rect 18680 -580 18690 -550
rect 18720 -580 18730 -550
rect 18680 -600 18730 -580
rect 18680 -630 18690 -600
rect 18720 -630 18730 -600
rect 18680 -650 18730 -630
rect 18680 -680 18690 -650
rect 18720 -680 18730 -650
rect 18680 -690 18730 -680
rect 18765 -500 18815 -490
rect 18765 -530 18775 -500
rect 18805 -530 18815 -500
rect 18765 -550 18815 -530
rect 18765 -580 18775 -550
rect 18805 -580 18815 -550
rect 18765 -600 18815 -580
rect 18765 -630 18775 -600
rect 18805 -630 18815 -600
rect 18765 -650 18815 -630
rect 18765 -680 18775 -650
rect 18805 -680 18815 -650
rect 18765 -690 18815 -680
rect 18850 -500 18900 -490
rect 18850 -530 18860 -500
rect 18890 -530 18900 -500
rect 18850 -550 18900 -530
rect 18850 -580 18860 -550
rect 18890 -580 18900 -550
rect 18850 -600 18900 -580
rect 18850 -630 18860 -600
rect 18890 -630 18900 -600
rect 18850 -650 18900 -630
rect 18850 -680 18860 -650
rect 18890 -680 18900 -650
rect 18850 -690 18900 -680
rect 18935 -500 18985 -490
rect 18935 -530 18945 -500
rect 18975 -530 18985 -500
rect 18935 -550 18985 -530
rect 18935 -580 18945 -550
rect 18975 -580 18985 -550
rect 18935 -600 18985 -580
rect 18935 -630 18945 -600
rect 18975 -630 18985 -600
rect 18935 -650 18985 -630
rect 18935 -680 18945 -650
rect 18975 -680 18985 -650
rect 18935 -690 18985 -680
rect 19020 -500 19070 -490
rect 19020 -530 19030 -500
rect 19060 -530 19070 -500
rect 19020 -550 19070 -530
rect 19020 -580 19030 -550
rect 19060 -580 19070 -550
rect 19020 -600 19070 -580
rect 19020 -630 19030 -600
rect 19060 -630 19070 -600
rect 19020 -650 19070 -630
rect 19020 -680 19030 -650
rect 19060 -680 19070 -650
rect 19020 -690 19070 -680
rect 19105 -500 19155 -490
rect 19105 -530 19115 -500
rect 19145 -530 19155 -500
rect 19105 -550 19155 -530
rect 19105 -580 19115 -550
rect 19145 -580 19155 -550
rect 19105 -600 19155 -580
rect 19105 -630 19115 -600
rect 19145 -630 19155 -600
rect 19105 -650 19155 -630
rect 19105 -680 19115 -650
rect 19145 -680 19155 -650
rect 19105 -690 19155 -680
rect 19190 -500 19240 -490
rect 19190 -530 19200 -500
rect 19230 -530 19240 -500
rect 19190 -550 19240 -530
rect 19190 -580 19200 -550
rect 19230 -580 19240 -550
rect 19190 -600 19240 -580
rect 19190 -630 19200 -600
rect 19230 -630 19240 -600
rect 19190 -650 19240 -630
rect 19190 -680 19200 -650
rect 19230 -680 19240 -650
rect 19190 -690 19240 -680
rect 19275 -500 19325 -490
rect 19275 -530 19285 -500
rect 19315 -530 19325 -500
rect 19275 -550 19325 -530
rect 19275 -580 19285 -550
rect 19315 -580 19325 -550
rect 19275 -600 19325 -580
rect 19275 -630 19285 -600
rect 19315 -630 19325 -600
rect 19275 -650 19325 -630
rect 19275 -680 19285 -650
rect 19315 -680 19325 -650
rect 19275 -690 19325 -680
rect 19360 -500 19410 -490
rect 19360 -530 19370 -500
rect 19400 -530 19410 -500
rect 19360 -550 19410 -530
rect 19360 -580 19370 -550
rect 19400 -580 19410 -550
rect 19360 -600 19410 -580
rect 19360 -630 19370 -600
rect 19400 -630 19410 -600
rect 19360 -650 19410 -630
rect 19360 -680 19370 -650
rect 19400 -680 19410 -650
rect 19360 -690 19410 -680
rect 19445 -500 19495 -490
rect 19445 -530 19455 -500
rect 19485 -530 19495 -500
rect 19445 -550 19495 -530
rect 19445 -580 19455 -550
rect 19485 -580 19495 -550
rect 19445 -600 19495 -580
rect 19445 -630 19455 -600
rect 19485 -630 19495 -600
rect 19445 -650 19495 -630
rect 19445 -680 19455 -650
rect 19485 -680 19495 -650
rect 19445 -690 19495 -680
rect 19530 -500 19580 -490
rect 19530 -530 19540 -500
rect 19570 -530 19580 -500
rect 19530 -550 19580 -530
rect 19530 -580 19540 -550
rect 19570 -580 19580 -550
rect 19530 -600 19580 -580
rect 19530 -630 19540 -600
rect 19570 -630 19580 -600
rect 19530 -650 19580 -630
rect 19530 -680 19540 -650
rect 19570 -680 19580 -650
rect 19530 -690 19580 -680
rect 19615 -500 19665 -490
rect 19615 -530 19625 -500
rect 19655 -530 19665 -500
rect 19615 -550 19665 -530
rect 19615 -580 19625 -550
rect 19655 -580 19665 -550
rect 19615 -600 19665 -580
rect 19615 -630 19625 -600
rect 19655 -630 19665 -600
rect 19615 -650 19665 -630
rect 19615 -680 19625 -650
rect 19655 -680 19665 -650
rect 19615 -690 19665 -680
rect 19700 -500 19750 -490
rect 19700 -530 19710 -500
rect 19740 -530 19750 -500
rect 19700 -550 19750 -530
rect 19700 -580 19710 -550
rect 19740 -580 19750 -550
rect 19700 -600 19750 -580
rect 19700 -630 19710 -600
rect 19740 -630 19750 -600
rect 19700 -650 19750 -630
rect 19700 -680 19710 -650
rect 19740 -680 19750 -650
rect 19700 -690 19750 -680
rect 19785 -500 19835 -490
rect 19785 -530 19795 -500
rect 19825 -530 19835 -500
rect 19785 -550 19835 -530
rect 19785 -580 19795 -550
rect 19825 -580 19835 -550
rect 19785 -600 19835 -580
rect 19785 -630 19795 -600
rect 19825 -630 19835 -600
rect 19785 -650 19835 -630
rect 19785 -680 19795 -650
rect 19825 -680 19835 -650
rect 19785 -690 19835 -680
rect 19870 -500 19920 -490
rect 19870 -530 19880 -500
rect 19910 -530 19920 -500
rect 19870 -550 19920 -530
rect 19870 -580 19880 -550
rect 19910 -580 19920 -550
rect 19870 -600 19920 -580
rect 19870 -630 19880 -600
rect 19910 -630 19920 -600
rect 19870 -650 19920 -630
rect 19870 -680 19880 -650
rect 19910 -680 19920 -650
rect 19870 -690 19920 -680
rect 19955 -500 20005 -490
rect 19955 -530 19965 -500
rect 19995 -530 20005 -500
rect 19955 -550 20005 -530
rect 19955 -580 19965 -550
rect 19995 -580 20005 -550
rect 19955 -600 20005 -580
rect 19955 -630 19965 -600
rect 19995 -630 20005 -600
rect 19955 -650 20005 -630
rect 19955 -680 19965 -650
rect 19995 -680 20005 -650
rect 19955 -690 20005 -680
rect 20040 -500 20090 -490
rect 20040 -530 20050 -500
rect 20080 -530 20090 -500
rect 20040 -550 20090 -530
rect 20040 -580 20050 -550
rect 20080 -580 20090 -550
rect 20040 -600 20090 -580
rect 20040 -630 20050 -600
rect 20080 -630 20090 -600
rect 20040 -650 20090 -630
rect 20040 -680 20050 -650
rect 20080 -680 20090 -650
rect 20040 -690 20090 -680
rect 20125 -500 20175 -490
rect 20125 -530 20135 -500
rect 20165 -530 20175 -500
rect 20125 -550 20175 -530
rect 20125 -580 20135 -550
rect 20165 -580 20175 -550
rect 20125 -600 20175 -580
rect 20125 -630 20135 -600
rect 20165 -630 20175 -600
rect 20125 -650 20175 -630
rect 20125 -680 20135 -650
rect 20165 -680 20175 -650
rect 20125 -690 20175 -680
rect 20210 -500 20260 -490
rect 20210 -530 20220 -500
rect 20250 -530 20260 -500
rect 20210 -550 20260 -530
rect 20210 -580 20220 -550
rect 20250 -580 20260 -550
rect 20210 -600 20260 -580
rect 20210 -630 20220 -600
rect 20250 -630 20260 -600
rect 20210 -650 20260 -630
rect 20210 -680 20220 -650
rect 20250 -680 20260 -650
rect 20210 -690 20260 -680
rect 20295 -500 20345 -490
rect 20295 -530 20305 -500
rect 20335 -530 20345 -500
rect 20295 -550 20345 -530
rect 20295 -580 20305 -550
rect 20335 -580 20345 -550
rect 20295 -600 20345 -580
rect 20295 -630 20305 -600
rect 20335 -630 20345 -600
rect 20295 -650 20345 -630
rect 20295 -680 20305 -650
rect 20335 -680 20345 -650
rect 20295 -690 20345 -680
rect 20380 -500 20430 -490
rect 20380 -530 20390 -500
rect 20420 -530 20430 -500
rect 20380 -550 20430 -530
rect 20380 -580 20390 -550
rect 20420 -580 20430 -550
rect 20380 -600 20430 -580
rect 20380 -630 20390 -600
rect 20420 -630 20430 -600
rect 20380 -650 20430 -630
rect 20380 -680 20390 -650
rect 20420 -680 20430 -650
rect 20380 -690 20430 -680
rect 20465 -500 20515 -490
rect 20465 -530 20475 -500
rect 20505 -530 20515 -500
rect 20465 -550 20515 -530
rect 20465 -580 20475 -550
rect 20505 -580 20515 -550
rect 20465 -600 20515 -580
rect 20465 -630 20475 -600
rect 20505 -630 20515 -600
rect 20465 -650 20515 -630
rect 20465 -680 20475 -650
rect 20505 -680 20515 -650
rect 20465 -690 20515 -680
rect 20550 -500 20600 -490
rect 20550 -530 20560 -500
rect 20590 -530 20600 -500
rect 20550 -550 20600 -530
rect 20550 -580 20560 -550
rect 20590 -580 20600 -550
rect 20550 -600 20600 -580
rect 20550 -630 20560 -600
rect 20590 -630 20600 -600
rect 20550 -650 20600 -630
rect 20550 -680 20560 -650
rect 20590 -680 20600 -650
rect 20550 -690 20600 -680
rect 20635 -500 20685 -490
rect 20635 -530 20645 -500
rect 20675 -530 20685 -500
rect 20635 -550 20685 -530
rect 20635 -580 20645 -550
rect 20675 -580 20685 -550
rect 20635 -600 20685 -580
rect 20635 -630 20645 -600
rect 20675 -630 20685 -600
rect 20635 -650 20685 -630
rect 20635 -680 20645 -650
rect 20675 -680 20685 -650
rect 20635 -690 20685 -680
rect 20720 -500 20770 -490
rect 20720 -530 20730 -500
rect 20760 -530 20770 -500
rect 20720 -550 20770 -530
rect 20720 -580 20730 -550
rect 20760 -580 20770 -550
rect 20720 -600 20770 -580
rect 20720 -630 20730 -600
rect 20760 -630 20770 -600
rect 20720 -650 20770 -630
rect 20720 -680 20730 -650
rect 20760 -680 20770 -650
rect 20720 -690 20770 -680
rect 20805 -500 20855 -490
rect 20805 -530 20815 -500
rect 20845 -530 20855 -500
rect 20805 -550 20855 -530
rect 20805 -580 20815 -550
rect 20845 -580 20855 -550
rect 20805 -600 20855 -580
rect 20805 -630 20815 -600
rect 20845 -630 20855 -600
rect 20805 -650 20855 -630
rect 20805 -680 20815 -650
rect 20845 -680 20855 -650
rect 20805 -690 20855 -680
rect 20890 -500 20940 -490
rect 20890 -530 20900 -500
rect 20930 -530 20940 -500
rect 20890 -550 20940 -530
rect 20890 -580 20900 -550
rect 20930 -580 20940 -550
rect 20890 -600 20940 -580
rect 20890 -630 20900 -600
rect 20930 -630 20940 -600
rect 20890 -650 20940 -630
rect 20890 -680 20900 -650
rect 20930 -680 20940 -650
rect 20890 -690 20940 -680
rect 20975 -500 21025 -490
rect 20975 -530 20985 -500
rect 21015 -530 21025 -500
rect 20975 -550 21025 -530
rect 20975 -580 20985 -550
rect 21015 -580 21025 -550
rect 20975 -600 21025 -580
rect 20975 -630 20985 -600
rect 21015 -630 21025 -600
rect 20975 -650 21025 -630
rect 20975 -680 20985 -650
rect 21015 -680 21025 -650
rect 20975 -690 21025 -680
rect 21060 -500 21110 -490
rect 21060 -530 21070 -500
rect 21100 -530 21110 -500
rect 21060 -550 21110 -530
rect 21060 -580 21070 -550
rect 21100 -580 21110 -550
rect 21060 -600 21110 -580
rect 21060 -630 21070 -600
rect 21100 -630 21110 -600
rect 21060 -650 21110 -630
rect 21060 -680 21070 -650
rect 21100 -680 21110 -650
rect 21060 -690 21110 -680
rect 21145 -500 21195 -490
rect 21145 -530 21155 -500
rect 21185 -530 21195 -500
rect 21145 -550 21195 -530
rect 21145 -580 21155 -550
rect 21185 -580 21195 -550
rect 21145 -600 21195 -580
rect 21145 -630 21155 -600
rect 21185 -630 21195 -600
rect 21145 -650 21195 -630
rect 21145 -680 21155 -650
rect 21185 -680 21195 -650
rect 21145 -690 21195 -680
rect 21230 -500 21280 -490
rect 21230 -530 21240 -500
rect 21270 -530 21280 -500
rect 21230 -550 21280 -530
rect 21230 -580 21240 -550
rect 21270 -580 21280 -550
rect 21230 -600 21280 -580
rect 21230 -630 21240 -600
rect 21270 -630 21280 -600
rect 21230 -650 21280 -630
rect 21230 -680 21240 -650
rect 21270 -680 21280 -650
rect 21230 -690 21280 -680
rect 21315 -500 21365 -490
rect 21315 -530 21325 -500
rect 21355 -530 21365 -500
rect 21315 -550 21365 -530
rect 21315 -580 21325 -550
rect 21355 -580 21365 -550
rect 21315 -600 21365 -580
rect 21315 -630 21325 -600
rect 21355 -630 21365 -600
rect 21315 -650 21365 -630
rect 21315 -680 21325 -650
rect 21355 -680 21365 -650
rect 21315 -690 21365 -680
rect 21400 -500 21450 -490
rect 21400 -530 21410 -500
rect 21440 -530 21450 -500
rect 21400 -550 21450 -530
rect 21400 -580 21410 -550
rect 21440 -580 21450 -550
rect 21400 -600 21450 -580
rect 21400 -630 21410 -600
rect 21440 -630 21450 -600
rect 21400 -650 21450 -630
rect 21400 -680 21410 -650
rect 21440 -680 21450 -650
rect 21400 -690 21450 -680
rect 21485 -500 21535 -490
rect 21485 -530 21495 -500
rect 21525 -530 21535 -500
rect 21485 -550 21535 -530
rect 21485 -580 21495 -550
rect 21525 -580 21535 -550
rect 21485 -600 21535 -580
rect 21485 -630 21495 -600
rect 21525 -630 21535 -600
rect 21485 -650 21535 -630
rect 21485 -680 21495 -650
rect 21525 -680 21535 -650
rect 21485 -690 21535 -680
rect 21570 -500 21620 -490
rect 21570 -530 21580 -500
rect 21610 -530 21620 -500
rect 21570 -550 21620 -530
rect 21570 -580 21580 -550
rect 21610 -580 21620 -550
rect 21570 -600 21620 -580
rect 21570 -630 21580 -600
rect 21610 -630 21620 -600
rect 21570 -650 21620 -630
rect 21570 -680 21580 -650
rect 21610 -680 21620 -650
rect 21570 -690 21620 -680
rect 21655 -500 21705 -490
rect 21655 -530 21665 -500
rect 21695 -530 21705 -500
rect 21655 -550 21705 -530
rect 21655 -580 21665 -550
rect 21695 -580 21705 -550
rect 21655 -600 21705 -580
rect 21655 -630 21665 -600
rect 21695 -630 21705 -600
rect 21655 -650 21705 -630
rect 21655 -680 21665 -650
rect 21695 -680 21705 -650
rect 21655 -690 21705 -680
rect 21740 -500 21790 -490
rect 21740 -530 21750 -500
rect 21780 -530 21790 -500
rect 21740 -550 21790 -530
rect 21740 -580 21750 -550
rect 21780 -580 21790 -550
rect 21740 -600 21790 -580
rect 21740 -630 21750 -600
rect 21780 -630 21790 -600
rect 21740 -650 21790 -630
rect 21740 -680 21750 -650
rect 21780 -680 21790 -650
rect 21740 -690 21790 -680
rect 21825 -500 21875 -490
rect 21825 -530 21835 -500
rect 21865 -530 21875 -500
rect 21825 -550 21875 -530
rect 21825 -580 21835 -550
rect 21865 -580 21875 -550
rect 21825 -600 21875 -580
rect 21825 -630 21835 -600
rect 21865 -630 21875 -600
rect 21825 -650 21875 -630
rect 21825 -680 21835 -650
rect 21865 -680 21875 -650
rect 21825 -690 21875 -680
rect 21910 -500 21960 -490
rect 21910 -530 21920 -500
rect 21950 -530 21960 -500
rect 21910 -550 21960 -530
rect 21910 -580 21920 -550
rect 21950 -580 21960 -550
rect 21910 -600 21960 -580
rect 21910 -630 21920 -600
rect 21950 -630 21960 -600
rect 21910 -650 21960 -630
rect 21910 -680 21920 -650
rect 21950 -680 21960 -650
rect 21910 -690 21960 -680
rect 21995 -500 22045 -490
rect 21995 -530 22005 -500
rect 22035 -530 22045 -500
rect 21995 -550 22045 -530
rect 21995 -580 22005 -550
rect 22035 -580 22045 -550
rect 21995 -600 22045 -580
rect 21995 -630 22005 -600
rect 22035 -630 22045 -600
rect 21995 -650 22045 -630
rect 21995 -680 22005 -650
rect 22035 -680 22045 -650
rect 21995 -690 22045 -680
rect 22080 -500 22130 -490
rect 22080 -530 22090 -500
rect 22120 -530 22130 -500
rect 22080 -550 22130 -530
rect 22080 -580 22090 -550
rect 22120 -580 22130 -550
rect 22080 -600 22130 -580
rect 22080 -630 22090 -600
rect 22120 -630 22130 -600
rect 22080 -650 22130 -630
rect 22080 -680 22090 -650
rect 22120 -680 22130 -650
rect 22080 -690 22130 -680
rect 22165 -500 22215 -490
rect 22165 -530 22175 -500
rect 22205 -530 22215 -500
rect 22165 -550 22215 -530
rect 22165 -580 22175 -550
rect 22205 -580 22215 -550
rect 22165 -600 22215 -580
rect 22165 -630 22175 -600
rect 22205 -630 22215 -600
rect 22165 -650 22215 -630
rect 22165 -680 22175 -650
rect 22205 -680 22215 -650
rect 22165 -690 22215 -680
rect 22250 -500 22300 -490
rect 22250 -530 22260 -500
rect 22290 -530 22300 -500
rect 22250 -550 22300 -530
rect 22250 -580 22260 -550
rect 22290 -580 22300 -550
rect 22250 -600 22300 -580
rect 22250 -630 22260 -600
rect 22290 -630 22300 -600
rect 22250 -650 22300 -630
rect 22250 -680 22260 -650
rect 22290 -680 22300 -650
rect 22250 -690 22300 -680
rect 22335 -500 22385 -490
rect 22335 -530 22345 -500
rect 22375 -530 22385 -500
rect 22335 -550 22385 -530
rect 22335 -580 22345 -550
rect 22375 -580 22385 -550
rect 22335 -600 22385 -580
rect 22335 -630 22345 -600
rect 22375 -630 22385 -600
rect 22335 -650 22385 -630
rect 22335 -680 22345 -650
rect 22375 -680 22385 -650
rect 22335 -690 22385 -680
rect 22420 -500 22470 -490
rect 22420 -530 22430 -500
rect 22460 -530 22470 -500
rect 22420 -550 22470 -530
rect 22420 -580 22430 -550
rect 22460 -580 22470 -550
rect 22420 -600 22470 -580
rect 22420 -630 22430 -600
rect 22460 -630 22470 -600
rect 22420 -650 22470 -630
rect 22420 -680 22430 -650
rect 22460 -680 22470 -650
rect 22420 -690 22470 -680
rect 22505 -500 22555 -490
rect 22505 -530 22515 -500
rect 22545 -530 22555 -500
rect 22505 -550 22555 -530
rect 22505 -580 22515 -550
rect 22545 -580 22555 -550
rect 22505 -600 22555 -580
rect 22505 -630 22515 -600
rect 22545 -630 22555 -600
rect 22505 -650 22555 -630
rect 22505 -680 22515 -650
rect 22545 -680 22555 -650
rect 22505 -690 22555 -680
rect 22590 -500 22640 -490
rect 22590 -530 22600 -500
rect 22630 -530 22640 -500
rect 22590 -550 22640 -530
rect 22590 -580 22600 -550
rect 22630 -580 22640 -550
rect 22590 -600 22640 -580
rect 22590 -630 22600 -600
rect 22630 -630 22640 -600
rect 22590 -650 22640 -630
rect 22590 -680 22600 -650
rect 22630 -680 22640 -650
rect 22590 -690 22640 -680
rect 22675 -500 22725 -490
rect 22675 -530 22685 -500
rect 22715 -530 22725 -500
rect 22675 -550 22725 -530
rect 22675 -580 22685 -550
rect 22715 -580 22725 -550
rect 22675 -600 22725 -580
rect 22675 -630 22685 -600
rect 22715 -630 22725 -600
rect 22675 -650 22725 -630
rect 22675 -680 22685 -650
rect 22715 -680 22725 -650
rect 22675 -690 22725 -680
rect 22760 -500 22810 -490
rect 22760 -530 22770 -500
rect 22800 -530 22810 -500
rect 22760 -550 22810 -530
rect 22760 -580 22770 -550
rect 22800 -580 22810 -550
rect 22760 -600 22810 -580
rect 22760 -630 22770 -600
rect 22800 -630 22810 -600
rect 22760 -650 22810 -630
rect 22760 -680 22770 -650
rect 22800 -680 22810 -650
rect 22760 -690 22810 -680
rect 22845 -500 22895 -490
rect 22845 -530 22855 -500
rect 22885 -530 22895 -500
rect 22845 -550 22895 -530
rect 22845 -580 22855 -550
rect 22885 -580 22895 -550
rect 22845 -600 22895 -580
rect 22845 -630 22855 -600
rect 22885 -630 22895 -600
rect 22845 -650 22895 -630
rect 22845 -680 22855 -650
rect 22885 -680 22895 -650
rect 22845 -690 22895 -680
rect 22930 -500 22980 -490
rect 22930 -530 22940 -500
rect 22970 -530 22980 -500
rect 22930 -550 22980 -530
rect 22930 -580 22940 -550
rect 22970 -580 22980 -550
rect 22930 -600 22980 -580
rect 22930 -630 22940 -600
rect 22970 -630 22980 -600
rect 22930 -650 22980 -630
rect 22930 -680 22940 -650
rect 22970 -680 22980 -650
rect 22930 -690 22980 -680
rect 23015 -500 23065 -490
rect 23015 -530 23025 -500
rect 23055 -530 23065 -500
rect 23015 -550 23065 -530
rect 23015 -580 23025 -550
rect 23055 -580 23065 -550
rect 23015 -600 23065 -580
rect 23015 -630 23025 -600
rect 23055 -630 23065 -600
rect 23015 -650 23065 -630
rect 23015 -680 23025 -650
rect 23055 -680 23065 -650
rect 23015 -690 23065 -680
rect 23100 -500 23150 -490
rect 23100 -530 23110 -500
rect 23140 -530 23150 -500
rect 23100 -550 23150 -530
rect 23100 -580 23110 -550
rect 23140 -580 23150 -550
rect 23100 -600 23150 -580
rect 23100 -630 23110 -600
rect 23140 -630 23150 -600
rect 23100 -650 23150 -630
rect 23100 -680 23110 -650
rect 23140 -680 23150 -650
rect 23100 -690 23150 -680
rect 23185 -500 23235 -490
rect 23185 -530 23195 -500
rect 23225 -530 23235 -500
rect 23185 -550 23235 -530
rect 23185 -580 23195 -550
rect 23225 -580 23235 -550
rect 23185 -600 23235 -580
rect 23185 -630 23195 -600
rect 23225 -630 23235 -600
rect 23185 -650 23235 -630
rect 23185 -680 23195 -650
rect 23225 -680 23235 -650
rect 23185 -690 23235 -680
rect 23270 -500 23320 -490
rect 23270 -530 23280 -500
rect 23310 -530 23320 -500
rect 23270 -550 23320 -530
rect 23270 -580 23280 -550
rect 23310 -580 23320 -550
rect 23270 -600 23320 -580
rect 23270 -630 23280 -600
rect 23310 -630 23320 -600
rect 23270 -650 23320 -630
rect 23270 -680 23280 -650
rect 23310 -680 23320 -650
rect 23270 -690 23320 -680
rect 23355 -500 23405 -490
rect 23355 -530 23365 -500
rect 23395 -530 23405 -500
rect 23355 -550 23405 -530
rect 23355 -580 23365 -550
rect 23395 -580 23405 -550
rect 23355 -600 23405 -580
rect 23355 -630 23365 -600
rect 23395 -630 23405 -600
rect 23355 -650 23405 -630
rect 23355 -680 23365 -650
rect 23395 -680 23405 -650
rect 23355 -690 23405 -680
rect 23440 -500 23490 -490
rect 23440 -530 23450 -500
rect 23480 -530 23490 -500
rect 23440 -550 23490 -530
rect 23440 -580 23450 -550
rect 23480 -580 23490 -550
rect 23440 -600 23490 -580
rect 23440 -630 23450 -600
rect 23480 -630 23490 -600
rect 23440 -650 23490 -630
rect 23440 -680 23450 -650
rect 23480 -680 23490 -650
rect 23440 -690 23490 -680
rect 23525 -500 23575 -490
rect 23525 -530 23535 -500
rect 23565 -530 23575 -500
rect 23525 -550 23575 -530
rect 23525 -580 23535 -550
rect 23565 -580 23575 -550
rect 23525 -600 23575 -580
rect 23525 -630 23535 -600
rect 23565 -630 23575 -600
rect 23525 -650 23575 -630
rect 23525 -680 23535 -650
rect 23565 -680 23575 -650
rect 23525 -690 23575 -680
rect 23610 -500 23660 -490
rect 23610 -530 23620 -500
rect 23650 -530 23660 -500
rect 23610 -550 23660 -530
rect 23610 -580 23620 -550
rect 23650 -580 23660 -550
rect 23610 -600 23660 -580
rect 23610 -630 23620 -600
rect 23650 -630 23660 -600
rect 23610 -650 23660 -630
rect 23610 -680 23620 -650
rect 23650 -680 23660 -650
rect 23610 -690 23660 -680
rect 23695 -500 23745 -490
rect 23695 -530 23705 -500
rect 23735 -530 23745 -500
rect 23695 -550 23745 -530
rect 23695 -580 23705 -550
rect 23735 -580 23745 -550
rect 23695 -600 23745 -580
rect 23695 -630 23705 -600
rect 23735 -630 23745 -600
rect 23695 -650 23745 -630
rect 23695 -680 23705 -650
rect 23735 -680 23745 -650
rect 23695 -690 23745 -680
rect 23780 -500 23830 -490
rect 23780 -530 23790 -500
rect 23820 -530 23830 -500
rect 23780 -550 23830 -530
rect 23780 -580 23790 -550
rect 23820 -580 23830 -550
rect 23780 -600 23830 -580
rect 23780 -630 23790 -600
rect 23820 -630 23830 -600
rect 23780 -650 23830 -630
rect 23780 -680 23790 -650
rect 23820 -680 23830 -650
rect 23780 -690 23830 -680
rect 23865 -500 23915 -490
rect 23865 -530 23875 -500
rect 23905 -530 23915 -500
rect 23865 -550 23915 -530
rect 23865 -580 23875 -550
rect 23905 -580 23915 -550
rect 23865 -600 23915 -580
rect 23865 -630 23875 -600
rect 23905 -630 23915 -600
rect 23865 -650 23915 -630
rect 23865 -680 23875 -650
rect 23905 -680 23915 -650
rect 23865 -690 23915 -680
rect 23950 -500 24000 -490
rect 23950 -530 23960 -500
rect 23990 -530 24000 -500
rect 23950 -550 24000 -530
rect 23950 -580 23960 -550
rect 23990 -580 24000 -550
rect 23950 -600 24000 -580
rect 23950 -630 23960 -600
rect 23990 -630 24000 -600
rect 23950 -650 24000 -630
rect 23950 -680 23960 -650
rect 23990 -680 24000 -650
rect 23950 -690 24000 -680
rect 24035 -500 24085 -490
rect 24035 -530 24045 -500
rect 24075 -530 24085 -500
rect 24035 -550 24085 -530
rect 24035 -580 24045 -550
rect 24075 -580 24085 -550
rect 24035 -600 24085 -580
rect 24035 -630 24045 -600
rect 24075 -630 24085 -600
rect 24035 -650 24085 -630
rect 24035 -680 24045 -650
rect 24075 -680 24085 -650
rect 24035 -690 24085 -680
rect 24120 -500 24170 -490
rect 24120 -530 24130 -500
rect 24160 -530 24170 -500
rect 24120 -550 24170 -530
rect 24120 -580 24130 -550
rect 24160 -580 24170 -550
rect 24120 -600 24170 -580
rect 24120 -630 24130 -600
rect 24160 -630 24170 -600
rect 24120 -650 24170 -630
rect 24120 -680 24130 -650
rect 24160 -680 24170 -650
rect 24120 -690 24170 -680
rect 24205 -500 24255 -490
rect 24205 -530 24215 -500
rect 24245 -530 24255 -500
rect 24205 -550 24255 -530
rect 24205 -580 24215 -550
rect 24245 -580 24255 -550
rect 24205 -600 24255 -580
rect 24205 -630 24215 -600
rect 24245 -630 24255 -600
rect 24205 -650 24255 -630
rect 24205 -680 24215 -650
rect 24245 -680 24255 -650
rect 24205 -690 24255 -680
rect 24290 -500 24340 -490
rect 24290 -530 24300 -500
rect 24330 -530 24340 -500
rect 24290 -550 24340 -530
rect 24290 -580 24300 -550
rect 24330 -580 24340 -550
rect 24290 -600 24340 -580
rect 24290 -630 24300 -600
rect 24330 -630 24340 -600
rect 24290 -650 24340 -630
rect 24290 -680 24300 -650
rect 24330 -680 24340 -650
rect 24290 -690 24340 -680
rect 24375 -500 24425 -490
rect 24375 -530 24385 -500
rect 24415 -530 24425 -500
rect 24375 -550 24425 -530
rect 24375 -580 24385 -550
rect 24415 -580 24425 -550
rect 24375 -600 24425 -580
rect 24375 -630 24385 -600
rect 24415 -630 24425 -600
rect 24375 -650 24425 -630
rect 24375 -680 24385 -650
rect 24415 -680 24425 -650
rect 24375 -690 24425 -680
rect 24460 -500 24510 -490
rect 24460 -530 24470 -500
rect 24500 -530 24510 -500
rect 24460 -550 24510 -530
rect 24460 -580 24470 -550
rect 24500 -580 24510 -550
rect 24460 -600 24510 -580
rect 24460 -630 24470 -600
rect 24500 -630 24510 -600
rect 24460 -650 24510 -630
rect 24460 -680 24470 -650
rect 24500 -680 24510 -650
rect 24460 -690 24510 -680
rect 24545 -500 24595 -490
rect 24545 -530 24555 -500
rect 24585 -530 24595 -500
rect 24545 -550 24595 -530
rect 24545 -580 24555 -550
rect 24585 -580 24595 -550
rect 24545 -600 24595 -580
rect 24545 -630 24555 -600
rect 24585 -630 24595 -600
rect 24545 -650 24595 -630
rect 24545 -680 24555 -650
rect 24585 -680 24595 -650
rect 24545 -690 24595 -680
rect 24630 -500 24680 -490
rect 24630 -530 24640 -500
rect 24670 -530 24680 -500
rect 24630 -550 24680 -530
rect 24630 -580 24640 -550
rect 24670 -580 24680 -550
rect 24630 -600 24680 -580
rect 24630 -630 24640 -600
rect 24670 -630 24680 -600
rect 24630 -650 24680 -630
rect 24630 -680 24640 -650
rect 24670 -680 24680 -650
rect 24630 -690 24680 -680
rect 24715 -500 24765 -490
rect 24715 -530 24725 -500
rect 24755 -530 24765 -500
rect 24715 -550 24765 -530
rect 24715 -580 24725 -550
rect 24755 -580 24765 -550
rect 24715 -600 24765 -580
rect 24715 -630 24725 -600
rect 24755 -630 24765 -600
rect 24715 -650 24765 -630
rect 24715 -680 24725 -650
rect 24755 -680 24765 -650
rect 24715 -690 24765 -680
rect 24800 -500 24850 -490
rect 24800 -530 24810 -500
rect 24840 -530 24850 -500
rect 24800 -550 24850 -530
rect 24800 -580 24810 -550
rect 24840 -580 24850 -550
rect 24800 -600 24850 -580
rect 24800 -630 24810 -600
rect 24840 -630 24850 -600
rect 24800 -650 24850 -630
rect 24800 -680 24810 -650
rect 24840 -680 24850 -650
rect 24800 -690 24850 -680
rect 24885 -500 24935 -490
rect 24885 -530 24895 -500
rect 24925 -530 24935 -500
rect 24885 -550 24935 -530
rect 24885 -580 24895 -550
rect 24925 -580 24935 -550
rect 24885 -600 24935 -580
rect 24885 -630 24895 -600
rect 24925 -630 24935 -600
rect 24885 -650 24935 -630
rect 24885 -680 24895 -650
rect 24925 -680 24935 -650
rect 24885 -690 24935 -680
rect 24970 -500 25020 -490
rect 24970 -530 24980 -500
rect 25010 -530 25020 -500
rect 24970 -550 25020 -530
rect 24970 -580 24980 -550
rect 25010 -580 25020 -550
rect 24970 -600 25020 -580
rect 24970 -630 24980 -600
rect 25010 -630 25020 -600
rect 24970 -650 25020 -630
rect 24970 -680 24980 -650
rect 25010 -680 25020 -650
rect 24970 -690 25020 -680
rect 25055 -500 25105 -490
rect 25055 -530 25065 -500
rect 25095 -530 25105 -500
rect 25055 -550 25105 -530
rect 25055 -580 25065 -550
rect 25095 -580 25105 -550
rect 25055 -600 25105 -580
rect 25055 -630 25065 -600
rect 25095 -630 25105 -600
rect 25055 -650 25105 -630
rect 25055 -680 25065 -650
rect 25095 -680 25105 -650
rect 25055 -690 25105 -680
rect 25140 -500 25190 -490
rect 25140 -530 25150 -500
rect 25180 -530 25190 -500
rect 25140 -550 25190 -530
rect 25140 -580 25150 -550
rect 25180 -580 25190 -550
rect 25140 -600 25190 -580
rect 25140 -630 25150 -600
rect 25180 -630 25190 -600
rect 25140 -650 25190 -630
rect 25140 -680 25150 -650
rect 25180 -680 25190 -650
rect 25140 -690 25190 -680
rect 25225 -500 25275 -490
rect 25225 -530 25235 -500
rect 25265 -530 25275 -500
rect 25225 -550 25275 -530
rect 25225 -580 25235 -550
rect 25265 -580 25275 -550
rect 25225 -600 25275 -580
rect 25225 -630 25235 -600
rect 25265 -630 25275 -600
rect 25225 -650 25275 -630
rect 25225 -680 25235 -650
rect 25265 -680 25275 -650
rect 25225 -690 25275 -680
rect 25310 -500 25360 -490
rect 25310 -530 25320 -500
rect 25350 -530 25360 -500
rect 25310 -550 25360 -530
rect 25310 -580 25320 -550
rect 25350 -580 25360 -550
rect 25310 -600 25360 -580
rect 25310 -630 25320 -600
rect 25350 -630 25360 -600
rect 25310 -650 25360 -630
rect 25310 -680 25320 -650
rect 25350 -680 25360 -650
rect 25310 -690 25360 -680
rect 25395 -500 25445 -490
rect 25395 -530 25405 -500
rect 25435 -530 25445 -500
rect 25395 -550 25445 -530
rect 25395 -580 25405 -550
rect 25435 -580 25445 -550
rect 25395 -600 25445 -580
rect 25395 -630 25405 -600
rect 25435 -630 25445 -600
rect 25395 -650 25445 -630
rect 25395 -680 25405 -650
rect 25435 -680 25445 -650
rect 25395 -690 25445 -680
rect 25480 -500 25530 -490
rect 25480 -530 25490 -500
rect 25520 -530 25530 -500
rect 25480 -550 25530 -530
rect 25480 -580 25490 -550
rect 25520 -580 25530 -550
rect 25480 -600 25530 -580
rect 25480 -630 25490 -600
rect 25520 -630 25530 -600
rect 25480 -650 25530 -630
rect 25480 -680 25490 -650
rect 25520 -680 25530 -650
rect 25480 -690 25530 -680
rect 25565 -500 25615 -490
rect 25565 -530 25575 -500
rect 25605 -530 25615 -500
rect 25565 -550 25615 -530
rect 25565 -580 25575 -550
rect 25605 -580 25615 -550
rect 25565 -600 25615 -580
rect 25565 -630 25575 -600
rect 25605 -630 25615 -600
rect 25565 -650 25615 -630
rect 25565 -680 25575 -650
rect 25605 -680 25615 -650
rect 25565 -690 25615 -680
rect 25650 -500 25700 -490
rect 25650 -530 25660 -500
rect 25690 -530 25700 -500
rect 25650 -550 25700 -530
rect 25650 -580 25660 -550
rect 25690 -580 25700 -550
rect 25650 -600 25700 -580
rect 25650 -630 25660 -600
rect 25690 -630 25700 -600
rect 25650 -650 25700 -630
rect 25650 -680 25660 -650
rect 25690 -680 25700 -650
rect 25650 -690 25700 -680
rect 25735 -500 25785 -490
rect 25735 -530 25745 -500
rect 25775 -530 25785 -500
rect 25735 -550 25785 -530
rect 25735 -580 25745 -550
rect 25775 -580 25785 -550
rect 25735 -600 25785 -580
rect 25735 -630 25745 -600
rect 25775 -630 25785 -600
rect 25735 -650 25785 -630
rect 25735 -680 25745 -650
rect 25775 -680 25785 -650
rect 25735 -690 25785 -680
rect 25820 -500 25870 -490
rect 25820 -530 25830 -500
rect 25860 -530 25870 -500
rect 25820 -550 25870 -530
rect 25820 -580 25830 -550
rect 25860 -580 25870 -550
rect 25820 -600 25870 -580
rect 25820 -630 25830 -600
rect 25860 -630 25870 -600
rect 25820 -650 25870 -630
rect 25820 -680 25830 -650
rect 25860 -680 25870 -650
rect 25820 -690 25870 -680
rect 25905 -500 25955 -490
rect 25905 -530 25915 -500
rect 25945 -530 25955 -500
rect 25905 -550 25955 -530
rect 25905 -580 25915 -550
rect 25945 -580 25955 -550
rect 25905 -600 25955 -580
rect 25905 -630 25915 -600
rect 25945 -630 25955 -600
rect 25905 -650 25955 -630
rect 25905 -680 25915 -650
rect 25945 -680 25955 -650
rect 25905 -690 25955 -680
rect 25990 -500 26040 -490
rect 25990 -530 26000 -500
rect 26030 -530 26040 -500
rect 25990 -550 26040 -530
rect 25990 -580 26000 -550
rect 26030 -580 26040 -550
rect 25990 -600 26040 -580
rect 25990 -630 26000 -600
rect 26030 -630 26040 -600
rect 25990 -650 26040 -630
rect 25990 -680 26000 -650
rect 26030 -680 26040 -650
rect 25990 -690 26040 -680
rect 26075 -500 26125 -490
rect 26075 -530 26085 -500
rect 26115 -530 26125 -500
rect 26075 -550 26125 -530
rect 26075 -580 26085 -550
rect 26115 -580 26125 -550
rect 26075 -600 26125 -580
rect 26075 -630 26085 -600
rect 26115 -630 26125 -600
rect 26075 -650 26125 -630
rect 26075 -680 26085 -650
rect 26115 -680 26125 -650
rect 26075 -690 26125 -680
rect 26160 -500 26210 -490
rect 26160 -530 26170 -500
rect 26200 -530 26210 -500
rect 26160 -550 26210 -530
rect 26160 -580 26170 -550
rect 26200 -580 26210 -550
rect 26160 -600 26210 -580
rect 26160 -630 26170 -600
rect 26200 -630 26210 -600
rect 26160 -650 26210 -630
rect 26160 -680 26170 -650
rect 26200 -680 26210 -650
rect 26160 -690 26210 -680
rect 26245 -500 26295 -490
rect 26245 -530 26255 -500
rect 26285 -530 26295 -500
rect 26245 -550 26295 -530
rect 26245 -580 26255 -550
rect 26285 -580 26295 -550
rect 26245 -600 26295 -580
rect 26245 -630 26255 -600
rect 26285 -630 26295 -600
rect 26245 -650 26295 -630
rect 26245 -680 26255 -650
rect 26285 -680 26295 -650
rect 26245 -690 26295 -680
rect 26330 -500 26380 -490
rect 26330 -530 26340 -500
rect 26370 -530 26380 -500
rect 26330 -550 26380 -530
rect 26330 -580 26340 -550
rect 26370 -580 26380 -550
rect 26330 -600 26380 -580
rect 26330 -630 26340 -600
rect 26370 -630 26380 -600
rect 26330 -650 26380 -630
rect 26330 -680 26340 -650
rect 26370 -680 26380 -650
rect 26330 -690 26380 -680
rect 26415 -500 26465 -490
rect 26415 -530 26425 -500
rect 26455 -530 26465 -500
rect 26415 -550 26465 -530
rect 26415 -580 26425 -550
rect 26455 -580 26465 -550
rect 26415 -600 26465 -580
rect 26415 -630 26425 -600
rect 26455 -630 26465 -600
rect 26415 -650 26465 -630
rect 26415 -680 26425 -650
rect 26455 -680 26465 -650
rect 26415 -690 26465 -680
rect 26500 -500 26550 -490
rect 26500 -530 26510 -500
rect 26540 -530 26550 -500
rect 26500 -550 26550 -530
rect 26500 -580 26510 -550
rect 26540 -580 26550 -550
rect 26500 -600 26550 -580
rect 26500 -630 26510 -600
rect 26540 -630 26550 -600
rect 26500 -650 26550 -630
rect 26500 -680 26510 -650
rect 26540 -680 26550 -650
rect 26500 -690 26550 -680
rect 26585 -500 26635 -490
rect 26585 -530 26595 -500
rect 26625 -530 26635 -500
rect 26585 -550 26635 -530
rect 26585 -580 26595 -550
rect 26625 -580 26635 -550
rect 26585 -600 26635 -580
rect 26585 -630 26595 -600
rect 26625 -630 26635 -600
rect 26585 -650 26635 -630
rect 26585 -680 26595 -650
rect 26625 -680 26635 -650
rect 26585 -690 26635 -680
rect 26670 -500 26720 -490
rect 26670 -530 26680 -500
rect 26710 -530 26720 -500
rect 26670 -550 26720 -530
rect 26670 -580 26680 -550
rect 26710 -580 26720 -550
rect 26670 -600 26720 -580
rect 26670 -630 26680 -600
rect 26710 -630 26720 -600
rect 26670 -650 26720 -630
rect 26670 -680 26680 -650
rect 26710 -680 26720 -650
rect 26670 -690 26720 -680
rect 26755 -500 26805 -490
rect 26755 -530 26765 -500
rect 26795 -530 26805 -500
rect 26755 -550 26805 -530
rect 26755 -580 26765 -550
rect 26795 -580 26805 -550
rect 26755 -600 26805 -580
rect 26755 -630 26765 -600
rect 26795 -630 26805 -600
rect 26755 -650 26805 -630
rect 26755 -680 26765 -650
rect 26795 -680 26805 -650
rect 26755 -690 26805 -680
rect 26840 -500 26890 -490
rect 26840 -530 26850 -500
rect 26880 -530 26890 -500
rect 26840 -550 26890 -530
rect 26840 -580 26850 -550
rect 26880 -580 26890 -550
rect 26840 -600 26890 -580
rect 26840 -630 26850 -600
rect 26880 -630 26890 -600
rect 26840 -650 26890 -630
rect 26840 -680 26850 -650
rect 26880 -680 26890 -650
rect 26840 -690 26890 -680
rect 26925 -500 26975 -490
rect 26925 -530 26935 -500
rect 26965 -530 26975 -500
rect 26925 -550 26975 -530
rect 26925 -580 26935 -550
rect 26965 -580 26975 -550
rect 26925 -600 26975 -580
rect 26925 -630 26935 -600
rect 26965 -630 26975 -600
rect 26925 -650 26975 -630
rect 26925 -680 26935 -650
rect 26965 -680 26975 -650
rect 26925 -690 26975 -680
rect 27010 -500 27060 -490
rect 27010 -530 27020 -500
rect 27050 -530 27060 -500
rect 27010 -550 27060 -530
rect 27010 -580 27020 -550
rect 27050 -580 27060 -550
rect 27010 -600 27060 -580
rect 27010 -630 27020 -600
rect 27050 -630 27060 -600
rect 27010 -650 27060 -630
rect 27010 -680 27020 -650
rect 27050 -680 27060 -650
rect 27010 -690 27060 -680
rect 27095 -500 27145 -490
rect 27095 -530 27105 -500
rect 27135 -530 27145 -500
rect 27095 -550 27145 -530
rect 27095 -580 27105 -550
rect 27135 -580 27145 -550
rect 27095 -600 27145 -580
rect 27095 -630 27105 -600
rect 27135 -630 27145 -600
rect 27095 -650 27145 -630
rect 27095 -680 27105 -650
rect 27135 -680 27145 -650
rect 27095 -690 27145 -680
rect 27180 -500 27230 -490
rect 27180 -530 27190 -500
rect 27220 -530 27230 -500
rect 27180 -550 27230 -530
rect 27180 -580 27190 -550
rect 27220 -580 27230 -550
rect 27180 -600 27230 -580
rect 27180 -630 27190 -600
rect 27220 -630 27230 -600
rect 27180 -650 27230 -630
rect 27180 -680 27190 -650
rect 27220 -680 27230 -650
rect 27180 -690 27230 -680
rect 27265 -500 27315 -490
rect 27265 -530 27275 -500
rect 27305 -530 27315 -500
rect 27265 -550 27315 -530
rect 27265 -580 27275 -550
rect 27305 -580 27315 -550
rect 27265 -600 27315 -580
rect 27265 -630 27275 -600
rect 27305 -630 27315 -600
rect 27265 -650 27315 -630
rect 27265 -680 27275 -650
rect 27305 -680 27315 -650
rect 27265 -690 27315 -680
rect 27350 -500 27400 -490
rect 27350 -530 27360 -500
rect 27390 -530 27400 -500
rect 27350 -550 27400 -530
rect 27350 -580 27360 -550
rect 27390 -580 27400 -550
rect 27350 -600 27400 -580
rect 27350 -630 27360 -600
rect 27390 -630 27400 -600
rect 27350 -650 27400 -630
rect 27350 -680 27360 -650
rect 27390 -680 27400 -650
rect 27350 -690 27400 -680
rect 27435 -500 27485 -490
rect 27435 -530 27445 -500
rect 27475 -530 27485 -500
rect 27435 -550 27485 -530
rect 27435 -580 27445 -550
rect 27475 -580 27485 -550
rect 27435 -600 27485 -580
rect 27435 -630 27445 -600
rect 27475 -630 27485 -600
rect 27435 -650 27485 -630
rect 27435 -680 27445 -650
rect 27475 -680 27485 -650
rect 27435 -690 27485 -680
rect 27520 -500 27570 -490
rect 27520 -530 27530 -500
rect 27560 -530 27570 -500
rect 27520 -550 27570 -530
rect 27520 -580 27530 -550
rect 27560 -580 27570 -550
rect 27520 -600 27570 -580
rect 27520 -630 27530 -600
rect 27560 -630 27570 -600
rect 27520 -650 27570 -630
rect 27520 -680 27530 -650
rect 27560 -680 27570 -650
rect 27520 -690 27570 -680
rect 27605 -500 27655 -490
rect 27605 -530 27615 -500
rect 27645 -530 27655 -500
rect 27605 -550 27655 -530
rect 27605 -580 27615 -550
rect 27645 -580 27655 -550
rect 27605 -600 27655 -580
rect 27605 -630 27615 -600
rect 27645 -630 27655 -600
rect 27605 -650 27655 -630
rect 27605 -680 27615 -650
rect 27645 -680 27655 -650
rect 27605 -690 27655 -680
rect 27690 -500 27740 -490
rect 27690 -530 27700 -500
rect 27730 -530 27740 -500
rect 27690 -550 27740 -530
rect 27690 -580 27700 -550
rect 27730 -580 27740 -550
rect 27690 -600 27740 -580
rect 27690 -630 27700 -600
rect 27730 -630 27740 -600
rect 27690 -650 27740 -630
rect 27690 -680 27700 -650
rect 27730 -680 27740 -650
rect 27690 -690 27740 -680
rect 27775 -500 27825 -490
rect 27775 -530 27785 -500
rect 27815 -530 27825 -500
rect 27775 -550 27825 -530
rect 27775 -580 27785 -550
rect 27815 -580 27825 -550
rect 27775 -600 27825 -580
rect 27775 -630 27785 -600
rect 27815 -630 27825 -600
rect 27775 -650 27825 -630
rect 27775 -680 27785 -650
rect 27815 -680 27825 -650
rect 27775 -690 27825 -680
rect 27860 -500 27910 -490
rect 27860 -530 27870 -500
rect 27900 -530 27910 -500
rect 27860 -550 27910 -530
rect 27860 -580 27870 -550
rect 27900 -580 27910 -550
rect 27860 -600 27910 -580
rect 27860 -630 27870 -600
rect 27900 -630 27910 -600
rect 27860 -650 27910 -630
rect 27860 -680 27870 -650
rect 27900 -680 27910 -650
rect 27860 -690 27910 -680
rect 27945 -500 27995 -490
rect 27945 -530 27955 -500
rect 27985 -530 27995 -500
rect 27945 -550 27995 -530
rect 27945 -580 27955 -550
rect 27985 -580 27995 -550
rect 27945 -600 27995 -580
rect 27945 -630 27955 -600
rect 27985 -630 27995 -600
rect 27945 -650 27995 -630
rect 27945 -680 27955 -650
rect 27985 -680 27995 -650
rect 27945 -690 27995 -680
rect 28030 -500 28080 -490
rect 28030 -530 28040 -500
rect 28070 -530 28080 -500
rect 28030 -550 28080 -530
rect 28030 -580 28040 -550
rect 28070 -580 28080 -550
rect 28030 -600 28080 -580
rect 28030 -630 28040 -600
rect 28070 -630 28080 -600
rect 28030 -650 28080 -630
rect 28030 -680 28040 -650
rect 28070 -680 28080 -650
rect 28030 -690 28080 -680
rect 28115 -500 28165 -490
rect 28115 -530 28125 -500
rect 28155 -530 28165 -500
rect 28115 -550 28165 -530
rect 28115 -580 28125 -550
rect 28155 -580 28165 -550
rect 28115 -600 28165 -580
rect 28115 -630 28125 -600
rect 28155 -630 28165 -600
rect 28115 -650 28165 -630
rect 28115 -680 28125 -650
rect 28155 -680 28165 -650
rect 28115 -690 28165 -680
rect 28200 -500 28250 -490
rect 28200 -530 28210 -500
rect 28240 -530 28250 -500
rect 28200 -550 28250 -530
rect 28200 -580 28210 -550
rect 28240 -580 28250 -550
rect 28200 -600 28250 -580
rect 28200 -630 28210 -600
rect 28240 -630 28250 -600
rect 28200 -650 28250 -630
rect 28200 -680 28210 -650
rect 28240 -680 28250 -650
rect 28200 -690 28250 -680
rect 28285 -500 28335 -490
rect 28285 -530 28295 -500
rect 28325 -530 28335 -500
rect 28285 -550 28335 -530
rect 28285 -580 28295 -550
rect 28325 -580 28335 -550
rect 28285 -600 28335 -580
rect 28285 -630 28295 -600
rect 28325 -630 28335 -600
rect 28285 -650 28335 -630
rect 28285 -680 28295 -650
rect 28325 -680 28335 -650
rect 28285 -690 28335 -680
rect 28370 -500 28420 -490
rect 28370 -530 28380 -500
rect 28410 -530 28420 -500
rect 28370 -550 28420 -530
rect 28370 -580 28380 -550
rect 28410 -580 28420 -550
rect 28370 -600 28420 -580
rect 28370 -630 28380 -600
rect 28410 -630 28420 -600
rect 28370 -650 28420 -630
rect 28370 -680 28380 -650
rect 28410 -680 28420 -650
rect 28370 -690 28420 -680
rect 28455 -500 28505 -490
rect 28455 -530 28465 -500
rect 28495 -530 28505 -500
rect 28455 -550 28505 -530
rect 28455 -580 28465 -550
rect 28495 -580 28505 -550
rect 28455 -600 28505 -580
rect 28455 -630 28465 -600
rect 28495 -630 28505 -600
rect 28455 -650 28505 -630
rect 28455 -680 28465 -650
rect 28495 -680 28505 -650
rect 28455 -690 28505 -680
rect 28540 -500 28590 -490
rect 28540 -530 28550 -500
rect 28580 -530 28590 -500
rect 28540 -550 28590 -530
rect 28540 -580 28550 -550
rect 28580 -580 28590 -550
rect 28540 -600 28590 -580
rect 28540 -630 28550 -600
rect 28580 -630 28590 -600
rect 28540 -650 28590 -630
rect 28540 -680 28550 -650
rect 28580 -680 28590 -650
rect 28540 -690 28590 -680
rect 28625 -500 28675 -490
rect 28625 -530 28635 -500
rect 28665 -530 28675 -500
rect 28625 -550 28675 -530
rect 28625 -580 28635 -550
rect 28665 -580 28675 -550
rect 28625 -600 28675 -580
rect 28625 -630 28635 -600
rect 28665 -630 28675 -600
rect 28625 -650 28675 -630
rect 28625 -680 28635 -650
rect 28665 -680 28675 -650
rect 28625 -690 28675 -680
rect 28710 -500 28760 -490
rect 28710 -530 28720 -500
rect 28750 -530 28760 -500
rect 28710 -550 28760 -530
rect 28710 -580 28720 -550
rect 28750 -580 28760 -550
rect 28710 -600 28760 -580
rect 28710 -630 28720 -600
rect 28750 -630 28760 -600
rect 28710 -650 28760 -630
rect 28710 -680 28720 -650
rect 28750 -680 28760 -650
rect 28710 -690 28760 -680
rect 28795 -500 28845 -490
rect 28795 -530 28805 -500
rect 28835 -530 28845 -500
rect 28795 -550 28845 -530
rect 28795 -580 28805 -550
rect 28835 -580 28845 -550
rect 28795 -600 28845 -580
rect 28795 -630 28805 -600
rect 28835 -630 28845 -600
rect 28795 -650 28845 -630
rect 28795 -680 28805 -650
rect 28835 -680 28845 -650
rect 28795 -690 28845 -680
rect 28880 -500 28930 -490
rect 28880 -530 28890 -500
rect 28920 -530 28930 -500
rect 28880 -550 28930 -530
rect 28880 -580 28890 -550
rect 28920 -580 28930 -550
rect 28880 -600 28930 -580
rect 28880 -630 28890 -600
rect 28920 -630 28930 -600
rect 28880 -650 28930 -630
rect 28880 -680 28890 -650
rect 28920 -680 28930 -650
rect 28880 -690 28930 -680
rect 28965 -500 29015 -490
rect 28965 -530 28975 -500
rect 29005 -530 29015 -500
rect 28965 -550 29015 -530
rect 28965 -580 28975 -550
rect 29005 -580 29015 -550
rect 28965 -600 29015 -580
rect 28965 -630 28975 -600
rect 29005 -630 29015 -600
rect 28965 -650 29015 -630
rect 28965 -680 28975 -650
rect 29005 -680 29015 -650
rect 28965 -690 29015 -680
rect 29050 -500 29100 -490
rect 29050 -530 29060 -500
rect 29090 -530 29100 -500
rect 29050 -550 29100 -530
rect 29050 -580 29060 -550
rect 29090 -580 29100 -550
rect 29050 -600 29100 -580
rect 29050 -630 29060 -600
rect 29090 -630 29100 -600
rect 29050 -650 29100 -630
rect 29050 -680 29060 -650
rect 29090 -680 29100 -650
rect 29050 -690 29100 -680
rect 29135 -500 29185 -490
rect 29135 -530 29145 -500
rect 29175 -530 29185 -500
rect 29135 -550 29185 -530
rect 29135 -580 29145 -550
rect 29175 -580 29185 -550
rect 29135 -600 29185 -580
rect 29135 -630 29145 -600
rect 29175 -630 29185 -600
rect 29135 -650 29185 -630
rect 29135 -680 29145 -650
rect 29175 -680 29185 -650
rect 29135 -690 29185 -680
rect 29220 -500 29270 -490
rect 29220 -530 29230 -500
rect 29260 -530 29270 -500
rect 29220 -550 29270 -530
rect 29220 -580 29230 -550
rect 29260 -580 29270 -550
rect 29220 -600 29270 -580
rect 29220 -630 29230 -600
rect 29260 -630 29270 -600
rect 29220 -650 29270 -630
rect 29220 -680 29230 -650
rect 29260 -680 29270 -650
rect 29220 -690 29270 -680
rect 29305 -500 29355 -490
rect 29305 -530 29315 -500
rect 29345 -530 29355 -500
rect 29305 -550 29355 -530
rect 29305 -580 29315 -550
rect 29345 -580 29355 -550
rect 29305 -600 29355 -580
rect 29305 -630 29315 -600
rect 29345 -630 29355 -600
rect 29305 -650 29355 -630
rect 29305 -680 29315 -650
rect 29345 -680 29355 -650
rect 29305 -690 29355 -680
rect 29390 -500 29440 -490
rect 29390 -530 29400 -500
rect 29430 -530 29440 -500
rect 29390 -550 29440 -530
rect 29390 -580 29400 -550
rect 29430 -580 29440 -550
rect 29390 -600 29440 -580
rect 29390 -630 29400 -600
rect 29430 -630 29440 -600
rect 29390 -650 29440 -630
rect 29390 -680 29400 -650
rect 29430 -680 29440 -650
rect 29390 -690 29440 -680
rect 29475 -500 29525 -490
rect 29475 -530 29485 -500
rect 29515 -530 29525 -500
rect 29475 -550 29525 -530
rect 29475 -580 29485 -550
rect 29515 -580 29525 -550
rect 29475 -600 29525 -580
rect 29475 -630 29485 -600
rect 29515 -630 29525 -600
rect 29475 -650 29525 -630
rect 29475 -680 29485 -650
rect 29515 -680 29525 -650
rect 29475 -690 29525 -680
rect 29560 -500 29610 -490
rect 29560 -530 29570 -500
rect 29600 -530 29610 -500
rect 29560 -550 29610 -530
rect 29560 -580 29570 -550
rect 29600 -580 29610 -550
rect 29560 -600 29610 -580
rect 29560 -630 29570 -600
rect 29600 -630 29610 -600
rect 29560 -650 29610 -630
rect 29560 -680 29570 -650
rect 29600 -680 29610 -650
rect 29560 -690 29610 -680
rect 29645 -500 29695 -490
rect 29645 -530 29655 -500
rect 29685 -530 29695 -500
rect 29645 -550 29695 -530
rect 29645 -580 29655 -550
rect 29685 -580 29695 -550
rect 29645 -600 29695 -580
rect 29645 -630 29655 -600
rect 29685 -630 29695 -600
rect 29645 -650 29695 -630
rect 29645 -680 29655 -650
rect 29685 -680 29695 -650
rect 29645 -690 29695 -680
rect 29730 -500 29780 -490
rect 29730 -530 29740 -500
rect 29770 -530 29780 -500
rect 29730 -550 29780 -530
rect 29730 -580 29740 -550
rect 29770 -580 29780 -550
rect 29730 -600 29780 -580
rect 29730 -630 29740 -600
rect 29770 -630 29780 -600
rect 29730 -650 29780 -630
rect 29730 -680 29740 -650
rect 29770 -680 29780 -650
rect 29730 -690 29780 -680
rect 29815 -500 29865 -490
rect 29815 -530 29825 -500
rect 29855 -530 29865 -500
rect 29815 -550 29865 -530
rect 29815 -580 29825 -550
rect 29855 -580 29865 -550
rect 29815 -600 29865 -580
rect 29815 -630 29825 -600
rect 29855 -630 29865 -600
rect 29815 -650 29865 -630
rect 29815 -680 29825 -650
rect 29855 -680 29865 -650
rect 29815 -690 29865 -680
rect 29900 -500 29950 -490
rect 29900 -530 29910 -500
rect 29940 -530 29950 -500
rect 29900 -550 29950 -530
rect 29900 -580 29910 -550
rect 29940 -580 29950 -550
rect 29900 -600 29950 -580
rect 29900 -630 29910 -600
rect 29940 -630 29950 -600
rect 29900 -650 29950 -630
rect 29900 -680 29910 -650
rect 29940 -680 29950 -650
rect 29900 -690 29950 -680
rect 29985 -500 30035 -490
rect 29985 -530 29995 -500
rect 30025 -530 30035 -500
rect 29985 -550 30035 -530
rect 29985 -580 29995 -550
rect 30025 -580 30035 -550
rect 29985 -600 30035 -580
rect 29985 -630 29995 -600
rect 30025 -630 30035 -600
rect 29985 -650 30035 -630
rect 29985 -680 29995 -650
rect 30025 -680 30035 -650
rect 29985 -690 30035 -680
rect 30070 -500 30120 -490
rect 30070 -530 30080 -500
rect 30110 -530 30120 -500
rect 30070 -550 30120 -530
rect 30070 -580 30080 -550
rect 30110 -580 30120 -550
rect 30070 -600 30120 -580
rect 30070 -630 30080 -600
rect 30110 -630 30120 -600
rect 30070 -650 30120 -630
rect 30070 -680 30080 -650
rect 30110 -680 30120 -650
rect 30070 -690 30120 -680
rect 30155 -500 30205 -490
rect 30155 -530 30165 -500
rect 30195 -530 30205 -500
rect 30155 -550 30205 -530
rect 30155 -580 30165 -550
rect 30195 -580 30205 -550
rect 30155 -600 30205 -580
rect 30155 -630 30165 -600
rect 30195 -630 30205 -600
rect 30155 -650 30205 -630
rect 30155 -680 30165 -650
rect 30195 -680 30205 -650
rect 30155 -690 30205 -680
rect 30240 -500 30290 -490
rect 30240 -530 30250 -500
rect 30280 -530 30290 -500
rect 30240 -550 30290 -530
rect 30240 -580 30250 -550
rect 30280 -580 30290 -550
rect 30240 -600 30290 -580
rect 30240 -630 30250 -600
rect 30280 -630 30290 -600
rect 30240 -650 30290 -630
rect 30240 -680 30250 -650
rect 30280 -680 30290 -650
rect 30240 -690 30290 -680
rect 30325 -500 30375 -490
rect 30325 -530 30335 -500
rect 30365 -530 30375 -500
rect 30325 -550 30375 -530
rect 30325 -580 30335 -550
rect 30365 -580 30375 -550
rect 30325 -600 30375 -580
rect 30325 -630 30335 -600
rect 30365 -630 30375 -600
rect 30325 -650 30375 -630
rect 30325 -680 30335 -650
rect 30365 -680 30375 -650
rect 30325 -690 30375 -680
rect 30410 -500 30460 -490
rect 30410 -530 30420 -500
rect 30450 -530 30460 -500
rect 30410 -550 30460 -530
rect 30410 -580 30420 -550
rect 30450 -580 30460 -550
rect 30410 -600 30460 -580
rect 30410 -630 30420 -600
rect 30450 -630 30460 -600
rect 30410 -650 30460 -630
rect 30410 -680 30420 -650
rect 30450 -680 30460 -650
rect 30410 -690 30460 -680
rect 30495 -500 30545 -490
rect 30495 -530 30505 -500
rect 30535 -530 30545 -500
rect 30495 -550 30545 -530
rect 30495 -580 30505 -550
rect 30535 -580 30545 -550
rect 30495 -600 30545 -580
rect 30495 -630 30505 -600
rect 30535 -630 30545 -600
rect 30495 -650 30545 -630
rect 30495 -680 30505 -650
rect 30535 -680 30545 -650
rect 30495 -690 30545 -680
rect 30580 -500 30630 -490
rect 30580 -530 30590 -500
rect 30620 -530 30630 -500
rect 30580 -550 30630 -530
rect 30580 -580 30590 -550
rect 30620 -580 30630 -550
rect 30580 -600 30630 -580
rect 30580 -630 30590 -600
rect 30620 -630 30630 -600
rect 30580 -650 30630 -630
rect 30580 -680 30590 -650
rect 30620 -680 30630 -650
rect 30580 -690 30630 -680
rect 30665 -500 30715 -490
rect 30665 -530 30675 -500
rect 30705 -530 30715 -500
rect 30665 -550 30715 -530
rect 30665 -580 30675 -550
rect 30705 -580 30715 -550
rect 30665 -600 30715 -580
rect 30665 -630 30675 -600
rect 30705 -630 30715 -600
rect 30665 -650 30715 -630
rect 30665 -680 30675 -650
rect 30705 -680 30715 -650
rect 30665 -690 30715 -680
rect 30750 -500 30800 -490
rect 30750 -530 30760 -500
rect 30790 -530 30800 -500
rect 30750 -550 30800 -530
rect 30750 -580 30760 -550
rect 30790 -580 30800 -550
rect 30750 -600 30800 -580
rect 30750 -630 30760 -600
rect 30790 -630 30800 -600
rect 30750 -650 30800 -630
rect 30750 -680 30760 -650
rect 30790 -680 30800 -650
rect 30750 -690 30800 -680
rect 30835 -500 30885 -490
rect 30835 -530 30845 -500
rect 30875 -530 30885 -500
rect 30835 -550 30885 -530
rect 30835 -580 30845 -550
rect 30875 -580 30885 -550
rect 30835 -600 30885 -580
rect 30835 -630 30845 -600
rect 30875 -630 30885 -600
rect 30835 -650 30885 -630
rect 30835 -680 30845 -650
rect 30875 -680 30885 -650
rect 30835 -690 30885 -680
rect 30920 -500 30970 -490
rect 30920 -530 30930 -500
rect 30960 -530 30970 -500
rect 30920 -550 30970 -530
rect 30920 -580 30930 -550
rect 30960 -580 30970 -550
rect 30920 -600 30970 -580
rect 30920 -630 30930 -600
rect 30960 -630 30970 -600
rect 30920 -650 30970 -630
rect 30920 -680 30930 -650
rect 30960 -680 30970 -650
rect 30920 -690 30970 -680
rect 31005 -500 31055 -490
rect 31005 -530 31015 -500
rect 31045 -530 31055 -500
rect 31005 -550 31055 -530
rect 31005 -580 31015 -550
rect 31045 -580 31055 -550
rect 31005 -600 31055 -580
rect 31005 -630 31015 -600
rect 31045 -630 31055 -600
rect 31005 -650 31055 -630
rect 31005 -680 31015 -650
rect 31045 -680 31055 -650
rect 31005 -690 31055 -680
rect 31090 -500 31140 -490
rect 31090 -530 31100 -500
rect 31130 -530 31140 -500
rect 31090 -550 31140 -530
rect 31090 -580 31100 -550
rect 31130 -580 31140 -550
rect 31090 -600 31140 -580
rect 31090 -630 31100 -600
rect 31130 -630 31140 -600
rect 31090 -650 31140 -630
rect 31090 -680 31100 -650
rect 31130 -680 31140 -650
rect 31090 -690 31140 -680
rect 31175 -500 31225 -490
rect 31175 -530 31185 -500
rect 31215 -530 31225 -500
rect 31175 -550 31225 -530
rect 31175 -580 31185 -550
rect 31215 -580 31225 -550
rect 31175 -600 31225 -580
rect 31175 -630 31185 -600
rect 31215 -630 31225 -600
rect 31175 -650 31225 -630
rect 31175 -680 31185 -650
rect 31215 -680 31225 -650
rect 31175 -690 31225 -680
rect 31260 -500 31310 -490
rect 31260 -530 31270 -500
rect 31300 -530 31310 -500
rect 31260 -550 31310 -530
rect 31260 -580 31270 -550
rect 31300 -580 31310 -550
rect 31260 -600 31310 -580
rect 31260 -630 31270 -600
rect 31300 -630 31310 -600
rect 31260 -650 31310 -630
rect 31260 -680 31270 -650
rect 31300 -680 31310 -650
rect 31260 -690 31310 -680
rect 31345 -500 31395 -490
rect 31345 -530 31355 -500
rect 31385 -530 31395 -500
rect 31345 -550 31395 -530
rect 31345 -580 31355 -550
rect 31385 -580 31395 -550
rect 31345 -600 31395 -580
rect 31345 -630 31355 -600
rect 31385 -630 31395 -600
rect 31345 -650 31395 -630
rect 31345 -680 31355 -650
rect 31385 -680 31395 -650
rect 31345 -690 31395 -680
rect 31430 -500 31480 -490
rect 31430 -530 31440 -500
rect 31470 -530 31480 -500
rect 31430 -550 31480 -530
rect 31430 -580 31440 -550
rect 31470 -580 31480 -550
rect 31430 -600 31480 -580
rect 31430 -630 31440 -600
rect 31470 -630 31480 -600
rect 31430 -650 31480 -630
rect 31430 -680 31440 -650
rect 31470 -680 31480 -650
rect 31430 -690 31480 -680
rect 31515 -500 31565 -490
rect 31515 -530 31525 -500
rect 31555 -530 31565 -500
rect 31515 -550 31565 -530
rect 31515 -580 31525 -550
rect 31555 -580 31565 -550
rect 31515 -600 31565 -580
rect 31515 -630 31525 -600
rect 31555 -630 31565 -600
rect 31515 -650 31565 -630
rect 31515 -680 31525 -650
rect 31555 -680 31565 -650
rect 31515 -690 31565 -680
rect 31600 -500 31650 -490
rect 31600 -530 31610 -500
rect 31640 -530 31650 -500
rect 31600 -550 31650 -530
rect 31600 -580 31610 -550
rect 31640 -580 31650 -550
rect 31600 -600 31650 -580
rect 31600 -630 31610 -600
rect 31640 -630 31650 -600
rect 31600 -650 31650 -630
rect 31600 -680 31610 -650
rect 31640 -680 31650 -650
rect 31600 -690 31650 -680
rect 31685 -500 31735 -490
rect 31685 -530 31695 -500
rect 31725 -530 31735 -500
rect 31685 -550 31735 -530
rect 31685 -580 31695 -550
rect 31725 -580 31735 -550
rect 31685 -600 31735 -580
rect 31685 -630 31695 -600
rect 31725 -630 31735 -600
rect 31685 -650 31735 -630
rect 31685 -680 31695 -650
rect 31725 -680 31735 -650
rect 31685 -690 31735 -680
rect 31770 -500 31820 -490
rect 31770 -530 31780 -500
rect 31810 -530 31820 -500
rect 31770 -550 31820 -530
rect 31770 -580 31780 -550
rect 31810 -580 31820 -550
rect 31770 -600 31820 -580
rect 31770 -630 31780 -600
rect 31810 -630 31820 -600
rect 31770 -650 31820 -630
rect 31770 -680 31780 -650
rect 31810 -680 31820 -650
rect 31770 -690 31820 -680
rect 31855 -500 31905 -490
rect 31855 -530 31865 -500
rect 31895 -530 31905 -500
rect 31855 -550 31905 -530
rect 31855 -580 31865 -550
rect 31895 -580 31905 -550
rect 31855 -600 31905 -580
rect 31855 -630 31865 -600
rect 31895 -630 31905 -600
rect 31855 -650 31905 -630
rect 31855 -680 31865 -650
rect 31895 -680 31905 -650
rect 31855 -690 31905 -680
rect 31940 -500 31990 -490
rect 31940 -530 31950 -500
rect 31980 -530 31990 -500
rect 31940 -550 31990 -530
rect 31940 -580 31950 -550
rect 31980 -580 31990 -550
rect 31940 -600 31990 -580
rect 31940 -630 31950 -600
rect 31980 -630 31990 -600
rect 31940 -650 31990 -630
rect 31940 -680 31950 -650
rect 31980 -680 31990 -650
rect 31940 -690 31990 -680
rect 32025 -500 32075 -490
rect 32025 -530 32035 -500
rect 32065 -530 32075 -500
rect 32025 -550 32075 -530
rect 32025 -580 32035 -550
rect 32065 -580 32075 -550
rect 32025 -600 32075 -580
rect 32025 -630 32035 -600
rect 32065 -630 32075 -600
rect 32025 -650 32075 -630
rect 32025 -680 32035 -650
rect 32065 -680 32075 -650
rect 32025 -690 32075 -680
rect 32110 -500 32160 -490
rect 32110 -530 32120 -500
rect 32150 -530 32160 -500
rect 32110 -550 32160 -530
rect 32110 -580 32120 -550
rect 32150 -580 32160 -550
rect 32110 -600 32160 -580
rect 32110 -630 32120 -600
rect 32150 -630 32160 -600
rect 32110 -650 32160 -630
rect 32110 -680 32120 -650
rect 32150 -680 32160 -650
rect 32110 -690 32160 -680
rect 32195 -500 32245 -490
rect 32195 -530 32205 -500
rect 32235 -530 32245 -500
rect 32195 -550 32245 -530
rect 32195 -580 32205 -550
rect 32235 -580 32245 -550
rect 32195 -600 32245 -580
rect 32195 -630 32205 -600
rect 32235 -630 32245 -600
rect 32195 -650 32245 -630
rect 32195 -680 32205 -650
rect 32235 -680 32245 -650
rect 32195 -690 32245 -680
rect 32280 -500 32330 -490
rect 32280 -530 32290 -500
rect 32320 -530 32330 -500
rect 32280 -550 32330 -530
rect 32280 -580 32290 -550
rect 32320 -580 32330 -550
rect 32280 -600 32330 -580
rect 32280 -630 32290 -600
rect 32320 -630 32330 -600
rect 32280 -650 32330 -630
rect 32280 -680 32290 -650
rect 32320 -680 32330 -650
rect 32280 -690 32330 -680
rect 32365 -500 32415 -490
rect 32365 -530 32375 -500
rect 32405 -530 32415 -500
rect 32365 -550 32415 -530
rect 32365 -580 32375 -550
rect 32405 -580 32415 -550
rect 32365 -600 32415 -580
rect 32365 -630 32375 -600
rect 32405 -630 32415 -600
rect 32365 -650 32415 -630
rect 32365 -680 32375 -650
rect 32405 -680 32415 -650
rect 32365 -690 32415 -680
rect 32450 -500 32500 -490
rect 32450 -530 32460 -500
rect 32490 -530 32500 -500
rect 32450 -550 32500 -530
rect 32450 -580 32460 -550
rect 32490 -580 32500 -550
rect 32450 -600 32500 -580
rect 32450 -630 32460 -600
rect 32490 -630 32500 -600
rect 32450 -650 32500 -630
rect 32450 -680 32460 -650
rect 32490 -680 32500 -650
rect 32450 -690 32500 -680
rect 32535 -500 32585 -490
rect 32535 -530 32545 -500
rect 32575 -530 32585 -500
rect 32535 -550 32585 -530
rect 32535 -580 32545 -550
rect 32575 -580 32585 -550
rect 32535 -600 32585 -580
rect 32535 -630 32545 -600
rect 32575 -630 32585 -600
rect 32535 -650 32585 -630
rect 32535 -680 32545 -650
rect 32575 -680 32585 -650
rect 32535 -690 32585 -680
rect 32620 -500 32670 -490
rect 32620 -530 32630 -500
rect 32660 -530 32670 -500
rect 32620 -550 32670 -530
rect 32620 -580 32630 -550
rect 32660 -580 32670 -550
rect 32620 -600 32670 -580
rect 32620 -630 32630 -600
rect 32660 -630 32670 -600
rect 32620 -650 32670 -630
rect 32620 -680 32630 -650
rect 32660 -680 32670 -650
rect 32620 -690 32670 -680
rect 32705 -500 32755 -490
rect 32705 -530 32715 -500
rect 32745 -530 32755 -500
rect 32705 -550 32755 -530
rect 32705 -580 32715 -550
rect 32745 -580 32755 -550
rect 32705 -600 32755 -580
rect 32705 -630 32715 -600
rect 32745 -630 32755 -600
rect 32705 -650 32755 -630
rect 32705 -680 32715 -650
rect 32745 -680 32755 -650
rect 32705 -690 32755 -680
rect 32790 -500 32840 -490
rect 32790 -530 32800 -500
rect 32830 -530 32840 -500
rect 32790 -550 32840 -530
rect 32790 -580 32800 -550
rect 32830 -580 32840 -550
rect 32790 -600 32840 -580
rect 32790 -630 32800 -600
rect 32830 -630 32840 -600
rect 32790 -650 32840 -630
rect 32790 -680 32800 -650
rect 32830 -680 32840 -650
rect 32790 -690 32840 -680
rect 32875 -500 32925 -490
rect 32875 -530 32885 -500
rect 32915 -530 32925 -500
rect 32875 -550 32925 -530
rect 32875 -580 32885 -550
rect 32915 -580 32925 -550
rect 32875 -600 32925 -580
rect 32875 -630 32885 -600
rect 32915 -630 32925 -600
rect 32875 -650 32925 -630
rect 32875 -680 32885 -650
rect 32915 -680 32925 -650
rect 32875 -690 32925 -680
rect 32960 -500 33010 -490
rect 32960 -530 32970 -500
rect 33000 -530 33010 -500
rect 32960 -550 33010 -530
rect 32960 -580 32970 -550
rect 33000 -580 33010 -550
rect 32960 -600 33010 -580
rect 32960 -630 32970 -600
rect 33000 -630 33010 -600
rect 32960 -650 33010 -630
rect 32960 -680 32970 -650
rect 33000 -680 33010 -650
rect 32960 -690 33010 -680
rect 33045 -500 33095 -490
rect 33045 -530 33055 -500
rect 33085 -530 33095 -500
rect 33045 -550 33095 -530
rect 33045 -580 33055 -550
rect 33085 -580 33095 -550
rect 33045 -600 33095 -580
rect 33045 -630 33055 -600
rect 33085 -630 33095 -600
rect 33045 -650 33095 -630
rect 33045 -680 33055 -650
rect 33085 -680 33095 -650
rect 33045 -690 33095 -680
rect 33130 -500 33180 -490
rect 33130 -530 33140 -500
rect 33170 -530 33180 -500
rect 33130 -550 33180 -530
rect 33130 -580 33140 -550
rect 33170 -580 33180 -550
rect 33130 -600 33180 -580
rect 33130 -630 33140 -600
rect 33170 -630 33180 -600
rect 33130 -650 33180 -630
rect 33130 -680 33140 -650
rect 33170 -680 33180 -650
rect 33130 -690 33180 -680
rect 33215 -500 33265 -490
rect 33215 -530 33225 -500
rect 33255 -530 33265 -500
rect 33215 -550 33265 -530
rect 33215 -580 33225 -550
rect 33255 -580 33265 -550
rect 33215 -600 33265 -580
rect 33215 -630 33225 -600
rect 33255 -630 33265 -600
rect 33215 -650 33265 -630
rect 33215 -680 33225 -650
rect 33255 -680 33265 -650
rect 33215 -690 33265 -680
rect 33300 -500 33350 -490
rect 33300 -530 33310 -500
rect 33340 -530 33350 -500
rect 33300 -550 33350 -530
rect 33300 -580 33310 -550
rect 33340 -580 33350 -550
rect 33300 -600 33350 -580
rect 33300 -630 33310 -600
rect 33340 -630 33350 -600
rect 33300 -650 33350 -630
rect 33300 -680 33310 -650
rect 33340 -680 33350 -650
rect 33300 -690 33350 -680
rect 33385 -500 33435 -490
rect 33385 -530 33395 -500
rect 33425 -530 33435 -500
rect 33385 -550 33435 -530
rect 33385 -580 33395 -550
rect 33425 -580 33435 -550
rect 33385 -600 33435 -580
rect 33385 -630 33395 -600
rect 33425 -630 33435 -600
rect 33385 -650 33435 -630
rect 33385 -680 33395 -650
rect 33425 -680 33435 -650
rect 33385 -690 33435 -680
rect 33470 -500 33520 -490
rect 33470 -530 33480 -500
rect 33510 -530 33520 -500
rect 33470 -550 33520 -530
rect 33470 -580 33480 -550
rect 33510 -580 33520 -550
rect 33470 -600 33520 -580
rect 33470 -630 33480 -600
rect 33510 -630 33520 -600
rect 33470 -650 33520 -630
rect 33470 -680 33480 -650
rect 33510 -680 33520 -650
rect 33470 -690 33520 -680
rect 33555 -500 33605 -490
rect 33555 -530 33565 -500
rect 33595 -530 33605 -500
rect 33555 -550 33605 -530
rect 33555 -580 33565 -550
rect 33595 -580 33605 -550
rect 33555 -600 33605 -580
rect 33555 -630 33565 -600
rect 33595 -630 33605 -600
rect 33555 -650 33605 -630
rect 33555 -680 33565 -650
rect 33595 -680 33605 -650
rect 33555 -690 33605 -680
rect 33640 -500 33690 -490
rect 33640 -530 33650 -500
rect 33680 -530 33690 -500
rect 33640 -550 33690 -530
rect 33640 -580 33650 -550
rect 33680 -580 33690 -550
rect 33640 -600 33690 -580
rect 33640 -630 33650 -600
rect 33680 -630 33690 -600
rect 33640 -650 33690 -630
rect 33640 -680 33650 -650
rect 33680 -680 33690 -650
rect 33640 -690 33690 -680
rect 33725 -500 33775 -490
rect 33725 -530 33735 -500
rect 33765 -530 33775 -500
rect 33725 -550 33775 -530
rect 33725 -580 33735 -550
rect 33765 -580 33775 -550
rect 33725 -600 33775 -580
rect 33725 -630 33735 -600
rect 33765 -630 33775 -600
rect 33725 -650 33775 -630
rect 33725 -680 33735 -650
rect 33765 -680 33775 -650
rect 33725 -690 33775 -680
rect 33810 -500 33860 -490
rect 33810 -530 33820 -500
rect 33850 -530 33860 -500
rect 33810 -550 33860 -530
rect 33810 -580 33820 -550
rect 33850 -580 33860 -550
rect 33810 -600 33860 -580
rect 33810 -630 33820 -600
rect 33850 -630 33860 -600
rect 33810 -650 33860 -630
rect 33810 -680 33820 -650
rect 33850 -680 33860 -650
rect 33810 -690 33860 -680
rect 33895 -500 33945 -490
rect 33895 -530 33905 -500
rect 33935 -530 33945 -500
rect 33895 -550 33945 -530
rect 33895 -580 33905 -550
rect 33935 -580 33945 -550
rect 33895 -600 33945 -580
rect 33895 -630 33905 -600
rect 33935 -630 33945 -600
rect 33895 -650 33945 -630
rect 33895 -680 33905 -650
rect 33935 -680 33945 -650
rect 33895 -690 33945 -680
rect 33980 -500 34030 -490
rect 33980 -530 33990 -500
rect 34020 -530 34030 -500
rect 33980 -550 34030 -530
rect 33980 -580 33990 -550
rect 34020 -580 34030 -550
rect 33980 -600 34030 -580
rect 33980 -630 33990 -600
rect 34020 -630 34030 -600
rect 33980 -650 34030 -630
rect 33980 -680 33990 -650
rect 34020 -680 34030 -650
rect 33980 -690 34030 -680
rect 34065 -500 34115 -490
rect 34065 -530 34075 -500
rect 34105 -530 34115 -500
rect 34065 -550 34115 -530
rect 34065 -580 34075 -550
rect 34105 -580 34115 -550
rect 34065 -600 34115 -580
rect 34065 -630 34075 -600
rect 34105 -630 34115 -600
rect 34065 -650 34115 -630
rect 34065 -680 34075 -650
rect 34105 -680 34115 -650
rect 34065 -690 34115 -680
rect 34150 -500 34200 -490
rect 34150 -530 34160 -500
rect 34190 -530 34200 -500
rect 34150 -550 34200 -530
rect 34150 -580 34160 -550
rect 34190 -580 34200 -550
rect 34150 -600 34200 -580
rect 34150 -630 34160 -600
rect 34190 -630 34200 -600
rect 34150 -650 34200 -630
rect 34150 -680 34160 -650
rect 34190 -680 34200 -650
rect 34150 -690 34200 -680
rect 34235 -500 34285 -490
rect 34235 -530 34245 -500
rect 34275 -530 34285 -500
rect 34235 -550 34285 -530
rect 34235 -580 34245 -550
rect 34275 -580 34285 -550
rect 34235 -600 34285 -580
rect 34235 -630 34245 -600
rect 34275 -630 34285 -600
rect 34235 -650 34285 -630
rect 34235 -680 34245 -650
rect 34275 -680 34285 -650
rect 34235 -690 34285 -680
rect 34320 -500 34370 -490
rect 34320 -530 34330 -500
rect 34360 -530 34370 -500
rect 34320 -550 34370 -530
rect 34320 -580 34330 -550
rect 34360 -580 34370 -550
rect 34320 -600 34370 -580
rect 34320 -630 34330 -600
rect 34360 -630 34370 -600
rect 34320 -650 34370 -630
rect 34320 -680 34330 -650
rect 34360 -680 34370 -650
rect 34320 -690 34370 -680
rect 34405 -500 34455 -490
rect 34405 -530 34415 -500
rect 34445 -530 34455 -500
rect 34405 -550 34455 -530
rect 34405 -580 34415 -550
rect 34445 -580 34455 -550
rect 34405 -600 34455 -580
rect 34405 -630 34415 -600
rect 34445 -630 34455 -600
rect 34405 -650 34455 -630
rect 34405 -680 34415 -650
rect 34445 -680 34455 -650
rect 34405 -690 34455 -680
rect 34490 -500 34540 -490
rect 34490 -530 34500 -500
rect 34530 -530 34540 -500
rect 34490 -550 34540 -530
rect 34490 -580 34500 -550
rect 34530 -580 34540 -550
rect 34490 -600 34540 -580
rect 34490 -630 34500 -600
rect 34530 -630 34540 -600
rect 34490 -650 34540 -630
rect 34490 -680 34500 -650
rect 34530 -680 34540 -650
rect 34490 -690 34540 -680
rect 34575 -500 34625 -490
rect 34575 -530 34585 -500
rect 34615 -530 34625 -500
rect 34575 -550 34625 -530
rect 34575 -580 34585 -550
rect 34615 -580 34625 -550
rect 34575 -600 34625 -580
rect 34575 -630 34585 -600
rect 34615 -630 34625 -600
rect 34575 -650 34625 -630
rect 34575 -680 34585 -650
rect 34615 -680 34625 -650
rect 34575 -690 34625 -680
rect 34660 -500 34710 -490
rect 34660 -530 34670 -500
rect 34700 -530 34710 -500
rect 34660 -550 34710 -530
rect 34660 -580 34670 -550
rect 34700 -580 34710 -550
rect 34660 -600 34710 -580
rect 34660 -630 34670 -600
rect 34700 -630 34710 -600
rect 34660 -650 34710 -630
rect 34660 -680 34670 -650
rect 34700 -680 34710 -650
rect 34660 -690 34710 -680
rect 34745 -500 34795 -490
rect 34745 -530 34755 -500
rect 34785 -530 34795 -500
rect 34745 -550 34795 -530
rect 34745 -580 34755 -550
rect 34785 -580 34795 -550
rect 34745 -600 34795 -580
rect 34745 -630 34755 -600
rect 34785 -630 34795 -600
rect 34745 -650 34795 -630
rect 34745 -680 34755 -650
rect 34785 -680 34795 -650
rect 34745 -690 34795 -680
rect 34830 -500 34880 -490
rect 34830 -530 34840 -500
rect 34870 -530 34880 -500
rect 34830 -550 34880 -530
rect 34830 -580 34840 -550
rect 34870 -580 34880 -550
rect 34830 -600 34880 -580
rect 34830 -630 34840 -600
rect 34870 -630 34880 -600
rect 34830 -650 34880 -630
rect 34830 -680 34840 -650
rect 34870 -680 34880 -650
rect 34830 -690 34880 -680
rect 34915 -500 34965 -490
rect 34915 -530 34925 -500
rect 34955 -530 34965 -500
rect 34915 -550 34965 -530
rect 34915 -580 34925 -550
rect 34955 -580 34965 -550
rect 34915 -600 34965 -580
rect 34915 -630 34925 -600
rect 34955 -630 34965 -600
rect 34915 -650 34965 -630
rect 34915 -680 34925 -650
rect 34955 -680 34965 -650
rect 34915 -690 34965 -680
rect 35000 -500 35050 -490
rect 35000 -530 35010 -500
rect 35040 -530 35050 -500
rect 35000 -550 35050 -530
rect 35000 -580 35010 -550
rect 35040 -580 35050 -550
rect 35000 -600 35050 -580
rect 35000 -630 35010 -600
rect 35040 -630 35050 -600
rect 35000 -650 35050 -630
rect 35000 -680 35010 -650
rect 35040 -680 35050 -650
rect 35000 -690 35050 -680
rect 35085 -500 35135 -490
rect 35085 -530 35095 -500
rect 35125 -530 35135 -500
rect 35085 -550 35135 -530
rect 35085 -580 35095 -550
rect 35125 -580 35135 -550
rect 35085 -600 35135 -580
rect 35085 -630 35095 -600
rect 35125 -630 35135 -600
rect 35085 -650 35135 -630
rect 35085 -680 35095 -650
rect 35125 -680 35135 -650
rect 35085 -690 35135 -680
rect 35170 -500 35220 -490
rect 35170 -530 35180 -500
rect 35210 -530 35220 -500
rect 35170 -550 35220 -530
rect 35170 -580 35180 -550
rect 35210 -580 35220 -550
rect 35170 -600 35220 -580
rect 35170 -630 35180 -600
rect 35210 -630 35220 -600
rect 35170 -650 35220 -630
rect 35170 -680 35180 -650
rect 35210 -680 35220 -650
rect 35170 -690 35220 -680
rect 35255 -500 35305 -490
rect 35255 -530 35265 -500
rect 35295 -530 35305 -500
rect 35255 -550 35305 -530
rect 35255 -580 35265 -550
rect 35295 -580 35305 -550
rect 35255 -600 35305 -580
rect 35255 -630 35265 -600
rect 35295 -630 35305 -600
rect 35255 -650 35305 -630
rect 35255 -680 35265 -650
rect 35295 -680 35305 -650
rect 35255 -690 35305 -680
rect 35340 -500 35390 -490
rect 35340 -530 35350 -500
rect 35380 -530 35390 -500
rect 35340 -550 35390 -530
rect 35340 -580 35350 -550
rect 35380 -580 35390 -550
rect 35340 -600 35390 -580
rect 35340 -630 35350 -600
rect 35380 -630 35390 -600
rect 35340 -650 35390 -630
rect 35340 -680 35350 -650
rect 35380 -680 35390 -650
rect 35340 -690 35390 -680
rect 35425 -500 35475 -490
rect 35425 -530 35435 -500
rect 35465 -530 35475 -500
rect 35425 -550 35475 -530
rect 35425 -580 35435 -550
rect 35465 -580 35475 -550
rect 35425 -600 35475 -580
rect 35425 -630 35435 -600
rect 35465 -630 35475 -600
rect 35425 -650 35475 -630
rect 35425 -680 35435 -650
rect 35465 -680 35475 -650
rect 35425 -690 35475 -680
rect 35510 -500 35560 -490
rect 35510 -530 35520 -500
rect 35550 -530 35560 -500
rect 35510 -550 35560 -530
rect 35510 -580 35520 -550
rect 35550 -580 35560 -550
rect 35510 -600 35560 -580
rect 35510 -630 35520 -600
rect 35550 -630 35560 -600
rect 35510 -650 35560 -630
rect 35510 -680 35520 -650
rect 35550 -680 35560 -650
rect 35510 -690 35560 -680
rect 35595 -500 35645 -490
rect 35595 -530 35605 -500
rect 35635 -530 35645 -500
rect 35595 -550 35645 -530
rect 35595 -580 35605 -550
rect 35635 -580 35645 -550
rect 35595 -600 35645 -580
rect 35595 -630 35605 -600
rect 35635 -630 35645 -600
rect 35595 -650 35645 -630
rect 35595 -680 35605 -650
rect 35635 -680 35645 -650
rect 35595 -690 35645 -680
rect 35680 -500 35730 -490
rect 35680 -530 35690 -500
rect 35720 -530 35730 -500
rect 35680 -550 35730 -530
rect 35680 -580 35690 -550
rect 35720 -580 35730 -550
rect 35680 -600 35730 -580
rect 35680 -630 35690 -600
rect 35720 -630 35730 -600
rect 35680 -650 35730 -630
rect 35680 -680 35690 -650
rect 35720 -680 35730 -650
rect 35680 -690 35730 -680
rect 35765 -500 35815 -490
rect 35765 -530 35775 -500
rect 35805 -530 35815 -500
rect 35765 -550 35815 -530
rect 35765 -580 35775 -550
rect 35805 -580 35815 -550
rect 35765 -600 35815 -580
rect 35765 -630 35775 -600
rect 35805 -630 35815 -600
rect 35765 -650 35815 -630
rect 35765 -680 35775 -650
rect 35805 -680 35815 -650
rect 35765 -690 35815 -680
rect 35850 -500 35900 -490
rect 35850 -530 35860 -500
rect 35890 -530 35900 -500
rect 35850 -550 35900 -530
rect 35850 -580 35860 -550
rect 35890 -580 35900 -550
rect 35850 -600 35900 -580
rect 35850 -630 35860 -600
rect 35890 -630 35900 -600
rect 35850 -650 35900 -630
rect 35850 -680 35860 -650
rect 35890 -680 35900 -650
rect 35850 -690 35900 -680
rect 35935 -500 35985 -490
rect 35935 -530 35945 -500
rect 35975 -530 35985 -500
rect 35935 -550 35985 -530
rect 35935 -580 35945 -550
rect 35975 -580 35985 -550
rect 35935 -600 35985 -580
rect 35935 -630 35945 -600
rect 35975 -630 35985 -600
rect 35935 -650 35985 -630
rect 35935 -680 35945 -650
rect 35975 -680 35985 -650
rect 35935 -690 35985 -680
rect 36020 -500 36070 -490
rect 36020 -530 36030 -500
rect 36060 -530 36070 -500
rect 36020 -550 36070 -530
rect 36020 -580 36030 -550
rect 36060 -580 36070 -550
rect 36020 -600 36070 -580
rect 36020 -630 36030 -600
rect 36060 -630 36070 -600
rect 36020 -650 36070 -630
rect 36020 -680 36030 -650
rect 36060 -680 36070 -650
rect 36020 -690 36070 -680
rect 36105 -500 36155 -490
rect 36105 -530 36115 -500
rect 36145 -530 36155 -500
rect 36105 -550 36155 -530
rect 36105 -580 36115 -550
rect 36145 -580 36155 -550
rect 36105 -600 36155 -580
rect 36105 -630 36115 -600
rect 36145 -630 36155 -600
rect 36105 -650 36155 -630
rect 36105 -680 36115 -650
rect 36145 -680 36155 -650
rect 36105 -690 36155 -680
rect 36190 -500 36240 -490
rect 36190 -530 36200 -500
rect 36230 -530 36240 -500
rect 36190 -550 36240 -530
rect 36190 -580 36200 -550
rect 36230 -580 36240 -550
rect 36190 -600 36240 -580
rect 36190 -630 36200 -600
rect 36230 -630 36240 -600
rect 36190 -650 36240 -630
rect 36190 -680 36200 -650
rect 36230 -680 36240 -650
rect 36190 -690 36240 -680
rect 36275 -500 36325 -490
rect 36275 -530 36285 -500
rect 36315 -530 36325 -500
rect 36275 -550 36325 -530
rect 36275 -580 36285 -550
rect 36315 -580 36325 -550
rect 36275 -600 36325 -580
rect 36275 -630 36285 -600
rect 36315 -630 36325 -600
rect 36275 -650 36325 -630
rect 36275 -680 36285 -650
rect 36315 -680 36325 -650
rect 36275 -690 36325 -680
rect 36360 -500 36410 -490
rect 36360 -530 36370 -500
rect 36400 -530 36410 -500
rect 36360 -550 36410 -530
rect 36360 -580 36370 -550
rect 36400 -580 36410 -550
rect 36360 -600 36410 -580
rect 36360 -630 36370 -600
rect 36400 -630 36410 -600
rect 36360 -650 36410 -630
rect 36360 -680 36370 -650
rect 36400 -680 36410 -650
rect 36360 -690 36410 -680
rect 36445 -500 36495 -490
rect 36445 -530 36455 -500
rect 36485 -530 36495 -500
rect 36445 -550 36495 -530
rect 36445 -580 36455 -550
rect 36485 -580 36495 -550
rect 36445 -600 36495 -580
rect 36445 -630 36455 -600
rect 36485 -630 36495 -600
rect 36445 -650 36495 -630
rect 36445 -680 36455 -650
rect 36485 -680 36495 -650
rect 36445 -690 36495 -680
rect 36530 -500 36580 -490
rect 36530 -530 36540 -500
rect 36570 -530 36580 -500
rect 36530 -550 36580 -530
rect 36530 -580 36540 -550
rect 36570 -580 36580 -550
rect 36530 -600 36580 -580
rect 36530 -630 36540 -600
rect 36570 -630 36580 -600
rect 36530 -650 36580 -630
rect 36530 -680 36540 -650
rect 36570 -680 36580 -650
rect 36530 -690 36580 -680
rect 36615 -500 36665 -490
rect 36615 -530 36625 -500
rect 36655 -530 36665 -500
rect 36615 -550 36665 -530
rect 36615 -580 36625 -550
rect 36655 -580 36665 -550
rect 36615 -600 36665 -580
rect 36615 -630 36625 -600
rect 36655 -630 36665 -600
rect 36615 -650 36665 -630
rect 36615 -680 36625 -650
rect 36655 -680 36665 -650
rect 36615 -690 36665 -680
rect 36700 -500 36750 -490
rect 36700 -530 36710 -500
rect 36740 -530 36750 -500
rect 36700 -550 36750 -530
rect 36700 -580 36710 -550
rect 36740 -580 36750 -550
rect 36700 -600 36750 -580
rect 36700 -630 36710 -600
rect 36740 -630 36750 -600
rect 36700 -650 36750 -630
rect 36700 -680 36710 -650
rect 36740 -680 36750 -650
rect 36700 -690 36750 -680
rect 36785 -500 36835 -490
rect 36785 -530 36795 -500
rect 36825 -530 36835 -500
rect 36785 -550 36835 -530
rect 36785 -580 36795 -550
rect 36825 -580 36835 -550
rect 36785 -600 36835 -580
rect 36785 -630 36795 -600
rect 36825 -630 36835 -600
rect 36785 -650 36835 -630
rect 36785 -680 36795 -650
rect 36825 -680 36835 -650
rect 36785 -690 36835 -680
rect 36870 -500 36920 -490
rect 36870 -530 36880 -500
rect 36910 -530 36920 -500
rect 36870 -550 36920 -530
rect 36870 -580 36880 -550
rect 36910 -580 36920 -550
rect 36870 -600 36920 -580
rect 36870 -630 36880 -600
rect 36910 -630 36920 -600
rect 36870 -650 36920 -630
rect 36870 -680 36880 -650
rect 36910 -680 36920 -650
rect 36870 -690 36920 -680
rect 36955 -500 37005 -490
rect 36955 -530 36965 -500
rect 36995 -530 37005 -500
rect 36955 -550 37005 -530
rect 36955 -580 36965 -550
rect 36995 -580 37005 -550
rect 36955 -600 37005 -580
rect 36955 -630 36965 -600
rect 36995 -630 37005 -600
rect 36955 -650 37005 -630
rect 36955 -680 36965 -650
rect 36995 -680 37005 -650
rect 36955 -690 37005 -680
rect 37040 -500 37090 -490
rect 37040 -530 37050 -500
rect 37080 -530 37090 -500
rect 37040 -550 37090 -530
rect 37040 -580 37050 -550
rect 37080 -580 37090 -550
rect 37040 -600 37090 -580
rect 37040 -630 37050 -600
rect 37080 -630 37090 -600
rect 37040 -650 37090 -630
rect 37040 -680 37050 -650
rect 37080 -680 37090 -650
rect 37040 -690 37090 -680
rect 37125 -500 37175 -490
rect 37125 -530 37135 -500
rect 37165 -530 37175 -500
rect 37125 -550 37175 -530
rect 37125 -580 37135 -550
rect 37165 -580 37175 -550
rect 37125 -600 37175 -580
rect 37125 -630 37135 -600
rect 37165 -630 37175 -600
rect 37125 -650 37175 -630
rect 37125 -680 37135 -650
rect 37165 -680 37175 -650
rect 37125 -690 37175 -680
rect 37210 -500 37260 -490
rect 37210 -530 37220 -500
rect 37250 -530 37260 -500
rect 37210 -550 37260 -530
rect 37210 -580 37220 -550
rect 37250 -580 37260 -550
rect 37210 -600 37260 -580
rect 37210 -630 37220 -600
rect 37250 -630 37260 -600
rect 37210 -650 37260 -630
rect 37210 -680 37220 -650
rect 37250 -680 37260 -650
rect 37210 -690 37260 -680
rect 37295 -500 37345 -490
rect 37295 -530 37305 -500
rect 37335 -530 37345 -500
rect 37295 -550 37345 -530
rect 37295 -580 37305 -550
rect 37335 -580 37345 -550
rect 37295 -600 37345 -580
rect 37295 -630 37305 -600
rect 37335 -630 37345 -600
rect 37295 -650 37345 -630
rect 37295 -680 37305 -650
rect 37335 -680 37345 -650
rect 37295 -690 37345 -680
rect 37380 -500 37430 -490
rect 37380 -530 37390 -500
rect 37420 -530 37430 -500
rect 37380 -550 37430 -530
rect 37380 -580 37390 -550
rect 37420 -580 37430 -550
rect 37380 -600 37430 -580
rect 37380 -630 37390 -600
rect 37420 -630 37430 -600
rect 37380 -650 37430 -630
rect 37380 -680 37390 -650
rect 37420 -680 37430 -650
rect 37380 -690 37430 -680
rect 37465 -500 37515 -490
rect 37465 -530 37475 -500
rect 37505 -530 37515 -500
rect 37465 -550 37515 -530
rect 37465 -580 37475 -550
rect 37505 -580 37515 -550
rect 37465 -600 37515 -580
rect 37465 -630 37475 -600
rect 37505 -630 37515 -600
rect 37465 -650 37515 -630
rect 37465 -680 37475 -650
rect 37505 -680 37515 -650
rect 37465 -690 37515 -680
rect 37550 -500 37600 -490
rect 37550 -530 37560 -500
rect 37590 -530 37600 -500
rect 37550 -550 37600 -530
rect 37550 -580 37560 -550
rect 37590 -580 37600 -550
rect 37550 -600 37600 -580
rect 37550 -630 37560 -600
rect 37590 -630 37600 -600
rect 37550 -650 37600 -630
rect 37550 -680 37560 -650
rect 37590 -680 37600 -650
rect 37550 -690 37600 -680
rect 37635 -500 37685 -490
rect 37635 -530 37645 -500
rect 37675 -530 37685 -500
rect 37635 -550 37685 -530
rect 37635 -580 37645 -550
rect 37675 -580 37685 -550
rect 37635 -600 37685 -580
rect 37635 -630 37645 -600
rect 37675 -630 37685 -600
rect 37635 -650 37685 -630
rect 37635 -680 37645 -650
rect 37675 -680 37685 -650
rect 37635 -690 37685 -680
rect 37720 -500 37770 -490
rect 37720 -530 37730 -500
rect 37760 -530 37770 -500
rect 37720 -550 37770 -530
rect 37720 -580 37730 -550
rect 37760 -580 37770 -550
rect 37720 -600 37770 -580
rect 37720 -630 37730 -600
rect 37760 -630 37770 -600
rect 37720 -650 37770 -630
rect 37720 -680 37730 -650
rect 37760 -680 37770 -650
rect 37720 -690 37770 -680
rect 37805 -500 37855 -490
rect 37805 -530 37815 -500
rect 37845 -530 37855 -500
rect 37805 -550 37855 -530
rect 37805 -580 37815 -550
rect 37845 -580 37855 -550
rect 37805 -600 37855 -580
rect 37805 -630 37815 -600
rect 37845 -630 37855 -600
rect 37805 -650 37855 -630
rect 37805 -680 37815 -650
rect 37845 -680 37855 -650
rect 37805 -690 37855 -680
rect 37890 -500 37940 -490
rect 37890 -530 37900 -500
rect 37930 -530 37940 -500
rect 37890 -550 37940 -530
rect 37890 -580 37900 -550
rect 37930 -580 37940 -550
rect 37890 -600 37940 -580
rect 37890 -630 37900 -600
rect 37930 -630 37940 -600
rect 37890 -650 37940 -630
rect 37890 -680 37900 -650
rect 37930 -680 37940 -650
rect 37890 -690 37940 -680
rect 37975 -500 38025 -490
rect 37975 -530 37985 -500
rect 38015 -530 38025 -500
rect 37975 -550 38025 -530
rect 37975 -580 37985 -550
rect 38015 -580 38025 -550
rect 37975 -600 38025 -580
rect 37975 -630 37985 -600
rect 38015 -630 38025 -600
rect 37975 -650 38025 -630
rect 37975 -680 37985 -650
rect 38015 -680 38025 -650
rect 37975 -690 38025 -680
rect 38060 -500 38110 -490
rect 38060 -530 38070 -500
rect 38100 -530 38110 -500
rect 38060 -550 38110 -530
rect 38060 -580 38070 -550
rect 38100 -580 38110 -550
rect 38060 -600 38110 -580
rect 38060 -630 38070 -600
rect 38100 -630 38110 -600
rect 38060 -650 38110 -630
rect 38060 -680 38070 -650
rect 38100 -680 38110 -650
rect 38060 -690 38110 -680
rect 38145 -500 38195 -490
rect 38145 -530 38155 -500
rect 38185 -530 38195 -500
rect 38145 -550 38195 -530
rect 38145 -580 38155 -550
rect 38185 -580 38195 -550
rect 38145 -600 38195 -580
rect 38145 -630 38155 -600
rect 38185 -630 38195 -600
rect 38145 -650 38195 -630
rect 38145 -680 38155 -650
rect 38185 -680 38195 -650
rect 38145 -690 38195 -680
rect 38230 -500 38280 -490
rect 38230 -530 38240 -500
rect 38270 -530 38280 -500
rect 38230 -550 38280 -530
rect 38230 -580 38240 -550
rect 38270 -580 38280 -550
rect 38230 -600 38280 -580
rect 38230 -630 38240 -600
rect 38270 -630 38280 -600
rect 38230 -650 38280 -630
rect 38230 -680 38240 -650
rect 38270 -680 38280 -650
rect 38230 -690 38280 -680
rect 38315 -500 38365 -490
rect 38315 -530 38325 -500
rect 38355 -530 38365 -500
rect 38315 -550 38365 -530
rect 38315 -580 38325 -550
rect 38355 -580 38365 -550
rect 38315 -600 38365 -580
rect 38315 -630 38325 -600
rect 38355 -630 38365 -600
rect 38315 -650 38365 -630
rect 38315 -680 38325 -650
rect 38355 -680 38365 -650
rect 38315 -690 38365 -680
rect 38400 -500 38450 -490
rect 38400 -530 38410 -500
rect 38440 -530 38450 -500
rect 38400 -550 38450 -530
rect 38400 -580 38410 -550
rect 38440 -580 38450 -550
rect 38400 -600 38450 -580
rect 38400 -630 38410 -600
rect 38440 -630 38450 -600
rect 38400 -650 38450 -630
rect 38400 -680 38410 -650
rect 38440 -680 38450 -650
rect 38400 -690 38450 -680
rect 38485 -500 38535 -490
rect 38485 -530 38495 -500
rect 38525 -530 38535 -500
rect 38485 -550 38535 -530
rect 38485 -580 38495 -550
rect 38525 -580 38535 -550
rect 38485 -600 38535 -580
rect 38485 -630 38495 -600
rect 38525 -630 38535 -600
rect 38485 -650 38535 -630
rect 38485 -680 38495 -650
rect 38525 -680 38535 -650
rect 38485 -690 38535 -680
rect 38570 -500 38620 -490
rect 38570 -530 38580 -500
rect 38610 -530 38620 -500
rect 38570 -550 38620 -530
rect 38570 -580 38580 -550
rect 38610 -580 38620 -550
rect 38570 -600 38620 -580
rect 38570 -630 38580 -600
rect 38610 -630 38620 -600
rect 38570 -650 38620 -630
rect 38570 -680 38580 -650
rect 38610 -680 38620 -650
rect 38570 -690 38620 -680
rect 38655 -500 38705 -490
rect 38655 -530 38665 -500
rect 38695 -530 38705 -500
rect 38655 -550 38705 -530
rect 38655 -580 38665 -550
rect 38695 -580 38705 -550
rect 38655 -600 38705 -580
rect 38655 -630 38665 -600
rect 38695 -630 38705 -600
rect 38655 -650 38705 -630
rect 38655 -680 38665 -650
rect 38695 -680 38705 -650
rect 38655 -690 38705 -680
rect 38740 -500 38790 -490
rect 38740 -530 38750 -500
rect 38780 -530 38790 -500
rect 38740 -550 38790 -530
rect 38740 -580 38750 -550
rect 38780 -580 38790 -550
rect 38740 -600 38790 -580
rect 38740 -630 38750 -600
rect 38780 -630 38790 -600
rect 38740 -650 38790 -630
rect 38740 -680 38750 -650
rect 38780 -680 38790 -650
rect 38740 -690 38790 -680
rect 38825 -500 38875 -490
rect 38825 -530 38835 -500
rect 38865 -530 38875 -500
rect 38825 -550 38875 -530
rect 38825 -580 38835 -550
rect 38865 -580 38875 -550
rect 38825 -600 38875 -580
rect 38825 -630 38835 -600
rect 38865 -630 38875 -600
rect 38825 -650 38875 -630
rect 38825 -680 38835 -650
rect 38865 -680 38875 -650
rect 38825 -690 38875 -680
rect 38910 -500 38960 -490
rect 38910 -530 38920 -500
rect 38950 -530 38960 -500
rect 38910 -550 38960 -530
rect 38910 -580 38920 -550
rect 38950 -580 38960 -550
rect 38910 -600 38960 -580
rect 38910 -630 38920 -600
rect 38950 -630 38960 -600
rect 38910 -650 38960 -630
rect 38910 -680 38920 -650
rect 38950 -680 38960 -650
rect 38910 -690 38960 -680
rect 38995 -500 39045 -490
rect 38995 -530 39005 -500
rect 39035 -530 39045 -500
rect 38995 -550 39045 -530
rect 38995 -580 39005 -550
rect 39035 -580 39045 -550
rect 38995 -600 39045 -580
rect 38995 -630 39005 -600
rect 39035 -630 39045 -600
rect 38995 -650 39045 -630
rect 38995 -680 39005 -650
rect 39035 -680 39045 -650
rect 38995 -690 39045 -680
rect 39080 -500 39130 -490
rect 39080 -530 39090 -500
rect 39120 -530 39130 -500
rect 39080 -550 39130 -530
rect 39080 -580 39090 -550
rect 39120 -580 39130 -550
rect 39080 -600 39130 -580
rect 39080 -630 39090 -600
rect 39120 -630 39130 -600
rect 39080 -650 39130 -630
rect 39080 -680 39090 -650
rect 39120 -680 39130 -650
rect 39080 -690 39130 -680
rect 39165 -500 39215 -490
rect 39165 -530 39175 -500
rect 39205 -530 39215 -500
rect 39165 -550 39215 -530
rect 39165 -580 39175 -550
rect 39205 -580 39215 -550
rect 39165 -600 39215 -580
rect 39165 -630 39175 -600
rect 39205 -630 39215 -600
rect 39165 -650 39215 -630
rect 39165 -680 39175 -650
rect 39205 -680 39215 -650
rect 39165 -690 39215 -680
rect 39250 -500 39300 -490
rect 39250 -530 39260 -500
rect 39290 -530 39300 -500
rect 39250 -550 39300 -530
rect 39250 -580 39260 -550
rect 39290 -580 39300 -550
rect 39250 -600 39300 -580
rect 39250 -630 39260 -600
rect 39290 -630 39300 -600
rect 39250 -650 39300 -630
rect 39250 -680 39260 -650
rect 39290 -680 39300 -650
rect 39250 -690 39300 -680
rect 39335 -500 39385 -490
rect 39335 -530 39345 -500
rect 39375 -530 39385 -500
rect 39335 -550 39385 -530
rect 39335 -580 39345 -550
rect 39375 -580 39385 -550
rect 39335 -600 39385 -580
rect 39335 -630 39345 -600
rect 39375 -630 39385 -600
rect 39335 -650 39385 -630
rect 39335 -680 39345 -650
rect 39375 -680 39385 -650
rect 39335 -690 39385 -680
rect 39420 -500 39470 -490
rect 39420 -530 39430 -500
rect 39460 -530 39470 -500
rect 39420 -550 39470 -530
rect 39420 -580 39430 -550
rect 39460 -580 39470 -550
rect 39420 -600 39470 -580
rect 39420 -630 39430 -600
rect 39460 -630 39470 -600
rect 39420 -650 39470 -630
rect 39420 -680 39430 -650
rect 39460 -680 39470 -650
rect 39420 -690 39470 -680
rect 39505 -500 39555 -490
rect 39505 -530 39515 -500
rect 39545 -530 39555 -500
rect 39505 -550 39555 -530
rect 39505 -580 39515 -550
rect 39545 -580 39555 -550
rect 39505 -600 39555 -580
rect 39505 -630 39515 -600
rect 39545 -630 39555 -600
rect 39505 -650 39555 -630
rect 39505 -680 39515 -650
rect 39545 -680 39555 -650
rect 39505 -690 39555 -680
rect 39590 -500 39640 -490
rect 39590 -530 39600 -500
rect 39630 -530 39640 -500
rect 39590 -550 39640 -530
rect 39590 -580 39600 -550
rect 39630 -580 39640 -550
rect 39590 -600 39640 -580
rect 39590 -630 39600 -600
rect 39630 -630 39640 -600
rect 39590 -650 39640 -630
rect 39590 -680 39600 -650
rect 39630 -680 39640 -650
rect 39590 -690 39640 -680
rect 39675 -500 39725 -490
rect 39675 -530 39685 -500
rect 39715 -530 39725 -500
rect 39675 -550 39725 -530
rect 39675 -580 39685 -550
rect 39715 -580 39725 -550
rect 39675 -600 39725 -580
rect 39675 -630 39685 -600
rect 39715 -630 39725 -600
rect 39675 -650 39725 -630
rect 39675 -680 39685 -650
rect 39715 -680 39725 -650
rect 39675 -690 39725 -680
rect 39760 -500 39810 -490
rect 39760 -530 39770 -500
rect 39800 -530 39810 -500
rect 39760 -550 39810 -530
rect 39760 -580 39770 -550
rect 39800 -580 39810 -550
rect 39760 -600 39810 -580
rect 39760 -630 39770 -600
rect 39800 -630 39810 -600
rect 39760 -650 39810 -630
rect 39760 -680 39770 -650
rect 39800 -680 39810 -650
rect 39760 -690 39810 -680
rect 39845 -500 39895 -490
rect 39845 -530 39855 -500
rect 39885 -530 39895 -500
rect 39845 -550 39895 -530
rect 39845 -580 39855 -550
rect 39885 -580 39895 -550
rect 39845 -600 39895 -580
rect 39845 -630 39855 -600
rect 39885 -630 39895 -600
rect 39845 -650 39895 -630
rect 39845 -680 39855 -650
rect 39885 -680 39895 -650
rect 39845 -690 39895 -680
rect 39930 -500 39980 -490
rect 39930 -530 39940 -500
rect 39970 -530 39980 -500
rect 39930 -550 39980 -530
rect 39930 -580 39940 -550
rect 39970 -580 39980 -550
rect 39930 -600 39980 -580
rect 39930 -630 39940 -600
rect 39970 -630 39980 -600
rect 39930 -650 39980 -630
rect 39930 -680 39940 -650
rect 39970 -680 39980 -650
rect 39930 -690 39980 -680
rect 40015 -500 40065 -490
rect 40015 -530 40025 -500
rect 40055 -530 40065 -500
rect 40015 -550 40065 -530
rect 40015 -580 40025 -550
rect 40055 -580 40065 -550
rect 40015 -600 40065 -580
rect 40015 -630 40025 -600
rect 40055 -630 40065 -600
rect 40015 -650 40065 -630
rect 40015 -680 40025 -650
rect 40055 -680 40065 -650
rect 40015 -690 40065 -680
rect 40100 -500 40150 -490
rect 40100 -530 40110 -500
rect 40140 -530 40150 -500
rect 40100 -550 40150 -530
rect 40100 -580 40110 -550
rect 40140 -580 40150 -550
rect 40100 -600 40150 -580
rect 40100 -630 40110 -600
rect 40140 -630 40150 -600
rect 40100 -650 40150 -630
rect 40100 -680 40110 -650
rect 40140 -680 40150 -650
rect 40100 -690 40150 -680
rect 40185 -500 40235 -490
rect 40185 -530 40195 -500
rect 40225 -530 40235 -500
rect 40185 -550 40235 -530
rect 40185 -580 40195 -550
rect 40225 -580 40235 -550
rect 40185 -600 40235 -580
rect 40185 -630 40195 -600
rect 40225 -630 40235 -600
rect 40185 -650 40235 -630
rect 40185 -680 40195 -650
rect 40225 -680 40235 -650
rect 40185 -690 40235 -680
rect 40270 -500 40320 -490
rect 40270 -530 40280 -500
rect 40310 -530 40320 -500
rect 40270 -550 40320 -530
rect 40270 -580 40280 -550
rect 40310 -580 40320 -550
rect 40270 -600 40320 -580
rect 40270 -630 40280 -600
rect 40310 -630 40320 -600
rect 40270 -650 40320 -630
rect 40270 -680 40280 -650
rect 40310 -680 40320 -650
rect 40270 -690 40320 -680
rect 40355 -500 40405 -490
rect 40355 -530 40365 -500
rect 40395 -530 40405 -500
rect 40355 -550 40405 -530
rect 40355 -580 40365 -550
rect 40395 -580 40405 -550
rect 40355 -600 40405 -580
rect 40355 -630 40365 -600
rect 40395 -630 40405 -600
rect 40355 -650 40405 -630
rect 40355 -680 40365 -650
rect 40395 -680 40405 -650
rect 40355 -690 40405 -680
rect 40440 -500 40490 -490
rect 40440 -530 40450 -500
rect 40480 -530 40490 -500
rect 40440 -550 40490 -530
rect 40440 -580 40450 -550
rect 40480 -580 40490 -550
rect 40440 -600 40490 -580
rect 40440 -630 40450 -600
rect 40480 -630 40490 -600
rect 40440 -650 40490 -630
rect 40440 -680 40450 -650
rect 40480 -680 40490 -650
rect 40440 -690 40490 -680
rect 40525 -500 40575 -490
rect 40525 -530 40535 -500
rect 40565 -530 40575 -500
rect 40525 -550 40575 -530
rect 40525 -580 40535 -550
rect 40565 -580 40575 -550
rect 40525 -600 40575 -580
rect 40525 -630 40535 -600
rect 40565 -630 40575 -600
rect 40525 -650 40575 -630
rect 40525 -680 40535 -650
rect 40565 -680 40575 -650
rect 40525 -690 40575 -680
rect 40610 -500 40660 -490
rect 40610 -530 40620 -500
rect 40650 -530 40660 -500
rect 40610 -550 40660 -530
rect 40610 -580 40620 -550
rect 40650 -580 40660 -550
rect 40610 -600 40660 -580
rect 40610 -630 40620 -600
rect 40650 -630 40660 -600
rect 40610 -650 40660 -630
rect 40610 -680 40620 -650
rect 40650 -680 40660 -650
rect 40610 -690 40660 -680
rect 40695 -500 40745 -490
rect 40695 -530 40705 -500
rect 40735 -530 40745 -500
rect 40695 -550 40745 -530
rect 40695 -580 40705 -550
rect 40735 -580 40745 -550
rect 40695 -600 40745 -580
rect 40695 -630 40705 -600
rect 40735 -630 40745 -600
rect 40695 -650 40745 -630
rect 40695 -680 40705 -650
rect 40735 -680 40745 -650
rect 40695 -690 40745 -680
rect 40780 -500 40830 -490
rect 40780 -530 40790 -500
rect 40820 -530 40830 -500
rect 40780 -550 40830 -530
rect 40780 -580 40790 -550
rect 40820 -580 40830 -550
rect 40780 -600 40830 -580
rect 40780 -630 40790 -600
rect 40820 -630 40830 -600
rect 40780 -650 40830 -630
rect 40780 -680 40790 -650
rect 40820 -680 40830 -650
rect 40780 -690 40830 -680
rect 40865 -500 40915 -490
rect 40865 -530 40875 -500
rect 40905 -530 40915 -500
rect 40865 -550 40915 -530
rect 40865 -580 40875 -550
rect 40905 -580 40915 -550
rect 40865 -600 40915 -580
rect 40865 -630 40875 -600
rect 40905 -630 40915 -600
rect 40865 -650 40915 -630
rect 40865 -680 40875 -650
rect 40905 -680 40915 -650
rect 40865 -690 40915 -680
rect 40950 -500 41000 -490
rect 40950 -530 40960 -500
rect 40990 -530 41000 -500
rect 40950 -550 41000 -530
rect 40950 -580 40960 -550
rect 40990 -580 41000 -550
rect 40950 -600 41000 -580
rect 40950 -630 40960 -600
rect 40990 -630 41000 -600
rect 40950 -650 41000 -630
rect 40950 -680 40960 -650
rect 40990 -680 41000 -650
rect 40950 -690 41000 -680
rect 41035 -500 41085 -490
rect 41035 -530 41045 -500
rect 41075 -530 41085 -500
rect 41035 -550 41085 -530
rect 41035 -580 41045 -550
rect 41075 -580 41085 -550
rect 41035 -600 41085 -580
rect 41035 -630 41045 -600
rect 41075 -630 41085 -600
rect 41035 -650 41085 -630
rect 41035 -680 41045 -650
rect 41075 -680 41085 -650
rect 41035 -690 41085 -680
rect 41120 -500 41170 -490
rect 41120 -530 41130 -500
rect 41160 -530 41170 -500
rect 41120 -550 41170 -530
rect 41120 -580 41130 -550
rect 41160 -580 41170 -550
rect 41120 -600 41170 -580
rect 41120 -630 41130 -600
rect 41160 -630 41170 -600
rect 41120 -650 41170 -630
rect 41120 -680 41130 -650
rect 41160 -680 41170 -650
rect 41120 -690 41170 -680
rect 41205 -500 41255 -490
rect 41205 -530 41215 -500
rect 41245 -530 41255 -500
rect 41205 -550 41255 -530
rect 41205 -580 41215 -550
rect 41245 -580 41255 -550
rect 41205 -600 41255 -580
rect 41205 -630 41215 -600
rect 41245 -630 41255 -600
rect 41205 -650 41255 -630
rect 41205 -680 41215 -650
rect 41245 -680 41255 -650
rect 41205 -690 41255 -680
rect 41290 -500 41340 -490
rect 41290 -530 41300 -500
rect 41330 -530 41340 -500
rect 41290 -550 41340 -530
rect 41290 -580 41300 -550
rect 41330 -580 41340 -550
rect 41290 -600 41340 -580
rect 41290 -630 41300 -600
rect 41330 -630 41340 -600
rect 41290 -650 41340 -630
rect 41290 -680 41300 -650
rect 41330 -680 41340 -650
rect 41290 -690 41340 -680
rect 41375 -500 41425 -490
rect 41375 -530 41385 -500
rect 41415 -530 41425 -500
rect 41375 -550 41425 -530
rect 41375 -580 41385 -550
rect 41415 -580 41425 -550
rect 41375 -600 41425 -580
rect 41375 -630 41385 -600
rect 41415 -630 41425 -600
rect 41375 -650 41425 -630
rect 41375 -680 41385 -650
rect 41415 -680 41425 -650
rect 41375 -690 41425 -680
rect 41460 -500 41510 -490
rect 41460 -530 41470 -500
rect 41500 -530 41510 -500
rect 41460 -550 41510 -530
rect 41460 -580 41470 -550
rect 41500 -580 41510 -550
rect 41460 -600 41510 -580
rect 41460 -630 41470 -600
rect 41500 -630 41510 -600
rect 41460 -650 41510 -630
rect 41460 -680 41470 -650
rect 41500 -680 41510 -650
rect 41460 -690 41510 -680
rect 41545 -500 41595 -490
rect 41545 -530 41555 -500
rect 41585 -530 41595 -500
rect 41545 -550 41595 -530
rect 41545 -580 41555 -550
rect 41585 -580 41595 -550
rect 41545 -600 41595 -580
rect 41545 -630 41555 -600
rect 41585 -630 41595 -600
rect 41545 -650 41595 -630
rect 41545 -680 41555 -650
rect 41585 -680 41595 -650
rect 41545 -690 41595 -680
rect 41630 -500 41680 -490
rect 41630 -530 41640 -500
rect 41670 -530 41680 -500
rect 41630 -550 41680 -530
rect 41630 -580 41640 -550
rect 41670 -580 41680 -550
rect 41630 -600 41680 -580
rect 41630 -630 41640 -600
rect 41670 -630 41680 -600
rect 41630 -650 41680 -630
rect 41630 -680 41640 -650
rect 41670 -680 41680 -650
rect 41630 -690 41680 -680
rect 41715 -500 41765 -490
rect 41715 -530 41725 -500
rect 41755 -530 41765 -500
rect 41715 -550 41765 -530
rect 41715 -580 41725 -550
rect 41755 -580 41765 -550
rect 41715 -600 41765 -580
rect 41715 -630 41725 -600
rect 41755 -630 41765 -600
rect 41715 -650 41765 -630
rect 41715 -680 41725 -650
rect 41755 -680 41765 -650
rect 41715 -690 41765 -680
rect 41800 -500 41850 -490
rect 41800 -530 41810 -500
rect 41840 -530 41850 -500
rect 41800 -550 41850 -530
rect 41800 -580 41810 -550
rect 41840 -580 41850 -550
rect 41800 -600 41850 -580
rect 41800 -630 41810 -600
rect 41840 -630 41850 -600
rect 41800 -650 41850 -630
rect 41800 -680 41810 -650
rect 41840 -680 41850 -650
rect 41800 -690 41850 -680
rect 41885 -500 41935 -490
rect 41885 -530 41895 -500
rect 41925 -530 41935 -500
rect 41885 -550 41935 -530
rect 41885 -580 41895 -550
rect 41925 -580 41935 -550
rect 41885 -600 41935 -580
rect 41885 -630 41895 -600
rect 41925 -630 41935 -600
rect 41885 -650 41935 -630
rect 41885 -680 41895 -650
rect 41925 -680 41935 -650
rect 41885 -690 41935 -680
rect 41970 -500 42020 -490
rect 41970 -530 41980 -500
rect 42010 -530 42020 -500
rect 41970 -550 42020 -530
rect 41970 -580 41980 -550
rect 42010 -580 42020 -550
rect 41970 -600 42020 -580
rect 41970 -630 41980 -600
rect 42010 -630 42020 -600
rect 41970 -650 42020 -630
rect 41970 -680 41980 -650
rect 42010 -680 42020 -650
rect 41970 -690 42020 -680
rect 42055 -500 42105 -490
rect 42055 -530 42065 -500
rect 42095 -530 42105 -500
rect 42055 -550 42105 -530
rect 42055 -580 42065 -550
rect 42095 -580 42105 -550
rect 42055 -600 42105 -580
rect 42055 -630 42065 -600
rect 42095 -630 42105 -600
rect 42055 -650 42105 -630
rect 42055 -680 42065 -650
rect 42095 -680 42105 -650
rect 42055 -690 42105 -680
rect 42140 -500 42190 -490
rect 42140 -530 42150 -500
rect 42180 -530 42190 -500
rect 42140 -550 42190 -530
rect 42140 -580 42150 -550
rect 42180 -580 42190 -550
rect 42140 -600 42190 -580
rect 42140 -630 42150 -600
rect 42180 -630 42190 -600
rect 42140 -650 42190 -630
rect 42140 -680 42150 -650
rect 42180 -680 42190 -650
rect 42140 -690 42190 -680
rect 42225 -500 42275 -490
rect 42225 -530 42235 -500
rect 42265 -530 42275 -500
rect 42225 -550 42275 -530
rect 42225 -580 42235 -550
rect 42265 -580 42275 -550
rect 42225 -600 42275 -580
rect 42225 -630 42235 -600
rect 42265 -630 42275 -600
rect 42225 -650 42275 -630
rect 42225 -680 42235 -650
rect 42265 -680 42275 -650
rect 42225 -690 42275 -680
rect 42310 -500 42360 -490
rect 42310 -530 42320 -500
rect 42350 -530 42360 -500
rect 42310 -550 42360 -530
rect 42310 -580 42320 -550
rect 42350 -580 42360 -550
rect 42310 -600 42360 -580
rect 42310 -630 42320 -600
rect 42350 -630 42360 -600
rect 42310 -650 42360 -630
rect 42310 -680 42320 -650
rect 42350 -680 42360 -650
rect 42310 -690 42360 -680
rect 42395 -500 42445 -490
rect 42395 -530 42405 -500
rect 42435 -530 42445 -500
rect 42395 -550 42445 -530
rect 42395 -580 42405 -550
rect 42435 -580 42445 -550
rect 42395 -600 42445 -580
rect 42395 -630 42405 -600
rect 42435 -630 42445 -600
rect 42395 -650 42445 -630
rect 42395 -680 42405 -650
rect 42435 -680 42445 -650
rect 42395 -690 42445 -680
rect 42480 -500 42530 -490
rect 42480 -530 42490 -500
rect 42520 -530 42530 -500
rect 42480 -550 42530 -530
rect 42480 -580 42490 -550
rect 42520 -580 42530 -550
rect 42480 -600 42530 -580
rect 42480 -630 42490 -600
rect 42520 -630 42530 -600
rect 42480 -650 42530 -630
rect 42480 -680 42490 -650
rect 42520 -680 42530 -650
rect 42480 -690 42530 -680
rect 42565 -500 42615 -490
rect 42565 -530 42575 -500
rect 42605 -530 42615 -500
rect 42565 -550 42615 -530
rect 42565 -580 42575 -550
rect 42605 -580 42615 -550
rect 42565 -600 42615 -580
rect 42565 -630 42575 -600
rect 42605 -630 42615 -600
rect 42565 -650 42615 -630
rect 42565 -680 42575 -650
rect 42605 -680 42615 -650
rect 42565 -690 42615 -680
rect 42650 -500 42700 -490
rect 42650 -530 42660 -500
rect 42690 -530 42700 -500
rect 42650 -550 42700 -530
rect 42650 -580 42660 -550
rect 42690 -580 42700 -550
rect 42650 -600 42700 -580
rect 42650 -630 42660 -600
rect 42690 -630 42700 -600
rect 42650 -650 42700 -630
rect 42650 -680 42660 -650
rect 42690 -680 42700 -650
rect 42650 -690 42700 -680
rect 42735 -500 42785 -490
rect 42735 -530 42745 -500
rect 42775 -530 42785 -500
rect 42735 -550 42785 -530
rect 42735 -580 42745 -550
rect 42775 -580 42785 -550
rect 42735 -600 42785 -580
rect 42735 -630 42745 -600
rect 42775 -630 42785 -600
rect 42735 -650 42785 -630
rect 42735 -680 42745 -650
rect 42775 -680 42785 -650
rect 42735 -690 42785 -680
rect 42820 -500 42870 -490
rect 42820 -530 42830 -500
rect 42860 -530 42870 -500
rect 42820 -550 42870 -530
rect 42820 -580 42830 -550
rect 42860 -580 42870 -550
rect 42820 -600 42870 -580
rect 42820 -630 42830 -600
rect 42860 -630 42870 -600
rect 42820 -650 42870 -630
rect 42820 -680 42830 -650
rect 42860 -680 42870 -650
rect 42820 -690 42870 -680
rect 42905 -500 42955 -490
rect 42905 -530 42915 -500
rect 42945 -530 42955 -500
rect 42905 -550 42955 -530
rect 42905 -580 42915 -550
rect 42945 -580 42955 -550
rect 42905 -600 42955 -580
rect 42905 -630 42915 -600
rect 42945 -630 42955 -600
rect 42905 -650 42955 -630
rect 42905 -680 42915 -650
rect 42945 -680 42955 -650
rect 42905 -690 42955 -680
rect 42990 -500 43040 -490
rect 42990 -530 43000 -500
rect 43030 -530 43040 -500
rect 42990 -550 43040 -530
rect 42990 -580 43000 -550
rect 43030 -580 43040 -550
rect 42990 -600 43040 -580
rect 42990 -630 43000 -600
rect 43030 -630 43040 -600
rect 42990 -650 43040 -630
rect 42990 -680 43000 -650
rect 43030 -680 43040 -650
rect 42990 -690 43040 -680
rect 43075 -500 43125 -490
rect 43075 -530 43085 -500
rect 43115 -530 43125 -500
rect 43075 -550 43125 -530
rect 43075 -580 43085 -550
rect 43115 -580 43125 -550
rect 43075 -600 43125 -580
rect 43075 -630 43085 -600
rect 43115 -630 43125 -600
rect 43075 -650 43125 -630
rect 43075 -680 43085 -650
rect 43115 -680 43125 -650
rect 43075 -690 43125 -680
rect 43160 -500 43210 -490
rect 43160 -530 43170 -500
rect 43200 -530 43210 -500
rect 43160 -550 43210 -530
rect 43160 -580 43170 -550
rect 43200 -580 43210 -550
rect 43160 -600 43210 -580
rect 43160 -630 43170 -600
rect 43200 -630 43210 -600
rect 43160 -650 43210 -630
rect 43160 -680 43170 -650
rect 43200 -680 43210 -650
rect 43160 -690 43210 -680
rect 43245 -500 43295 -490
rect 43245 -530 43255 -500
rect 43285 -530 43295 -500
rect 43245 -550 43295 -530
rect 43245 -580 43255 -550
rect 43285 -580 43295 -550
rect 43245 -600 43295 -580
rect 43245 -630 43255 -600
rect 43285 -630 43295 -600
rect 43245 -650 43295 -630
rect 43245 -680 43255 -650
rect 43285 -680 43295 -650
rect 43245 -690 43295 -680
rect 43330 -500 43380 -490
rect 43330 -530 43340 -500
rect 43370 -530 43380 -500
rect 43330 -550 43380 -530
rect 43330 -580 43340 -550
rect 43370 -580 43380 -550
rect 43330 -600 43380 -580
rect 43330 -630 43340 -600
rect 43370 -630 43380 -600
rect 43330 -650 43380 -630
rect 43330 -680 43340 -650
rect 43370 -680 43380 -650
rect 43330 -690 43380 -680
rect 43415 -500 43465 -490
rect 43415 -530 43425 -500
rect 43455 -530 43465 -500
rect 43415 -550 43465 -530
rect 43415 -580 43425 -550
rect 43455 -580 43465 -550
rect 43415 -600 43465 -580
rect 43415 -630 43425 -600
rect 43455 -630 43465 -600
rect 43415 -650 43465 -630
rect 43415 -680 43425 -650
rect 43455 -680 43465 -650
rect 43415 -690 43465 -680
rect 43500 -500 43550 -490
rect 43500 -530 43510 -500
rect 43540 -530 43550 -500
rect 43500 -550 43550 -530
rect 43500 -580 43510 -550
rect 43540 -580 43550 -550
rect 43500 -600 43550 -580
rect 43500 -630 43510 -600
rect 43540 -630 43550 -600
rect 43500 -650 43550 -630
rect 43500 -680 43510 -650
rect 43540 -680 43550 -650
rect 43500 -690 43550 -680
rect 43585 -500 43635 -490
rect 43585 -530 43595 -500
rect 43625 -530 43635 -500
rect 43585 -550 43635 -530
rect 43585 -580 43595 -550
rect 43625 -580 43635 -550
rect 43585 -600 43635 -580
rect 43585 -630 43595 -600
rect 43625 -630 43635 -600
rect 43585 -650 43635 -630
rect 43585 -680 43595 -650
rect 43625 -680 43635 -650
rect 43585 -690 43635 -680
<< viali >>
rect 225 175 255 205
rect 310 125 340 155
rect 395 175 425 205
rect 480 125 510 155
rect 565 175 595 205
rect 760 175 790 205
rect 845 125 875 155
rect 930 175 960 205
rect 1015 125 1045 155
rect 1100 175 1130 205
rect 1185 125 1215 155
rect 1270 175 1300 205
rect 1355 125 1385 155
rect 1440 175 1470 205
rect 1525 125 1555 155
rect 1610 175 1640 205
rect 1695 125 1725 155
rect 1780 175 1810 205
rect 1865 125 1895 155
rect 1950 175 1980 205
rect 2035 125 2065 155
rect 2120 175 2150 205
rect 2270 175 2300 205
rect 2355 125 2385 155
rect 2440 175 2470 205
rect 2525 125 2555 155
rect 2610 175 2640 205
rect 2695 125 2725 155
rect 2780 175 2810 205
rect 2865 125 2895 155
rect 2950 175 2980 205
rect 3035 125 3065 155
rect 3120 175 3150 205
rect 3205 125 3235 155
rect 3290 175 3320 205
rect 3375 125 3405 155
rect 3460 175 3490 205
rect 3545 125 3575 155
rect 3630 175 3660 205
rect 3715 125 3745 155
rect 3800 175 3830 205
rect 3885 125 3915 155
rect 3970 175 4000 205
rect 4055 125 4085 155
rect 4140 175 4170 205
rect 4225 125 4255 155
rect 4310 175 4340 205
rect 4395 125 4425 155
rect 4480 175 4510 205
rect 4565 125 4595 155
rect 4650 175 4680 205
rect 4735 125 4765 155
rect 4820 175 4850 205
rect 4905 125 4935 155
rect 4990 175 5020 205
rect 5075 125 5105 155
rect 5160 175 5190 205
rect 5245 125 5275 155
rect 5330 175 5360 205
rect 5415 125 5445 155
rect 5500 175 5530 205
rect 5585 125 5615 155
rect 5670 175 5700 205
rect 5755 125 5785 155
rect 5840 175 5870 205
rect 5925 125 5955 155
rect 6010 175 6040 205
rect 6095 125 6125 155
rect 6180 175 6210 205
rect 6265 125 6295 155
rect 6350 175 6380 205
rect 6435 125 6465 155
rect 6520 175 6550 205
rect 6605 125 6635 155
rect 6690 175 6720 205
rect 6775 125 6805 155
rect 6860 175 6890 205
rect 6945 125 6975 155
rect 7030 175 7060 205
rect 7115 125 7145 155
rect 7200 175 7230 205
rect 7285 125 7315 155
rect 7370 175 7400 205
rect 7455 125 7485 155
rect 7540 175 7570 205
rect 7625 125 7655 155
rect 7710 175 7740 205
rect 7860 175 7890 205
rect 7945 125 7975 155
rect 8030 175 8060 205
rect 8115 125 8145 155
rect 8200 175 8230 205
rect 8285 125 8315 155
rect 8370 175 8400 205
rect 8455 125 8485 155
rect 8540 175 8570 205
rect 8625 125 8655 155
rect 8710 175 8740 205
rect 8795 125 8825 155
rect 8880 175 8910 205
rect 8965 125 8995 155
rect 9050 175 9080 205
rect 9135 125 9165 155
rect 9220 175 9250 205
rect 9305 125 9335 155
rect 9390 175 9420 205
rect 9475 125 9505 155
rect 9560 175 9590 205
rect 9645 125 9675 155
rect 9730 175 9760 205
rect 9815 125 9845 155
rect 9900 175 9930 205
rect 9985 125 10015 155
rect 10070 175 10100 205
rect 10155 125 10185 155
rect 10240 175 10270 205
rect 10325 125 10355 155
rect 10410 175 10440 205
rect 10495 125 10525 155
rect 10580 175 10610 205
rect 10665 125 10695 155
rect 10750 175 10780 205
rect 10835 125 10865 155
rect 10920 175 10950 205
rect 11005 125 11035 155
rect 11090 175 11120 205
rect 11175 125 11205 155
rect 11260 175 11290 205
rect 11345 125 11375 155
rect 11430 175 11460 205
rect 11515 125 11545 155
rect 11600 175 11630 205
rect 11685 125 11715 155
rect 11770 175 11800 205
rect 11855 125 11885 155
rect 11940 175 11970 205
rect 12025 125 12055 155
rect 12110 175 12140 205
rect 12195 125 12225 155
rect 12280 175 12310 205
rect 12365 125 12395 155
rect 12450 175 12480 205
rect 12535 125 12565 155
rect 12620 175 12650 205
rect 12705 125 12735 155
rect 12790 175 12820 205
rect 12875 125 12905 155
rect 12960 175 12990 205
rect 13045 125 13075 155
rect 13130 175 13160 205
rect 13215 125 13245 155
rect 13300 175 13330 205
rect 13385 125 13415 155
rect 13470 175 13500 205
rect 13555 125 13585 155
rect 13640 175 13670 205
rect 13725 125 13755 155
rect 13810 175 13840 205
rect 13895 125 13925 155
rect 13980 175 14010 205
rect 14065 125 14095 155
rect 14150 175 14180 205
rect 14235 125 14265 155
rect 14320 175 14350 205
rect 14405 125 14435 155
rect 14490 175 14520 205
rect 14575 125 14605 155
rect 14660 175 14690 205
rect 14745 125 14775 155
rect 14830 175 14860 205
rect 14915 125 14945 155
rect 15000 175 15030 205
rect 15085 125 15115 155
rect 15170 175 15200 205
rect 15255 125 15285 155
rect 15340 175 15370 205
rect 15425 125 15455 155
rect 15510 175 15540 205
rect 15595 125 15625 155
rect 15680 175 15710 205
rect 15765 125 15795 155
rect 15850 175 15880 205
rect 15935 125 15965 155
rect 16020 175 16050 205
rect 16105 125 16135 155
rect 16190 175 16220 205
rect 16275 125 16305 155
rect 16360 175 16390 205
rect 16445 125 16475 155
rect 16530 175 16560 205
rect 16615 125 16645 155
rect 16700 175 16730 205
rect 16785 125 16815 155
rect 16870 175 16900 205
rect 16955 125 16985 155
rect 17040 175 17070 205
rect 17125 125 17155 155
rect 17210 175 17240 205
rect 17295 125 17325 155
rect 17380 175 17410 205
rect 17465 125 17495 155
rect 17550 175 17580 205
rect 17635 125 17665 155
rect 17720 175 17750 205
rect 17805 125 17835 155
rect 17890 175 17920 205
rect 17975 125 18005 155
rect 18060 175 18090 205
rect 18145 125 18175 155
rect 18230 175 18260 205
rect 18315 125 18345 155
rect 18400 175 18430 205
rect 18485 125 18515 155
rect 18570 175 18600 205
rect 18655 125 18685 155
rect 18740 175 18770 205
rect 18825 125 18855 155
rect 18910 175 18940 205
rect 18995 125 19025 155
rect 19080 175 19110 205
rect 19165 125 19195 155
rect 19250 175 19280 205
rect 19335 125 19365 155
rect 19420 175 19450 205
rect 19505 125 19535 155
rect 19590 175 19620 205
rect 19675 125 19705 155
rect 19760 175 19790 205
rect 19845 125 19875 155
rect 19930 175 19960 205
rect 20015 125 20045 155
rect 20100 175 20130 205
rect 20185 125 20215 155
rect 20270 175 20300 205
rect 20355 125 20385 155
rect 20440 175 20470 205
rect 20525 125 20555 155
rect 20610 175 20640 205
rect 20695 125 20725 155
rect 20780 175 20810 205
rect 20865 125 20895 155
rect 20950 175 20980 205
rect 21035 125 21065 155
rect 21120 175 21150 205
rect 21205 125 21235 155
rect 21290 175 21320 205
rect 21375 125 21405 155
rect 21460 175 21490 205
rect 21545 125 21575 155
rect 21630 175 21660 205
rect 21715 125 21745 155
rect 21800 175 21830 205
rect 21885 125 21915 155
rect 21970 175 22000 205
rect 22055 125 22085 155
rect 22140 175 22170 205
rect 22225 125 22255 155
rect 22310 175 22340 205
rect 22395 125 22425 155
rect 22480 175 22510 205
rect 22565 125 22595 155
rect 22650 175 22680 205
rect 22735 125 22765 155
rect 22820 175 22850 205
rect 22905 125 22935 155
rect 22990 175 23020 205
rect 23075 125 23105 155
rect 23160 175 23190 205
rect 23245 125 23275 155
rect 23330 175 23360 205
rect 23415 125 23445 155
rect 23500 175 23530 205
rect 23585 125 23615 155
rect 23670 175 23700 205
rect 23755 125 23785 155
rect 23840 175 23870 205
rect 23925 125 23955 155
rect 24010 175 24040 205
rect 24095 125 24125 155
rect 24180 175 24210 205
rect 24265 125 24295 155
rect 24350 175 24380 205
rect 24435 125 24465 155
rect 24520 175 24550 205
rect 24605 125 24635 155
rect 24690 175 24720 205
rect 24775 125 24805 155
rect 24860 175 24890 205
rect 24945 125 24975 155
rect 25030 175 25060 205
rect 25115 125 25145 155
rect 25200 175 25230 205
rect 25285 125 25315 155
rect 25370 175 25400 205
rect 25455 125 25485 155
rect 25540 175 25570 205
rect 25625 125 25655 155
rect 25710 175 25740 205
rect 25795 125 25825 155
rect 25880 175 25910 205
rect 25965 125 25995 155
rect 26050 175 26080 205
rect 26135 125 26165 155
rect 26220 175 26250 205
rect 26305 125 26335 155
rect 26390 175 26420 205
rect 26475 125 26505 155
rect 26560 175 26590 205
rect 26645 125 26675 155
rect 26730 175 26760 205
rect 26815 125 26845 155
rect 26900 175 26930 205
rect 26985 125 27015 155
rect 27070 175 27100 205
rect 27155 125 27185 155
rect 27240 175 27270 205
rect 27325 125 27355 155
rect 27410 175 27440 205
rect 27495 125 27525 155
rect 27580 175 27610 205
rect 27665 125 27695 155
rect 27750 175 27780 205
rect 27835 125 27865 155
rect 27920 175 27950 205
rect 28005 125 28035 155
rect 28090 175 28120 205
rect 28175 125 28205 155
rect 28260 175 28290 205
rect 28345 125 28375 155
rect 28430 175 28460 205
rect 28515 125 28545 155
rect 28600 175 28630 205
rect 28685 125 28715 155
rect 28770 175 28800 205
rect 28855 125 28885 155
rect 28940 175 28970 205
rect 29025 125 29055 155
rect 29110 175 29140 205
rect 29195 125 29225 155
rect 29280 175 29310 205
rect 29365 125 29395 155
rect 29450 175 29480 205
rect 29535 125 29565 155
rect 29620 175 29650 205
rect 35 15 65 55
rect 225 10 255 40
rect 310 10 340 40
rect 395 10 425 40
rect 480 10 510 40
rect 565 10 595 40
rect 760 10 790 40
rect 845 10 875 40
rect 930 10 960 40
rect 1015 10 1045 40
rect 1100 10 1130 40
rect 1185 10 1215 40
rect 1270 10 1300 40
rect 1355 10 1385 40
rect 1440 10 1470 40
rect 1525 10 1555 40
rect 1610 10 1640 40
rect 1695 10 1725 40
rect 1780 10 1810 40
rect 1865 10 1895 40
rect 1950 10 1980 40
rect 2035 10 2065 40
rect 2120 10 2150 40
rect 2270 10 2300 40
rect 2355 10 2385 40
rect 2440 10 2470 40
rect 2525 10 2555 40
rect 2610 10 2640 40
rect 2695 10 2725 40
rect 2780 10 2810 40
rect 2865 10 2895 40
rect 2950 10 2980 40
rect 3035 10 3065 40
rect 3120 10 3150 40
rect 3205 10 3235 40
rect 3290 10 3320 40
rect 3375 10 3405 40
rect 3460 10 3490 40
rect 3545 10 3575 40
rect 3630 10 3660 40
rect 3715 10 3745 40
rect 3800 10 3830 40
rect 3885 10 3915 40
rect 3970 10 4000 40
rect 4055 10 4085 40
rect 4140 10 4170 40
rect 4225 10 4255 40
rect 4310 10 4340 40
rect 4395 10 4425 40
rect 4480 10 4510 40
rect 4565 10 4595 40
rect 4650 10 4680 40
rect 4735 10 4765 40
rect 4820 10 4850 40
rect 4905 10 4935 40
rect 4990 10 5020 40
rect 5075 10 5105 40
rect 5160 10 5190 40
rect 5245 10 5275 40
rect 5330 10 5360 40
rect 5415 10 5445 40
rect 5500 10 5530 40
rect 5585 10 5615 40
rect 5670 10 5700 40
rect 5755 10 5785 40
rect 5840 10 5870 40
rect 5925 10 5955 40
rect 6010 10 6040 40
rect 6095 10 6125 40
rect 6180 10 6210 40
rect 6265 10 6295 40
rect 6350 10 6380 40
rect 6435 10 6465 40
rect 6520 10 6550 40
rect 6605 10 6635 40
rect 6690 10 6720 40
rect 6775 10 6805 40
rect 6860 10 6890 40
rect 6945 10 6975 40
rect 7030 10 7060 40
rect 7115 10 7145 40
rect 7200 10 7230 40
rect 7285 10 7315 40
rect 7370 10 7400 40
rect 7455 10 7485 40
rect 7540 10 7570 40
rect 7625 10 7655 40
rect 7710 10 7740 40
rect 7860 10 7890 40
rect 7945 10 7975 40
rect 8030 10 8060 40
rect 8115 10 8145 40
rect 8200 10 8230 40
rect 8285 10 8315 40
rect 8370 10 8400 40
rect 8455 10 8485 40
rect 8540 10 8570 40
rect 8625 10 8655 40
rect 8710 10 8740 40
rect 8795 10 8825 40
rect 8880 10 8910 40
rect 8965 10 8995 40
rect 9050 10 9080 40
rect 9135 10 9165 40
rect 9220 10 9250 40
rect 9305 10 9335 40
rect 9390 10 9420 40
rect 9475 10 9505 40
rect 9560 10 9590 40
rect 9645 10 9675 40
rect 9730 10 9760 40
rect 9815 10 9845 40
rect 9900 10 9930 40
rect 9985 10 10015 40
rect 10070 10 10100 40
rect 10155 10 10185 40
rect 10240 10 10270 40
rect 10325 10 10355 40
rect 10410 10 10440 40
rect 10495 10 10525 40
rect 10580 10 10610 40
rect 10665 10 10695 40
rect 10750 10 10780 40
rect 10835 10 10865 40
rect 10920 10 10950 40
rect 11005 10 11035 40
rect 11090 10 11120 40
rect 11175 10 11205 40
rect 11260 10 11290 40
rect 11345 10 11375 40
rect 11430 10 11460 40
rect 11515 10 11545 40
rect 11600 10 11630 40
rect 11685 10 11715 40
rect 11770 10 11800 40
rect 11855 10 11885 40
rect 11940 10 11970 40
rect 12025 10 12055 40
rect 12110 10 12140 40
rect 12195 10 12225 40
rect 12280 10 12310 40
rect 12365 10 12395 40
rect 12450 10 12480 40
rect 12535 10 12565 40
rect 12620 10 12650 40
rect 12705 10 12735 40
rect 12790 10 12820 40
rect 12875 10 12905 40
rect 12960 10 12990 40
rect 13045 10 13075 40
rect 13130 10 13160 40
rect 13215 10 13245 40
rect 13300 10 13330 40
rect 13385 10 13415 40
rect 13470 10 13500 40
rect 13555 10 13585 40
rect 13640 10 13670 40
rect 13725 10 13755 40
rect 13810 10 13840 40
rect 13895 10 13925 40
rect 13980 10 14010 40
rect 14065 10 14095 40
rect 14150 10 14180 40
rect 14235 10 14265 40
rect 14320 10 14350 40
rect 14405 10 14435 40
rect 14490 10 14520 40
rect 14575 10 14605 40
rect 14660 10 14690 40
rect 14745 10 14775 40
rect 14830 10 14860 40
rect 14915 10 14945 40
rect 15000 10 15030 40
rect 15085 10 15115 40
rect 15170 10 15200 40
rect 15255 10 15285 40
rect 15340 10 15370 40
rect 15425 10 15455 40
rect 15510 10 15540 40
rect 15595 10 15625 40
rect 15680 10 15710 40
rect 15765 10 15795 40
rect 15850 10 15880 40
rect 15935 10 15965 40
rect 16020 10 16050 40
rect 16105 10 16135 40
rect 16190 10 16220 40
rect 16275 10 16305 40
rect 16360 10 16390 40
rect 16445 10 16475 40
rect 16530 10 16560 40
rect 16615 10 16645 40
rect 16700 10 16730 40
rect 16785 10 16815 40
rect 16870 10 16900 40
rect 16955 10 16985 40
rect 17040 10 17070 40
rect 17125 10 17155 40
rect 17210 10 17240 40
rect 17295 10 17325 40
rect 17380 10 17410 40
rect 17465 10 17495 40
rect 17550 10 17580 40
rect 17635 10 17665 40
rect 17720 10 17750 40
rect 17805 10 17835 40
rect 17890 10 17920 40
rect 17975 10 18005 40
rect 18060 10 18090 40
rect 18145 10 18175 40
rect 18230 10 18260 40
rect 18315 10 18345 40
rect 18400 10 18430 40
rect 18485 10 18515 40
rect 18570 10 18600 40
rect 18655 10 18685 40
rect 18740 10 18770 40
rect 18825 10 18855 40
rect 18910 10 18940 40
rect 18995 10 19025 40
rect 19080 10 19110 40
rect 19165 10 19195 40
rect 19250 10 19280 40
rect 19335 10 19365 40
rect 19420 10 19450 40
rect 19505 10 19535 40
rect 19590 10 19620 40
rect 19675 10 19705 40
rect 19760 10 19790 40
rect 19845 10 19875 40
rect 19930 10 19960 40
rect 20015 10 20045 40
rect 20100 10 20130 40
rect 20185 10 20215 40
rect 20270 10 20300 40
rect 20355 10 20385 40
rect 20440 10 20470 40
rect 20525 10 20555 40
rect 20610 10 20640 40
rect 20695 10 20725 40
rect 20780 10 20810 40
rect 20865 10 20895 40
rect 20950 10 20980 40
rect 21035 10 21065 40
rect 21120 10 21150 40
rect 21205 10 21235 40
rect 21290 10 21320 40
rect 21375 10 21405 40
rect 21460 10 21490 40
rect 21545 10 21575 40
rect 21630 10 21660 40
rect 21715 10 21745 40
rect 21800 10 21830 40
rect 21885 10 21915 40
rect 21970 10 22000 40
rect 22055 10 22085 40
rect 22140 10 22170 40
rect 22225 10 22255 40
rect 22310 10 22340 40
rect 22395 10 22425 40
rect 22480 10 22510 40
rect 22565 10 22595 40
rect 22650 10 22680 40
rect 22735 10 22765 40
rect 22820 10 22850 40
rect 22905 10 22935 40
rect 22990 10 23020 40
rect 23075 10 23105 40
rect 23160 10 23190 40
rect 23245 10 23275 40
rect 23330 10 23360 40
rect 23415 10 23445 40
rect 23500 10 23530 40
rect 23585 10 23615 40
rect 23670 10 23700 40
rect 23755 10 23785 40
rect 23840 10 23870 40
rect 23925 10 23955 40
rect 24010 10 24040 40
rect 24095 10 24125 40
rect 24180 10 24210 40
rect 24265 10 24295 40
rect 24350 10 24380 40
rect 24435 10 24465 40
rect 24520 10 24550 40
rect 24605 10 24635 40
rect 24690 10 24720 40
rect 24775 10 24805 40
rect 24860 10 24890 40
rect 24945 10 24975 40
rect 25030 10 25060 40
rect 25115 10 25145 40
rect 25200 10 25230 40
rect 25285 10 25315 40
rect 25370 10 25400 40
rect 25455 10 25485 40
rect 25540 10 25570 40
rect 25625 10 25655 40
rect 25710 10 25740 40
rect 25795 10 25825 40
rect 25880 10 25910 40
rect 25965 10 25995 40
rect 26050 10 26080 40
rect 26135 10 26165 40
rect 26220 10 26250 40
rect 26305 10 26335 40
rect 26390 10 26420 40
rect 26475 10 26505 40
rect 26560 10 26590 40
rect 26645 10 26675 40
rect 26730 10 26760 40
rect 26815 10 26845 40
rect 26900 10 26930 40
rect 26985 10 27015 40
rect 27070 10 27100 40
rect 27155 10 27185 40
rect 27240 10 27270 40
rect 27325 10 27355 40
rect 27410 10 27440 40
rect 27495 10 27525 40
rect 27580 10 27610 40
rect 27665 10 27695 40
rect 27750 10 27780 40
rect 27835 10 27865 40
rect 27920 10 27950 40
rect 28005 10 28035 40
rect 28090 10 28120 40
rect 28175 10 28205 40
rect 28260 10 28290 40
rect 28345 10 28375 40
rect 28430 10 28460 40
rect 28515 10 28545 40
rect 28600 10 28630 40
rect 28685 10 28715 40
rect 28770 10 28800 40
rect 28855 10 28885 40
rect 28940 10 28970 40
rect 29025 10 29055 40
rect 29110 10 29140 40
rect 29195 10 29225 40
rect 29280 10 29310 40
rect 29365 10 29395 40
rect 29450 10 29480 40
rect 29535 10 29565 40
rect 29620 10 29650 40
rect 100 -60 130 -30
rect 265 -60 300 -30
rect 350 -60 385 -30
rect 435 -60 470 -30
rect 520 -60 555 -30
rect 800 -60 835 -30
rect 885 -60 920 -30
rect 970 -60 1005 -30
rect 1055 -60 1090 -30
rect 1140 -60 1175 -30
rect 1225 -60 1260 -30
rect 1310 -60 1345 -30
rect 1395 -60 1430 -30
rect 1480 -60 1515 -30
rect 1565 -60 1600 -30
rect 1650 -60 1685 -30
rect 1735 -60 1770 -30
rect 1820 -60 1855 -30
rect 1905 -60 1940 -30
rect 1990 -60 2025 -30
rect 2075 -60 2110 -30
rect 2310 -60 2345 -30
rect 2395 -60 2430 -30
rect 2480 -60 2515 -30
rect 2565 -60 2600 -30
rect 2650 -60 2685 -30
rect 2735 -60 2770 -30
rect 2820 -60 2855 -30
rect 2905 -60 2940 -30
rect 2990 -60 3025 -30
rect 3075 -60 3110 -30
rect 3160 -60 3195 -30
rect 3245 -60 3280 -30
rect 3330 -60 3365 -30
rect 3415 -60 3450 -30
rect 3500 -60 3535 -30
rect 3585 -60 3620 -30
rect 3670 -60 3705 -30
rect 3755 -60 3790 -30
rect 3840 -60 3875 -30
rect 3925 -60 3960 -30
rect 4010 -60 4045 -30
rect 4095 -60 4130 -30
rect 4180 -60 4215 -30
rect 4265 -60 4300 -30
rect 4350 -60 4385 -30
rect 4435 -60 4470 -30
rect 4520 -60 4555 -30
rect 4605 -60 4640 -30
rect 4690 -60 4725 -30
rect 4775 -60 4810 -30
rect 4860 -60 4895 -30
rect 4945 -60 4980 -30
rect 5030 -60 5065 -30
rect 5115 -60 5150 -30
rect 5200 -60 5235 -30
rect 5285 -60 5320 -30
rect 5370 -60 5405 -30
rect 5455 -60 5490 -30
rect 5540 -60 5575 -30
rect 5625 -60 5660 -30
rect 5710 -60 5745 -30
rect 5795 -60 5830 -30
rect 5880 -60 5915 -30
rect 5965 -60 6000 -30
rect 6050 -60 6085 -30
rect 6135 -60 6170 -30
rect 6220 -60 6255 -30
rect 6305 -60 6340 -30
rect 6390 -60 6425 -30
rect 6475 -60 6510 -30
rect 6560 -60 6595 -30
rect 6645 -60 6680 -30
rect 6730 -60 6765 -30
rect 6815 -60 6850 -30
rect 6900 -60 6935 -30
rect 6985 -60 7020 -30
rect 7070 -60 7105 -30
rect 7155 -60 7190 -30
rect 7240 -60 7275 -30
rect 7325 -60 7360 -30
rect 7410 -60 7445 -30
rect 7495 -60 7530 -30
rect 7580 -60 7615 -30
rect 7665 -60 7700 -30
rect 7900 -60 7935 -30
rect 7985 -60 8020 -30
rect 8070 -60 8105 -30
rect 8155 -60 8190 -30
rect 8240 -60 8275 -30
rect 8325 -60 8360 -30
rect 8410 -60 8445 -30
rect 8495 -60 8530 -30
rect 8580 -60 8615 -30
rect 8665 -60 8700 -30
rect 8750 -60 8785 -30
rect 8835 -60 8870 -30
rect 8920 -60 8955 -30
rect 9005 -60 9040 -30
rect 9090 -60 9125 -30
rect 9175 -60 9210 -30
rect 9260 -60 9295 -30
rect 9345 -60 9380 -30
rect 9430 -60 9465 -30
rect 9515 -60 9550 -30
rect 9600 -60 9635 -30
rect 9685 -60 9720 -30
rect 9770 -60 9805 -30
rect 9855 -60 9890 -30
rect 9940 -60 9975 -30
rect 10025 -60 10060 -30
rect 10110 -60 10145 -30
rect 10195 -60 10230 -30
rect 10280 -60 10315 -30
rect 10365 -60 10400 -30
rect 10450 -60 10485 -30
rect 10535 -60 10570 -30
rect 10620 -60 10655 -30
rect 10705 -60 10740 -30
rect 10790 -60 10825 -30
rect 10875 -60 10910 -30
rect 10960 -60 10995 -30
rect 11045 -60 11080 -30
rect 11130 -60 11165 -30
rect 11215 -60 11250 -30
rect 11300 -60 11335 -30
rect 11385 -60 11420 -30
rect 11470 -60 11505 -30
rect 11555 -60 11590 -30
rect 11640 -60 11675 -30
rect 11725 -60 11760 -30
rect 11810 -60 11845 -30
rect 11895 -60 11930 -30
rect 11980 -60 12015 -30
rect 12065 -60 12100 -30
rect 12150 -60 12185 -30
rect 12235 -60 12270 -30
rect 12320 -60 12355 -30
rect 12405 -60 12440 -30
rect 12490 -60 12525 -30
rect 12575 -60 12610 -30
rect 12660 -60 12695 -30
rect 12745 -60 12780 -30
rect 12830 -60 12865 -30
rect 12915 -60 12950 -30
rect 13000 -60 13035 -30
rect 13085 -60 13120 -30
rect 13170 -60 13205 -30
rect 13255 -60 13290 -30
rect 13340 -60 13375 -30
rect 13425 -60 13460 -30
rect 13510 -60 13545 -30
rect 13595 -60 13630 -30
rect 13680 -60 13715 -30
rect 13765 -60 13800 -30
rect 13850 -60 13885 -30
rect 13935 -60 13970 -30
rect 14020 -60 14055 -30
rect 14105 -60 14140 -30
rect 14190 -60 14225 -30
rect 14275 -60 14310 -30
rect 14360 -60 14395 -30
rect 14445 -60 14480 -30
rect 14530 -60 14565 -30
rect 14615 -60 14650 -30
rect 14700 -60 14735 -30
rect 14785 -60 14820 -30
rect 14870 -60 14905 -30
rect 14955 -60 14990 -30
rect 15040 -60 15075 -30
rect 15125 -60 15160 -30
rect 15210 -60 15245 -30
rect 15295 -60 15330 -30
rect 15380 -60 15415 -30
rect 15465 -60 15500 -30
rect 15550 -60 15585 -30
rect 15635 -60 15670 -30
rect 15720 -60 15755 -30
rect 15805 -60 15840 -30
rect 15890 -60 15925 -30
rect 15975 -60 16010 -30
rect 16060 -60 16095 -30
rect 16145 -60 16180 -30
rect 16230 -60 16265 -30
rect 16315 -60 16350 -30
rect 16400 -60 16435 -30
rect 16485 -60 16520 -30
rect 16570 -60 16605 -30
rect 16655 -60 16690 -30
rect 16740 -60 16775 -30
rect 16825 -60 16860 -30
rect 16910 -60 16945 -30
rect 16995 -60 17030 -30
rect 17080 -60 17115 -30
rect 17165 -60 17200 -30
rect 17250 -60 17285 -30
rect 17335 -60 17370 -30
rect 17420 -60 17455 -30
rect 17505 -60 17540 -30
rect 17590 -60 17625 -30
rect 17675 -60 17710 -30
rect 17760 -60 17795 -30
rect 17845 -60 17880 -30
rect 17930 -60 17965 -30
rect 18015 -60 18050 -30
rect 18100 -60 18135 -30
rect 18185 -60 18220 -30
rect 18270 -60 18305 -30
rect 18355 -60 18390 -30
rect 18440 -60 18475 -30
rect 18525 -60 18560 -30
rect 18610 -60 18645 -30
rect 18695 -60 18730 -30
rect 18780 -60 18815 -30
rect 18865 -60 18900 -30
rect 18950 -60 18985 -30
rect 19035 -60 19070 -30
rect 19120 -60 19155 -30
rect 19205 -60 19240 -30
rect 19290 -60 19325 -30
rect 19375 -60 19410 -30
rect 19460 -60 19495 -30
rect 19545 -60 19580 -30
rect 19630 -60 19665 -30
rect 19715 -60 19750 -30
rect 19800 -60 19835 -30
rect 19885 -60 19920 -30
rect 19970 -60 20005 -30
rect 20055 -60 20090 -30
rect 20140 -60 20175 -30
rect 20225 -60 20260 -30
rect 20310 -60 20345 -30
rect 20395 -60 20430 -30
rect 20480 -60 20515 -30
rect 20565 -60 20600 -30
rect 20650 -60 20685 -30
rect 20735 -60 20770 -30
rect 20820 -60 20855 -30
rect 20905 -60 20940 -30
rect 20990 -60 21025 -30
rect 21075 -60 21110 -30
rect 21160 -60 21195 -30
rect 21245 -60 21280 -30
rect 21330 -60 21365 -30
rect 21415 -60 21450 -30
rect 21500 -60 21535 -30
rect 21585 -60 21620 -30
rect 21670 -60 21705 -30
rect 21755 -60 21790 -30
rect 21840 -60 21875 -30
rect 21925 -60 21960 -30
rect 22010 -60 22045 -30
rect 22095 -60 22130 -30
rect 22180 -60 22215 -30
rect 22265 -60 22300 -30
rect 22350 -60 22385 -30
rect 22435 -60 22470 -30
rect 22520 -60 22555 -30
rect 22605 -60 22640 -30
rect 22690 -60 22725 -30
rect 22775 -60 22810 -30
rect 22860 -60 22895 -30
rect 22945 -60 22980 -30
rect 23030 -60 23065 -30
rect 23115 -60 23150 -30
rect 23200 -60 23235 -30
rect 23285 -60 23320 -30
rect 23370 -60 23405 -30
rect 23455 -60 23490 -30
rect 23540 -60 23575 -30
rect 23625 -60 23660 -30
rect 23710 -60 23745 -30
rect 23795 -60 23830 -30
rect 23880 -60 23915 -30
rect 23965 -60 24000 -30
rect 24050 -60 24085 -30
rect 24135 -60 24170 -30
rect 24220 -60 24255 -30
rect 24305 -60 24340 -30
rect 24390 -60 24425 -30
rect 24475 -60 24510 -30
rect 24560 -60 24595 -30
rect 24645 -60 24680 -30
rect 24730 -60 24765 -30
rect 24815 -60 24850 -30
rect 24900 -60 24935 -30
rect 24985 -60 25020 -30
rect 25070 -60 25105 -30
rect 25155 -60 25190 -30
rect 25240 -60 25275 -30
rect 25325 -60 25360 -30
rect 25410 -60 25445 -30
rect 25495 -60 25530 -30
rect 25580 -60 25615 -30
rect 25665 -60 25700 -30
rect 25750 -60 25785 -30
rect 25835 -60 25870 -30
rect 25920 -60 25955 -30
rect 26005 -60 26040 -30
rect 26090 -60 26125 -30
rect 26175 -60 26210 -30
rect 26260 -60 26295 -30
rect 26345 -60 26380 -30
rect 26430 -60 26465 -30
rect 26515 -60 26550 -30
rect 26600 -60 26635 -30
rect 26685 -60 26720 -30
rect 26770 -60 26805 -30
rect 26855 -60 26890 -30
rect 26940 -60 26975 -30
rect 27025 -60 27060 -30
rect 27110 -60 27145 -30
rect 27195 -60 27230 -30
rect 27280 -60 27315 -30
rect 27365 -60 27400 -30
rect 27450 -60 27485 -30
rect 27535 -60 27570 -30
rect 27620 -60 27655 -30
rect 27705 -60 27740 -30
rect 27790 -60 27825 -30
rect 27875 -60 27910 -30
rect 27960 -60 27995 -30
rect 28045 -60 28080 -30
rect 28130 -60 28165 -30
rect 28215 -60 28250 -30
rect 28300 -60 28335 -30
rect 28385 -60 28420 -30
rect 28470 -60 28505 -30
rect 28555 -60 28590 -30
rect 28640 -60 28675 -30
rect 28725 -60 28760 -30
rect 28810 -60 28845 -30
rect 28895 -60 28930 -30
rect 28980 -60 29015 -30
rect 29065 -60 29100 -30
rect 29150 -60 29185 -30
rect 29235 -60 29270 -30
rect 29320 -60 29355 -30
rect 29405 -60 29440 -30
rect 29490 -60 29525 -30
rect 29575 -60 29610 -30
rect 115 -295 150 -265
rect 200 -295 235 -265
rect 285 -295 320 -265
rect 370 -295 405 -265
rect 455 -295 490 -265
rect 540 -295 575 -265
rect 625 -295 660 -265
rect 710 -295 745 -265
rect 795 -295 830 -265
rect 880 -295 915 -265
rect 965 -295 1000 -265
rect 1050 -295 1085 -265
rect 1135 -295 1170 -265
rect 1220 -295 1255 -265
rect 1305 -295 1340 -265
rect 1390 -295 1425 -265
rect 1475 -295 1510 -265
rect 1560 -295 1595 -265
rect 1645 -295 1680 -265
rect 1730 -295 1765 -265
rect 1815 -295 1850 -265
rect 1900 -295 1935 -265
rect 1985 -295 2020 -265
rect 2070 -295 2105 -265
rect 2155 -295 2190 -265
rect 2240 -295 2275 -265
rect 2325 -295 2360 -265
rect 2410 -295 2445 -265
rect 2495 -295 2530 -265
rect 2580 -295 2615 -265
rect 2665 -295 2700 -265
rect 2750 -295 2785 -265
rect 2835 -295 2870 -265
rect 2920 -295 2955 -265
rect 3005 -295 3040 -265
rect 3090 -295 3125 -265
rect 3175 -295 3210 -265
rect 3260 -295 3295 -265
rect 3345 -295 3380 -265
rect 3430 -295 3465 -265
rect 3515 -295 3550 -265
rect 3600 -295 3635 -265
rect 3685 -295 3720 -265
rect 3770 -295 3805 -265
rect 3855 -295 3890 -265
rect 3940 -295 3975 -265
rect 4025 -295 4060 -265
rect 4110 -295 4145 -265
rect 4195 -295 4230 -265
rect 4280 -295 4315 -265
rect 4365 -295 4400 -265
rect 4450 -295 4485 -265
rect 4535 -295 4570 -265
rect 4620 -295 4655 -265
rect 4705 -295 4740 -265
rect 4790 -295 4825 -265
rect 4875 -295 4910 -265
rect 4960 -295 4995 -265
rect 5045 -295 5080 -265
rect 5130 -295 5165 -265
rect 5215 -295 5250 -265
rect 5300 -295 5335 -265
rect 5385 -295 5420 -265
rect 5470 -295 5505 -265
rect 5555 -295 5590 -265
rect 5640 -295 5675 -265
rect 5725 -295 5760 -265
rect 5810 -295 5845 -265
rect 5895 -295 5930 -265
rect 5980 -295 6015 -265
rect 6065 -295 6100 -265
rect 6150 -295 6185 -265
rect 6235 -295 6270 -265
rect 6320 -295 6355 -265
rect 6405 -295 6440 -265
rect 6490 -295 6525 -265
rect 6575 -295 6610 -265
rect 6660 -295 6695 -265
rect 6745 -295 6780 -265
rect 6830 -295 6865 -265
rect 6915 -295 6950 -265
rect 7000 -295 7035 -265
rect 7085 -295 7120 -265
rect 7170 -295 7205 -265
rect 7255 -295 7290 -265
rect 7340 -295 7375 -265
rect 7425 -295 7460 -265
rect 7510 -295 7545 -265
rect 7595 -295 7630 -265
rect 7680 -295 7715 -265
rect 7765 -295 7800 -265
rect 7850 -295 7885 -265
rect 7935 -295 7970 -265
rect 8020 -295 8055 -265
rect 8105 -295 8140 -265
rect 8190 -295 8225 -265
rect 8275 -295 8310 -265
rect 8360 -295 8395 -265
rect 8445 -295 8480 -265
rect 8530 -295 8565 -265
rect 8615 -295 8650 -265
rect 8700 -295 8735 -265
rect 8785 -295 8820 -265
rect 8870 -295 8905 -265
rect 8955 -295 8990 -265
rect 9040 -295 9075 -265
rect 9125 -295 9160 -265
rect 9210 -295 9245 -265
rect 9295 -295 9330 -265
rect 9380 -295 9415 -265
rect 9465 -295 9500 -265
rect 9550 -295 9585 -265
rect 9635 -295 9670 -265
rect 9720 -295 9755 -265
rect 9805 -295 9840 -265
rect 9890 -295 9925 -265
rect 9975 -295 10010 -265
rect 10060 -295 10095 -265
rect 10145 -295 10180 -265
rect 10230 -295 10265 -265
rect 10315 -295 10350 -265
rect 10400 -295 10435 -265
rect 10485 -295 10520 -265
rect 10570 -295 10605 -265
rect 10655 -295 10690 -265
rect 10740 -295 10775 -265
rect 10825 -295 10860 -265
rect 10910 -295 10945 -265
rect 10995 -295 11030 -265
rect 11080 -295 11115 -265
rect 11165 -295 11200 -265
rect 11250 -295 11285 -265
rect 11335 -295 11370 -265
rect 11420 -295 11455 -265
rect 11505 -295 11540 -265
rect 11590 -295 11625 -265
rect 11675 -295 11710 -265
rect 11760 -295 11795 -265
rect 11845 -295 11880 -265
rect 11930 -295 11965 -265
rect 12015 -295 12050 -265
rect 12100 -295 12135 -265
rect 12185 -295 12220 -265
rect 12270 -295 12305 -265
rect 12355 -295 12390 -265
rect 12440 -295 12475 -265
rect 12525 -295 12560 -265
rect 12610 -295 12645 -265
rect 12695 -295 12730 -265
rect 12780 -295 12815 -265
rect 12865 -295 12900 -265
rect 12950 -295 12985 -265
rect 13035 -295 13070 -265
rect 13120 -295 13155 -265
rect 13205 -295 13240 -265
rect 13290 -295 13325 -265
rect 13375 -295 13410 -265
rect 13460 -295 13495 -265
rect 13545 -295 13580 -265
rect 13630 -295 13665 -265
rect 13715 -295 13750 -265
rect 13800 -295 13835 -265
rect 13885 -295 13920 -265
rect 13970 -295 14005 -265
rect 14055 -295 14090 -265
rect 14140 -295 14175 -265
rect 14225 -295 14260 -265
rect 14310 -295 14345 -265
rect 14395 -295 14430 -265
rect 14480 -295 14515 -265
rect 14565 -295 14600 -265
rect 14650 -295 14685 -265
rect 14735 -295 14770 -265
rect 14820 -295 14855 -265
rect 14905 -295 14940 -265
rect 14990 -295 15025 -265
rect 15075 -295 15110 -265
rect 15160 -295 15195 -265
rect 15245 -295 15280 -265
rect 15330 -295 15365 -265
rect 15415 -295 15450 -265
rect 15500 -295 15535 -265
rect 15585 -295 15620 -265
rect 15670 -295 15705 -265
rect 15755 -295 15790 -265
rect 15840 -295 15875 -265
rect 15925 -295 15960 -265
rect 16010 -295 16045 -265
rect 16095 -295 16130 -265
rect 16180 -295 16215 -265
rect 16265 -295 16300 -265
rect 16350 -295 16385 -265
rect 16435 -295 16470 -265
rect 16520 -295 16555 -265
rect 16605 -295 16640 -265
rect 16690 -295 16725 -265
rect 16775 -295 16810 -265
rect 16860 -295 16895 -265
rect 16945 -295 16980 -265
rect 17030 -295 17065 -265
rect 17115 -295 17150 -265
rect 17200 -295 17235 -265
rect 17285 -295 17320 -265
rect 17370 -295 17405 -265
rect 17455 -295 17490 -265
rect 17540 -295 17575 -265
rect 17625 -295 17660 -265
rect 17710 -295 17745 -265
rect 17795 -295 17830 -265
rect 17880 -295 17915 -265
rect 17965 -295 18000 -265
rect 18050 -295 18085 -265
rect 18135 -295 18170 -265
rect 18220 -295 18255 -265
rect 18305 -295 18340 -265
rect 18390 -295 18425 -265
rect 18475 -295 18510 -265
rect 18560 -295 18595 -265
rect 18645 -295 18680 -265
rect 18730 -295 18765 -265
rect 18815 -295 18850 -265
rect 18900 -295 18935 -265
rect 18985 -295 19020 -265
rect 19070 -295 19105 -265
rect 19155 -295 19190 -265
rect 19240 -295 19275 -265
rect 19325 -295 19360 -265
rect 19410 -295 19445 -265
rect 19495 -295 19530 -265
rect 19580 -295 19615 -265
rect 19665 -295 19700 -265
rect 19750 -295 19785 -265
rect 19835 -295 19870 -265
rect 19920 -295 19955 -265
rect 20005 -295 20040 -265
rect 20090 -295 20125 -265
rect 20175 -295 20210 -265
rect 20260 -295 20295 -265
rect 20345 -295 20380 -265
rect 20430 -295 20465 -265
rect 20515 -295 20550 -265
rect 20600 -295 20635 -265
rect 20685 -295 20720 -265
rect 20770 -295 20805 -265
rect 20855 -295 20890 -265
rect 20940 -295 20975 -265
rect 21025 -295 21060 -265
rect 21110 -295 21145 -265
rect 21195 -295 21230 -265
rect 21280 -295 21315 -265
rect 21365 -295 21400 -265
rect 21450 -295 21485 -265
rect 21535 -295 21570 -265
rect 21620 -295 21655 -265
rect 21705 -295 21740 -265
rect 21790 -295 21825 -265
rect 21875 -295 21910 -265
rect 21960 -295 21995 -265
rect 22045 -295 22080 -265
rect 22130 -295 22165 -265
rect 22215 -295 22250 -265
rect 22300 -295 22335 -265
rect 22385 -295 22420 -265
rect 22470 -295 22505 -265
rect 22555 -295 22590 -265
rect 22640 -295 22675 -265
rect 22725 -295 22760 -265
rect 22810 -295 22845 -265
rect 22895 -295 22930 -265
rect 22980 -295 23015 -265
rect 23065 -295 23100 -265
rect 23150 -295 23185 -265
rect 23235 -295 23270 -265
rect 23320 -295 23355 -265
rect 23405 -295 23440 -265
rect 23490 -295 23525 -265
rect 23575 -295 23610 -265
rect 23660 -295 23695 -265
rect 23745 -295 23780 -265
rect 23830 -295 23865 -265
rect 23915 -295 23950 -265
rect 24000 -295 24035 -265
rect 24085 -295 24120 -265
rect 24170 -295 24205 -265
rect 24255 -295 24290 -265
rect 24340 -295 24375 -265
rect 24425 -295 24460 -265
rect 24510 -295 24545 -265
rect 24595 -295 24630 -265
rect 24680 -295 24715 -265
rect 24765 -295 24800 -265
rect 24850 -295 24885 -265
rect 24935 -295 24970 -265
rect 25020 -295 25055 -265
rect 25105 -295 25140 -265
rect 25190 -295 25225 -265
rect 25275 -295 25310 -265
rect 25360 -295 25395 -265
rect 25445 -295 25480 -265
rect 25530 -295 25565 -265
rect 25615 -295 25650 -265
rect 25700 -295 25735 -265
rect 25785 -295 25820 -265
rect 25870 -295 25905 -265
rect 25955 -295 25990 -265
rect 26040 -295 26075 -265
rect 26125 -295 26160 -265
rect 26210 -295 26245 -265
rect 26295 -295 26330 -265
rect 26380 -295 26415 -265
rect 26465 -295 26500 -265
rect 26550 -295 26585 -265
rect 26635 -295 26670 -265
rect 26720 -295 26755 -265
rect 26805 -295 26840 -265
rect 26890 -295 26925 -265
rect 26975 -295 27010 -265
rect 27060 -295 27095 -265
rect 27145 -295 27180 -265
rect 27230 -295 27265 -265
rect 27315 -295 27350 -265
rect 27400 -295 27435 -265
rect 27485 -295 27520 -265
rect 27570 -295 27605 -265
rect 27655 -295 27690 -265
rect 27740 -295 27775 -265
rect 27825 -295 27860 -265
rect 27910 -295 27945 -265
rect 27995 -295 28030 -265
rect 28080 -295 28115 -265
rect 28165 -295 28200 -265
rect 28250 -295 28285 -265
rect 28335 -295 28370 -265
rect 28420 -295 28455 -265
rect 28505 -295 28540 -265
rect 28590 -295 28625 -265
rect 28675 -295 28710 -265
rect 28760 -295 28795 -265
rect 28845 -295 28880 -265
rect 28930 -295 28965 -265
rect 29015 -295 29050 -265
rect 29100 -295 29135 -265
rect 29185 -295 29220 -265
rect 29270 -295 29305 -265
rect 29355 -295 29390 -265
rect 29440 -295 29475 -265
rect 29525 -295 29560 -265
rect 29610 -295 29645 -265
rect 29695 -295 29730 -265
rect 29780 -295 29815 -265
rect 29865 -295 29900 -265
rect 29950 -295 29985 -265
rect 30035 -295 30070 -265
rect 30120 -295 30155 -265
rect 30205 -295 30240 -265
rect 30290 -295 30325 -265
rect 30375 -295 30410 -265
rect 30460 -295 30495 -265
rect 30545 -295 30580 -265
rect 30630 -295 30665 -265
rect 30715 -295 30750 -265
rect 30800 -295 30835 -265
rect 30885 -295 30920 -265
rect 30970 -295 31005 -265
rect 31055 -295 31090 -265
rect 31140 -295 31175 -265
rect 31225 -295 31260 -265
rect 31310 -295 31345 -265
rect 31395 -295 31430 -265
rect 31480 -295 31515 -265
rect 31565 -295 31600 -265
rect 31650 -295 31685 -265
rect 31735 -295 31770 -265
rect 31820 -295 31855 -265
rect 31905 -295 31940 -265
rect 31990 -295 32025 -265
rect 32075 -295 32110 -265
rect 32160 -295 32195 -265
rect 32245 -295 32280 -265
rect 32330 -295 32365 -265
rect 32415 -295 32450 -265
rect 32500 -295 32535 -265
rect 32585 -295 32620 -265
rect 32670 -295 32705 -265
rect 32755 -295 32790 -265
rect 32840 -295 32875 -265
rect 32925 -295 32960 -265
rect 33010 -295 33045 -265
rect 33095 -295 33130 -265
rect 33180 -295 33215 -265
rect 33265 -295 33300 -265
rect 33350 -295 33385 -265
rect 33435 -295 33470 -265
rect 33520 -295 33555 -265
rect 33605 -295 33640 -265
rect 33690 -295 33725 -265
rect 33775 -295 33810 -265
rect 33860 -295 33895 -265
rect 33945 -295 33980 -265
rect 34030 -295 34065 -265
rect 34115 -295 34150 -265
rect 34200 -295 34235 -265
rect 34285 -295 34320 -265
rect 34370 -295 34405 -265
rect 34455 -295 34490 -265
rect 34540 -295 34575 -265
rect 34625 -295 34660 -265
rect 34710 -295 34745 -265
rect 34795 -295 34830 -265
rect 34880 -295 34915 -265
rect 34965 -295 35000 -265
rect 35050 -295 35085 -265
rect 35135 -295 35170 -265
rect 35220 -295 35255 -265
rect 35305 -295 35340 -265
rect 35390 -295 35425 -265
rect 35475 -295 35510 -265
rect 35560 -295 35595 -265
rect 35645 -295 35680 -265
rect 35730 -295 35765 -265
rect 35815 -295 35850 -265
rect 35900 -295 35935 -265
rect 35985 -295 36020 -265
rect 36070 -295 36105 -265
rect 36155 -295 36190 -265
rect 36240 -295 36275 -265
rect 36325 -295 36360 -265
rect 36410 -295 36445 -265
rect 36495 -295 36530 -265
rect 36580 -295 36615 -265
rect 36665 -295 36700 -265
rect 36750 -295 36785 -265
rect 36835 -295 36870 -265
rect 36920 -295 36955 -265
rect 37005 -295 37040 -265
rect 37090 -295 37125 -265
rect 37175 -295 37210 -265
rect 37260 -295 37295 -265
rect 37345 -295 37380 -265
rect 37430 -295 37465 -265
rect 37515 -295 37550 -265
rect 37600 -295 37635 -265
rect 37685 -295 37720 -265
rect 37770 -295 37805 -265
rect 37855 -295 37890 -265
rect 37940 -295 37975 -265
rect 38025 -295 38060 -265
rect 38110 -295 38145 -265
rect 38195 -295 38230 -265
rect 38280 -295 38315 -265
rect 38365 -295 38400 -265
rect 38450 -295 38485 -265
rect 38535 -295 38570 -265
rect 38620 -295 38655 -265
rect 38705 -295 38740 -265
rect 38790 -295 38825 -265
rect 38875 -295 38910 -265
rect 38960 -295 38995 -265
rect 39045 -295 39080 -265
rect 39130 -295 39165 -265
rect 39215 -295 39250 -265
rect 39300 -295 39335 -265
rect 39385 -295 39420 -265
rect 39470 -295 39505 -265
rect 39555 -295 39590 -265
rect 39640 -295 39675 -265
rect 39725 -295 39760 -265
rect 39810 -295 39845 -265
rect 39895 -295 39930 -265
rect 39980 -295 40015 -265
rect 40065 -295 40100 -265
rect 40150 -295 40185 -265
rect 40235 -295 40270 -265
rect 40320 -295 40355 -265
rect 40405 -295 40440 -265
rect 40490 -295 40525 -265
rect 40575 -295 40610 -265
rect 40660 -295 40695 -265
rect 40745 -295 40780 -265
rect 40830 -295 40865 -265
rect 40915 -295 40950 -265
rect 41000 -295 41035 -265
rect 41085 -295 41120 -265
rect 41170 -295 41205 -265
rect 41255 -295 41290 -265
rect 41340 -295 41375 -265
rect 41425 -295 41460 -265
rect 41510 -295 41545 -265
rect 41595 -295 41630 -265
rect 41680 -295 41715 -265
rect 41765 -295 41800 -265
rect 41850 -295 41885 -265
rect 41935 -295 41970 -265
rect 42020 -295 42055 -265
rect 42105 -295 42140 -265
rect 42190 -295 42225 -265
rect 42275 -295 42310 -265
rect 42360 -295 42395 -265
rect 42445 -295 42480 -265
rect 42530 -295 42565 -265
rect 42615 -295 42650 -265
rect 42700 -295 42735 -265
rect 42785 -295 42820 -265
rect 42870 -295 42905 -265
rect 42955 -295 42990 -265
rect 43040 -295 43075 -265
rect 43125 -295 43160 -265
rect 43210 -295 43245 -265
rect 43295 -295 43330 -265
rect 43380 -295 43415 -265
rect 43465 -295 43500 -265
rect 43550 -295 43585 -265
rect 75 -365 105 -335
rect 160 -415 190 -385
rect 245 -365 275 -335
rect 330 -415 360 -385
rect 415 -365 445 -335
rect 500 -415 530 -385
rect 585 -365 615 -335
rect 670 -415 700 -385
rect 755 -365 785 -335
rect 840 -415 870 -385
rect 925 -365 955 -335
rect 1010 -415 1040 -385
rect 1095 -365 1125 -335
rect 1180 -415 1210 -385
rect 1265 -365 1295 -335
rect 1350 -415 1380 -385
rect 1435 -365 1465 -335
rect 1520 -415 1550 -385
rect 1605 -365 1635 -335
rect 1690 -415 1720 -385
rect 1775 -365 1805 -335
rect 1860 -415 1890 -385
rect 1945 -365 1975 -335
rect 2030 -415 2060 -385
rect 2115 -365 2145 -335
rect 2200 -415 2230 -385
rect 2285 -365 2315 -335
rect 2370 -415 2400 -385
rect 2455 -365 2485 -335
rect 2540 -415 2570 -385
rect 2625 -365 2655 -335
rect 2710 -415 2740 -385
rect 2795 -365 2825 -335
rect 2880 -415 2910 -385
rect 2965 -365 2995 -335
rect 3050 -415 3080 -385
rect 3135 -365 3165 -335
rect 3220 -415 3250 -385
rect 3305 -365 3335 -335
rect 3390 -415 3420 -385
rect 3475 -365 3505 -335
rect 3560 -415 3590 -385
rect 3645 -365 3675 -335
rect 3730 -415 3760 -385
rect 3815 -365 3845 -335
rect 3900 -415 3930 -385
rect 3985 -365 4015 -335
rect 4070 -415 4100 -385
rect 4155 -365 4185 -335
rect 4240 -415 4270 -385
rect 4325 -365 4355 -335
rect 4410 -415 4440 -385
rect 4495 -365 4525 -335
rect 4580 -415 4610 -385
rect 4665 -365 4695 -335
rect 4750 -415 4780 -385
rect 4835 -365 4865 -335
rect 4920 -415 4950 -385
rect 5005 -365 5035 -335
rect 5090 -415 5120 -385
rect 5175 -365 5205 -335
rect 5260 -415 5290 -385
rect 5345 -365 5375 -335
rect 5430 -415 5460 -385
rect 5515 -365 5545 -335
rect 5600 -415 5630 -385
rect 5685 -365 5715 -335
rect 5770 -415 5800 -385
rect 5855 -365 5885 -335
rect 5940 -415 5970 -385
rect 6025 -365 6055 -335
rect 6110 -415 6140 -385
rect 6195 -365 6225 -335
rect 6280 -415 6310 -385
rect 6365 -365 6395 -335
rect 6450 -415 6480 -385
rect 6535 -365 6565 -335
rect 6620 -415 6650 -385
rect 6705 -365 6735 -335
rect 6790 -415 6820 -385
rect 6875 -365 6905 -335
rect 6960 -415 6990 -385
rect 7045 -365 7075 -335
rect 7130 -415 7160 -385
rect 7215 -365 7245 -335
rect 7300 -415 7330 -385
rect 7385 -365 7415 -335
rect 7470 -415 7500 -385
rect 7555 -365 7585 -335
rect 7640 -415 7670 -385
rect 7725 -365 7755 -335
rect 7810 -415 7840 -385
rect 7895 -365 7925 -335
rect 7980 -415 8010 -385
rect 8065 -365 8095 -335
rect 8150 -415 8180 -385
rect 8235 -365 8265 -335
rect 8320 -415 8350 -385
rect 8405 -365 8435 -335
rect 8490 -415 8520 -385
rect 8575 -365 8605 -335
rect 8660 -415 8690 -385
rect 8745 -365 8775 -335
rect 8830 -415 8860 -385
rect 8915 -365 8945 -335
rect 9000 -415 9030 -385
rect 9085 -365 9115 -335
rect 9170 -415 9200 -385
rect 9255 -365 9285 -335
rect 9340 -415 9370 -385
rect 9425 -365 9455 -335
rect 9510 -415 9540 -385
rect 9595 -365 9625 -335
rect 9680 -415 9710 -385
rect 9765 -365 9795 -335
rect 9850 -415 9880 -385
rect 9935 -365 9965 -335
rect 10020 -415 10050 -385
rect 10105 -365 10135 -335
rect 10190 -415 10220 -385
rect 10275 -365 10305 -335
rect 10360 -415 10390 -385
rect 10445 -365 10475 -335
rect 10530 -415 10560 -385
rect 10615 -365 10645 -335
rect 10700 -415 10730 -385
rect 10785 -365 10815 -335
rect 10870 -415 10900 -385
rect 10955 -365 10985 -335
rect 11040 -415 11070 -385
rect 11125 -365 11155 -335
rect 11210 -415 11240 -385
rect 11295 -365 11325 -335
rect 11380 -415 11410 -385
rect 11465 -365 11495 -335
rect 11550 -415 11580 -385
rect 11635 -365 11665 -335
rect 11720 -415 11750 -385
rect 11805 -365 11835 -335
rect 11890 -415 11920 -385
rect 11975 -365 12005 -335
rect 12060 -415 12090 -385
rect 12145 -365 12175 -335
rect 12230 -415 12260 -385
rect 12315 -365 12345 -335
rect 12400 -415 12430 -385
rect 12485 -365 12515 -335
rect 12570 -415 12600 -385
rect 12655 -365 12685 -335
rect 12740 -415 12770 -385
rect 12825 -365 12855 -335
rect 12910 -415 12940 -385
rect 12995 -365 13025 -335
rect 13080 -415 13110 -385
rect 13165 -365 13195 -335
rect 13250 -415 13280 -385
rect 13335 -365 13365 -335
rect 13420 -415 13450 -385
rect 13505 -365 13535 -335
rect 13590 -415 13620 -385
rect 13675 -365 13705 -335
rect 13760 -415 13790 -385
rect 13845 -365 13875 -335
rect 13930 -415 13960 -385
rect 14015 -365 14045 -335
rect 14100 -415 14130 -385
rect 14185 -365 14215 -335
rect 14270 -415 14300 -385
rect 14355 -365 14385 -335
rect 14440 -415 14470 -385
rect 14525 -365 14555 -335
rect 14610 -415 14640 -385
rect 14695 -365 14725 -335
rect 14780 -415 14810 -385
rect 14865 -365 14895 -335
rect 14950 -415 14980 -385
rect 15035 -365 15065 -335
rect 15120 -415 15150 -385
rect 15205 -365 15235 -335
rect 15290 -415 15320 -385
rect 15375 -365 15405 -335
rect 15460 -415 15490 -385
rect 15545 -365 15575 -335
rect 15630 -415 15660 -385
rect 15715 -365 15745 -335
rect 15800 -415 15830 -385
rect 15885 -365 15915 -335
rect 15970 -415 16000 -385
rect 16055 -365 16085 -335
rect 16140 -415 16170 -385
rect 16225 -365 16255 -335
rect 16310 -415 16340 -385
rect 16395 -365 16425 -335
rect 16480 -415 16510 -385
rect 16565 -365 16595 -335
rect 16650 -415 16680 -385
rect 16735 -365 16765 -335
rect 16820 -415 16850 -385
rect 16905 -365 16935 -335
rect 16990 -415 17020 -385
rect 17075 -365 17105 -335
rect 17160 -415 17190 -385
rect 17245 -365 17275 -335
rect 17330 -415 17360 -385
rect 17415 -365 17445 -335
rect 17500 -415 17530 -385
rect 17585 -365 17615 -335
rect 17670 -415 17700 -385
rect 17755 -365 17785 -335
rect 17840 -415 17870 -385
rect 17925 -365 17955 -335
rect 18010 -415 18040 -385
rect 18095 -365 18125 -335
rect 18180 -415 18210 -385
rect 18265 -365 18295 -335
rect 18350 -415 18380 -385
rect 18435 -365 18465 -335
rect 18520 -415 18550 -385
rect 18605 -365 18635 -335
rect 18690 -415 18720 -385
rect 18775 -365 18805 -335
rect 18860 -415 18890 -385
rect 18945 -365 18975 -335
rect 19030 -415 19060 -385
rect 19115 -365 19145 -335
rect 19200 -415 19230 -385
rect 19285 -365 19315 -335
rect 19370 -415 19400 -385
rect 19455 -365 19485 -335
rect 19540 -415 19570 -385
rect 19625 -365 19655 -335
rect 19710 -415 19740 -385
rect 19795 -365 19825 -335
rect 19880 -415 19910 -385
rect 19965 -365 19995 -335
rect 20050 -415 20080 -385
rect 20135 -365 20165 -335
rect 20220 -415 20250 -385
rect 20305 -365 20335 -335
rect 20390 -415 20420 -385
rect 20475 -365 20505 -335
rect 20560 -415 20590 -385
rect 20645 -365 20675 -335
rect 20730 -415 20760 -385
rect 20815 -365 20845 -335
rect 20900 -415 20930 -385
rect 20985 -365 21015 -335
rect 21070 -415 21100 -385
rect 21155 -365 21185 -335
rect 21240 -415 21270 -385
rect 21325 -365 21355 -335
rect 21410 -415 21440 -385
rect 21495 -365 21525 -335
rect 21580 -415 21610 -385
rect 21665 -365 21695 -335
rect 21750 -415 21780 -385
rect 21835 -365 21865 -335
rect 21920 -415 21950 -385
rect 22005 -365 22035 -335
rect 22090 -415 22120 -385
rect 22175 -365 22205 -335
rect 22260 -415 22290 -385
rect 22345 -365 22375 -335
rect 22430 -415 22460 -385
rect 22515 -365 22545 -335
rect 22600 -415 22630 -385
rect 22685 -365 22715 -335
rect 22770 -415 22800 -385
rect 22855 -365 22885 -335
rect 22940 -415 22970 -385
rect 23025 -365 23055 -335
rect 23110 -415 23140 -385
rect 23195 -365 23225 -335
rect 23280 -415 23310 -385
rect 23365 -365 23395 -335
rect 23450 -415 23480 -385
rect 23535 -365 23565 -335
rect 23620 -415 23650 -385
rect 23705 -365 23735 -335
rect 23790 -415 23820 -385
rect 23875 -365 23905 -335
rect 23960 -415 23990 -385
rect 24045 -365 24075 -335
rect 24130 -415 24160 -385
rect 24215 -365 24245 -335
rect 24300 -415 24330 -385
rect 24385 -365 24415 -335
rect 24470 -415 24500 -385
rect 24555 -365 24585 -335
rect 24640 -415 24670 -385
rect 24725 -365 24755 -335
rect 24810 -415 24840 -385
rect 24895 -365 24925 -335
rect 24980 -415 25010 -385
rect 25065 -365 25095 -335
rect 25150 -415 25180 -385
rect 25235 -365 25265 -335
rect 25320 -415 25350 -385
rect 25405 -365 25435 -335
rect 25490 -415 25520 -385
rect 25575 -365 25605 -335
rect 25660 -415 25690 -385
rect 25745 -365 25775 -335
rect 25830 -415 25860 -385
rect 25915 -365 25945 -335
rect 26000 -415 26030 -385
rect 26085 -365 26115 -335
rect 26170 -415 26200 -385
rect 26255 -365 26285 -335
rect 26340 -415 26370 -385
rect 26425 -365 26455 -335
rect 26510 -415 26540 -385
rect 26595 -365 26625 -335
rect 26680 -415 26710 -385
rect 26765 -365 26795 -335
rect 26850 -415 26880 -385
rect 26935 -365 26965 -335
rect 27020 -415 27050 -385
rect 27105 -365 27135 -335
rect 27190 -415 27220 -385
rect 27275 -365 27305 -335
rect 27360 -415 27390 -385
rect 27445 -365 27475 -335
rect 27530 -415 27560 -385
rect 27615 -365 27645 -335
rect 27700 -415 27730 -385
rect 27785 -365 27815 -335
rect 27870 -415 27900 -385
rect 27955 -365 27985 -335
rect 28040 -415 28070 -385
rect 28125 -365 28155 -335
rect 28210 -415 28240 -385
rect 28295 -365 28325 -335
rect 28380 -415 28410 -385
rect 28465 -365 28495 -335
rect 28550 -415 28580 -385
rect 28635 -365 28665 -335
rect 28720 -415 28750 -385
rect 28805 -365 28835 -335
rect 28890 -415 28920 -385
rect 28975 -365 29005 -335
rect 29060 -415 29090 -385
rect 29145 -365 29175 -335
rect 29230 -415 29260 -385
rect 29315 -365 29345 -335
rect 29400 -415 29430 -385
rect 29485 -365 29515 -335
rect 29570 -415 29600 -385
rect 29655 -365 29685 -335
rect 29740 -415 29770 -385
rect 29825 -365 29855 -335
rect 29910 -415 29940 -385
rect 29995 -365 30025 -335
rect 30080 -415 30110 -385
rect 30165 -365 30195 -335
rect 30250 -415 30280 -385
rect 30335 -365 30365 -335
rect 30420 -415 30450 -385
rect 30505 -365 30535 -335
rect 30590 -415 30620 -385
rect 30675 -365 30705 -335
rect 30760 -415 30790 -385
rect 30845 -365 30875 -335
rect 30930 -415 30960 -385
rect 31015 -365 31045 -335
rect 31100 -415 31130 -385
rect 31185 -365 31215 -335
rect 31270 -415 31300 -385
rect 31355 -365 31385 -335
rect 31440 -415 31470 -385
rect 31525 -365 31555 -335
rect 31610 -415 31640 -385
rect 31695 -365 31725 -335
rect 31780 -415 31810 -385
rect 31865 -365 31895 -335
rect 31950 -415 31980 -385
rect 32035 -365 32065 -335
rect 32120 -415 32150 -385
rect 32205 -365 32235 -335
rect 32290 -415 32320 -385
rect 32375 -365 32405 -335
rect 32460 -415 32490 -385
rect 32545 -365 32575 -335
rect 32630 -415 32660 -385
rect 32715 -365 32745 -335
rect 32800 -415 32830 -385
rect 32885 -365 32915 -335
rect 32970 -415 33000 -385
rect 33055 -365 33085 -335
rect 33140 -415 33170 -385
rect 33225 -365 33255 -335
rect 33310 -415 33340 -385
rect 33395 -365 33425 -335
rect 33480 -415 33510 -385
rect 33565 -365 33595 -335
rect 33650 -415 33680 -385
rect 33735 -365 33765 -335
rect 33820 -415 33850 -385
rect 33905 -365 33935 -335
rect 33990 -415 34020 -385
rect 34075 -365 34105 -335
rect 34160 -415 34190 -385
rect 34245 -365 34275 -335
rect 34330 -415 34360 -385
rect 34415 -365 34445 -335
rect 34500 -415 34530 -385
rect 34585 -365 34615 -335
rect 34670 -415 34700 -385
rect 34755 -365 34785 -335
rect 34840 -415 34870 -385
rect 34925 -365 34955 -335
rect 35010 -415 35040 -385
rect 35095 -365 35125 -335
rect 35180 -415 35210 -385
rect 35265 -365 35295 -335
rect 35350 -415 35380 -385
rect 35435 -365 35465 -335
rect 35520 -415 35550 -385
rect 35605 -365 35635 -335
rect 35690 -415 35720 -385
rect 35775 -365 35805 -335
rect 35860 -415 35890 -385
rect 35945 -365 35975 -335
rect 36030 -415 36060 -385
rect 36115 -365 36145 -335
rect 36200 -415 36230 -385
rect 36285 -365 36315 -335
rect 36370 -415 36400 -385
rect 36455 -365 36485 -335
rect 36540 -415 36570 -385
rect 36625 -365 36655 -335
rect 36710 -415 36740 -385
rect 36795 -365 36825 -335
rect 36880 -415 36910 -385
rect 36965 -365 36995 -335
rect 37050 -415 37080 -385
rect 37135 -365 37165 -335
rect 37220 -415 37250 -385
rect 37305 -365 37335 -335
rect 37390 -415 37420 -385
rect 37475 -365 37505 -335
rect 37560 -415 37590 -385
rect 37645 -365 37675 -335
rect 37730 -415 37760 -385
rect 37815 -365 37845 -335
rect 37900 -415 37930 -385
rect 37985 -365 38015 -335
rect 38070 -415 38100 -385
rect 38155 -365 38185 -335
rect 38240 -415 38270 -385
rect 38325 -365 38355 -335
rect 38410 -415 38440 -385
rect 38495 -365 38525 -335
rect 38580 -415 38610 -385
rect 38665 -365 38695 -335
rect 38750 -415 38780 -385
rect 38835 -365 38865 -335
rect 38920 -415 38950 -385
rect 39005 -365 39035 -335
rect 39090 -415 39120 -385
rect 39175 -365 39205 -335
rect 39260 -415 39290 -385
rect 39345 -365 39375 -335
rect 39430 -415 39460 -385
rect 39515 -365 39545 -335
rect 39600 -415 39630 -385
rect 39685 -365 39715 -335
rect 39770 -415 39800 -385
rect 39855 -365 39885 -335
rect 39940 -415 39970 -385
rect 40025 -365 40055 -335
rect 40110 -415 40140 -385
rect 40195 -365 40225 -335
rect 40280 -415 40310 -385
rect 40365 -365 40395 -335
rect 40450 -415 40480 -385
rect 40535 -365 40565 -335
rect 40620 -415 40650 -385
rect 40705 -365 40735 -335
rect 40790 -415 40820 -385
rect 40875 -365 40905 -335
rect 40960 -415 40990 -385
rect 41045 -365 41075 -335
rect 41130 -415 41160 -385
rect 41215 -365 41245 -335
rect 41300 -415 41330 -385
rect 41385 -365 41415 -335
rect 41470 -415 41500 -385
rect 41555 -365 41585 -335
rect 41640 -415 41670 -385
rect 41725 -365 41755 -335
rect 41810 -415 41840 -385
rect 41895 -365 41925 -335
rect 41980 -415 42010 -385
rect 42065 -365 42095 -335
rect 42150 -415 42180 -385
rect 42235 -365 42265 -335
rect 42320 -415 42350 -385
rect 42405 -365 42435 -335
rect 42490 -415 42520 -385
rect 42575 -365 42605 -335
rect 42660 -415 42690 -385
rect 42745 -365 42775 -335
rect 42830 -415 42860 -385
rect 42915 -365 42945 -335
rect 43000 -415 43030 -385
rect 43085 -365 43115 -335
rect 43170 -415 43200 -385
rect 43255 -365 43285 -335
rect 43340 -415 43370 -385
rect 43425 -365 43455 -335
rect 43510 -415 43540 -385
rect 43595 -365 43625 -335
rect 75 -580 105 -550
rect 75 -680 105 -650
rect 160 -530 190 -500
rect 160 -630 190 -600
rect 245 -580 275 -550
rect 245 -680 275 -650
rect 330 -530 360 -500
rect 330 -630 360 -600
rect 415 -580 445 -550
rect 415 -680 445 -650
rect 500 -530 530 -500
rect 500 -630 530 -600
rect 585 -580 615 -550
rect 585 -680 615 -650
rect 670 -530 700 -500
rect 670 -630 700 -600
rect 755 -580 785 -550
rect 755 -680 785 -650
rect 840 -530 870 -500
rect 840 -630 870 -600
rect 925 -580 955 -550
rect 925 -680 955 -650
rect 1010 -530 1040 -500
rect 1010 -630 1040 -600
rect 1095 -580 1125 -550
rect 1095 -680 1125 -650
rect 1180 -530 1210 -500
rect 1180 -630 1210 -600
rect 1265 -580 1295 -550
rect 1265 -680 1295 -650
rect 1350 -530 1380 -500
rect 1350 -630 1380 -600
rect 1435 -580 1465 -550
rect 1435 -680 1465 -650
rect 1520 -530 1550 -500
rect 1520 -630 1550 -600
rect 1605 -580 1635 -550
rect 1605 -680 1635 -650
rect 1690 -530 1720 -500
rect 1690 -630 1720 -600
rect 1775 -580 1805 -550
rect 1775 -680 1805 -650
rect 1860 -530 1890 -500
rect 1860 -630 1890 -600
rect 1945 -580 1975 -550
rect 1945 -680 1975 -650
rect 2030 -530 2060 -500
rect 2030 -630 2060 -600
rect 2115 -580 2145 -550
rect 2115 -680 2145 -650
rect 2200 -530 2230 -500
rect 2200 -630 2230 -600
rect 2285 -580 2315 -550
rect 2285 -680 2315 -650
rect 2370 -530 2400 -500
rect 2370 -630 2400 -600
rect 2455 -580 2485 -550
rect 2455 -680 2485 -650
rect 2540 -530 2570 -500
rect 2540 -630 2570 -600
rect 2625 -580 2655 -550
rect 2625 -680 2655 -650
rect 2710 -530 2740 -500
rect 2710 -630 2740 -600
rect 2795 -580 2825 -550
rect 2795 -680 2825 -650
rect 2880 -530 2910 -500
rect 2880 -630 2910 -600
rect 2965 -580 2995 -550
rect 2965 -680 2995 -650
rect 3050 -530 3080 -500
rect 3050 -630 3080 -600
rect 3135 -580 3165 -550
rect 3135 -680 3165 -650
rect 3220 -530 3250 -500
rect 3220 -630 3250 -600
rect 3305 -580 3335 -550
rect 3305 -680 3335 -650
rect 3390 -530 3420 -500
rect 3390 -630 3420 -600
rect 3475 -580 3505 -550
rect 3475 -680 3505 -650
rect 3560 -530 3590 -500
rect 3560 -630 3590 -600
rect 3645 -580 3675 -550
rect 3645 -680 3675 -650
rect 3730 -530 3760 -500
rect 3730 -630 3760 -600
rect 3815 -580 3845 -550
rect 3815 -680 3845 -650
rect 3900 -530 3930 -500
rect 3900 -630 3930 -600
rect 3985 -580 4015 -550
rect 3985 -680 4015 -650
rect 4070 -530 4100 -500
rect 4070 -630 4100 -600
rect 4155 -580 4185 -550
rect 4155 -680 4185 -650
rect 4240 -530 4270 -500
rect 4240 -630 4270 -600
rect 4325 -580 4355 -550
rect 4325 -680 4355 -650
rect 4410 -530 4440 -500
rect 4410 -630 4440 -600
rect 4495 -580 4525 -550
rect 4495 -680 4525 -650
rect 4580 -530 4610 -500
rect 4580 -630 4610 -600
rect 4665 -580 4695 -550
rect 4665 -680 4695 -650
rect 4750 -530 4780 -500
rect 4750 -630 4780 -600
rect 4835 -580 4865 -550
rect 4835 -680 4865 -650
rect 4920 -530 4950 -500
rect 4920 -630 4950 -600
rect 5005 -580 5035 -550
rect 5005 -680 5035 -650
rect 5090 -530 5120 -500
rect 5090 -630 5120 -600
rect 5175 -580 5205 -550
rect 5175 -680 5205 -650
rect 5260 -530 5290 -500
rect 5260 -630 5290 -600
rect 5345 -580 5375 -550
rect 5345 -680 5375 -650
rect 5430 -530 5460 -500
rect 5430 -630 5460 -600
rect 5515 -580 5545 -550
rect 5515 -680 5545 -650
rect 5600 -530 5630 -500
rect 5600 -630 5630 -600
rect 5685 -580 5715 -550
rect 5685 -680 5715 -650
rect 5770 -530 5800 -500
rect 5770 -630 5800 -600
rect 5855 -580 5885 -550
rect 5855 -680 5885 -650
rect 5940 -530 5970 -500
rect 5940 -630 5970 -600
rect 6025 -580 6055 -550
rect 6025 -680 6055 -650
rect 6110 -530 6140 -500
rect 6110 -630 6140 -600
rect 6195 -580 6225 -550
rect 6195 -680 6225 -650
rect 6280 -530 6310 -500
rect 6280 -630 6310 -600
rect 6365 -580 6395 -550
rect 6365 -680 6395 -650
rect 6450 -530 6480 -500
rect 6450 -630 6480 -600
rect 6535 -580 6565 -550
rect 6535 -680 6565 -650
rect 6620 -530 6650 -500
rect 6620 -630 6650 -600
rect 6705 -580 6735 -550
rect 6705 -680 6735 -650
rect 6790 -530 6820 -500
rect 6790 -630 6820 -600
rect 6875 -580 6905 -550
rect 6875 -680 6905 -650
rect 6960 -530 6990 -500
rect 6960 -630 6990 -600
rect 7045 -580 7075 -550
rect 7045 -680 7075 -650
rect 7130 -530 7160 -500
rect 7130 -630 7160 -600
rect 7215 -580 7245 -550
rect 7215 -680 7245 -650
rect 7300 -530 7330 -500
rect 7300 -630 7330 -600
rect 7385 -580 7415 -550
rect 7385 -680 7415 -650
rect 7470 -530 7500 -500
rect 7470 -630 7500 -600
rect 7555 -580 7585 -550
rect 7555 -680 7585 -650
rect 7640 -530 7670 -500
rect 7640 -630 7670 -600
rect 7725 -580 7755 -550
rect 7725 -680 7755 -650
rect 7810 -530 7840 -500
rect 7810 -630 7840 -600
rect 7895 -580 7925 -550
rect 7895 -680 7925 -650
rect 7980 -530 8010 -500
rect 7980 -630 8010 -600
rect 8065 -580 8095 -550
rect 8065 -680 8095 -650
rect 8150 -530 8180 -500
rect 8150 -630 8180 -600
rect 8235 -580 8265 -550
rect 8235 -680 8265 -650
rect 8320 -530 8350 -500
rect 8320 -630 8350 -600
rect 8405 -580 8435 -550
rect 8405 -680 8435 -650
rect 8490 -530 8520 -500
rect 8490 -630 8520 -600
rect 8575 -580 8605 -550
rect 8575 -680 8605 -650
rect 8660 -530 8690 -500
rect 8660 -630 8690 -600
rect 8745 -580 8775 -550
rect 8745 -680 8775 -650
rect 8830 -530 8860 -500
rect 8830 -630 8860 -600
rect 8915 -580 8945 -550
rect 8915 -680 8945 -650
rect 9000 -530 9030 -500
rect 9000 -630 9030 -600
rect 9085 -580 9115 -550
rect 9085 -680 9115 -650
rect 9170 -530 9200 -500
rect 9170 -630 9200 -600
rect 9255 -580 9285 -550
rect 9255 -680 9285 -650
rect 9340 -530 9370 -500
rect 9340 -630 9370 -600
rect 9425 -580 9455 -550
rect 9425 -680 9455 -650
rect 9510 -530 9540 -500
rect 9510 -630 9540 -600
rect 9595 -580 9625 -550
rect 9595 -680 9625 -650
rect 9680 -530 9710 -500
rect 9680 -630 9710 -600
rect 9765 -580 9795 -550
rect 9765 -680 9795 -650
rect 9850 -530 9880 -500
rect 9850 -630 9880 -600
rect 9935 -580 9965 -550
rect 9935 -680 9965 -650
rect 10020 -530 10050 -500
rect 10020 -630 10050 -600
rect 10105 -580 10135 -550
rect 10105 -680 10135 -650
rect 10190 -530 10220 -500
rect 10190 -630 10220 -600
rect 10275 -580 10305 -550
rect 10275 -680 10305 -650
rect 10360 -530 10390 -500
rect 10360 -630 10390 -600
rect 10445 -580 10475 -550
rect 10445 -680 10475 -650
rect 10530 -530 10560 -500
rect 10530 -630 10560 -600
rect 10615 -580 10645 -550
rect 10615 -680 10645 -650
rect 10700 -530 10730 -500
rect 10700 -630 10730 -600
rect 10785 -580 10815 -550
rect 10785 -680 10815 -650
rect 10870 -530 10900 -500
rect 10870 -630 10900 -600
rect 10955 -580 10985 -550
rect 10955 -680 10985 -650
rect 11040 -530 11070 -500
rect 11040 -630 11070 -600
rect 11125 -580 11155 -550
rect 11125 -680 11155 -650
rect 11210 -530 11240 -500
rect 11210 -630 11240 -600
rect 11295 -580 11325 -550
rect 11295 -680 11325 -650
rect 11380 -530 11410 -500
rect 11380 -630 11410 -600
rect 11465 -580 11495 -550
rect 11465 -680 11495 -650
rect 11550 -530 11580 -500
rect 11550 -630 11580 -600
rect 11635 -580 11665 -550
rect 11635 -680 11665 -650
rect 11720 -530 11750 -500
rect 11720 -630 11750 -600
rect 11805 -580 11835 -550
rect 11805 -680 11835 -650
rect 11890 -530 11920 -500
rect 11890 -630 11920 -600
rect 11975 -580 12005 -550
rect 11975 -680 12005 -650
rect 12060 -530 12090 -500
rect 12060 -630 12090 -600
rect 12145 -580 12175 -550
rect 12145 -680 12175 -650
rect 12230 -530 12260 -500
rect 12230 -630 12260 -600
rect 12315 -580 12345 -550
rect 12315 -680 12345 -650
rect 12400 -530 12430 -500
rect 12400 -630 12430 -600
rect 12485 -580 12515 -550
rect 12485 -680 12515 -650
rect 12570 -530 12600 -500
rect 12570 -630 12600 -600
rect 12655 -580 12685 -550
rect 12655 -680 12685 -650
rect 12740 -530 12770 -500
rect 12740 -630 12770 -600
rect 12825 -580 12855 -550
rect 12825 -680 12855 -650
rect 12910 -530 12940 -500
rect 12910 -630 12940 -600
rect 12995 -580 13025 -550
rect 12995 -680 13025 -650
rect 13080 -530 13110 -500
rect 13080 -630 13110 -600
rect 13165 -580 13195 -550
rect 13165 -680 13195 -650
rect 13250 -530 13280 -500
rect 13250 -630 13280 -600
rect 13335 -580 13365 -550
rect 13335 -680 13365 -650
rect 13420 -530 13450 -500
rect 13420 -630 13450 -600
rect 13505 -580 13535 -550
rect 13505 -680 13535 -650
rect 13590 -530 13620 -500
rect 13590 -630 13620 -600
rect 13675 -580 13705 -550
rect 13675 -680 13705 -650
rect 13760 -530 13790 -500
rect 13760 -630 13790 -600
rect 13845 -580 13875 -550
rect 13845 -680 13875 -650
rect 13930 -530 13960 -500
rect 13930 -630 13960 -600
rect 14015 -580 14045 -550
rect 14015 -680 14045 -650
rect 14100 -530 14130 -500
rect 14100 -630 14130 -600
rect 14185 -580 14215 -550
rect 14185 -680 14215 -650
rect 14270 -530 14300 -500
rect 14270 -630 14300 -600
rect 14355 -580 14385 -550
rect 14355 -680 14385 -650
rect 14440 -530 14470 -500
rect 14440 -630 14470 -600
rect 14525 -580 14555 -550
rect 14525 -680 14555 -650
rect 14610 -530 14640 -500
rect 14610 -630 14640 -600
rect 14695 -580 14725 -550
rect 14695 -680 14725 -650
rect 14780 -530 14810 -500
rect 14780 -630 14810 -600
rect 14865 -580 14895 -550
rect 14865 -680 14895 -650
rect 14950 -530 14980 -500
rect 14950 -630 14980 -600
rect 15035 -580 15065 -550
rect 15035 -680 15065 -650
rect 15120 -530 15150 -500
rect 15120 -630 15150 -600
rect 15205 -580 15235 -550
rect 15205 -680 15235 -650
rect 15290 -530 15320 -500
rect 15290 -630 15320 -600
rect 15375 -580 15405 -550
rect 15375 -680 15405 -650
rect 15460 -530 15490 -500
rect 15460 -630 15490 -600
rect 15545 -580 15575 -550
rect 15545 -680 15575 -650
rect 15630 -530 15660 -500
rect 15630 -630 15660 -600
rect 15715 -580 15745 -550
rect 15715 -680 15745 -650
rect 15800 -530 15830 -500
rect 15800 -630 15830 -600
rect 15885 -580 15915 -550
rect 15885 -680 15915 -650
rect 15970 -530 16000 -500
rect 15970 -630 16000 -600
rect 16055 -580 16085 -550
rect 16055 -680 16085 -650
rect 16140 -530 16170 -500
rect 16140 -630 16170 -600
rect 16225 -580 16255 -550
rect 16225 -680 16255 -650
rect 16310 -530 16340 -500
rect 16310 -630 16340 -600
rect 16395 -580 16425 -550
rect 16395 -680 16425 -650
rect 16480 -530 16510 -500
rect 16480 -630 16510 -600
rect 16565 -580 16595 -550
rect 16565 -680 16595 -650
rect 16650 -530 16680 -500
rect 16650 -630 16680 -600
rect 16735 -580 16765 -550
rect 16735 -680 16765 -650
rect 16820 -530 16850 -500
rect 16820 -630 16850 -600
rect 16905 -580 16935 -550
rect 16905 -680 16935 -650
rect 16990 -530 17020 -500
rect 16990 -630 17020 -600
rect 17075 -580 17105 -550
rect 17075 -680 17105 -650
rect 17160 -530 17190 -500
rect 17160 -630 17190 -600
rect 17245 -580 17275 -550
rect 17245 -680 17275 -650
rect 17330 -530 17360 -500
rect 17330 -630 17360 -600
rect 17415 -580 17445 -550
rect 17415 -680 17445 -650
rect 17500 -530 17530 -500
rect 17500 -630 17530 -600
rect 17585 -580 17615 -550
rect 17585 -680 17615 -650
rect 17670 -530 17700 -500
rect 17670 -630 17700 -600
rect 17755 -580 17785 -550
rect 17755 -680 17785 -650
rect 17840 -530 17870 -500
rect 17840 -630 17870 -600
rect 17925 -580 17955 -550
rect 17925 -680 17955 -650
rect 18010 -530 18040 -500
rect 18010 -630 18040 -600
rect 18095 -580 18125 -550
rect 18095 -680 18125 -650
rect 18180 -530 18210 -500
rect 18180 -630 18210 -600
rect 18265 -580 18295 -550
rect 18265 -680 18295 -650
rect 18350 -530 18380 -500
rect 18350 -630 18380 -600
rect 18435 -580 18465 -550
rect 18435 -680 18465 -650
rect 18520 -530 18550 -500
rect 18520 -630 18550 -600
rect 18605 -580 18635 -550
rect 18605 -680 18635 -650
rect 18690 -530 18720 -500
rect 18690 -630 18720 -600
rect 18775 -580 18805 -550
rect 18775 -680 18805 -650
rect 18860 -530 18890 -500
rect 18860 -630 18890 -600
rect 18945 -580 18975 -550
rect 18945 -680 18975 -650
rect 19030 -530 19060 -500
rect 19030 -630 19060 -600
rect 19115 -580 19145 -550
rect 19115 -680 19145 -650
rect 19200 -530 19230 -500
rect 19200 -630 19230 -600
rect 19285 -580 19315 -550
rect 19285 -680 19315 -650
rect 19370 -530 19400 -500
rect 19370 -630 19400 -600
rect 19455 -580 19485 -550
rect 19455 -680 19485 -650
rect 19540 -530 19570 -500
rect 19540 -630 19570 -600
rect 19625 -580 19655 -550
rect 19625 -680 19655 -650
rect 19710 -530 19740 -500
rect 19710 -630 19740 -600
rect 19795 -580 19825 -550
rect 19795 -680 19825 -650
rect 19880 -530 19910 -500
rect 19880 -630 19910 -600
rect 19965 -580 19995 -550
rect 19965 -680 19995 -650
rect 20050 -530 20080 -500
rect 20050 -630 20080 -600
rect 20135 -580 20165 -550
rect 20135 -680 20165 -650
rect 20220 -530 20250 -500
rect 20220 -630 20250 -600
rect 20305 -580 20335 -550
rect 20305 -680 20335 -650
rect 20390 -530 20420 -500
rect 20390 -630 20420 -600
rect 20475 -580 20505 -550
rect 20475 -680 20505 -650
rect 20560 -530 20590 -500
rect 20560 -630 20590 -600
rect 20645 -580 20675 -550
rect 20645 -680 20675 -650
rect 20730 -530 20760 -500
rect 20730 -630 20760 -600
rect 20815 -580 20845 -550
rect 20815 -680 20845 -650
rect 20900 -530 20930 -500
rect 20900 -630 20930 -600
rect 20985 -580 21015 -550
rect 20985 -680 21015 -650
rect 21070 -530 21100 -500
rect 21070 -630 21100 -600
rect 21155 -580 21185 -550
rect 21155 -680 21185 -650
rect 21240 -530 21270 -500
rect 21240 -630 21270 -600
rect 21325 -580 21355 -550
rect 21325 -680 21355 -650
rect 21410 -530 21440 -500
rect 21410 -630 21440 -600
rect 21495 -580 21525 -550
rect 21495 -680 21525 -650
rect 21580 -530 21610 -500
rect 21580 -630 21610 -600
rect 21665 -580 21695 -550
rect 21665 -680 21695 -650
rect 21750 -530 21780 -500
rect 21750 -630 21780 -600
rect 21835 -580 21865 -550
rect 21835 -680 21865 -650
rect 21920 -530 21950 -500
rect 21920 -630 21950 -600
rect 22005 -580 22035 -550
rect 22005 -680 22035 -650
rect 22090 -530 22120 -500
rect 22090 -630 22120 -600
rect 22175 -580 22205 -550
rect 22175 -680 22205 -650
rect 22260 -530 22290 -500
rect 22260 -630 22290 -600
rect 22345 -580 22375 -550
rect 22345 -680 22375 -650
rect 22430 -530 22460 -500
rect 22430 -630 22460 -600
rect 22515 -580 22545 -550
rect 22515 -680 22545 -650
rect 22600 -530 22630 -500
rect 22600 -630 22630 -600
rect 22685 -580 22715 -550
rect 22685 -680 22715 -650
rect 22770 -530 22800 -500
rect 22770 -630 22800 -600
rect 22855 -580 22885 -550
rect 22855 -680 22885 -650
rect 22940 -530 22970 -500
rect 22940 -630 22970 -600
rect 23025 -580 23055 -550
rect 23025 -680 23055 -650
rect 23110 -530 23140 -500
rect 23110 -630 23140 -600
rect 23195 -580 23225 -550
rect 23195 -680 23225 -650
rect 23280 -530 23310 -500
rect 23280 -630 23310 -600
rect 23365 -580 23395 -550
rect 23365 -680 23395 -650
rect 23450 -530 23480 -500
rect 23450 -630 23480 -600
rect 23535 -580 23565 -550
rect 23535 -680 23565 -650
rect 23620 -530 23650 -500
rect 23620 -630 23650 -600
rect 23705 -580 23735 -550
rect 23705 -680 23735 -650
rect 23790 -530 23820 -500
rect 23790 -630 23820 -600
rect 23875 -580 23905 -550
rect 23875 -680 23905 -650
rect 23960 -530 23990 -500
rect 23960 -630 23990 -600
rect 24045 -580 24075 -550
rect 24045 -680 24075 -650
rect 24130 -530 24160 -500
rect 24130 -630 24160 -600
rect 24215 -580 24245 -550
rect 24215 -680 24245 -650
rect 24300 -530 24330 -500
rect 24300 -630 24330 -600
rect 24385 -580 24415 -550
rect 24385 -680 24415 -650
rect 24470 -530 24500 -500
rect 24470 -630 24500 -600
rect 24555 -580 24585 -550
rect 24555 -680 24585 -650
rect 24640 -530 24670 -500
rect 24640 -630 24670 -600
rect 24725 -580 24755 -550
rect 24725 -680 24755 -650
rect 24810 -530 24840 -500
rect 24810 -630 24840 -600
rect 24895 -580 24925 -550
rect 24895 -680 24925 -650
rect 24980 -530 25010 -500
rect 24980 -630 25010 -600
rect 25065 -580 25095 -550
rect 25065 -680 25095 -650
rect 25150 -530 25180 -500
rect 25150 -630 25180 -600
rect 25235 -580 25265 -550
rect 25235 -680 25265 -650
rect 25320 -530 25350 -500
rect 25320 -630 25350 -600
rect 25405 -580 25435 -550
rect 25405 -680 25435 -650
rect 25490 -530 25520 -500
rect 25490 -630 25520 -600
rect 25575 -580 25605 -550
rect 25575 -680 25605 -650
rect 25660 -530 25690 -500
rect 25660 -630 25690 -600
rect 25745 -580 25775 -550
rect 25745 -680 25775 -650
rect 25830 -530 25860 -500
rect 25830 -630 25860 -600
rect 25915 -580 25945 -550
rect 25915 -680 25945 -650
rect 26000 -530 26030 -500
rect 26000 -630 26030 -600
rect 26085 -580 26115 -550
rect 26085 -680 26115 -650
rect 26170 -530 26200 -500
rect 26170 -630 26200 -600
rect 26255 -580 26285 -550
rect 26255 -680 26285 -650
rect 26340 -530 26370 -500
rect 26340 -630 26370 -600
rect 26425 -580 26455 -550
rect 26425 -680 26455 -650
rect 26510 -530 26540 -500
rect 26510 -630 26540 -600
rect 26595 -580 26625 -550
rect 26595 -680 26625 -650
rect 26680 -530 26710 -500
rect 26680 -630 26710 -600
rect 26765 -580 26795 -550
rect 26765 -680 26795 -650
rect 26850 -530 26880 -500
rect 26850 -630 26880 -600
rect 26935 -580 26965 -550
rect 26935 -680 26965 -650
rect 27020 -530 27050 -500
rect 27020 -630 27050 -600
rect 27105 -580 27135 -550
rect 27105 -680 27135 -650
rect 27190 -530 27220 -500
rect 27190 -630 27220 -600
rect 27275 -580 27305 -550
rect 27275 -680 27305 -650
rect 27360 -530 27390 -500
rect 27360 -630 27390 -600
rect 27445 -580 27475 -550
rect 27445 -680 27475 -650
rect 27530 -530 27560 -500
rect 27530 -630 27560 -600
rect 27615 -580 27645 -550
rect 27615 -680 27645 -650
rect 27700 -530 27730 -500
rect 27700 -630 27730 -600
rect 27785 -580 27815 -550
rect 27785 -680 27815 -650
rect 27870 -530 27900 -500
rect 27870 -630 27900 -600
rect 27955 -580 27985 -550
rect 27955 -680 27985 -650
rect 28040 -530 28070 -500
rect 28040 -630 28070 -600
rect 28125 -580 28155 -550
rect 28125 -680 28155 -650
rect 28210 -530 28240 -500
rect 28210 -630 28240 -600
rect 28295 -580 28325 -550
rect 28295 -680 28325 -650
rect 28380 -530 28410 -500
rect 28380 -630 28410 -600
rect 28465 -580 28495 -550
rect 28465 -680 28495 -650
rect 28550 -530 28580 -500
rect 28550 -630 28580 -600
rect 28635 -580 28665 -550
rect 28635 -680 28665 -650
rect 28720 -530 28750 -500
rect 28720 -630 28750 -600
rect 28805 -580 28835 -550
rect 28805 -680 28835 -650
rect 28890 -530 28920 -500
rect 28890 -630 28920 -600
rect 28975 -580 29005 -550
rect 28975 -680 29005 -650
rect 29060 -530 29090 -500
rect 29060 -630 29090 -600
rect 29145 -580 29175 -550
rect 29145 -680 29175 -650
rect 29230 -530 29260 -500
rect 29230 -630 29260 -600
rect 29315 -580 29345 -550
rect 29315 -680 29345 -650
rect 29400 -530 29430 -500
rect 29400 -630 29430 -600
rect 29485 -580 29515 -550
rect 29485 -680 29515 -650
rect 29570 -530 29600 -500
rect 29570 -630 29600 -600
rect 29655 -580 29685 -550
rect 29655 -680 29685 -650
rect 29740 -530 29770 -500
rect 29740 -630 29770 -600
rect 29825 -580 29855 -550
rect 29825 -680 29855 -650
rect 29910 -530 29940 -500
rect 29910 -630 29940 -600
rect 29995 -580 30025 -550
rect 29995 -680 30025 -650
rect 30080 -530 30110 -500
rect 30080 -630 30110 -600
rect 30165 -580 30195 -550
rect 30165 -680 30195 -650
rect 30250 -530 30280 -500
rect 30250 -630 30280 -600
rect 30335 -580 30365 -550
rect 30335 -680 30365 -650
rect 30420 -530 30450 -500
rect 30420 -630 30450 -600
rect 30505 -580 30535 -550
rect 30505 -680 30535 -650
rect 30590 -530 30620 -500
rect 30590 -630 30620 -600
rect 30675 -580 30705 -550
rect 30675 -680 30705 -650
rect 30760 -530 30790 -500
rect 30760 -630 30790 -600
rect 30845 -580 30875 -550
rect 30845 -680 30875 -650
rect 30930 -530 30960 -500
rect 30930 -630 30960 -600
rect 31015 -580 31045 -550
rect 31015 -680 31045 -650
rect 31100 -530 31130 -500
rect 31100 -630 31130 -600
rect 31185 -580 31215 -550
rect 31185 -680 31215 -650
rect 31270 -530 31300 -500
rect 31270 -630 31300 -600
rect 31355 -580 31385 -550
rect 31355 -680 31385 -650
rect 31440 -530 31470 -500
rect 31440 -630 31470 -600
rect 31525 -580 31555 -550
rect 31525 -680 31555 -650
rect 31610 -530 31640 -500
rect 31610 -630 31640 -600
rect 31695 -580 31725 -550
rect 31695 -680 31725 -650
rect 31780 -530 31810 -500
rect 31780 -630 31810 -600
rect 31865 -580 31895 -550
rect 31865 -680 31895 -650
rect 31950 -530 31980 -500
rect 31950 -630 31980 -600
rect 32035 -580 32065 -550
rect 32035 -680 32065 -650
rect 32120 -530 32150 -500
rect 32120 -630 32150 -600
rect 32205 -580 32235 -550
rect 32205 -680 32235 -650
rect 32290 -530 32320 -500
rect 32290 -630 32320 -600
rect 32375 -580 32405 -550
rect 32375 -680 32405 -650
rect 32460 -530 32490 -500
rect 32460 -630 32490 -600
rect 32545 -580 32575 -550
rect 32545 -680 32575 -650
rect 32630 -530 32660 -500
rect 32630 -630 32660 -600
rect 32715 -580 32745 -550
rect 32715 -680 32745 -650
rect 32800 -530 32830 -500
rect 32800 -630 32830 -600
rect 32885 -580 32915 -550
rect 32885 -680 32915 -650
rect 32970 -530 33000 -500
rect 32970 -630 33000 -600
rect 33055 -580 33085 -550
rect 33055 -680 33085 -650
rect 33140 -530 33170 -500
rect 33140 -630 33170 -600
rect 33225 -580 33255 -550
rect 33225 -680 33255 -650
rect 33310 -530 33340 -500
rect 33310 -630 33340 -600
rect 33395 -580 33425 -550
rect 33395 -680 33425 -650
rect 33480 -530 33510 -500
rect 33480 -630 33510 -600
rect 33565 -580 33595 -550
rect 33565 -680 33595 -650
rect 33650 -530 33680 -500
rect 33650 -630 33680 -600
rect 33735 -580 33765 -550
rect 33735 -680 33765 -650
rect 33820 -530 33850 -500
rect 33820 -630 33850 -600
rect 33905 -580 33935 -550
rect 33905 -680 33935 -650
rect 33990 -530 34020 -500
rect 33990 -630 34020 -600
rect 34075 -580 34105 -550
rect 34075 -680 34105 -650
rect 34160 -530 34190 -500
rect 34160 -630 34190 -600
rect 34245 -580 34275 -550
rect 34245 -680 34275 -650
rect 34330 -530 34360 -500
rect 34330 -630 34360 -600
rect 34415 -580 34445 -550
rect 34415 -680 34445 -650
rect 34500 -530 34530 -500
rect 34500 -630 34530 -600
rect 34585 -580 34615 -550
rect 34585 -680 34615 -650
rect 34670 -530 34700 -500
rect 34670 -630 34700 -600
rect 34755 -580 34785 -550
rect 34755 -680 34785 -650
rect 34840 -530 34870 -500
rect 34840 -630 34870 -600
rect 34925 -580 34955 -550
rect 34925 -680 34955 -650
rect 35010 -530 35040 -500
rect 35010 -630 35040 -600
rect 35095 -580 35125 -550
rect 35095 -680 35125 -650
rect 35180 -530 35210 -500
rect 35180 -630 35210 -600
rect 35265 -580 35295 -550
rect 35265 -680 35295 -650
rect 35350 -530 35380 -500
rect 35350 -630 35380 -600
rect 35435 -580 35465 -550
rect 35435 -680 35465 -650
rect 35520 -530 35550 -500
rect 35520 -630 35550 -600
rect 35605 -580 35635 -550
rect 35605 -680 35635 -650
rect 35690 -530 35720 -500
rect 35690 -630 35720 -600
rect 35775 -580 35805 -550
rect 35775 -680 35805 -650
rect 35860 -530 35890 -500
rect 35860 -630 35890 -600
rect 35945 -580 35975 -550
rect 35945 -680 35975 -650
rect 36030 -530 36060 -500
rect 36030 -630 36060 -600
rect 36115 -580 36145 -550
rect 36115 -680 36145 -650
rect 36200 -530 36230 -500
rect 36200 -630 36230 -600
rect 36285 -580 36315 -550
rect 36285 -680 36315 -650
rect 36370 -530 36400 -500
rect 36370 -630 36400 -600
rect 36455 -580 36485 -550
rect 36455 -680 36485 -650
rect 36540 -530 36570 -500
rect 36540 -630 36570 -600
rect 36625 -580 36655 -550
rect 36625 -680 36655 -650
rect 36710 -530 36740 -500
rect 36710 -630 36740 -600
rect 36795 -580 36825 -550
rect 36795 -680 36825 -650
rect 36880 -530 36910 -500
rect 36880 -630 36910 -600
rect 36965 -580 36995 -550
rect 36965 -680 36995 -650
rect 37050 -530 37080 -500
rect 37050 -630 37080 -600
rect 37135 -580 37165 -550
rect 37135 -680 37165 -650
rect 37220 -530 37250 -500
rect 37220 -630 37250 -600
rect 37305 -580 37335 -550
rect 37305 -680 37335 -650
rect 37390 -530 37420 -500
rect 37390 -630 37420 -600
rect 37475 -580 37505 -550
rect 37475 -680 37505 -650
rect 37560 -530 37590 -500
rect 37560 -630 37590 -600
rect 37645 -580 37675 -550
rect 37645 -680 37675 -650
rect 37730 -530 37760 -500
rect 37730 -630 37760 -600
rect 37815 -580 37845 -550
rect 37815 -680 37845 -650
rect 37900 -530 37930 -500
rect 37900 -630 37930 -600
rect 37985 -580 38015 -550
rect 37985 -680 38015 -650
rect 38070 -530 38100 -500
rect 38070 -630 38100 -600
rect 38155 -580 38185 -550
rect 38155 -680 38185 -650
rect 38240 -530 38270 -500
rect 38240 -630 38270 -600
rect 38325 -580 38355 -550
rect 38325 -680 38355 -650
rect 38410 -530 38440 -500
rect 38410 -630 38440 -600
rect 38495 -580 38525 -550
rect 38495 -680 38525 -650
rect 38580 -530 38610 -500
rect 38580 -630 38610 -600
rect 38665 -580 38695 -550
rect 38665 -680 38695 -650
rect 38750 -530 38780 -500
rect 38750 -630 38780 -600
rect 38835 -580 38865 -550
rect 38835 -680 38865 -650
rect 38920 -530 38950 -500
rect 38920 -630 38950 -600
rect 39005 -580 39035 -550
rect 39005 -680 39035 -650
rect 39090 -530 39120 -500
rect 39090 -630 39120 -600
rect 39175 -580 39205 -550
rect 39175 -680 39205 -650
rect 39260 -530 39290 -500
rect 39260 -630 39290 -600
rect 39345 -580 39375 -550
rect 39345 -680 39375 -650
rect 39430 -530 39460 -500
rect 39430 -630 39460 -600
rect 39515 -580 39545 -550
rect 39515 -680 39545 -650
rect 39600 -530 39630 -500
rect 39600 -630 39630 -600
rect 39685 -580 39715 -550
rect 39685 -680 39715 -650
rect 39770 -530 39800 -500
rect 39770 -630 39800 -600
rect 39855 -580 39885 -550
rect 39855 -680 39885 -650
rect 39940 -530 39970 -500
rect 39940 -630 39970 -600
rect 40025 -580 40055 -550
rect 40025 -680 40055 -650
rect 40110 -530 40140 -500
rect 40110 -630 40140 -600
rect 40195 -580 40225 -550
rect 40195 -680 40225 -650
rect 40280 -530 40310 -500
rect 40280 -630 40310 -600
rect 40365 -580 40395 -550
rect 40365 -680 40395 -650
rect 40450 -530 40480 -500
rect 40450 -630 40480 -600
rect 40535 -580 40565 -550
rect 40535 -680 40565 -650
rect 40620 -530 40650 -500
rect 40620 -630 40650 -600
rect 40705 -580 40735 -550
rect 40705 -680 40735 -650
rect 40790 -530 40820 -500
rect 40790 -630 40820 -600
rect 40875 -580 40905 -550
rect 40875 -680 40905 -650
rect 40960 -530 40990 -500
rect 40960 -630 40990 -600
rect 41045 -580 41075 -550
rect 41045 -680 41075 -650
rect 41130 -530 41160 -500
rect 41130 -630 41160 -600
rect 41215 -580 41245 -550
rect 41215 -680 41245 -650
rect 41300 -530 41330 -500
rect 41300 -630 41330 -600
rect 41385 -580 41415 -550
rect 41385 -680 41415 -650
rect 41470 -530 41500 -500
rect 41470 -630 41500 -600
rect 41555 -580 41585 -550
rect 41555 -680 41585 -650
rect 41640 -530 41670 -500
rect 41640 -630 41670 -600
rect 41725 -580 41755 -550
rect 41725 -680 41755 -650
rect 41810 -530 41840 -500
rect 41810 -630 41840 -600
rect 41895 -580 41925 -550
rect 41895 -680 41925 -650
rect 41980 -530 42010 -500
rect 41980 -630 42010 -600
rect 42065 -580 42095 -550
rect 42065 -680 42095 -650
rect 42150 -530 42180 -500
rect 42150 -630 42180 -600
rect 42235 -580 42265 -550
rect 42235 -680 42265 -650
rect 42320 -530 42350 -500
rect 42320 -630 42350 -600
rect 42405 -580 42435 -550
rect 42405 -680 42435 -650
rect 42490 -530 42520 -500
rect 42490 -630 42520 -600
rect 42575 -580 42605 -550
rect 42575 -680 42605 -650
rect 42660 -530 42690 -500
rect 42660 -630 42690 -600
rect 42745 -580 42775 -550
rect 42745 -680 42775 -650
rect 42830 -530 42860 -500
rect 42830 -630 42860 -600
rect 42915 -580 42945 -550
rect 42915 -680 42945 -650
rect 43000 -530 43030 -500
rect 43000 -630 43030 -600
rect 43085 -580 43115 -550
rect 43085 -680 43115 -650
rect 43170 -530 43200 -500
rect 43170 -630 43200 -600
rect 43255 -580 43285 -550
rect 43255 -680 43285 -650
rect 43340 -530 43370 -500
rect 43340 -630 43370 -600
rect 43425 -580 43455 -550
rect 43425 -680 43455 -650
rect 43510 -530 43540 -500
rect 43510 -630 43540 -600
rect 43595 -580 43625 -550
rect 43595 -680 43625 -650
<< metal1 >>
rect 25 55 75 65
rect 25 15 35 55
rect 65 15 75 55
rect 25 5 75 15
rect 90 -30 140 215
rect 215 205 265 215
rect 215 175 225 205
rect 255 175 265 205
rect 215 165 265 175
rect 385 205 435 215
rect 385 175 395 205
rect 425 175 435 205
rect 385 165 435 175
rect 555 205 605 215
rect 555 175 565 205
rect 595 175 605 205
rect 555 165 605 175
rect 750 205 800 215
rect 750 175 760 205
rect 790 175 800 205
rect 750 165 800 175
rect 920 205 970 215
rect 920 175 930 205
rect 960 175 970 205
rect 920 165 970 175
rect 1090 205 1140 215
rect 1090 175 1100 205
rect 1130 175 1140 205
rect 1090 165 1140 175
rect 1260 205 1310 215
rect 1260 175 1270 205
rect 1300 175 1310 205
rect 1260 165 1310 175
rect 1430 205 1480 215
rect 1430 175 1440 205
rect 1470 175 1480 205
rect 1430 165 1480 175
rect 1600 205 1650 215
rect 1600 175 1610 205
rect 1640 175 1650 205
rect 1600 165 1650 175
rect 1770 205 1820 215
rect 1770 175 1780 205
rect 1810 175 1820 205
rect 1770 165 1820 175
rect 1940 205 1990 215
rect 1940 175 1950 205
rect 1980 175 1990 205
rect 1940 165 1990 175
rect 2110 205 2160 215
rect 2110 175 2120 205
rect 2150 175 2160 205
rect 2110 165 2160 175
rect 2260 205 2310 215
rect 2260 175 2270 205
rect 2300 175 2310 205
rect 2260 165 2310 175
rect 2430 205 2480 215
rect 2430 175 2440 205
rect 2470 175 2480 205
rect 2430 165 2480 175
rect 2600 205 2650 215
rect 2600 175 2610 205
rect 2640 175 2650 205
rect 2600 165 2650 175
rect 2770 205 2820 215
rect 2770 175 2780 205
rect 2810 175 2820 205
rect 2770 165 2820 175
rect 2940 205 2990 215
rect 2940 175 2950 205
rect 2980 175 2990 205
rect 2940 165 2990 175
rect 3110 205 3160 215
rect 3110 175 3120 205
rect 3150 175 3160 205
rect 3110 165 3160 175
rect 3280 205 3330 215
rect 3280 175 3290 205
rect 3320 175 3330 205
rect 3280 165 3330 175
rect 3450 205 3500 215
rect 3450 175 3460 205
rect 3490 175 3500 205
rect 3450 165 3500 175
rect 3620 205 3670 215
rect 3620 175 3630 205
rect 3660 175 3670 205
rect 3620 165 3670 175
rect 3790 205 3840 215
rect 3790 175 3800 205
rect 3830 175 3840 205
rect 3790 165 3840 175
rect 3960 205 4010 215
rect 3960 175 3970 205
rect 4000 175 4010 205
rect 3960 165 4010 175
rect 4130 205 4180 215
rect 4130 175 4140 205
rect 4170 175 4180 205
rect 4130 165 4180 175
rect 4300 205 4350 215
rect 4300 175 4310 205
rect 4340 175 4350 205
rect 4300 165 4350 175
rect 4470 205 4520 215
rect 4470 175 4480 205
rect 4510 175 4520 205
rect 4470 165 4520 175
rect 4640 205 4690 215
rect 4640 175 4650 205
rect 4680 175 4690 205
rect 4640 165 4690 175
rect 4810 205 4860 215
rect 4810 175 4820 205
rect 4850 175 4860 205
rect 4810 165 4860 175
rect 4980 205 5030 215
rect 4980 175 4990 205
rect 5020 175 5030 205
rect 4980 165 5030 175
rect 5150 205 5200 215
rect 5150 175 5160 205
rect 5190 175 5200 205
rect 5150 165 5200 175
rect 5320 205 5370 215
rect 5320 175 5330 205
rect 5360 175 5370 205
rect 5320 165 5370 175
rect 5490 205 5540 215
rect 5490 175 5500 205
rect 5530 175 5540 205
rect 5490 165 5540 175
rect 5660 205 5710 215
rect 5660 175 5670 205
rect 5700 175 5710 205
rect 5660 165 5710 175
rect 5830 205 5880 215
rect 5830 175 5840 205
rect 5870 175 5880 205
rect 5830 165 5880 175
rect 6000 205 6050 215
rect 6000 175 6010 205
rect 6040 175 6050 205
rect 6000 165 6050 175
rect 6170 205 6220 215
rect 6170 175 6180 205
rect 6210 175 6220 205
rect 6170 165 6220 175
rect 6340 205 6390 215
rect 6340 175 6350 205
rect 6380 175 6390 205
rect 6340 165 6390 175
rect 6510 205 6560 215
rect 6510 175 6520 205
rect 6550 175 6560 205
rect 6510 165 6560 175
rect 6680 205 6730 215
rect 6680 175 6690 205
rect 6720 175 6730 205
rect 6680 165 6730 175
rect 6850 205 6900 215
rect 6850 175 6860 205
rect 6890 175 6900 205
rect 6850 165 6900 175
rect 7020 205 7070 215
rect 7020 175 7030 205
rect 7060 175 7070 205
rect 7020 165 7070 175
rect 7190 205 7240 215
rect 7190 175 7200 205
rect 7230 175 7240 205
rect 7190 165 7240 175
rect 7360 205 7410 215
rect 7360 175 7370 205
rect 7400 175 7410 205
rect 7360 165 7410 175
rect 7530 205 7580 215
rect 7530 175 7540 205
rect 7570 175 7580 205
rect 7530 165 7580 175
rect 7700 205 7750 215
rect 7700 175 7710 205
rect 7740 175 7750 205
rect 7700 165 7750 175
rect 7850 205 7900 215
rect 7850 175 7860 205
rect 7890 175 7900 205
rect 7850 165 7900 175
rect 8020 205 8070 215
rect 8020 175 8030 205
rect 8060 175 8070 205
rect 8020 165 8070 175
rect 8190 205 8240 215
rect 8190 175 8200 205
rect 8230 175 8240 205
rect 8190 165 8240 175
rect 8360 205 8410 215
rect 8360 175 8370 205
rect 8400 175 8410 205
rect 8360 165 8410 175
rect 8530 205 8580 215
rect 8530 175 8540 205
rect 8570 175 8580 205
rect 8530 165 8580 175
rect 8700 205 8750 215
rect 8700 175 8710 205
rect 8740 175 8750 205
rect 8700 165 8750 175
rect 8870 205 8920 215
rect 8870 175 8880 205
rect 8910 175 8920 205
rect 8870 165 8920 175
rect 9040 205 9090 215
rect 9040 175 9050 205
rect 9080 175 9090 205
rect 9040 165 9090 175
rect 9210 205 9260 215
rect 9210 175 9220 205
rect 9250 175 9260 205
rect 9210 165 9260 175
rect 9380 205 9430 215
rect 9380 175 9390 205
rect 9420 175 9430 205
rect 9380 165 9430 175
rect 9550 205 9600 215
rect 9550 175 9560 205
rect 9590 175 9600 205
rect 9550 165 9600 175
rect 9720 205 9770 215
rect 9720 175 9730 205
rect 9760 175 9770 205
rect 9720 165 9770 175
rect 9890 205 9940 215
rect 9890 175 9900 205
rect 9930 175 9940 205
rect 9890 165 9940 175
rect 10060 205 10110 215
rect 10060 175 10070 205
rect 10100 175 10110 205
rect 10060 165 10110 175
rect 10230 205 10280 215
rect 10230 175 10240 205
rect 10270 175 10280 205
rect 10230 165 10280 175
rect 10400 205 10450 215
rect 10400 175 10410 205
rect 10440 175 10450 205
rect 10400 165 10450 175
rect 10570 205 10620 215
rect 10570 175 10580 205
rect 10610 175 10620 205
rect 10570 165 10620 175
rect 10740 205 10790 215
rect 10740 175 10750 205
rect 10780 175 10790 205
rect 10740 165 10790 175
rect 10910 205 10960 215
rect 10910 175 10920 205
rect 10950 175 10960 205
rect 10910 165 10960 175
rect 11080 205 11130 215
rect 11080 175 11090 205
rect 11120 175 11130 205
rect 11080 165 11130 175
rect 11250 205 11300 215
rect 11250 175 11260 205
rect 11290 175 11300 205
rect 11250 165 11300 175
rect 11420 205 11470 215
rect 11420 175 11430 205
rect 11460 175 11470 205
rect 11420 165 11470 175
rect 11590 205 11640 215
rect 11590 175 11600 205
rect 11630 175 11640 205
rect 11590 165 11640 175
rect 11760 205 11810 215
rect 11760 175 11770 205
rect 11800 175 11810 205
rect 11760 165 11810 175
rect 11930 205 11980 215
rect 11930 175 11940 205
rect 11970 175 11980 205
rect 11930 165 11980 175
rect 12100 205 12150 215
rect 12100 175 12110 205
rect 12140 175 12150 205
rect 12100 165 12150 175
rect 12270 205 12320 215
rect 12270 175 12280 205
rect 12310 175 12320 205
rect 12270 165 12320 175
rect 12440 205 12490 215
rect 12440 175 12450 205
rect 12480 175 12490 205
rect 12440 165 12490 175
rect 12610 205 12660 215
rect 12610 175 12620 205
rect 12650 175 12660 205
rect 12610 165 12660 175
rect 12780 205 12830 215
rect 12780 175 12790 205
rect 12820 175 12830 205
rect 12780 165 12830 175
rect 12950 205 13000 215
rect 12950 175 12960 205
rect 12990 175 13000 205
rect 12950 165 13000 175
rect 13120 205 13170 215
rect 13120 175 13130 205
rect 13160 175 13170 205
rect 13120 165 13170 175
rect 13290 205 13340 215
rect 13290 175 13300 205
rect 13330 175 13340 205
rect 13290 165 13340 175
rect 13460 205 13510 215
rect 13460 175 13470 205
rect 13500 175 13510 205
rect 13460 165 13510 175
rect 13630 205 13680 215
rect 13630 175 13640 205
rect 13670 175 13680 205
rect 13630 165 13680 175
rect 13800 205 13850 215
rect 13800 175 13810 205
rect 13840 175 13850 205
rect 13800 165 13850 175
rect 13970 205 14020 215
rect 13970 175 13980 205
rect 14010 175 14020 205
rect 13970 165 14020 175
rect 14140 205 14190 215
rect 14140 175 14150 205
rect 14180 175 14190 205
rect 14140 165 14190 175
rect 14310 205 14360 215
rect 14310 175 14320 205
rect 14350 175 14360 205
rect 14310 165 14360 175
rect 14480 205 14530 215
rect 14480 175 14490 205
rect 14520 175 14530 205
rect 14480 165 14530 175
rect 14650 205 14700 215
rect 14650 175 14660 205
rect 14690 175 14700 205
rect 14650 165 14700 175
rect 14820 205 14870 215
rect 14820 175 14830 205
rect 14860 175 14870 205
rect 14820 165 14870 175
rect 14990 205 15040 215
rect 14990 175 15000 205
rect 15030 175 15040 205
rect 14990 165 15040 175
rect 15160 205 15210 215
rect 15160 175 15170 205
rect 15200 175 15210 205
rect 15160 165 15210 175
rect 15330 205 15380 215
rect 15330 175 15340 205
rect 15370 175 15380 205
rect 15330 165 15380 175
rect 15500 205 15550 215
rect 15500 175 15510 205
rect 15540 175 15550 205
rect 15500 165 15550 175
rect 15670 205 15720 215
rect 15670 175 15680 205
rect 15710 175 15720 205
rect 15670 165 15720 175
rect 15840 205 15890 215
rect 15840 175 15850 205
rect 15880 175 15890 205
rect 15840 165 15890 175
rect 16010 205 16060 215
rect 16010 175 16020 205
rect 16050 175 16060 205
rect 16010 165 16060 175
rect 16180 205 16230 215
rect 16180 175 16190 205
rect 16220 175 16230 205
rect 16180 165 16230 175
rect 16350 205 16400 215
rect 16350 175 16360 205
rect 16390 175 16400 205
rect 16350 165 16400 175
rect 16520 205 16570 215
rect 16520 175 16530 205
rect 16560 175 16570 205
rect 16520 165 16570 175
rect 16690 205 16740 215
rect 16690 175 16700 205
rect 16730 175 16740 205
rect 16690 165 16740 175
rect 16860 205 16910 215
rect 16860 175 16870 205
rect 16900 175 16910 205
rect 16860 165 16910 175
rect 17030 205 17080 215
rect 17030 175 17040 205
rect 17070 175 17080 205
rect 17030 165 17080 175
rect 17200 205 17250 215
rect 17200 175 17210 205
rect 17240 175 17250 205
rect 17200 165 17250 175
rect 17370 205 17420 215
rect 17370 175 17380 205
rect 17410 175 17420 205
rect 17370 165 17420 175
rect 17540 205 17590 215
rect 17540 175 17550 205
rect 17580 175 17590 205
rect 17540 165 17590 175
rect 17710 205 17760 215
rect 17710 175 17720 205
rect 17750 175 17760 205
rect 17710 165 17760 175
rect 17880 205 17930 215
rect 17880 175 17890 205
rect 17920 175 17930 205
rect 17880 165 17930 175
rect 18050 205 18100 215
rect 18050 175 18060 205
rect 18090 175 18100 205
rect 18050 165 18100 175
rect 18220 205 18270 215
rect 18220 175 18230 205
rect 18260 175 18270 205
rect 18220 165 18270 175
rect 18390 205 18440 215
rect 18390 175 18400 205
rect 18430 175 18440 205
rect 18390 165 18440 175
rect 18560 205 18610 215
rect 18560 175 18570 205
rect 18600 175 18610 205
rect 18560 165 18610 175
rect 18730 205 18780 215
rect 18730 175 18740 205
rect 18770 175 18780 205
rect 18730 165 18780 175
rect 18900 205 18950 215
rect 18900 175 18910 205
rect 18940 175 18950 205
rect 18900 165 18950 175
rect 19070 205 19120 215
rect 19070 175 19080 205
rect 19110 175 19120 205
rect 19070 165 19120 175
rect 19240 205 19290 215
rect 19240 175 19250 205
rect 19280 175 19290 205
rect 19240 165 19290 175
rect 19410 205 19460 215
rect 19410 175 19420 205
rect 19450 175 19460 205
rect 19410 165 19460 175
rect 19580 205 19630 215
rect 19580 175 19590 205
rect 19620 175 19630 205
rect 19580 165 19630 175
rect 19750 205 19800 215
rect 19750 175 19760 205
rect 19790 175 19800 205
rect 19750 165 19800 175
rect 19920 205 19970 215
rect 19920 175 19930 205
rect 19960 175 19970 205
rect 19920 165 19970 175
rect 20090 205 20140 215
rect 20090 175 20100 205
rect 20130 175 20140 205
rect 20090 165 20140 175
rect 20260 205 20310 215
rect 20260 175 20270 205
rect 20300 175 20310 205
rect 20260 165 20310 175
rect 20430 205 20480 215
rect 20430 175 20440 205
rect 20470 175 20480 205
rect 20430 165 20480 175
rect 20600 205 20650 215
rect 20600 175 20610 205
rect 20640 175 20650 205
rect 20600 165 20650 175
rect 20770 205 20820 215
rect 20770 175 20780 205
rect 20810 175 20820 205
rect 20770 165 20820 175
rect 20940 205 20990 215
rect 20940 175 20950 205
rect 20980 175 20990 205
rect 20940 165 20990 175
rect 21110 205 21160 215
rect 21110 175 21120 205
rect 21150 175 21160 205
rect 21110 165 21160 175
rect 21280 205 21330 215
rect 21280 175 21290 205
rect 21320 175 21330 205
rect 21280 165 21330 175
rect 21450 205 21500 215
rect 21450 175 21460 205
rect 21490 175 21500 205
rect 21450 165 21500 175
rect 21620 205 21670 215
rect 21620 175 21630 205
rect 21660 175 21670 205
rect 21620 165 21670 175
rect 21790 205 21840 215
rect 21790 175 21800 205
rect 21830 175 21840 205
rect 21790 165 21840 175
rect 21960 205 22010 215
rect 21960 175 21970 205
rect 22000 175 22010 205
rect 21960 165 22010 175
rect 22130 205 22180 215
rect 22130 175 22140 205
rect 22170 175 22180 205
rect 22130 165 22180 175
rect 22300 205 22350 215
rect 22300 175 22310 205
rect 22340 175 22350 205
rect 22300 165 22350 175
rect 22470 205 22520 215
rect 22470 175 22480 205
rect 22510 175 22520 205
rect 22470 165 22520 175
rect 22640 205 22690 215
rect 22640 175 22650 205
rect 22680 175 22690 205
rect 22640 165 22690 175
rect 22810 205 22860 215
rect 22810 175 22820 205
rect 22850 175 22860 205
rect 22810 165 22860 175
rect 22980 205 23030 215
rect 22980 175 22990 205
rect 23020 175 23030 205
rect 22980 165 23030 175
rect 23150 205 23200 215
rect 23150 175 23160 205
rect 23190 175 23200 205
rect 23150 165 23200 175
rect 23320 205 23370 215
rect 23320 175 23330 205
rect 23360 175 23370 205
rect 23320 165 23370 175
rect 23490 205 23540 215
rect 23490 175 23500 205
rect 23530 175 23540 205
rect 23490 165 23540 175
rect 23660 205 23710 215
rect 23660 175 23670 205
rect 23700 175 23710 205
rect 23660 165 23710 175
rect 23830 205 23880 215
rect 23830 175 23840 205
rect 23870 175 23880 205
rect 23830 165 23880 175
rect 24000 205 24050 215
rect 24000 175 24010 205
rect 24040 175 24050 205
rect 24000 165 24050 175
rect 24170 205 24220 215
rect 24170 175 24180 205
rect 24210 175 24220 205
rect 24170 165 24220 175
rect 24340 205 24390 215
rect 24340 175 24350 205
rect 24380 175 24390 205
rect 24340 165 24390 175
rect 24510 205 24560 215
rect 24510 175 24520 205
rect 24550 175 24560 205
rect 24510 165 24560 175
rect 24680 205 24730 215
rect 24680 175 24690 205
rect 24720 175 24730 205
rect 24680 165 24730 175
rect 24850 205 24900 215
rect 24850 175 24860 205
rect 24890 175 24900 205
rect 24850 165 24900 175
rect 25020 205 25070 215
rect 25020 175 25030 205
rect 25060 175 25070 205
rect 25020 165 25070 175
rect 25190 205 25240 215
rect 25190 175 25200 205
rect 25230 175 25240 205
rect 25190 165 25240 175
rect 25360 205 25410 215
rect 25360 175 25370 205
rect 25400 175 25410 205
rect 25360 165 25410 175
rect 25530 205 25580 215
rect 25530 175 25540 205
rect 25570 175 25580 205
rect 25530 165 25580 175
rect 25700 205 25750 215
rect 25700 175 25710 205
rect 25740 175 25750 205
rect 25700 165 25750 175
rect 25870 205 25920 215
rect 25870 175 25880 205
rect 25910 175 25920 205
rect 25870 165 25920 175
rect 26040 205 26090 215
rect 26040 175 26050 205
rect 26080 175 26090 205
rect 26040 165 26090 175
rect 26210 205 26260 215
rect 26210 175 26220 205
rect 26250 175 26260 205
rect 26210 165 26260 175
rect 26380 205 26430 215
rect 26380 175 26390 205
rect 26420 175 26430 205
rect 26380 165 26430 175
rect 26550 205 26600 215
rect 26550 175 26560 205
rect 26590 175 26600 205
rect 26550 165 26600 175
rect 26720 205 26770 215
rect 26720 175 26730 205
rect 26760 175 26770 205
rect 26720 165 26770 175
rect 26890 205 26940 215
rect 26890 175 26900 205
rect 26930 175 26940 205
rect 26890 165 26940 175
rect 27060 205 27110 215
rect 27060 175 27070 205
rect 27100 175 27110 205
rect 27060 165 27110 175
rect 27230 205 27280 215
rect 27230 175 27240 205
rect 27270 175 27280 205
rect 27230 165 27280 175
rect 27400 205 27450 215
rect 27400 175 27410 205
rect 27440 175 27450 205
rect 27400 165 27450 175
rect 27570 205 27620 215
rect 27570 175 27580 205
rect 27610 175 27620 205
rect 27570 165 27620 175
rect 27740 205 27790 215
rect 27740 175 27750 205
rect 27780 175 27790 205
rect 27740 165 27790 175
rect 27910 205 27960 215
rect 27910 175 27920 205
rect 27950 175 27960 205
rect 27910 165 27960 175
rect 28080 205 28130 215
rect 28080 175 28090 205
rect 28120 175 28130 205
rect 28080 165 28130 175
rect 28250 205 28300 215
rect 28250 175 28260 205
rect 28290 175 28300 205
rect 28250 165 28300 175
rect 28420 205 28470 215
rect 28420 175 28430 205
rect 28460 175 28470 205
rect 28420 165 28470 175
rect 28590 205 28640 215
rect 28590 175 28600 205
rect 28630 175 28640 205
rect 28590 165 28640 175
rect 28760 205 28810 215
rect 28760 175 28770 205
rect 28800 175 28810 205
rect 28760 165 28810 175
rect 28930 205 28980 215
rect 28930 175 28940 205
rect 28970 175 28980 205
rect 28930 165 28980 175
rect 29100 205 29150 215
rect 29100 175 29110 205
rect 29140 175 29150 205
rect 29100 165 29150 175
rect 29270 205 29320 215
rect 29270 175 29280 205
rect 29310 175 29320 205
rect 29270 165 29320 175
rect 29440 205 29490 215
rect 29440 175 29450 205
rect 29480 175 29490 205
rect 29440 165 29490 175
rect 29610 205 29660 215
rect 29610 175 29620 205
rect 29650 175 29660 205
rect 29610 165 29660 175
rect 300 155 350 160
rect 300 125 310 155
rect 340 125 350 155
rect 300 100 350 125
rect 300 65 310 100
rect 340 65 350 100
rect 215 40 265 50
rect 215 10 225 40
rect 255 10 265 40
rect 215 0 265 10
rect 300 40 350 65
rect 470 155 520 160
rect 470 125 480 155
rect 510 125 520 155
rect 470 100 520 125
rect 470 65 480 100
rect 510 65 520 100
rect 300 10 310 40
rect 340 10 350 40
rect 300 0 350 10
rect 385 40 435 50
rect 385 10 395 40
rect 425 10 435 40
rect 385 0 435 10
rect 470 40 520 65
rect 835 155 885 160
rect 835 125 845 155
rect 875 125 885 155
rect 835 100 885 125
rect 835 65 845 100
rect 875 65 885 100
rect 470 10 480 40
rect 510 10 520 40
rect 470 0 520 10
rect 555 40 605 50
rect 555 10 565 40
rect 595 10 605 40
rect 555 0 605 10
rect 750 40 800 50
rect 750 10 760 40
rect 790 10 800 40
rect 750 0 800 10
rect 835 40 885 65
rect 1005 155 1055 160
rect 1005 125 1015 155
rect 1045 125 1055 155
rect 1005 100 1055 125
rect 1005 65 1015 100
rect 1045 65 1055 100
rect 835 10 845 40
rect 875 10 885 40
rect 835 0 885 10
rect 920 40 970 50
rect 920 10 930 40
rect 960 10 970 40
rect 920 0 970 10
rect 1005 40 1055 65
rect 1175 155 1225 160
rect 1175 125 1185 155
rect 1215 125 1225 155
rect 1175 100 1225 125
rect 1175 65 1185 100
rect 1215 65 1225 100
rect 1005 10 1015 40
rect 1045 10 1055 40
rect 1005 0 1055 10
rect 1090 40 1140 50
rect 1090 10 1100 40
rect 1130 10 1140 40
rect 1090 0 1140 10
rect 1175 40 1225 65
rect 1345 155 1395 160
rect 1345 125 1355 155
rect 1385 125 1395 155
rect 1345 100 1395 125
rect 1345 65 1355 100
rect 1385 65 1395 100
rect 1175 10 1185 40
rect 1215 10 1225 40
rect 1175 0 1225 10
rect 1260 40 1310 50
rect 1260 10 1270 40
rect 1300 10 1310 40
rect 1260 0 1310 10
rect 1345 40 1395 65
rect 1515 155 1565 160
rect 1515 125 1525 155
rect 1555 125 1565 155
rect 1515 100 1565 125
rect 1515 65 1525 100
rect 1555 65 1565 100
rect 1345 10 1355 40
rect 1385 10 1395 40
rect 1345 0 1395 10
rect 1430 40 1480 50
rect 1430 10 1440 40
rect 1470 10 1480 40
rect 1430 0 1480 10
rect 1515 40 1565 65
rect 1685 155 1735 160
rect 1685 125 1695 155
rect 1725 125 1735 155
rect 1685 100 1735 125
rect 1685 65 1695 100
rect 1725 65 1735 100
rect 1515 10 1525 40
rect 1555 10 1565 40
rect 1515 0 1565 10
rect 1600 40 1650 50
rect 1600 10 1610 40
rect 1640 10 1650 40
rect 1600 0 1650 10
rect 1685 40 1735 65
rect 1855 155 1905 160
rect 1855 125 1865 155
rect 1895 125 1905 155
rect 1855 100 1905 125
rect 1855 65 1865 100
rect 1895 65 1905 100
rect 1685 10 1695 40
rect 1725 10 1735 40
rect 1685 0 1735 10
rect 1770 40 1820 50
rect 1770 10 1780 40
rect 1810 10 1820 40
rect 1770 0 1820 10
rect 1855 40 1905 65
rect 2025 155 2075 160
rect 2025 125 2035 155
rect 2065 125 2075 155
rect 2025 100 2075 125
rect 2025 65 2035 100
rect 2065 65 2075 100
rect 1855 10 1865 40
rect 1895 10 1905 40
rect 1855 0 1905 10
rect 1940 40 1990 50
rect 1940 10 1950 40
rect 1980 10 1990 40
rect 1940 0 1990 10
rect 2025 40 2075 65
rect 2345 155 2395 160
rect 2345 125 2355 155
rect 2385 125 2395 155
rect 2345 100 2395 125
rect 2345 65 2355 100
rect 2385 65 2395 100
rect 2025 10 2035 40
rect 2065 10 2075 40
rect 2025 0 2075 10
rect 2110 40 2160 50
rect 2110 10 2120 40
rect 2150 10 2160 40
rect 2110 0 2160 10
rect 2260 40 2310 50
rect 2260 10 2270 40
rect 2300 10 2310 40
rect 2260 0 2310 10
rect 2345 40 2395 65
rect 2515 155 2565 160
rect 2515 125 2525 155
rect 2555 125 2565 155
rect 2515 100 2565 125
rect 2515 65 2525 100
rect 2555 65 2565 100
rect 2345 10 2355 40
rect 2385 10 2395 40
rect 2345 0 2395 10
rect 2430 40 2480 50
rect 2430 10 2440 40
rect 2470 10 2480 40
rect 2430 0 2480 10
rect 2515 40 2565 65
rect 2685 155 2735 160
rect 2685 125 2695 155
rect 2725 125 2735 155
rect 2685 100 2735 125
rect 2685 65 2695 100
rect 2725 65 2735 100
rect 2515 10 2525 40
rect 2555 10 2565 40
rect 2515 0 2565 10
rect 2600 40 2650 50
rect 2600 10 2610 40
rect 2640 10 2650 40
rect 2600 0 2650 10
rect 2685 40 2735 65
rect 2855 155 2905 160
rect 2855 125 2865 155
rect 2895 125 2905 155
rect 2855 100 2905 125
rect 2855 65 2865 100
rect 2895 65 2905 100
rect 2685 10 2695 40
rect 2725 10 2735 40
rect 2685 0 2735 10
rect 2770 40 2820 50
rect 2770 10 2780 40
rect 2810 10 2820 40
rect 2770 0 2820 10
rect 2855 40 2905 65
rect 3025 155 3075 160
rect 3025 125 3035 155
rect 3065 125 3075 155
rect 3025 100 3075 125
rect 3025 65 3035 100
rect 3065 65 3075 100
rect 2855 10 2865 40
rect 2895 10 2905 40
rect 2855 0 2905 10
rect 2940 40 2990 50
rect 2940 10 2950 40
rect 2980 10 2990 40
rect 2940 0 2990 10
rect 3025 40 3075 65
rect 3195 155 3245 160
rect 3195 125 3205 155
rect 3235 125 3245 155
rect 3195 100 3245 125
rect 3195 65 3205 100
rect 3235 65 3245 100
rect 3025 10 3035 40
rect 3065 10 3075 40
rect 3025 0 3075 10
rect 3110 40 3160 50
rect 3110 10 3120 40
rect 3150 10 3160 40
rect 3110 0 3160 10
rect 3195 40 3245 65
rect 3365 155 3415 160
rect 3365 125 3375 155
rect 3405 125 3415 155
rect 3365 100 3415 125
rect 3365 65 3375 100
rect 3405 65 3415 100
rect 3195 10 3205 40
rect 3235 10 3245 40
rect 3195 0 3245 10
rect 3280 40 3330 50
rect 3280 10 3290 40
rect 3320 10 3330 40
rect 3280 0 3330 10
rect 3365 40 3415 65
rect 3535 155 3585 160
rect 3535 125 3545 155
rect 3575 125 3585 155
rect 3535 100 3585 125
rect 3535 65 3545 100
rect 3575 65 3585 100
rect 3365 10 3375 40
rect 3405 10 3415 40
rect 3365 0 3415 10
rect 3450 40 3500 50
rect 3450 10 3460 40
rect 3490 10 3500 40
rect 3450 0 3500 10
rect 3535 40 3585 65
rect 3705 155 3755 160
rect 3705 125 3715 155
rect 3745 125 3755 155
rect 3705 100 3755 125
rect 3705 65 3715 100
rect 3745 65 3755 100
rect 3535 10 3545 40
rect 3575 10 3585 40
rect 3535 0 3585 10
rect 3620 40 3670 50
rect 3620 10 3630 40
rect 3660 10 3670 40
rect 3620 0 3670 10
rect 3705 40 3755 65
rect 3875 155 3925 160
rect 3875 125 3885 155
rect 3915 125 3925 155
rect 3875 100 3925 125
rect 3875 65 3885 100
rect 3915 65 3925 100
rect 3705 10 3715 40
rect 3745 10 3755 40
rect 3705 0 3755 10
rect 3790 40 3840 50
rect 3790 10 3800 40
rect 3830 10 3840 40
rect 3790 0 3840 10
rect 3875 40 3925 65
rect 4045 155 4095 160
rect 4045 125 4055 155
rect 4085 125 4095 155
rect 4045 100 4095 125
rect 4045 65 4055 100
rect 4085 65 4095 100
rect 3875 10 3885 40
rect 3915 10 3925 40
rect 3875 0 3925 10
rect 3960 40 4010 50
rect 3960 10 3970 40
rect 4000 10 4010 40
rect 3960 0 4010 10
rect 4045 40 4095 65
rect 4215 155 4265 160
rect 4215 125 4225 155
rect 4255 125 4265 155
rect 4215 100 4265 125
rect 4215 65 4225 100
rect 4255 65 4265 100
rect 4045 10 4055 40
rect 4085 10 4095 40
rect 4045 0 4095 10
rect 4130 40 4180 50
rect 4130 10 4140 40
rect 4170 10 4180 40
rect 4130 0 4180 10
rect 4215 40 4265 65
rect 4385 155 4435 160
rect 4385 125 4395 155
rect 4425 125 4435 155
rect 4385 100 4435 125
rect 4385 65 4395 100
rect 4425 65 4435 100
rect 4215 10 4225 40
rect 4255 10 4265 40
rect 4215 0 4265 10
rect 4300 40 4350 50
rect 4300 10 4310 40
rect 4340 10 4350 40
rect 4300 0 4350 10
rect 4385 40 4435 65
rect 4555 155 4605 160
rect 4555 125 4565 155
rect 4595 125 4605 155
rect 4555 100 4605 125
rect 4555 65 4565 100
rect 4595 65 4605 100
rect 4385 10 4395 40
rect 4425 10 4435 40
rect 4385 0 4435 10
rect 4470 40 4520 50
rect 4470 10 4480 40
rect 4510 10 4520 40
rect 4470 0 4520 10
rect 4555 40 4605 65
rect 4725 155 4775 160
rect 4725 125 4735 155
rect 4765 125 4775 155
rect 4725 100 4775 125
rect 4725 65 4735 100
rect 4765 65 4775 100
rect 4555 10 4565 40
rect 4595 10 4605 40
rect 4555 0 4605 10
rect 4640 40 4690 50
rect 4640 10 4650 40
rect 4680 10 4690 40
rect 4640 0 4690 10
rect 4725 40 4775 65
rect 4895 155 4945 160
rect 4895 125 4905 155
rect 4935 125 4945 155
rect 4895 100 4945 125
rect 4895 65 4905 100
rect 4935 65 4945 100
rect 4725 10 4735 40
rect 4765 10 4775 40
rect 4725 0 4775 10
rect 4810 40 4860 50
rect 4810 10 4820 40
rect 4850 10 4860 40
rect 4810 0 4860 10
rect 4895 40 4945 65
rect 5065 155 5115 160
rect 5065 125 5075 155
rect 5105 125 5115 155
rect 5065 100 5115 125
rect 5065 65 5075 100
rect 5105 65 5115 100
rect 4895 10 4905 40
rect 4935 10 4945 40
rect 4895 0 4945 10
rect 4980 40 5030 50
rect 4980 10 4990 40
rect 5020 10 5030 40
rect 4980 0 5030 10
rect 5065 40 5115 65
rect 5235 155 5285 160
rect 5235 125 5245 155
rect 5275 125 5285 155
rect 5235 100 5285 125
rect 5235 65 5245 100
rect 5275 65 5285 100
rect 5065 10 5075 40
rect 5105 10 5115 40
rect 5065 0 5115 10
rect 5150 40 5200 50
rect 5150 10 5160 40
rect 5190 10 5200 40
rect 5150 0 5200 10
rect 5235 40 5285 65
rect 5405 155 5455 160
rect 5405 125 5415 155
rect 5445 125 5455 155
rect 5405 100 5455 125
rect 5405 65 5415 100
rect 5445 65 5455 100
rect 5235 10 5245 40
rect 5275 10 5285 40
rect 5235 0 5285 10
rect 5320 40 5370 50
rect 5320 10 5330 40
rect 5360 10 5370 40
rect 5320 0 5370 10
rect 5405 40 5455 65
rect 5575 155 5625 160
rect 5575 125 5585 155
rect 5615 125 5625 155
rect 5575 100 5625 125
rect 5575 65 5585 100
rect 5615 65 5625 100
rect 5405 10 5415 40
rect 5445 10 5455 40
rect 5405 0 5455 10
rect 5490 40 5540 50
rect 5490 10 5500 40
rect 5530 10 5540 40
rect 5490 0 5540 10
rect 5575 40 5625 65
rect 5745 155 5795 160
rect 5745 125 5755 155
rect 5785 125 5795 155
rect 5745 100 5795 125
rect 5745 65 5755 100
rect 5785 65 5795 100
rect 5575 10 5585 40
rect 5615 10 5625 40
rect 5575 0 5625 10
rect 5660 40 5710 50
rect 5660 10 5670 40
rect 5700 10 5710 40
rect 5660 0 5710 10
rect 5745 40 5795 65
rect 5915 155 5965 160
rect 5915 125 5925 155
rect 5955 125 5965 155
rect 5915 100 5965 125
rect 5915 65 5925 100
rect 5955 65 5965 100
rect 5745 10 5755 40
rect 5785 10 5795 40
rect 5745 0 5795 10
rect 5830 40 5880 50
rect 5830 10 5840 40
rect 5870 10 5880 40
rect 5830 0 5880 10
rect 5915 40 5965 65
rect 6085 155 6135 160
rect 6085 125 6095 155
rect 6125 125 6135 155
rect 6085 100 6135 125
rect 6085 65 6095 100
rect 6125 65 6135 100
rect 5915 10 5925 40
rect 5955 10 5965 40
rect 5915 0 5965 10
rect 6000 40 6050 50
rect 6000 10 6010 40
rect 6040 10 6050 40
rect 6000 0 6050 10
rect 6085 40 6135 65
rect 6255 155 6305 160
rect 6255 125 6265 155
rect 6295 125 6305 155
rect 6255 100 6305 125
rect 6255 65 6265 100
rect 6295 65 6305 100
rect 6085 10 6095 40
rect 6125 10 6135 40
rect 6085 0 6135 10
rect 6170 40 6220 50
rect 6170 10 6180 40
rect 6210 10 6220 40
rect 6170 0 6220 10
rect 6255 40 6305 65
rect 6425 155 6475 160
rect 6425 125 6435 155
rect 6465 125 6475 155
rect 6425 100 6475 125
rect 6425 65 6435 100
rect 6465 65 6475 100
rect 6255 10 6265 40
rect 6295 10 6305 40
rect 6255 0 6305 10
rect 6340 40 6390 50
rect 6340 10 6350 40
rect 6380 10 6390 40
rect 6340 0 6390 10
rect 6425 40 6475 65
rect 6595 155 6645 160
rect 6595 125 6605 155
rect 6635 125 6645 155
rect 6595 100 6645 125
rect 6595 65 6605 100
rect 6635 65 6645 100
rect 6425 10 6435 40
rect 6465 10 6475 40
rect 6425 0 6475 10
rect 6510 40 6560 50
rect 6510 10 6520 40
rect 6550 10 6560 40
rect 6510 0 6560 10
rect 6595 40 6645 65
rect 6765 155 6815 160
rect 6765 125 6775 155
rect 6805 125 6815 155
rect 6765 100 6815 125
rect 6765 65 6775 100
rect 6805 65 6815 100
rect 6595 10 6605 40
rect 6635 10 6645 40
rect 6595 0 6645 10
rect 6680 40 6730 50
rect 6680 10 6690 40
rect 6720 10 6730 40
rect 6680 0 6730 10
rect 6765 40 6815 65
rect 6935 155 6985 160
rect 6935 125 6945 155
rect 6975 125 6985 155
rect 6935 100 6985 125
rect 6935 65 6945 100
rect 6975 65 6985 100
rect 6765 10 6775 40
rect 6805 10 6815 40
rect 6765 0 6815 10
rect 6850 40 6900 50
rect 6850 10 6860 40
rect 6890 10 6900 40
rect 6850 0 6900 10
rect 6935 40 6985 65
rect 7105 155 7155 160
rect 7105 125 7115 155
rect 7145 125 7155 155
rect 7105 100 7155 125
rect 7105 65 7115 100
rect 7145 65 7155 100
rect 6935 10 6945 40
rect 6975 10 6985 40
rect 6935 0 6985 10
rect 7020 40 7070 50
rect 7020 10 7030 40
rect 7060 10 7070 40
rect 7020 0 7070 10
rect 7105 40 7155 65
rect 7275 155 7325 160
rect 7275 125 7285 155
rect 7315 125 7325 155
rect 7275 100 7325 125
rect 7275 65 7285 100
rect 7315 65 7325 100
rect 7105 10 7115 40
rect 7145 10 7155 40
rect 7105 0 7155 10
rect 7190 40 7240 50
rect 7190 10 7200 40
rect 7230 10 7240 40
rect 7190 0 7240 10
rect 7275 40 7325 65
rect 7445 155 7495 160
rect 7445 125 7455 155
rect 7485 125 7495 155
rect 7445 100 7495 125
rect 7445 65 7455 100
rect 7485 65 7495 100
rect 7275 10 7285 40
rect 7315 10 7325 40
rect 7275 0 7325 10
rect 7360 40 7410 50
rect 7360 10 7370 40
rect 7400 10 7410 40
rect 7360 0 7410 10
rect 7445 40 7495 65
rect 7615 155 7665 160
rect 7615 125 7625 155
rect 7655 125 7665 155
rect 7615 100 7665 125
rect 7615 65 7625 100
rect 7655 65 7665 100
rect 7445 10 7455 40
rect 7485 10 7495 40
rect 7445 0 7495 10
rect 7530 40 7580 50
rect 7530 10 7540 40
rect 7570 10 7580 40
rect 7530 0 7580 10
rect 7615 40 7665 65
rect 7935 155 7985 160
rect 7935 125 7945 155
rect 7975 125 7985 155
rect 7935 100 7985 125
rect 7935 65 7945 100
rect 7975 65 7985 100
rect 7615 10 7625 40
rect 7655 10 7665 40
rect 7615 0 7665 10
rect 7700 40 7750 50
rect 7700 10 7710 40
rect 7740 10 7750 40
rect 7700 0 7750 10
rect 7850 40 7900 50
rect 7850 10 7860 40
rect 7890 10 7900 40
rect 7850 0 7900 10
rect 7935 40 7985 65
rect 8105 155 8155 160
rect 8105 125 8115 155
rect 8145 125 8155 155
rect 8105 100 8155 125
rect 8105 65 8115 100
rect 8145 65 8155 100
rect 7935 10 7945 40
rect 7975 10 7985 40
rect 7935 0 7985 10
rect 8020 40 8070 50
rect 8020 10 8030 40
rect 8060 10 8070 40
rect 8020 0 8070 10
rect 8105 40 8155 65
rect 8275 155 8325 160
rect 8275 125 8285 155
rect 8315 125 8325 155
rect 8275 100 8325 125
rect 8275 65 8285 100
rect 8315 65 8325 100
rect 8105 10 8115 40
rect 8145 10 8155 40
rect 8105 0 8155 10
rect 8190 40 8240 50
rect 8190 10 8200 40
rect 8230 10 8240 40
rect 8190 0 8240 10
rect 8275 40 8325 65
rect 8445 155 8495 160
rect 8445 125 8455 155
rect 8485 125 8495 155
rect 8445 100 8495 125
rect 8445 65 8455 100
rect 8485 65 8495 100
rect 8275 10 8285 40
rect 8315 10 8325 40
rect 8275 0 8325 10
rect 8360 40 8410 50
rect 8360 10 8370 40
rect 8400 10 8410 40
rect 8360 0 8410 10
rect 8445 40 8495 65
rect 8615 155 8665 160
rect 8615 125 8625 155
rect 8655 125 8665 155
rect 8615 100 8665 125
rect 8615 65 8625 100
rect 8655 65 8665 100
rect 8445 10 8455 40
rect 8485 10 8495 40
rect 8445 0 8495 10
rect 8530 40 8580 50
rect 8530 10 8540 40
rect 8570 10 8580 40
rect 8530 0 8580 10
rect 8615 40 8665 65
rect 8785 155 8835 160
rect 8785 125 8795 155
rect 8825 125 8835 155
rect 8785 100 8835 125
rect 8785 65 8795 100
rect 8825 65 8835 100
rect 8615 10 8625 40
rect 8655 10 8665 40
rect 8615 0 8665 10
rect 8700 40 8750 50
rect 8700 10 8710 40
rect 8740 10 8750 40
rect 8700 0 8750 10
rect 8785 40 8835 65
rect 8955 155 9005 160
rect 8955 125 8965 155
rect 8995 125 9005 155
rect 8955 100 9005 125
rect 8955 65 8965 100
rect 8995 65 9005 100
rect 8785 10 8795 40
rect 8825 10 8835 40
rect 8785 0 8835 10
rect 8870 40 8920 50
rect 8870 10 8880 40
rect 8910 10 8920 40
rect 8870 0 8920 10
rect 8955 40 9005 65
rect 9125 155 9175 160
rect 9125 125 9135 155
rect 9165 125 9175 155
rect 9125 100 9175 125
rect 9125 65 9135 100
rect 9165 65 9175 100
rect 8955 10 8965 40
rect 8995 10 9005 40
rect 8955 0 9005 10
rect 9040 40 9090 50
rect 9040 10 9050 40
rect 9080 10 9090 40
rect 9040 0 9090 10
rect 9125 40 9175 65
rect 9295 155 9345 160
rect 9295 125 9305 155
rect 9335 125 9345 155
rect 9295 100 9345 125
rect 9295 65 9305 100
rect 9335 65 9345 100
rect 9125 10 9135 40
rect 9165 10 9175 40
rect 9125 0 9175 10
rect 9210 40 9260 50
rect 9210 10 9220 40
rect 9250 10 9260 40
rect 9210 0 9260 10
rect 9295 40 9345 65
rect 9465 155 9515 160
rect 9465 125 9475 155
rect 9505 125 9515 155
rect 9465 100 9515 125
rect 9465 65 9475 100
rect 9505 65 9515 100
rect 9295 10 9305 40
rect 9335 10 9345 40
rect 9295 0 9345 10
rect 9380 40 9430 50
rect 9380 10 9390 40
rect 9420 10 9430 40
rect 9380 0 9430 10
rect 9465 40 9515 65
rect 9635 155 9685 160
rect 9635 125 9645 155
rect 9675 125 9685 155
rect 9635 100 9685 125
rect 9635 65 9645 100
rect 9675 65 9685 100
rect 9465 10 9475 40
rect 9505 10 9515 40
rect 9465 0 9515 10
rect 9550 40 9600 50
rect 9550 10 9560 40
rect 9590 10 9600 40
rect 9550 0 9600 10
rect 9635 40 9685 65
rect 9805 155 9855 160
rect 9805 125 9815 155
rect 9845 125 9855 155
rect 9805 100 9855 125
rect 9805 65 9815 100
rect 9845 65 9855 100
rect 9635 10 9645 40
rect 9675 10 9685 40
rect 9635 0 9685 10
rect 9720 40 9770 50
rect 9720 10 9730 40
rect 9760 10 9770 40
rect 9720 0 9770 10
rect 9805 40 9855 65
rect 9975 155 10025 160
rect 9975 125 9985 155
rect 10015 125 10025 155
rect 9975 100 10025 125
rect 9975 65 9985 100
rect 10015 65 10025 100
rect 9805 10 9815 40
rect 9845 10 9855 40
rect 9805 0 9855 10
rect 9890 40 9940 50
rect 9890 10 9900 40
rect 9930 10 9940 40
rect 9890 0 9940 10
rect 9975 40 10025 65
rect 10145 155 10195 160
rect 10145 125 10155 155
rect 10185 125 10195 155
rect 10145 100 10195 125
rect 10145 65 10155 100
rect 10185 65 10195 100
rect 9975 10 9985 40
rect 10015 10 10025 40
rect 9975 0 10025 10
rect 10060 40 10110 50
rect 10060 10 10070 40
rect 10100 10 10110 40
rect 10060 0 10110 10
rect 10145 40 10195 65
rect 10315 155 10365 160
rect 10315 125 10325 155
rect 10355 125 10365 155
rect 10315 100 10365 125
rect 10315 65 10325 100
rect 10355 65 10365 100
rect 10145 10 10155 40
rect 10185 10 10195 40
rect 10145 0 10195 10
rect 10230 40 10280 50
rect 10230 10 10240 40
rect 10270 10 10280 40
rect 10230 0 10280 10
rect 10315 40 10365 65
rect 10485 155 10535 160
rect 10485 125 10495 155
rect 10525 125 10535 155
rect 10485 100 10535 125
rect 10485 65 10495 100
rect 10525 65 10535 100
rect 10315 10 10325 40
rect 10355 10 10365 40
rect 10315 0 10365 10
rect 10400 40 10450 50
rect 10400 10 10410 40
rect 10440 10 10450 40
rect 10400 0 10450 10
rect 10485 40 10535 65
rect 10655 155 10705 160
rect 10655 125 10665 155
rect 10695 125 10705 155
rect 10655 100 10705 125
rect 10655 65 10665 100
rect 10695 65 10705 100
rect 10485 10 10495 40
rect 10525 10 10535 40
rect 10485 0 10535 10
rect 10570 40 10620 50
rect 10570 10 10580 40
rect 10610 10 10620 40
rect 10570 0 10620 10
rect 10655 40 10705 65
rect 10825 155 10875 160
rect 10825 125 10835 155
rect 10865 125 10875 155
rect 10825 100 10875 125
rect 10825 65 10835 100
rect 10865 65 10875 100
rect 10655 10 10665 40
rect 10695 10 10705 40
rect 10655 0 10705 10
rect 10740 40 10790 50
rect 10740 10 10750 40
rect 10780 10 10790 40
rect 10740 0 10790 10
rect 10825 40 10875 65
rect 10995 155 11045 160
rect 10995 125 11005 155
rect 11035 125 11045 155
rect 10995 100 11045 125
rect 10995 65 11005 100
rect 11035 65 11045 100
rect 10825 10 10835 40
rect 10865 10 10875 40
rect 10825 0 10875 10
rect 10910 40 10960 50
rect 10910 10 10920 40
rect 10950 10 10960 40
rect 10910 0 10960 10
rect 10995 40 11045 65
rect 11165 155 11215 160
rect 11165 125 11175 155
rect 11205 125 11215 155
rect 11165 100 11215 125
rect 11165 65 11175 100
rect 11205 65 11215 100
rect 10995 10 11005 40
rect 11035 10 11045 40
rect 10995 0 11045 10
rect 11080 40 11130 50
rect 11080 10 11090 40
rect 11120 10 11130 40
rect 11080 0 11130 10
rect 11165 40 11215 65
rect 11335 155 11385 160
rect 11335 125 11345 155
rect 11375 125 11385 155
rect 11335 100 11385 125
rect 11335 65 11345 100
rect 11375 65 11385 100
rect 11165 10 11175 40
rect 11205 10 11215 40
rect 11165 0 11215 10
rect 11250 40 11300 50
rect 11250 10 11260 40
rect 11290 10 11300 40
rect 11250 0 11300 10
rect 11335 40 11385 65
rect 11505 155 11555 160
rect 11505 125 11515 155
rect 11545 125 11555 155
rect 11505 100 11555 125
rect 11505 65 11515 100
rect 11545 65 11555 100
rect 11335 10 11345 40
rect 11375 10 11385 40
rect 11335 0 11385 10
rect 11420 40 11470 50
rect 11420 10 11430 40
rect 11460 10 11470 40
rect 11420 0 11470 10
rect 11505 40 11555 65
rect 11675 155 11725 160
rect 11675 125 11685 155
rect 11715 125 11725 155
rect 11675 100 11725 125
rect 11675 65 11685 100
rect 11715 65 11725 100
rect 11505 10 11515 40
rect 11545 10 11555 40
rect 11505 0 11555 10
rect 11590 40 11640 50
rect 11590 10 11600 40
rect 11630 10 11640 40
rect 11590 0 11640 10
rect 11675 40 11725 65
rect 11845 155 11895 160
rect 11845 125 11855 155
rect 11885 125 11895 155
rect 11845 100 11895 125
rect 11845 65 11855 100
rect 11885 65 11895 100
rect 11675 10 11685 40
rect 11715 10 11725 40
rect 11675 0 11725 10
rect 11760 40 11810 50
rect 11760 10 11770 40
rect 11800 10 11810 40
rect 11760 0 11810 10
rect 11845 40 11895 65
rect 12015 155 12065 160
rect 12015 125 12025 155
rect 12055 125 12065 155
rect 12015 100 12065 125
rect 12015 65 12025 100
rect 12055 65 12065 100
rect 11845 10 11855 40
rect 11885 10 11895 40
rect 11845 0 11895 10
rect 11930 40 11980 50
rect 11930 10 11940 40
rect 11970 10 11980 40
rect 11930 0 11980 10
rect 12015 40 12065 65
rect 12185 155 12235 160
rect 12185 125 12195 155
rect 12225 125 12235 155
rect 12185 100 12235 125
rect 12185 65 12195 100
rect 12225 65 12235 100
rect 12015 10 12025 40
rect 12055 10 12065 40
rect 12015 0 12065 10
rect 12100 40 12150 50
rect 12100 10 12110 40
rect 12140 10 12150 40
rect 12100 0 12150 10
rect 12185 40 12235 65
rect 12355 155 12405 160
rect 12355 125 12365 155
rect 12395 125 12405 155
rect 12355 100 12405 125
rect 12355 65 12365 100
rect 12395 65 12405 100
rect 12185 10 12195 40
rect 12225 10 12235 40
rect 12185 0 12235 10
rect 12270 40 12320 50
rect 12270 10 12280 40
rect 12310 10 12320 40
rect 12270 0 12320 10
rect 12355 40 12405 65
rect 12525 155 12575 160
rect 12525 125 12535 155
rect 12565 125 12575 155
rect 12525 100 12575 125
rect 12525 65 12535 100
rect 12565 65 12575 100
rect 12355 10 12365 40
rect 12395 10 12405 40
rect 12355 0 12405 10
rect 12440 40 12490 50
rect 12440 10 12450 40
rect 12480 10 12490 40
rect 12440 0 12490 10
rect 12525 40 12575 65
rect 12695 155 12745 160
rect 12695 125 12705 155
rect 12735 125 12745 155
rect 12695 100 12745 125
rect 12695 65 12705 100
rect 12735 65 12745 100
rect 12525 10 12535 40
rect 12565 10 12575 40
rect 12525 0 12575 10
rect 12610 40 12660 50
rect 12610 10 12620 40
rect 12650 10 12660 40
rect 12610 0 12660 10
rect 12695 40 12745 65
rect 12865 155 12915 160
rect 12865 125 12875 155
rect 12905 125 12915 155
rect 12865 100 12915 125
rect 12865 65 12875 100
rect 12905 65 12915 100
rect 12695 10 12705 40
rect 12735 10 12745 40
rect 12695 0 12745 10
rect 12780 40 12830 50
rect 12780 10 12790 40
rect 12820 10 12830 40
rect 12780 0 12830 10
rect 12865 40 12915 65
rect 13035 155 13085 160
rect 13035 125 13045 155
rect 13075 125 13085 155
rect 13035 100 13085 125
rect 13035 65 13045 100
rect 13075 65 13085 100
rect 12865 10 12875 40
rect 12905 10 12915 40
rect 12865 0 12915 10
rect 12950 40 13000 50
rect 12950 10 12960 40
rect 12990 10 13000 40
rect 12950 0 13000 10
rect 13035 40 13085 65
rect 13205 155 13255 160
rect 13205 125 13215 155
rect 13245 125 13255 155
rect 13205 100 13255 125
rect 13205 65 13215 100
rect 13245 65 13255 100
rect 13035 10 13045 40
rect 13075 10 13085 40
rect 13035 0 13085 10
rect 13120 40 13170 50
rect 13120 10 13130 40
rect 13160 10 13170 40
rect 13120 0 13170 10
rect 13205 40 13255 65
rect 13375 155 13425 160
rect 13375 125 13385 155
rect 13415 125 13425 155
rect 13375 100 13425 125
rect 13375 65 13385 100
rect 13415 65 13425 100
rect 13205 10 13215 40
rect 13245 10 13255 40
rect 13205 0 13255 10
rect 13290 40 13340 50
rect 13290 10 13300 40
rect 13330 10 13340 40
rect 13290 0 13340 10
rect 13375 40 13425 65
rect 13545 155 13595 160
rect 13545 125 13555 155
rect 13585 125 13595 155
rect 13545 100 13595 125
rect 13545 65 13555 100
rect 13585 65 13595 100
rect 13375 10 13385 40
rect 13415 10 13425 40
rect 13375 0 13425 10
rect 13460 40 13510 50
rect 13460 10 13470 40
rect 13500 10 13510 40
rect 13460 0 13510 10
rect 13545 40 13595 65
rect 13715 155 13765 160
rect 13715 125 13725 155
rect 13755 125 13765 155
rect 13715 100 13765 125
rect 13715 65 13725 100
rect 13755 65 13765 100
rect 13545 10 13555 40
rect 13585 10 13595 40
rect 13545 0 13595 10
rect 13630 40 13680 50
rect 13630 10 13640 40
rect 13670 10 13680 40
rect 13630 0 13680 10
rect 13715 40 13765 65
rect 13885 155 13935 160
rect 13885 125 13895 155
rect 13925 125 13935 155
rect 13885 100 13935 125
rect 13885 65 13895 100
rect 13925 65 13935 100
rect 13715 10 13725 40
rect 13755 10 13765 40
rect 13715 0 13765 10
rect 13800 40 13850 50
rect 13800 10 13810 40
rect 13840 10 13850 40
rect 13800 0 13850 10
rect 13885 40 13935 65
rect 14055 155 14105 160
rect 14055 125 14065 155
rect 14095 125 14105 155
rect 14055 100 14105 125
rect 14055 65 14065 100
rect 14095 65 14105 100
rect 13885 10 13895 40
rect 13925 10 13935 40
rect 13885 0 13935 10
rect 13970 40 14020 50
rect 13970 10 13980 40
rect 14010 10 14020 40
rect 13970 0 14020 10
rect 14055 40 14105 65
rect 14225 155 14275 160
rect 14225 125 14235 155
rect 14265 125 14275 155
rect 14225 100 14275 125
rect 14225 65 14235 100
rect 14265 65 14275 100
rect 14055 10 14065 40
rect 14095 10 14105 40
rect 14055 0 14105 10
rect 14140 40 14190 50
rect 14140 10 14150 40
rect 14180 10 14190 40
rect 14140 0 14190 10
rect 14225 40 14275 65
rect 14395 155 14445 160
rect 14395 125 14405 155
rect 14435 125 14445 155
rect 14395 100 14445 125
rect 14395 65 14405 100
rect 14435 65 14445 100
rect 14225 10 14235 40
rect 14265 10 14275 40
rect 14225 0 14275 10
rect 14310 40 14360 50
rect 14310 10 14320 40
rect 14350 10 14360 40
rect 14310 0 14360 10
rect 14395 40 14445 65
rect 14565 155 14615 160
rect 14565 125 14575 155
rect 14605 125 14615 155
rect 14565 100 14615 125
rect 14565 65 14575 100
rect 14605 65 14615 100
rect 14395 10 14405 40
rect 14435 10 14445 40
rect 14395 0 14445 10
rect 14480 40 14530 50
rect 14480 10 14490 40
rect 14520 10 14530 40
rect 14480 0 14530 10
rect 14565 40 14615 65
rect 14735 155 14785 160
rect 14735 125 14745 155
rect 14775 125 14785 155
rect 14735 100 14785 125
rect 14735 65 14745 100
rect 14775 65 14785 100
rect 14565 10 14575 40
rect 14605 10 14615 40
rect 14565 0 14615 10
rect 14650 40 14700 50
rect 14650 10 14660 40
rect 14690 10 14700 40
rect 14650 0 14700 10
rect 14735 40 14785 65
rect 14905 155 14955 160
rect 14905 125 14915 155
rect 14945 125 14955 155
rect 14905 100 14955 125
rect 14905 65 14915 100
rect 14945 65 14955 100
rect 14735 10 14745 40
rect 14775 10 14785 40
rect 14735 0 14785 10
rect 14820 40 14870 50
rect 14820 10 14830 40
rect 14860 10 14870 40
rect 14820 0 14870 10
rect 14905 40 14955 65
rect 15075 155 15125 160
rect 15075 125 15085 155
rect 15115 125 15125 155
rect 15075 100 15125 125
rect 15075 65 15085 100
rect 15115 65 15125 100
rect 14905 10 14915 40
rect 14945 10 14955 40
rect 14905 0 14955 10
rect 14990 40 15040 50
rect 14990 10 15000 40
rect 15030 10 15040 40
rect 14990 0 15040 10
rect 15075 40 15125 65
rect 15245 155 15295 160
rect 15245 125 15255 155
rect 15285 125 15295 155
rect 15245 100 15295 125
rect 15245 65 15255 100
rect 15285 65 15295 100
rect 15075 10 15085 40
rect 15115 10 15125 40
rect 15075 0 15125 10
rect 15160 40 15210 50
rect 15160 10 15170 40
rect 15200 10 15210 40
rect 15160 0 15210 10
rect 15245 40 15295 65
rect 15415 155 15465 160
rect 15415 125 15425 155
rect 15455 125 15465 155
rect 15415 100 15465 125
rect 15415 65 15425 100
rect 15455 65 15465 100
rect 15245 10 15255 40
rect 15285 10 15295 40
rect 15245 0 15295 10
rect 15330 40 15380 50
rect 15330 10 15340 40
rect 15370 10 15380 40
rect 15330 0 15380 10
rect 15415 40 15465 65
rect 15585 155 15635 160
rect 15585 125 15595 155
rect 15625 125 15635 155
rect 15585 100 15635 125
rect 15585 65 15595 100
rect 15625 65 15635 100
rect 15415 10 15425 40
rect 15455 10 15465 40
rect 15415 0 15465 10
rect 15500 40 15550 50
rect 15500 10 15510 40
rect 15540 10 15550 40
rect 15500 0 15550 10
rect 15585 40 15635 65
rect 15755 155 15805 160
rect 15755 125 15765 155
rect 15795 125 15805 155
rect 15755 100 15805 125
rect 15755 65 15765 100
rect 15795 65 15805 100
rect 15585 10 15595 40
rect 15625 10 15635 40
rect 15585 0 15635 10
rect 15670 40 15720 50
rect 15670 10 15680 40
rect 15710 10 15720 40
rect 15670 0 15720 10
rect 15755 40 15805 65
rect 15925 155 15975 160
rect 15925 125 15935 155
rect 15965 125 15975 155
rect 15925 100 15975 125
rect 15925 65 15935 100
rect 15965 65 15975 100
rect 15755 10 15765 40
rect 15795 10 15805 40
rect 15755 0 15805 10
rect 15840 40 15890 50
rect 15840 10 15850 40
rect 15880 10 15890 40
rect 15840 0 15890 10
rect 15925 40 15975 65
rect 16095 155 16145 160
rect 16095 125 16105 155
rect 16135 125 16145 155
rect 16095 100 16145 125
rect 16095 65 16105 100
rect 16135 65 16145 100
rect 15925 10 15935 40
rect 15965 10 15975 40
rect 15925 0 15975 10
rect 16010 40 16060 50
rect 16010 10 16020 40
rect 16050 10 16060 40
rect 16010 0 16060 10
rect 16095 40 16145 65
rect 16265 155 16315 160
rect 16265 125 16275 155
rect 16305 125 16315 155
rect 16265 100 16315 125
rect 16265 65 16275 100
rect 16305 65 16315 100
rect 16095 10 16105 40
rect 16135 10 16145 40
rect 16095 0 16145 10
rect 16180 40 16230 50
rect 16180 10 16190 40
rect 16220 10 16230 40
rect 16180 0 16230 10
rect 16265 40 16315 65
rect 16435 155 16485 160
rect 16435 125 16445 155
rect 16475 125 16485 155
rect 16435 100 16485 125
rect 16435 65 16445 100
rect 16475 65 16485 100
rect 16265 10 16275 40
rect 16305 10 16315 40
rect 16265 0 16315 10
rect 16350 40 16400 50
rect 16350 10 16360 40
rect 16390 10 16400 40
rect 16350 0 16400 10
rect 16435 40 16485 65
rect 16605 155 16655 160
rect 16605 125 16615 155
rect 16645 125 16655 155
rect 16605 100 16655 125
rect 16605 65 16615 100
rect 16645 65 16655 100
rect 16435 10 16445 40
rect 16475 10 16485 40
rect 16435 0 16485 10
rect 16520 40 16570 50
rect 16520 10 16530 40
rect 16560 10 16570 40
rect 16520 0 16570 10
rect 16605 40 16655 65
rect 16775 155 16825 160
rect 16775 125 16785 155
rect 16815 125 16825 155
rect 16775 100 16825 125
rect 16775 65 16785 100
rect 16815 65 16825 100
rect 16605 10 16615 40
rect 16645 10 16655 40
rect 16605 0 16655 10
rect 16690 40 16740 50
rect 16690 10 16700 40
rect 16730 10 16740 40
rect 16690 0 16740 10
rect 16775 40 16825 65
rect 16945 155 16995 160
rect 16945 125 16955 155
rect 16985 125 16995 155
rect 16945 100 16995 125
rect 16945 65 16955 100
rect 16985 65 16995 100
rect 16775 10 16785 40
rect 16815 10 16825 40
rect 16775 0 16825 10
rect 16860 40 16910 50
rect 16860 10 16870 40
rect 16900 10 16910 40
rect 16860 0 16910 10
rect 16945 40 16995 65
rect 17115 155 17165 160
rect 17115 125 17125 155
rect 17155 125 17165 155
rect 17115 100 17165 125
rect 17115 65 17125 100
rect 17155 65 17165 100
rect 16945 10 16955 40
rect 16985 10 16995 40
rect 16945 0 16995 10
rect 17030 40 17080 50
rect 17030 10 17040 40
rect 17070 10 17080 40
rect 17030 0 17080 10
rect 17115 40 17165 65
rect 17285 155 17335 160
rect 17285 125 17295 155
rect 17325 125 17335 155
rect 17285 100 17335 125
rect 17285 65 17295 100
rect 17325 65 17335 100
rect 17115 10 17125 40
rect 17155 10 17165 40
rect 17115 0 17165 10
rect 17200 40 17250 50
rect 17200 10 17210 40
rect 17240 10 17250 40
rect 17200 0 17250 10
rect 17285 40 17335 65
rect 17455 155 17505 160
rect 17455 125 17465 155
rect 17495 125 17505 155
rect 17455 100 17505 125
rect 17455 65 17465 100
rect 17495 65 17505 100
rect 17285 10 17295 40
rect 17325 10 17335 40
rect 17285 0 17335 10
rect 17370 40 17420 50
rect 17370 10 17380 40
rect 17410 10 17420 40
rect 17370 0 17420 10
rect 17455 40 17505 65
rect 17625 155 17675 160
rect 17625 125 17635 155
rect 17665 125 17675 155
rect 17625 100 17675 125
rect 17625 65 17635 100
rect 17665 65 17675 100
rect 17455 10 17465 40
rect 17495 10 17505 40
rect 17455 0 17505 10
rect 17540 40 17590 50
rect 17540 10 17550 40
rect 17580 10 17590 40
rect 17540 0 17590 10
rect 17625 40 17675 65
rect 17795 155 17845 160
rect 17795 125 17805 155
rect 17835 125 17845 155
rect 17795 100 17845 125
rect 17795 65 17805 100
rect 17835 65 17845 100
rect 17625 10 17635 40
rect 17665 10 17675 40
rect 17625 0 17675 10
rect 17710 40 17760 50
rect 17710 10 17720 40
rect 17750 10 17760 40
rect 17710 0 17760 10
rect 17795 40 17845 65
rect 17965 155 18015 160
rect 17965 125 17975 155
rect 18005 125 18015 155
rect 17965 100 18015 125
rect 17965 65 17975 100
rect 18005 65 18015 100
rect 17795 10 17805 40
rect 17835 10 17845 40
rect 17795 0 17845 10
rect 17880 40 17930 50
rect 17880 10 17890 40
rect 17920 10 17930 40
rect 17880 0 17930 10
rect 17965 40 18015 65
rect 18135 155 18185 160
rect 18135 125 18145 155
rect 18175 125 18185 155
rect 18135 100 18185 125
rect 18135 65 18145 100
rect 18175 65 18185 100
rect 17965 10 17975 40
rect 18005 10 18015 40
rect 17965 0 18015 10
rect 18050 40 18100 50
rect 18050 10 18060 40
rect 18090 10 18100 40
rect 18050 0 18100 10
rect 18135 40 18185 65
rect 18305 155 18355 160
rect 18305 125 18315 155
rect 18345 125 18355 155
rect 18305 100 18355 125
rect 18305 65 18315 100
rect 18345 65 18355 100
rect 18135 10 18145 40
rect 18175 10 18185 40
rect 18135 0 18185 10
rect 18220 40 18270 50
rect 18220 10 18230 40
rect 18260 10 18270 40
rect 18220 0 18270 10
rect 18305 40 18355 65
rect 18475 155 18525 160
rect 18475 125 18485 155
rect 18515 125 18525 155
rect 18475 100 18525 125
rect 18475 65 18485 100
rect 18515 65 18525 100
rect 18305 10 18315 40
rect 18345 10 18355 40
rect 18305 0 18355 10
rect 18390 40 18440 50
rect 18390 10 18400 40
rect 18430 10 18440 40
rect 18390 0 18440 10
rect 18475 40 18525 65
rect 18645 155 18695 160
rect 18645 125 18655 155
rect 18685 125 18695 155
rect 18645 100 18695 125
rect 18645 65 18655 100
rect 18685 65 18695 100
rect 18475 10 18485 40
rect 18515 10 18525 40
rect 18475 0 18525 10
rect 18560 40 18610 50
rect 18560 10 18570 40
rect 18600 10 18610 40
rect 18560 0 18610 10
rect 18645 40 18695 65
rect 18815 155 18865 160
rect 18815 125 18825 155
rect 18855 125 18865 155
rect 18815 100 18865 125
rect 18815 65 18825 100
rect 18855 65 18865 100
rect 18645 10 18655 40
rect 18685 10 18695 40
rect 18645 0 18695 10
rect 18730 40 18780 50
rect 18730 10 18740 40
rect 18770 10 18780 40
rect 18730 0 18780 10
rect 18815 40 18865 65
rect 18985 155 19035 160
rect 18985 125 18995 155
rect 19025 125 19035 155
rect 18985 100 19035 125
rect 18985 65 18995 100
rect 19025 65 19035 100
rect 18815 10 18825 40
rect 18855 10 18865 40
rect 18815 0 18865 10
rect 18900 40 18950 50
rect 18900 10 18910 40
rect 18940 10 18950 40
rect 18900 0 18950 10
rect 18985 40 19035 65
rect 19155 155 19205 160
rect 19155 125 19165 155
rect 19195 125 19205 155
rect 19155 100 19205 125
rect 19155 65 19165 100
rect 19195 65 19205 100
rect 18985 10 18995 40
rect 19025 10 19035 40
rect 18985 0 19035 10
rect 19070 40 19120 50
rect 19070 10 19080 40
rect 19110 10 19120 40
rect 19070 0 19120 10
rect 19155 40 19205 65
rect 19325 155 19375 160
rect 19325 125 19335 155
rect 19365 125 19375 155
rect 19325 100 19375 125
rect 19325 65 19335 100
rect 19365 65 19375 100
rect 19155 10 19165 40
rect 19195 10 19205 40
rect 19155 0 19205 10
rect 19240 40 19290 50
rect 19240 10 19250 40
rect 19280 10 19290 40
rect 19240 0 19290 10
rect 19325 40 19375 65
rect 19495 155 19545 160
rect 19495 125 19505 155
rect 19535 125 19545 155
rect 19495 100 19545 125
rect 19495 65 19505 100
rect 19535 65 19545 100
rect 19325 10 19335 40
rect 19365 10 19375 40
rect 19325 0 19375 10
rect 19410 40 19460 50
rect 19410 10 19420 40
rect 19450 10 19460 40
rect 19410 0 19460 10
rect 19495 40 19545 65
rect 19665 155 19715 160
rect 19665 125 19675 155
rect 19705 125 19715 155
rect 19665 100 19715 125
rect 19665 65 19675 100
rect 19705 65 19715 100
rect 19495 10 19505 40
rect 19535 10 19545 40
rect 19495 0 19545 10
rect 19580 40 19630 50
rect 19580 10 19590 40
rect 19620 10 19630 40
rect 19580 0 19630 10
rect 19665 40 19715 65
rect 19835 155 19885 160
rect 19835 125 19845 155
rect 19875 125 19885 155
rect 19835 100 19885 125
rect 19835 65 19845 100
rect 19875 65 19885 100
rect 19665 10 19675 40
rect 19705 10 19715 40
rect 19665 0 19715 10
rect 19750 40 19800 50
rect 19750 10 19760 40
rect 19790 10 19800 40
rect 19750 0 19800 10
rect 19835 40 19885 65
rect 20005 155 20055 160
rect 20005 125 20015 155
rect 20045 125 20055 155
rect 20005 100 20055 125
rect 20005 65 20015 100
rect 20045 65 20055 100
rect 19835 10 19845 40
rect 19875 10 19885 40
rect 19835 0 19885 10
rect 19920 40 19970 50
rect 19920 10 19930 40
rect 19960 10 19970 40
rect 19920 0 19970 10
rect 20005 40 20055 65
rect 20175 155 20225 160
rect 20175 125 20185 155
rect 20215 125 20225 155
rect 20175 100 20225 125
rect 20175 65 20185 100
rect 20215 65 20225 100
rect 20005 10 20015 40
rect 20045 10 20055 40
rect 20005 0 20055 10
rect 20090 40 20140 50
rect 20090 10 20100 40
rect 20130 10 20140 40
rect 20090 0 20140 10
rect 20175 40 20225 65
rect 20345 155 20395 160
rect 20345 125 20355 155
rect 20385 125 20395 155
rect 20345 100 20395 125
rect 20345 65 20355 100
rect 20385 65 20395 100
rect 20175 10 20185 40
rect 20215 10 20225 40
rect 20175 0 20225 10
rect 20260 40 20310 50
rect 20260 10 20270 40
rect 20300 10 20310 40
rect 20260 0 20310 10
rect 20345 40 20395 65
rect 20515 155 20565 160
rect 20515 125 20525 155
rect 20555 125 20565 155
rect 20515 100 20565 125
rect 20515 65 20525 100
rect 20555 65 20565 100
rect 20345 10 20355 40
rect 20385 10 20395 40
rect 20345 0 20395 10
rect 20430 40 20480 50
rect 20430 10 20440 40
rect 20470 10 20480 40
rect 20430 0 20480 10
rect 20515 40 20565 65
rect 20685 155 20735 160
rect 20685 125 20695 155
rect 20725 125 20735 155
rect 20685 100 20735 125
rect 20685 65 20695 100
rect 20725 65 20735 100
rect 20515 10 20525 40
rect 20555 10 20565 40
rect 20515 0 20565 10
rect 20600 40 20650 50
rect 20600 10 20610 40
rect 20640 10 20650 40
rect 20600 0 20650 10
rect 20685 40 20735 65
rect 20855 155 20905 160
rect 20855 125 20865 155
rect 20895 125 20905 155
rect 20855 100 20905 125
rect 20855 65 20865 100
rect 20895 65 20905 100
rect 20685 10 20695 40
rect 20725 10 20735 40
rect 20685 0 20735 10
rect 20770 40 20820 50
rect 20770 10 20780 40
rect 20810 10 20820 40
rect 20770 0 20820 10
rect 20855 40 20905 65
rect 21025 155 21075 160
rect 21025 125 21035 155
rect 21065 125 21075 155
rect 21025 100 21075 125
rect 21025 65 21035 100
rect 21065 65 21075 100
rect 20855 10 20865 40
rect 20895 10 20905 40
rect 20855 0 20905 10
rect 20940 40 20990 50
rect 20940 10 20950 40
rect 20980 10 20990 40
rect 20940 0 20990 10
rect 21025 40 21075 65
rect 21195 155 21245 160
rect 21195 125 21205 155
rect 21235 125 21245 155
rect 21195 100 21245 125
rect 21195 65 21205 100
rect 21235 65 21245 100
rect 21025 10 21035 40
rect 21065 10 21075 40
rect 21025 0 21075 10
rect 21110 40 21160 50
rect 21110 10 21120 40
rect 21150 10 21160 40
rect 21110 0 21160 10
rect 21195 40 21245 65
rect 21365 155 21415 160
rect 21365 125 21375 155
rect 21405 125 21415 155
rect 21365 100 21415 125
rect 21365 65 21375 100
rect 21405 65 21415 100
rect 21195 10 21205 40
rect 21235 10 21245 40
rect 21195 0 21245 10
rect 21280 40 21330 50
rect 21280 10 21290 40
rect 21320 10 21330 40
rect 21280 0 21330 10
rect 21365 40 21415 65
rect 21535 155 21585 160
rect 21535 125 21545 155
rect 21575 125 21585 155
rect 21535 100 21585 125
rect 21535 65 21545 100
rect 21575 65 21585 100
rect 21365 10 21375 40
rect 21405 10 21415 40
rect 21365 0 21415 10
rect 21450 40 21500 50
rect 21450 10 21460 40
rect 21490 10 21500 40
rect 21450 0 21500 10
rect 21535 40 21585 65
rect 21705 155 21755 160
rect 21705 125 21715 155
rect 21745 125 21755 155
rect 21705 100 21755 125
rect 21705 65 21715 100
rect 21745 65 21755 100
rect 21535 10 21545 40
rect 21575 10 21585 40
rect 21535 0 21585 10
rect 21620 40 21670 50
rect 21620 10 21630 40
rect 21660 10 21670 40
rect 21620 0 21670 10
rect 21705 40 21755 65
rect 21875 155 21925 160
rect 21875 125 21885 155
rect 21915 125 21925 155
rect 21875 100 21925 125
rect 21875 65 21885 100
rect 21915 65 21925 100
rect 21705 10 21715 40
rect 21745 10 21755 40
rect 21705 0 21755 10
rect 21790 40 21840 50
rect 21790 10 21800 40
rect 21830 10 21840 40
rect 21790 0 21840 10
rect 21875 40 21925 65
rect 22045 155 22095 160
rect 22045 125 22055 155
rect 22085 125 22095 155
rect 22045 100 22095 125
rect 22045 65 22055 100
rect 22085 65 22095 100
rect 21875 10 21885 40
rect 21915 10 21925 40
rect 21875 0 21925 10
rect 21960 40 22010 50
rect 21960 10 21970 40
rect 22000 10 22010 40
rect 21960 0 22010 10
rect 22045 40 22095 65
rect 22215 155 22265 160
rect 22215 125 22225 155
rect 22255 125 22265 155
rect 22215 100 22265 125
rect 22215 65 22225 100
rect 22255 65 22265 100
rect 22045 10 22055 40
rect 22085 10 22095 40
rect 22045 0 22095 10
rect 22130 40 22180 50
rect 22130 10 22140 40
rect 22170 10 22180 40
rect 22130 0 22180 10
rect 22215 40 22265 65
rect 22385 155 22435 160
rect 22385 125 22395 155
rect 22425 125 22435 155
rect 22385 100 22435 125
rect 22385 65 22395 100
rect 22425 65 22435 100
rect 22215 10 22225 40
rect 22255 10 22265 40
rect 22215 0 22265 10
rect 22300 40 22350 50
rect 22300 10 22310 40
rect 22340 10 22350 40
rect 22300 0 22350 10
rect 22385 40 22435 65
rect 22555 155 22605 160
rect 22555 125 22565 155
rect 22595 125 22605 155
rect 22555 100 22605 125
rect 22555 65 22565 100
rect 22595 65 22605 100
rect 22385 10 22395 40
rect 22425 10 22435 40
rect 22385 0 22435 10
rect 22470 40 22520 50
rect 22470 10 22480 40
rect 22510 10 22520 40
rect 22470 0 22520 10
rect 22555 40 22605 65
rect 22725 155 22775 160
rect 22725 125 22735 155
rect 22765 125 22775 155
rect 22725 100 22775 125
rect 22725 65 22735 100
rect 22765 65 22775 100
rect 22555 10 22565 40
rect 22595 10 22605 40
rect 22555 0 22605 10
rect 22640 40 22690 50
rect 22640 10 22650 40
rect 22680 10 22690 40
rect 22640 0 22690 10
rect 22725 40 22775 65
rect 22895 155 22945 160
rect 22895 125 22905 155
rect 22935 125 22945 155
rect 22895 100 22945 125
rect 22895 65 22905 100
rect 22935 65 22945 100
rect 22725 10 22735 40
rect 22765 10 22775 40
rect 22725 0 22775 10
rect 22810 40 22860 50
rect 22810 10 22820 40
rect 22850 10 22860 40
rect 22810 0 22860 10
rect 22895 40 22945 65
rect 23065 155 23115 160
rect 23065 125 23075 155
rect 23105 125 23115 155
rect 23065 100 23115 125
rect 23065 65 23075 100
rect 23105 65 23115 100
rect 22895 10 22905 40
rect 22935 10 22945 40
rect 22895 0 22945 10
rect 22980 40 23030 50
rect 22980 10 22990 40
rect 23020 10 23030 40
rect 22980 0 23030 10
rect 23065 40 23115 65
rect 23235 155 23285 160
rect 23235 125 23245 155
rect 23275 125 23285 155
rect 23235 100 23285 125
rect 23235 65 23245 100
rect 23275 65 23285 100
rect 23065 10 23075 40
rect 23105 10 23115 40
rect 23065 0 23115 10
rect 23150 40 23200 50
rect 23150 10 23160 40
rect 23190 10 23200 40
rect 23150 0 23200 10
rect 23235 40 23285 65
rect 23405 155 23455 160
rect 23405 125 23415 155
rect 23445 125 23455 155
rect 23405 100 23455 125
rect 23405 65 23415 100
rect 23445 65 23455 100
rect 23235 10 23245 40
rect 23275 10 23285 40
rect 23235 0 23285 10
rect 23320 40 23370 50
rect 23320 10 23330 40
rect 23360 10 23370 40
rect 23320 0 23370 10
rect 23405 40 23455 65
rect 23575 155 23625 160
rect 23575 125 23585 155
rect 23615 125 23625 155
rect 23575 100 23625 125
rect 23575 65 23585 100
rect 23615 65 23625 100
rect 23405 10 23415 40
rect 23445 10 23455 40
rect 23405 0 23455 10
rect 23490 40 23540 50
rect 23490 10 23500 40
rect 23530 10 23540 40
rect 23490 0 23540 10
rect 23575 40 23625 65
rect 23745 155 23795 160
rect 23745 125 23755 155
rect 23785 125 23795 155
rect 23745 100 23795 125
rect 23745 65 23755 100
rect 23785 65 23795 100
rect 23575 10 23585 40
rect 23615 10 23625 40
rect 23575 0 23625 10
rect 23660 40 23710 50
rect 23660 10 23670 40
rect 23700 10 23710 40
rect 23660 0 23710 10
rect 23745 40 23795 65
rect 23915 155 23965 160
rect 23915 125 23925 155
rect 23955 125 23965 155
rect 23915 100 23965 125
rect 23915 65 23925 100
rect 23955 65 23965 100
rect 23745 10 23755 40
rect 23785 10 23795 40
rect 23745 0 23795 10
rect 23830 40 23880 50
rect 23830 10 23840 40
rect 23870 10 23880 40
rect 23830 0 23880 10
rect 23915 40 23965 65
rect 24085 155 24135 160
rect 24085 125 24095 155
rect 24125 125 24135 155
rect 24085 100 24135 125
rect 24085 65 24095 100
rect 24125 65 24135 100
rect 23915 10 23925 40
rect 23955 10 23965 40
rect 23915 0 23965 10
rect 24000 40 24050 50
rect 24000 10 24010 40
rect 24040 10 24050 40
rect 24000 0 24050 10
rect 24085 40 24135 65
rect 24255 155 24305 160
rect 24255 125 24265 155
rect 24295 125 24305 155
rect 24255 100 24305 125
rect 24255 65 24265 100
rect 24295 65 24305 100
rect 24085 10 24095 40
rect 24125 10 24135 40
rect 24085 0 24135 10
rect 24170 40 24220 50
rect 24170 10 24180 40
rect 24210 10 24220 40
rect 24170 0 24220 10
rect 24255 40 24305 65
rect 24425 155 24475 160
rect 24425 125 24435 155
rect 24465 125 24475 155
rect 24425 100 24475 125
rect 24425 65 24435 100
rect 24465 65 24475 100
rect 24255 10 24265 40
rect 24295 10 24305 40
rect 24255 0 24305 10
rect 24340 40 24390 50
rect 24340 10 24350 40
rect 24380 10 24390 40
rect 24340 0 24390 10
rect 24425 40 24475 65
rect 24595 155 24645 160
rect 24595 125 24605 155
rect 24635 125 24645 155
rect 24595 100 24645 125
rect 24595 65 24605 100
rect 24635 65 24645 100
rect 24425 10 24435 40
rect 24465 10 24475 40
rect 24425 0 24475 10
rect 24510 40 24560 50
rect 24510 10 24520 40
rect 24550 10 24560 40
rect 24510 0 24560 10
rect 24595 40 24645 65
rect 24765 155 24815 160
rect 24765 125 24775 155
rect 24805 125 24815 155
rect 24765 100 24815 125
rect 24765 65 24775 100
rect 24805 65 24815 100
rect 24595 10 24605 40
rect 24635 10 24645 40
rect 24595 0 24645 10
rect 24680 40 24730 50
rect 24680 10 24690 40
rect 24720 10 24730 40
rect 24680 0 24730 10
rect 24765 40 24815 65
rect 24935 155 24985 160
rect 24935 125 24945 155
rect 24975 125 24985 155
rect 24935 100 24985 125
rect 24935 65 24945 100
rect 24975 65 24985 100
rect 24765 10 24775 40
rect 24805 10 24815 40
rect 24765 0 24815 10
rect 24850 40 24900 50
rect 24850 10 24860 40
rect 24890 10 24900 40
rect 24850 0 24900 10
rect 24935 40 24985 65
rect 25105 155 25155 160
rect 25105 125 25115 155
rect 25145 125 25155 155
rect 25105 100 25155 125
rect 25105 65 25115 100
rect 25145 65 25155 100
rect 24935 10 24945 40
rect 24975 10 24985 40
rect 24935 0 24985 10
rect 25020 40 25070 50
rect 25020 10 25030 40
rect 25060 10 25070 40
rect 25020 0 25070 10
rect 25105 40 25155 65
rect 25275 155 25325 160
rect 25275 125 25285 155
rect 25315 125 25325 155
rect 25275 100 25325 125
rect 25275 65 25285 100
rect 25315 65 25325 100
rect 25105 10 25115 40
rect 25145 10 25155 40
rect 25105 0 25155 10
rect 25190 40 25240 50
rect 25190 10 25200 40
rect 25230 10 25240 40
rect 25190 0 25240 10
rect 25275 40 25325 65
rect 25445 155 25495 160
rect 25445 125 25455 155
rect 25485 125 25495 155
rect 25445 100 25495 125
rect 25445 65 25455 100
rect 25485 65 25495 100
rect 25275 10 25285 40
rect 25315 10 25325 40
rect 25275 0 25325 10
rect 25360 40 25410 50
rect 25360 10 25370 40
rect 25400 10 25410 40
rect 25360 0 25410 10
rect 25445 40 25495 65
rect 25615 155 25665 160
rect 25615 125 25625 155
rect 25655 125 25665 155
rect 25615 100 25665 125
rect 25615 65 25625 100
rect 25655 65 25665 100
rect 25445 10 25455 40
rect 25485 10 25495 40
rect 25445 0 25495 10
rect 25530 40 25580 50
rect 25530 10 25540 40
rect 25570 10 25580 40
rect 25530 0 25580 10
rect 25615 40 25665 65
rect 25785 155 25835 160
rect 25785 125 25795 155
rect 25825 125 25835 155
rect 25785 100 25835 125
rect 25785 65 25795 100
rect 25825 65 25835 100
rect 25615 10 25625 40
rect 25655 10 25665 40
rect 25615 0 25665 10
rect 25700 40 25750 50
rect 25700 10 25710 40
rect 25740 10 25750 40
rect 25700 0 25750 10
rect 25785 40 25835 65
rect 25955 155 26005 160
rect 25955 125 25965 155
rect 25995 125 26005 155
rect 25955 100 26005 125
rect 25955 65 25965 100
rect 25995 65 26005 100
rect 25785 10 25795 40
rect 25825 10 25835 40
rect 25785 0 25835 10
rect 25870 40 25920 50
rect 25870 10 25880 40
rect 25910 10 25920 40
rect 25870 0 25920 10
rect 25955 40 26005 65
rect 26125 155 26175 160
rect 26125 125 26135 155
rect 26165 125 26175 155
rect 26125 100 26175 125
rect 26125 65 26135 100
rect 26165 65 26175 100
rect 25955 10 25965 40
rect 25995 10 26005 40
rect 25955 0 26005 10
rect 26040 40 26090 50
rect 26040 10 26050 40
rect 26080 10 26090 40
rect 26040 0 26090 10
rect 26125 40 26175 65
rect 26295 155 26345 160
rect 26295 125 26305 155
rect 26335 125 26345 155
rect 26295 100 26345 125
rect 26295 65 26305 100
rect 26335 65 26345 100
rect 26125 10 26135 40
rect 26165 10 26175 40
rect 26125 0 26175 10
rect 26210 40 26260 50
rect 26210 10 26220 40
rect 26250 10 26260 40
rect 26210 0 26260 10
rect 26295 40 26345 65
rect 26465 155 26515 160
rect 26465 125 26475 155
rect 26505 125 26515 155
rect 26465 100 26515 125
rect 26465 65 26475 100
rect 26505 65 26515 100
rect 26295 10 26305 40
rect 26335 10 26345 40
rect 26295 0 26345 10
rect 26380 40 26430 50
rect 26380 10 26390 40
rect 26420 10 26430 40
rect 26380 0 26430 10
rect 26465 40 26515 65
rect 26635 155 26685 160
rect 26635 125 26645 155
rect 26675 125 26685 155
rect 26635 100 26685 125
rect 26635 65 26645 100
rect 26675 65 26685 100
rect 26465 10 26475 40
rect 26505 10 26515 40
rect 26465 0 26515 10
rect 26550 40 26600 50
rect 26550 10 26560 40
rect 26590 10 26600 40
rect 26550 0 26600 10
rect 26635 40 26685 65
rect 26805 155 26855 160
rect 26805 125 26815 155
rect 26845 125 26855 155
rect 26805 100 26855 125
rect 26805 65 26815 100
rect 26845 65 26855 100
rect 26635 10 26645 40
rect 26675 10 26685 40
rect 26635 0 26685 10
rect 26720 40 26770 50
rect 26720 10 26730 40
rect 26760 10 26770 40
rect 26720 0 26770 10
rect 26805 40 26855 65
rect 26975 155 27025 160
rect 26975 125 26985 155
rect 27015 125 27025 155
rect 26975 100 27025 125
rect 26975 65 26985 100
rect 27015 65 27025 100
rect 26805 10 26815 40
rect 26845 10 26855 40
rect 26805 0 26855 10
rect 26890 40 26940 50
rect 26890 10 26900 40
rect 26930 10 26940 40
rect 26890 0 26940 10
rect 26975 40 27025 65
rect 27145 155 27195 160
rect 27145 125 27155 155
rect 27185 125 27195 155
rect 27145 100 27195 125
rect 27145 65 27155 100
rect 27185 65 27195 100
rect 26975 10 26985 40
rect 27015 10 27025 40
rect 26975 0 27025 10
rect 27060 40 27110 50
rect 27060 10 27070 40
rect 27100 10 27110 40
rect 27060 0 27110 10
rect 27145 40 27195 65
rect 27315 155 27365 160
rect 27315 125 27325 155
rect 27355 125 27365 155
rect 27315 100 27365 125
rect 27315 65 27325 100
rect 27355 65 27365 100
rect 27145 10 27155 40
rect 27185 10 27195 40
rect 27145 0 27195 10
rect 27230 40 27280 50
rect 27230 10 27240 40
rect 27270 10 27280 40
rect 27230 0 27280 10
rect 27315 40 27365 65
rect 27485 155 27535 160
rect 27485 125 27495 155
rect 27525 125 27535 155
rect 27485 100 27535 125
rect 27485 65 27495 100
rect 27525 65 27535 100
rect 27315 10 27325 40
rect 27355 10 27365 40
rect 27315 0 27365 10
rect 27400 40 27450 50
rect 27400 10 27410 40
rect 27440 10 27450 40
rect 27400 0 27450 10
rect 27485 40 27535 65
rect 27655 155 27705 160
rect 27655 125 27665 155
rect 27695 125 27705 155
rect 27655 100 27705 125
rect 27655 65 27665 100
rect 27695 65 27705 100
rect 27485 10 27495 40
rect 27525 10 27535 40
rect 27485 0 27535 10
rect 27570 40 27620 50
rect 27570 10 27580 40
rect 27610 10 27620 40
rect 27570 0 27620 10
rect 27655 40 27705 65
rect 27825 155 27875 160
rect 27825 125 27835 155
rect 27865 125 27875 155
rect 27825 100 27875 125
rect 27825 65 27835 100
rect 27865 65 27875 100
rect 27655 10 27665 40
rect 27695 10 27705 40
rect 27655 0 27705 10
rect 27740 40 27790 50
rect 27740 10 27750 40
rect 27780 10 27790 40
rect 27740 0 27790 10
rect 27825 40 27875 65
rect 27995 155 28045 160
rect 27995 125 28005 155
rect 28035 125 28045 155
rect 27995 100 28045 125
rect 27995 65 28005 100
rect 28035 65 28045 100
rect 27825 10 27835 40
rect 27865 10 27875 40
rect 27825 0 27875 10
rect 27910 40 27960 50
rect 27910 10 27920 40
rect 27950 10 27960 40
rect 27910 0 27960 10
rect 27995 40 28045 65
rect 28165 155 28215 160
rect 28165 125 28175 155
rect 28205 125 28215 155
rect 28165 100 28215 125
rect 28165 65 28175 100
rect 28205 65 28215 100
rect 27995 10 28005 40
rect 28035 10 28045 40
rect 27995 0 28045 10
rect 28080 40 28130 50
rect 28080 10 28090 40
rect 28120 10 28130 40
rect 28080 0 28130 10
rect 28165 40 28215 65
rect 28335 155 28385 160
rect 28335 125 28345 155
rect 28375 125 28385 155
rect 28335 100 28385 125
rect 28335 65 28345 100
rect 28375 65 28385 100
rect 28165 10 28175 40
rect 28205 10 28215 40
rect 28165 0 28215 10
rect 28250 40 28300 50
rect 28250 10 28260 40
rect 28290 10 28300 40
rect 28250 0 28300 10
rect 28335 40 28385 65
rect 28505 155 28555 160
rect 28505 125 28515 155
rect 28545 125 28555 155
rect 28505 100 28555 125
rect 28505 65 28515 100
rect 28545 65 28555 100
rect 28335 10 28345 40
rect 28375 10 28385 40
rect 28335 0 28385 10
rect 28420 40 28470 50
rect 28420 10 28430 40
rect 28460 10 28470 40
rect 28420 0 28470 10
rect 28505 40 28555 65
rect 28675 155 28725 160
rect 28675 125 28685 155
rect 28715 125 28725 155
rect 28675 100 28725 125
rect 28675 65 28685 100
rect 28715 65 28725 100
rect 28505 10 28515 40
rect 28545 10 28555 40
rect 28505 0 28555 10
rect 28590 40 28640 50
rect 28590 10 28600 40
rect 28630 10 28640 40
rect 28590 0 28640 10
rect 28675 40 28725 65
rect 28845 155 28895 160
rect 28845 125 28855 155
rect 28885 125 28895 155
rect 28845 100 28895 125
rect 28845 65 28855 100
rect 28885 65 28895 100
rect 28675 10 28685 40
rect 28715 10 28725 40
rect 28675 0 28725 10
rect 28760 40 28810 50
rect 28760 10 28770 40
rect 28800 10 28810 40
rect 28760 0 28810 10
rect 28845 40 28895 65
rect 29015 155 29065 160
rect 29015 125 29025 155
rect 29055 125 29065 155
rect 29015 100 29065 125
rect 29015 65 29025 100
rect 29055 65 29065 100
rect 28845 10 28855 40
rect 28885 10 28895 40
rect 28845 0 28895 10
rect 28930 40 28980 50
rect 28930 10 28940 40
rect 28970 10 28980 40
rect 28930 0 28980 10
rect 29015 40 29065 65
rect 29185 155 29235 160
rect 29185 125 29195 155
rect 29225 125 29235 155
rect 29185 100 29235 125
rect 29185 65 29195 100
rect 29225 65 29235 100
rect 29015 10 29025 40
rect 29055 10 29065 40
rect 29015 0 29065 10
rect 29100 40 29150 50
rect 29100 10 29110 40
rect 29140 10 29150 40
rect 29100 0 29150 10
rect 29185 40 29235 65
rect 29355 155 29405 160
rect 29355 125 29365 155
rect 29395 125 29405 155
rect 29355 100 29405 125
rect 29355 65 29365 100
rect 29395 65 29405 100
rect 29185 10 29195 40
rect 29225 10 29235 40
rect 29185 0 29235 10
rect 29270 40 29320 50
rect 29270 10 29280 40
rect 29310 10 29320 40
rect 29270 0 29320 10
rect 29355 40 29405 65
rect 29525 155 29575 160
rect 29525 125 29535 155
rect 29565 125 29575 155
rect 29525 100 29575 125
rect 29525 65 29535 100
rect 29565 65 29575 100
rect 29355 10 29365 40
rect 29395 10 29405 40
rect 29355 0 29405 10
rect 29440 40 29490 50
rect 29440 10 29450 40
rect 29480 10 29490 40
rect 29440 0 29490 10
rect 29525 40 29575 65
rect 29525 10 29535 40
rect 29565 10 29575 40
rect 29525 0 29575 10
rect 29610 40 29660 50
rect 29610 10 29620 40
rect 29650 10 29660 40
rect 29610 0 29660 10
rect 90 -60 100 -30
rect 130 -60 140 -30
rect 90 -90 140 -60
rect 255 -30 310 -20
rect 255 -60 265 -30
rect 300 -60 310 -30
rect 255 -70 310 -60
rect 340 -30 395 -20
rect 340 -60 350 -30
rect 385 -60 395 -30
rect 340 -70 395 -60
rect 425 -30 480 -20
rect 425 -60 435 -30
rect 470 -60 480 -30
rect 425 -70 480 -60
rect 510 -30 565 -20
rect 510 -60 520 -30
rect 555 -60 565 -30
rect 510 -70 565 -60
rect 790 -30 845 -20
rect 790 -60 800 -30
rect 835 -60 845 -30
rect 790 -70 845 -60
rect 875 -30 930 -20
rect 875 -60 885 -30
rect 920 -60 930 -30
rect 875 -70 930 -60
rect 960 -30 1015 -20
rect 960 -60 970 -30
rect 1005 -60 1015 -30
rect 960 -70 1015 -60
rect 1045 -30 1100 -20
rect 1045 -60 1055 -30
rect 1090 -60 1100 -30
rect 1045 -70 1100 -60
rect 1130 -30 1185 -20
rect 1130 -60 1140 -30
rect 1175 -60 1185 -30
rect 1130 -70 1185 -60
rect 1215 -30 1270 -20
rect 1215 -60 1225 -30
rect 1260 -60 1270 -30
rect 1215 -70 1270 -60
rect 1300 -30 1355 -20
rect 1300 -60 1310 -30
rect 1345 -60 1355 -30
rect 1300 -70 1355 -60
rect 1385 -30 1440 -20
rect 1385 -60 1395 -30
rect 1430 -60 1440 -30
rect 1385 -70 1440 -60
rect 1470 -30 1525 -20
rect 1470 -60 1480 -30
rect 1515 -60 1525 -30
rect 1470 -70 1525 -60
rect 1555 -30 1610 -20
rect 1555 -60 1565 -30
rect 1600 -60 1610 -30
rect 1555 -70 1610 -60
rect 1640 -30 1695 -20
rect 1640 -60 1650 -30
rect 1685 -60 1695 -30
rect 1640 -70 1695 -60
rect 1725 -30 1780 -20
rect 1725 -60 1735 -30
rect 1770 -60 1780 -30
rect 1725 -70 1780 -60
rect 1810 -30 1865 -20
rect 1810 -60 1820 -30
rect 1855 -60 1865 -30
rect 1810 -70 1865 -60
rect 1895 -30 1950 -20
rect 1895 -60 1905 -30
rect 1940 -60 1950 -30
rect 1895 -70 1950 -60
rect 1980 -30 2035 -20
rect 1980 -60 1990 -30
rect 2025 -60 2035 -30
rect 1980 -70 2035 -60
rect 2065 -30 2120 -20
rect 2065 -60 2075 -30
rect 2110 -60 2120 -30
rect 2065 -70 2120 -60
rect 2300 -30 2355 -20
rect 2300 -60 2310 -30
rect 2345 -60 2355 -30
rect 2300 -70 2355 -60
rect 2385 -30 2440 -20
rect 2385 -60 2395 -30
rect 2430 -60 2440 -30
rect 2385 -70 2440 -60
rect 2470 -30 2525 -20
rect 2470 -60 2480 -30
rect 2515 -60 2525 -30
rect 2470 -70 2525 -60
rect 2555 -30 2610 -20
rect 2555 -60 2565 -30
rect 2600 -60 2610 -30
rect 2555 -70 2610 -60
rect 2640 -30 2695 -20
rect 2640 -60 2650 -30
rect 2685 -60 2695 -30
rect 2640 -70 2695 -60
rect 2725 -30 2780 -20
rect 2725 -60 2735 -30
rect 2770 -60 2780 -30
rect 2725 -70 2780 -60
rect 2810 -30 2865 -20
rect 2810 -60 2820 -30
rect 2855 -60 2865 -30
rect 2810 -70 2865 -60
rect 2895 -30 2950 -20
rect 2895 -60 2905 -30
rect 2940 -60 2950 -30
rect 2895 -70 2950 -60
rect 2980 -30 3035 -20
rect 2980 -60 2990 -30
rect 3025 -60 3035 -30
rect 2980 -70 3035 -60
rect 3065 -30 3120 -20
rect 3065 -60 3075 -30
rect 3110 -60 3120 -30
rect 3065 -70 3120 -60
rect 3150 -30 3205 -20
rect 3150 -60 3160 -30
rect 3195 -60 3205 -30
rect 3150 -70 3205 -60
rect 3235 -30 3290 -20
rect 3235 -60 3245 -30
rect 3280 -60 3290 -30
rect 3235 -70 3290 -60
rect 3320 -30 3375 -20
rect 3320 -60 3330 -30
rect 3365 -60 3375 -30
rect 3320 -70 3375 -60
rect 3405 -30 3460 -20
rect 3405 -60 3415 -30
rect 3450 -60 3460 -30
rect 3405 -70 3460 -60
rect 3490 -30 3545 -20
rect 3490 -60 3500 -30
rect 3535 -60 3545 -30
rect 3490 -70 3545 -60
rect 3575 -30 3630 -20
rect 3575 -60 3585 -30
rect 3620 -60 3630 -30
rect 3575 -70 3630 -60
rect 3660 -30 3715 -20
rect 3660 -60 3670 -30
rect 3705 -60 3715 -30
rect 3660 -70 3715 -60
rect 3745 -30 3800 -20
rect 3745 -60 3755 -30
rect 3790 -60 3800 -30
rect 3745 -70 3800 -60
rect 3830 -30 3885 -20
rect 3830 -60 3840 -30
rect 3875 -60 3885 -30
rect 3830 -70 3885 -60
rect 3915 -30 3970 -20
rect 3915 -60 3925 -30
rect 3960 -60 3970 -30
rect 3915 -70 3970 -60
rect 4000 -30 4055 -20
rect 4000 -60 4010 -30
rect 4045 -60 4055 -30
rect 4000 -70 4055 -60
rect 4085 -30 4140 -20
rect 4085 -60 4095 -30
rect 4130 -60 4140 -30
rect 4085 -70 4140 -60
rect 4170 -30 4225 -20
rect 4170 -60 4180 -30
rect 4215 -60 4225 -30
rect 4170 -70 4225 -60
rect 4255 -30 4310 -20
rect 4255 -60 4265 -30
rect 4300 -60 4310 -30
rect 4255 -70 4310 -60
rect 4340 -30 4395 -20
rect 4340 -60 4350 -30
rect 4385 -60 4395 -30
rect 4340 -70 4395 -60
rect 4425 -30 4480 -20
rect 4425 -60 4435 -30
rect 4470 -60 4480 -30
rect 4425 -70 4480 -60
rect 4510 -30 4565 -20
rect 4510 -60 4520 -30
rect 4555 -60 4565 -30
rect 4510 -70 4565 -60
rect 4595 -30 4650 -20
rect 4595 -60 4605 -30
rect 4640 -60 4650 -30
rect 4595 -70 4650 -60
rect 4680 -30 4735 -20
rect 4680 -60 4690 -30
rect 4725 -60 4735 -30
rect 4680 -70 4735 -60
rect 4765 -30 4820 -20
rect 4765 -60 4775 -30
rect 4810 -60 4820 -30
rect 4765 -70 4820 -60
rect 4850 -30 4905 -20
rect 4850 -60 4860 -30
rect 4895 -60 4905 -30
rect 4850 -70 4905 -60
rect 4935 -30 4990 -20
rect 4935 -60 4945 -30
rect 4980 -60 4990 -30
rect 4935 -70 4990 -60
rect 5020 -30 5075 -20
rect 5020 -60 5030 -30
rect 5065 -60 5075 -30
rect 5020 -70 5075 -60
rect 5105 -30 5160 -20
rect 5105 -60 5115 -30
rect 5150 -60 5160 -30
rect 5105 -70 5160 -60
rect 5190 -30 5245 -20
rect 5190 -60 5200 -30
rect 5235 -60 5245 -30
rect 5190 -70 5245 -60
rect 5275 -30 5330 -20
rect 5275 -60 5285 -30
rect 5320 -60 5330 -30
rect 5275 -70 5330 -60
rect 5360 -30 5415 -20
rect 5360 -60 5370 -30
rect 5405 -60 5415 -30
rect 5360 -70 5415 -60
rect 5445 -30 5500 -20
rect 5445 -60 5455 -30
rect 5490 -60 5500 -30
rect 5445 -70 5500 -60
rect 5530 -30 5585 -20
rect 5530 -60 5540 -30
rect 5575 -60 5585 -30
rect 5530 -70 5585 -60
rect 5615 -30 5670 -20
rect 5615 -60 5625 -30
rect 5660 -60 5670 -30
rect 5615 -70 5670 -60
rect 5700 -30 5755 -20
rect 5700 -60 5710 -30
rect 5745 -60 5755 -30
rect 5700 -70 5755 -60
rect 5785 -30 5840 -20
rect 5785 -60 5795 -30
rect 5830 -60 5840 -30
rect 5785 -70 5840 -60
rect 5870 -30 5925 -20
rect 5870 -60 5880 -30
rect 5915 -60 5925 -30
rect 5870 -70 5925 -60
rect 5955 -30 6010 -20
rect 5955 -60 5965 -30
rect 6000 -60 6010 -30
rect 5955 -70 6010 -60
rect 6040 -30 6095 -20
rect 6040 -60 6050 -30
rect 6085 -60 6095 -30
rect 6040 -70 6095 -60
rect 6125 -30 6180 -20
rect 6125 -60 6135 -30
rect 6170 -60 6180 -30
rect 6125 -70 6180 -60
rect 6210 -30 6265 -20
rect 6210 -60 6220 -30
rect 6255 -60 6265 -30
rect 6210 -70 6265 -60
rect 6295 -30 6350 -20
rect 6295 -60 6305 -30
rect 6340 -60 6350 -30
rect 6295 -70 6350 -60
rect 6380 -30 6435 -20
rect 6380 -60 6390 -30
rect 6425 -60 6435 -30
rect 6380 -70 6435 -60
rect 6465 -30 6520 -20
rect 6465 -60 6475 -30
rect 6510 -60 6520 -30
rect 6465 -70 6520 -60
rect 6550 -30 6605 -20
rect 6550 -60 6560 -30
rect 6595 -60 6605 -30
rect 6550 -70 6605 -60
rect 6635 -30 6690 -20
rect 6635 -60 6645 -30
rect 6680 -60 6690 -30
rect 6635 -70 6690 -60
rect 6720 -30 6775 -20
rect 6720 -60 6730 -30
rect 6765 -60 6775 -30
rect 6720 -70 6775 -60
rect 6805 -30 6860 -20
rect 6805 -60 6815 -30
rect 6850 -60 6860 -30
rect 6805 -70 6860 -60
rect 6890 -30 6945 -20
rect 6890 -60 6900 -30
rect 6935 -60 6945 -30
rect 6890 -70 6945 -60
rect 6975 -30 7030 -20
rect 6975 -60 6985 -30
rect 7020 -60 7030 -30
rect 6975 -70 7030 -60
rect 7060 -30 7115 -20
rect 7060 -60 7070 -30
rect 7105 -60 7115 -30
rect 7060 -70 7115 -60
rect 7145 -30 7200 -20
rect 7145 -60 7155 -30
rect 7190 -60 7200 -30
rect 7145 -70 7200 -60
rect 7230 -30 7285 -20
rect 7230 -60 7240 -30
rect 7275 -60 7285 -30
rect 7230 -70 7285 -60
rect 7315 -30 7370 -20
rect 7315 -60 7325 -30
rect 7360 -60 7370 -30
rect 7315 -70 7370 -60
rect 7400 -30 7455 -20
rect 7400 -60 7410 -30
rect 7445 -60 7455 -30
rect 7400 -70 7455 -60
rect 7485 -30 7540 -20
rect 7485 -60 7495 -30
rect 7530 -60 7540 -30
rect 7485 -70 7540 -60
rect 7570 -30 7625 -20
rect 7570 -60 7580 -30
rect 7615 -60 7625 -30
rect 7570 -70 7625 -60
rect 7655 -30 7710 -20
rect 7655 -60 7665 -30
rect 7700 -60 7710 -30
rect 7655 -70 7710 -60
rect 7890 -30 7945 -20
rect 7890 -60 7900 -30
rect 7935 -60 7945 -30
rect 7890 -70 7945 -60
rect 7975 -30 8030 -20
rect 7975 -60 7985 -30
rect 8020 -60 8030 -30
rect 7975 -70 8030 -60
rect 8060 -30 8115 -20
rect 8060 -60 8070 -30
rect 8105 -60 8115 -30
rect 8060 -70 8115 -60
rect 8145 -30 8200 -20
rect 8145 -60 8155 -30
rect 8190 -60 8200 -30
rect 8145 -70 8200 -60
rect 8230 -30 8285 -20
rect 8230 -60 8240 -30
rect 8275 -60 8285 -30
rect 8230 -70 8285 -60
rect 8315 -30 8370 -20
rect 8315 -60 8325 -30
rect 8360 -60 8370 -30
rect 8315 -70 8370 -60
rect 8400 -30 8455 -20
rect 8400 -60 8410 -30
rect 8445 -60 8455 -30
rect 8400 -70 8455 -60
rect 8485 -30 8540 -20
rect 8485 -60 8495 -30
rect 8530 -60 8540 -30
rect 8485 -70 8540 -60
rect 8570 -30 8625 -20
rect 8570 -60 8580 -30
rect 8615 -60 8625 -30
rect 8570 -70 8625 -60
rect 8655 -30 8710 -20
rect 8655 -60 8665 -30
rect 8700 -60 8710 -30
rect 8655 -70 8710 -60
rect 8740 -30 8795 -20
rect 8740 -60 8750 -30
rect 8785 -60 8795 -30
rect 8740 -70 8795 -60
rect 8825 -30 8880 -20
rect 8825 -60 8835 -30
rect 8870 -60 8880 -30
rect 8825 -70 8880 -60
rect 8910 -30 8965 -20
rect 8910 -60 8920 -30
rect 8955 -60 8965 -30
rect 8910 -70 8965 -60
rect 8995 -30 9050 -20
rect 8995 -60 9005 -30
rect 9040 -60 9050 -30
rect 8995 -70 9050 -60
rect 9080 -30 9135 -20
rect 9080 -60 9090 -30
rect 9125 -60 9135 -30
rect 9080 -70 9135 -60
rect 9165 -30 9220 -20
rect 9165 -60 9175 -30
rect 9210 -60 9220 -30
rect 9165 -70 9220 -60
rect 9250 -30 9305 -20
rect 9250 -60 9260 -30
rect 9295 -60 9305 -30
rect 9250 -70 9305 -60
rect 9335 -30 9390 -20
rect 9335 -60 9345 -30
rect 9380 -60 9390 -30
rect 9335 -70 9390 -60
rect 9420 -30 9475 -20
rect 9420 -60 9430 -30
rect 9465 -60 9475 -30
rect 9420 -70 9475 -60
rect 9505 -30 9560 -20
rect 9505 -60 9515 -30
rect 9550 -60 9560 -30
rect 9505 -70 9560 -60
rect 9590 -30 9645 -20
rect 9590 -60 9600 -30
rect 9635 -60 9645 -30
rect 9590 -70 9645 -60
rect 9675 -30 9730 -20
rect 9675 -60 9685 -30
rect 9720 -60 9730 -30
rect 9675 -70 9730 -60
rect 9760 -30 9815 -20
rect 9760 -60 9770 -30
rect 9805 -60 9815 -30
rect 9760 -70 9815 -60
rect 9845 -30 9900 -20
rect 9845 -60 9855 -30
rect 9890 -60 9900 -30
rect 9845 -70 9900 -60
rect 9930 -30 9985 -20
rect 9930 -60 9940 -30
rect 9975 -60 9985 -30
rect 9930 -70 9985 -60
rect 10015 -30 10070 -20
rect 10015 -60 10025 -30
rect 10060 -60 10070 -30
rect 10015 -70 10070 -60
rect 10100 -30 10155 -20
rect 10100 -60 10110 -30
rect 10145 -60 10155 -30
rect 10100 -70 10155 -60
rect 10185 -30 10240 -20
rect 10185 -60 10195 -30
rect 10230 -60 10240 -30
rect 10185 -70 10240 -60
rect 10270 -30 10325 -20
rect 10270 -60 10280 -30
rect 10315 -60 10325 -30
rect 10270 -70 10325 -60
rect 10355 -30 10410 -20
rect 10355 -60 10365 -30
rect 10400 -60 10410 -30
rect 10355 -70 10410 -60
rect 10440 -30 10495 -20
rect 10440 -60 10450 -30
rect 10485 -60 10495 -30
rect 10440 -70 10495 -60
rect 10525 -30 10580 -20
rect 10525 -60 10535 -30
rect 10570 -60 10580 -30
rect 10525 -70 10580 -60
rect 10610 -30 10665 -20
rect 10610 -60 10620 -30
rect 10655 -60 10665 -30
rect 10610 -70 10665 -60
rect 10695 -30 10750 -20
rect 10695 -60 10705 -30
rect 10740 -60 10750 -30
rect 10695 -70 10750 -60
rect 10780 -30 10835 -20
rect 10780 -60 10790 -30
rect 10825 -60 10835 -30
rect 10780 -70 10835 -60
rect 10865 -30 10920 -20
rect 10865 -60 10875 -30
rect 10910 -60 10920 -30
rect 10865 -70 10920 -60
rect 10950 -30 11005 -20
rect 10950 -60 10960 -30
rect 10995 -60 11005 -30
rect 10950 -70 11005 -60
rect 11035 -30 11090 -20
rect 11035 -60 11045 -30
rect 11080 -60 11090 -30
rect 11035 -70 11090 -60
rect 11120 -30 11175 -20
rect 11120 -60 11130 -30
rect 11165 -60 11175 -30
rect 11120 -70 11175 -60
rect 11205 -30 11260 -20
rect 11205 -60 11215 -30
rect 11250 -60 11260 -30
rect 11205 -70 11260 -60
rect 11290 -30 11345 -20
rect 11290 -60 11300 -30
rect 11335 -60 11345 -30
rect 11290 -70 11345 -60
rect 11375 -30 11430 -20
rect 11375 -60 11385 -30
rect 11420 -60 11430 -30
rect 11375 -70 11430 -60
rect 11460 -30 11515 -20
rect 11460 -60 11470 -30
rect 11505 -60 11515 -30
rect 11460 -70 11515 -60
rect 11545 -30 11600 -20
rect 11545 -60 11555 -30
rect 11590 -60 11600 -30
rect 11545 -70 11600 -60
rect 11630 -30 11685 -20
rect 11630 -60 11640 -30
rect 11675 -60 11685 -30
rect 11630 -70 11685 -60
rect 11715 -30 11770 -20
rect 11715 -60 11725 -30
rect 11760 -60 11770 -30
rect 11715 -70 11770 -60
rect 11800 -30 11855 -20
rect 11800 -60 11810 -30
rect 11845 -60 11855 -30
rect 11800 -70 11855 -60
rect 11885 -30 11940 -20
rect 11885 -60 11895 -30
rect 11930 -60 11940 -30
rect 11885 -70 11940 -60
rect 11970 -30 12025 -20
rect 11970 -60 11980 -30
rect 12015 -60 12025 -30
rect 11970 -70 12025 -60
rect 12055 -30 12110 -20
rect 12055 -60 12065 -30
rect 12100 -60 12110 -30
rect 12055 -70 12110 -60
rect 12140 -30 12195 -20
rect 12140 -60 12150 -30
rect 12185 -60 12195 -30
rect 12140 -70 12195 -60
rect 12225 -30 12280 -20
rect 12225 -60 12235 -30
rect 12270 -60 12280 -30
rect 12225 -70 12280 -60
rect 12310 -30 12365 -20
rect 12310 -60 12320 -30
rect 12355 -60 12365 -30
rect 12310 -70 12365 -60
rect 12395 -30 12450 -20
rect 12395 -60 12405 -30
rect 12440 -60 12450 -30
rect 12395 -70 12450 -60
rect 12480 -30 12535 -20
rect 12480 -60 12490 -30
rect 12525 -60 12535 -30
rect 12480 -70 12535 -60
rect 12565 -30 12620 -20
rect 12565 -60 12575 -30
rect 12610 -60 12620 -30
rect 12565 -70 12620 -60
rect 12650 -30 12705 -20
rect 12650 -60 12660 -30
rect 12695 -60 12705 -30
rect 12650 -70 12705 -60
rect 12735 -30 12790 -20
rect 12735 -60 12745 -30
rect 12780 -60 12790 -30
rect 12735 -70 12790 -60
rect 12820 -30 12875 -20
rect 12820 -60 12830 -30
rect 12865 -60 12875 -30
rect 12820 -70 12875 -60
rect 12905 -30 12960 -20
rect 12905 -60 12915 -30
rect 12950 -60 12960 -30
rect 12905 -70 12960 -60
rect 12990 -30 13045 -20
rect 12990 -60 13000 -30
rect 13035 -60 13045 -30
rect 12990 -70 13045 -60
rect 13075 -30 13130 -20
rect 13075 -60 13085 -30
rect 13120 -60 13130 -30
rect 13075 -70 13130 -60
rect 13160 -30 13215 -20
rect 13160 -60 13170 -30
rect 13205 -60 13215 -30
rect 13160 -70 13215 -60
rect 13245 -30 13300 -20
rect 13245 -60 13255 -30
rect 13290 -60 13300 -30
rect 13245 -70 13300 -60
rect 13330 -30 13385 -20
rect 13330 -60 13340 -30
rect 13375 -60 13385 -30
rect 13330 -70 13385 -60
rect 13415 -30 13470 -20
rect 13415 -60 13425 -30
rect 13460 -60 13470 -30
rect 13415 -70 13470 -60
rect 13500 -30 13555 -20
rect 13500 -60 13510 -30
rect 13545 -60 13555 -30
rect 13500 -70 13555 -60
rect 13585 -30 13640 -20
rect 13585 -60 13595 -30
rect 13630 -60 13640 -30
rect 13585 -70 13640 -60
rect 13670 -30 13725 -20
rect 13670 -60 13680 -30
rect 13715 -60 13725 -30
rect 13670 -70 13725 -60
rect 13755 -30 13810 -20
rect 13755 -60 13765 -30
rect 13800 -60 13810 -30
rect 13755 -70 13810 -60
rect 13840 -30 13895 -20
rect 13840 -60 13850 -30
rect 13885 -60 13895 -30
rect 13840 -70 13895 -60
rect 13925 -30 13980 -20
rect 13925 -60 13935 -30
rect 13970 -60 13980 -30
rect 13925 -70 13980 -60
rect 14010 -30 14065 -20
rect 14010 -60 14020 -30
rect 14055 -60 14065 -30
rect 14010 -70 14065 -60
rect 14095 -30 14150 -20
rect 14095 -60 14105 -30
rect 14140 -60 14150 -30
rect 14095 -70 14150 -60
rect 14180 -30 14235 -20
rect 14180 -60 14190 -30
rect 14225 -60 14235 -30
rect 14180 -70 14235 -60
rect 14265 -30 14320 -20
rect 14265 -60 14275 -30
rect 14310 -60 14320 -30
rect 14265 -70 14320 -60
rect 14350 -30 14405 -20
rect 14350 -60 14360 -30
rect 14395 -60 14405 -30
rect 14350 -70 14405 -60
rect 14435 -30 14490 -20
rect 14435 -60 14445 -30
rect 14480 -60 14490 -30
rect 14435 -70 14490 -60
rect 14520 -30 14575 -20
rect 14520 -60 14530 -30
rect 14565 -60 14575 -30
rect 14520 -70 14575 -60
rect 14605 -30 14660 -20
rect 14605 -60 14615 -30
rect 14650 -60 14660 -30
rect 14605 -70 14660 -60
rect 14690 -30 14745 -20
rect 14690 -60 14700 -30
rect 14735 -60 14745 -30
rect 14690 -70 14745 -60
rect 14775 -30 14830 -20
rect 14775 -60 14785 -30
rect 14820 -60 14830 -30
rect 14775 -70 14830 -60
rect 14860 -30 14915 -20
rect 14860 -60 14870 -30
rect 14905 -60 14915 -30
rect 14860 -70 14915 -60
rect 14945 -30 15000 -20
rect 14945 -60 14955 -30
rect 14990 -60 15000 -30
rect 14945 -70 15000 -60
rect 15030 -30 15085 -20
rect 15030 -60 15040 -30
rect 15075 -60 15085 -30
rect 15030 -70 15085 -60
rect 15115 -30 15170 -20
rect 15115 -60 15125 -30
rect 15160 -60 15170 -30
rect 15115 -70 15170 -60
rect 15200 -30 15255 -20
rect 15200 -60 15210 -30
rect 15245 -60 15255 -30
rect 15200 -70 15255 -60
rect 15285 -30 15340 -20
rect 15285 -60 15295 -30
rect 15330 -60 15340 -30
rect 15285 -70 15340 -60
rect 15370 -30 15425 -20
rect 15370 -60 15380 -30
rect 15415 -60 15425 -30
rect 15370 -70 15425 -60
rect 15455 -30 15510 -20
rect 15455 -60 15465 -30
rect 15500 -60 15510 -30
rect 15455 -70 15510 -60
rect 15540 -30 15595 -20
rect 15540 -60 15550 -30
rect 15585 -60 15595 -30
rect 15540 -70 15595 -60
rect 15625 -30 15680 -20
rect 15625 -60 15635 -30
rect 15670 -60 15680 -30
rect 15625 -70 15680 -60
rect 15710 -30 15765 -20
rect 15710 -60 15720 -30
rect 15755 -60 15765 -30
rect 15710 -70 15765 -60
rect 15795 -30 15850 -20
rect 15795 -60 15805 -30
rect 15840 -60 15850 -30
rect 15795 -70 15850 -60
rect 15880 -30 15935 -20
rect 15880 -60 15890 -30
rect 15925 -60 15935 -30
rect 15880 -70 15935 -60
rect 15965 -30 16020 -20
rect 15965 -60 15975 -30
rect 16010 -60 16020 -30
rect 15965 -70 16020 -60
rect 16050 -30 16105 -20
rect 16050 -60 16060 -30
rect 16095 -60 16105 -30
rect 16050 -70 16105 -60
rect 16135 -30 16190 -20
rect 16135 -60 16145 -30
rect 16180 -60 16190 -30
rect 16135 -70 16190 -60
rect 16220 -30 16275 -20
rect 16220 -60 16230 -30
rect 16265 -60 16275 -30
rect 16220 -70 16275 -60
rect 16305 -30 16360 -20
rect 16305 -60 16315 -30
rect 16350 -60 16360 -30
rect 16305 -70 16360 -60
rect 16390 -30 16445 -20
rect 16390 -60 16400 -30
rect 16435 -60 16445 -30
rect 16390 -70 16445 -60
rect 16475 -30 16530 -20
rect 16475 -60 16485 -30
rect 16520 -60 16530 -30
rect 16475 -70 16530 -60
rect 16560 -30 16615 -20
rect 16560 -60 16570 -30
rect 16605 -60 16615 -30
rect 16560 -70 16615 -60
rect 16645 -30 16700 -20
rect 16645 -60 16655 -30
rect 16690 -60 16700 -30
rect 16645 -70 16700 -60
rect 16730 -30 16785 -20
rect 16730 -60 16740 -30
rect 16775 -60 16785 -30
rect 16730 -70 16785 -60
rect 16815 -30 16870 -20
rect 16815 -60 16825 -30
rect 16860 -60 16870 -30
rect 16815 -70 16870 -60
rect 16900 -30 16955 -20
rect 16900 -60 16910 -30
rect 16945 -60 16955 -30
rect 16900 -70 16955 -60
rect 16985 -30 17040 -20
rect 16985 -60 16995 -30
rect 17030 -60 17040 -30
rect 16985 -70 17040 -60
rect 17070 -30 17125 -20
rect 17070 -60 17080 -30
rect 17115 -60 17125 -30
rect 17070 -70 17125 -60
rect 17155 -30 17210 -20
rect 17155 -60 17165 -30
rect 17200 -60 17210 -30
rect 17155 -70 17210 -60
rect 17240 -30 17295 -20
rect 17240 -60 17250 -30
rect 17285 -60 17295 -30
rect 17240 -70 17295 -60
rect 17325 -30 17380 -20
rect 17325 -60 17335 -30
rect 17370 -60 17380 -30
rect 17325 -70 17380 -60
rect 17410 -30 17465 -20
rect 17410 -60 17420 -30
rect 17455 -60 17465 -30
rect 17410 -70 17465 -60
rect 17495 -30 17550 -20
rect 17495 -60 17505 -30
rect 17540 -60 17550 -30
rect 17495 -70 17550 -60
rect 17580 -30 17635 -20
rect 17580 -60 17590 -30
rect 17625 -60 17635 -30
rect 17580 -70 17635 -60
rect 17665 -30 17720 -20
rect 17665 -60 17675 -30
rect 17710 -60 17720 -30
rect 17665 -70 17720 -60
rect 17750 -30 17805 -20
rect 17750 -60 17760 -30
rect 17795 -60 17805 -30
rect 17750 -70 17805 -60
rect 17835 -30 17890 -20
rect 17835 -60 17845 -30
rect 17880 -60 17890 -30
rect 17835 -70 17890 -60
rect 17920 -30 17975 -20
rect 17920 -60 17930 -30
rect 17965 -60 17975 -30
rect 17920 -70 17975 -60
rect 18005 -30 18060 -20
rect 18005 -60 18015 -30
rect 18050 -60 18060 -30
rect 18005 -70 18060 -60
rect 18090 -30 18145 -20
rect 18090 -60 18100 -30
rect 18135 -60 18145 -30
rect 18090 -70 18145 -60
rect 18175 -30 18230 -20
rect 18175 -60 18185 -30
rect 18220 -60 18230 -30
rect 18175 -70 18230 -60
rect 18260 -30 18315 -20
rect 18260 -60 18270 -30
rect 18305 -60 18315 -30
rect 18260 -70 18315 -60
rect 18345 -30 18400 -20
rect 18345 -60 18355 -30
rect 18390 -60 18400 -30
rect 18345 -70 18400 -60
rect 18430 -30 18485 -20
rect 18430 -60 18440 -30
rect 18475 -60 18485 -30
rect 18430 -70 18485 -60
rect 18515 -30 18570 -20
rect 18515 -60 18525 -30
rect 18560 -60 18570 -30
rect 18515 -70 18570 -60
rect 18600 -30 18655 -20
rect 18600 -60 18610 -30
rect 18645 -60 18655 -30
rect 18600 -70 18655 -60
rect 18685 -30 18740 -20
rect 18685 -60 18695 -30
rect 18730 -60 18740 -30
rect 18685 -70 18740 -60
rect 18770 -30 18825 -20
rect 18770 -60 18780 -30
rect 18815 -60 18825 -30
rect 18770 -70 18825 -60
rect 18855 -30 18910 -20
rect 18855 -60 18865 -30
rect 18900 -60 18910 -30
rect 18855 -70 18910 -60
rect 18940 -30 18995 -20
rect 18940 -60 18950 -30
rect 18985 -60 18995 -30
rect 18940 -70 18995 -60
rect 19025 -30 19080 -20
rect 19025 -60 19035 -30
rect 19070 -60 19080 -30
rect 19025 -70 19080 -60
rect 19110 -30 19165 -20
rect 19110 -60 19120 -30
rect 19155 -60 19165 -30
rect 19110 -70 19165 -60
rect 19195 -30 19250 -20
rect 19195 -60 19205 -30
rect 19240 -60 19250 -30
rect 19195 -70 19250 -60
rect 19280 -30 19335 -20
rect 19280 -60 19290 -30
rect 19325 -60 19335 -30
rect 19280 -70 19335 -60
rect 19365 -30 19420 -20
rect 19365 -60 19375 -30
rect 19410 -60 19420 -30
rect 19365 -70 19420 -60
rect 19450 -30 19505 -20
rect 19450 -60 19460 -30
rect 19495 -60 19505 -30
rect 19450 -70 19505 -60
rect 19535 -30 19590 -20
rect 19535 -60 19545 -30
rect 19580 -60 19590 -30
rect 19535 -70 19590 -60
rect 19620 -30 19675 -20
rect 19620 -60 19630 -30
rect 19665 -60 19675 -30
rect 19620 -70 19675 -60
rect 19705 -30 19760 -20
rect 19705 -60 19715 -30
rect 19750 -60 19760 -30
rect 19705 -70 19760 -60
rect 19790 -30 19845 -20
rect 19790 -60 19800 -30
rect 19835 -60 19845 -30
rect 19790 -70 19845 -60
rect 19875 -30 19930 -20
rect 19875 -60 19885 -30
rect 19920 -60 19930 -30
rect 19875 -70 19930 -60
rect 19960 -30 20015 -20
rect 19960 -60 19970 -30
rect 20005 -60 20015 -30
rect 19960 -70 20015 -60
rect 20045 -30 20100 -20
rect 20045 -60 20055 -30
rect 20090 -60 20100 -30
rect 20045 -70 20100 -60
rect 20130 -30 20185 -20
rect 20130 -60 20140 -30
rect 20175 -60 20185 -30
rect 20130 -70 20185 -60
rect 20215 -30 20270 -20
rect 20215 -60 20225 -30
rect 20260 -60 20270 -30
rect 20215 -70 20270 -60
rect 20300 -30 20355 -20
rect 20300 -60 20310 -30
rect 20345 -60 20355 -30
rect 20300 -70 20355 -60
rect 20385 -30 20440 -20
rect 20385 -60 20395 -30
rect 20430 -60 20440 -30
rect 20385 -70 20440 -60
rect 20470 -30 20525 -20
rect 20470 -60 20480 -30
rect 20515 -60 20525 -30
rect 20470 -70 20525 -60
rect 20555 -30 20610 -20
rect 20555 -60 20565 -30
rect 20600 -60 20610 -30
rect 20555 -70 20610 -60
rect 20640 -30 20695 -20
rect 20640 -60 20650 -30
rect 20685 -60 20695 -30
rect 20640 -70 20695 -60
rect 20725 -30 20780 -20
rect 20725 -60 20735 -30
rect 20770 -60 20780 -30
rect 20725 -70 20780 -60
rect 20810 -30 20865 -20
rect 20810 -60 20820 -30
rect 20855 -60 20865 -30
rect 20810 -70 20865 -60
rect 20895 -30 20950 -20
rect 20895 -60 20905 -30
rect 20940 -60 20950 -30
rect 20895 -70 20950 -60
rect 20980 -30 21035 -20
rect 20980 -60 20990 -30
rect 21025 -60 21035 -30
rect 20980 -70 21035 -60
rect 21065 -30 21120 -20
rect 21065 -60 21075 -30
rect 21110 -60 21120 -30
rect 21065 -70 21120 -60
rect 21150 -30 21205 -20
rect 21150 -60 21160 -30
rect 21195 -60 21205 -30
rect 21150 -70 21205 -60
rect 21235 -30 21290 -20
rect 21235 -60 21245 -30
rect 21280 -60 21290 -30
rect 21235 -70 21290 -60
rect 21320 -30 21375 -20
rect 21320 -60 21330 -30
rect 21365 -60 21375 -30
rect 21320 -70 21375 -60
rect 21405 -30 21460 -20
rect 21405 -60 21415 -30
rect 21450 -60 21460 -30
rect 21405 -70 21460 -60
rect 21490 -30 21545 -20
rect 21490 -60 21500 -30
rect 21535 -60 21545 -30
rect 21490 -70 21545 -60
rect 21575 -30 21630 -20
rect 21575 -60 21585 -30
rect 21620 -60 21630 -30
rect 21575 -70 21630 -60
rect 21660 -30 21715 -20
rect 21660 -60 21670 -30
rect 21705 -60 21715 -30
rect 21660 -70 21715 -60
rect 21745 -30 21800 -20
rect 21745 -60 21755 -30
rect 21790 -60 21800 -30
rect 21745 -70 21800 -60
rect 21830 -30 21885 -20
rect 21830 -60 21840 -30
rect 21875 -60 21885 -30
rect 21830 -70 21885 -60
rect 21915 -30 21970 -20
rect 21915 -60 21925 -30
rect 21960 -60 21970 -30
rect 21915 -70 21970 -60
rect 22000 -30 22055 -20
rect 22000 -60 22010 -30
rect 22045 -60 22055 -30
rect 22000 -70 22055 -60
rect 22085 -30 22140 -20
rect 22085 -60 22095 -30
rect 22130 -60 22140 -30
rect 22085 -70 22140 -60
rect 22170 -30 22225 -20
rect 22170 -60 22180 -30
rect 22215 -60 22225 -30
rect 22170 -70 22225 -60
rect 22255 -30 22310 -20
rect 22255 -60 22265 -30
rect 22300 -60 22310 -30
rect 22255 -70 22310 -60
rect 22340 -30 22395 -20
rect 22340 -60 22350 -30
rect 22385 -60 22395 -30
rect 22340 -70 22395 -60
rect 22425 -30 22480 -20
rect 22425 -60 22435 -30
rect 22470 -60 22480 -30
rect 22425 -70 22480 -60
rect 22510 -30 22565 -20
rect 22510 -60 22520 -30
rect 22555 -60 22565 -30
rect 22510 -70 22565 -60
rect 22595 -30 22650 -20
rect 22595 -60 22605 -30
rect 22640 -60 22650 -30
rect 22595 -70 22650 -60
rect 22680 -30 22735 -20
rect 22680 -60 22690 -30
rect 22725 -60 22735 -30
rect 22680 -70 22735 -60
rect 22765 -30 22820 -20
rect 22765 -60 22775 -30
rect 22810 -60 22820 -30
rect 22765 -70 22820 -60
rect 22850 -30 22905 -20
rect 22850 -60 22860 -30
rect 22895 -60 22905 -30
rect 22850 -70 22905 -60
rect 22935 -30 22990 -20
rect 22935 -60 22945 -30
rect 22980 -60 22990 -30
rect 22935 -70 22990 -60
rect 23020 -30 23075 -20
rect 23020 -60 23030 -30
rect 23065 -60 23075 -30
rect 23020 -70 23075 -60
rect 23105 -30 23160 -20
rect 23105 -60 23115 -30
rect 23150 -60 23160 -30
rect 23105 -70 23160 -60
rect 23190 -30 23245 -20
rect 23190 -60 23200 -30
rect 23235 -60 23245 -30
rect 23190 -70 23245 -60
rect 23275 -30 23330 -20
rect 23275 -60 23285 -30
rect 23320 -60 23330 -30
rect 23275 -70 23330 -60
rect 23360 -30 23415 -20
rect 23360 -60 23370 -30
rect 23405 -60 23415 -30
rect 23360 -70 23415 -60
rect 23445 -30 23500 -20
rect 23445 -60 23455 -30
rect 23490 -60 23500 -30
rect 23445 -70 23500 -60
rect 23530 -30 23585 -20
rect 23530 -60 23540 -30
rect 23575 -60 23585 -30
rect 23530 -70 23585 -60
rect 23615 -30 23670 -20
rect 23615 -60 23625 -30
rect 23660 -60 23670 -30
rect 23615 -70 23670 -60
rect 23700 -30 23755 -20
rect 23700 -60 23710 -30
rect 23745 -60 23755 -30
rect 23700 -70 23755 -60
rect 23785 -30 23840 -20
rect 23785 -60 23795 -30
rect 23830 -60 23840 -30
rect 23785 -70 23840 -60
rect 23870 -30 23925 -20
rect 23870 -60 23880 -30
rect 23915 -60 23925 -30
rect 23870 -70 23925 -60
rect 23955 -30 24010 -20
rect 23955 -60 23965 -30
rect 24000 -60 24010 -30
rect 23955 -70 24010 -60
rect 24040 -30 24095 -20
rect 24040 -60 24050 -30
rect 24085 -60 24095 -30
rect 24040 -70 24095 -60
rect 24125 -30 24180 -20
rect 24125 -60 24135 -30
rect 24170 -60 24180 -30
rect 24125 -70 24180 -60
rect 24210 -30 24265 -20
rect 24210 -60 24220 -30
rect 24255 -60 24265 -30
rect 24210 -70 24265 -60
rect 24295 -30 24350 -20
rect 24295 -60 24305 -30
rect 24340 -60 24350 -30
rect 24295 -70 24350 -60
rect 24380 -30 24435 -20
rect 24380 -60 24390 -30
rect 24425 -60 24435 -30
rect 24380 -70 24435 -60
rect 24465 -30 24520 -20
rect 24465 -60 24475 -30
rect 24510 -60 24520 -30
rect 24465 -70 24520 -60
rect 24550 -30 24605 -20
rect 24550 -60 24560 -30
rect 24595 -60 24605 -30
rect 24550 -70 24605 -60
rect 24635 -30 24690 -20
rect 24635 -60 24645 -30
rect 24680 -60 24690 -30
rect 24635 -70 24690 -60
rect 24720 -30 24775 -20
rect 24720 -60 24730 -30
rect 24765 -60 24775 -30
rect 24720 -70 24775 -60
rect 24805 -30 24860 -20
rect 24805 -60 24815 -30
rect 24850 -60 24860 -30
rect 24805 -70 24860 -60
rect 24890 -30 24945 -20
rect 24890 -60 24900 -30
rect 24935 -60 24945 -30
rect 24890 -70 24945 -60
rect 24975 -30 25030 -20
rect 24975 -60 24985 -30
rect 25020 -60 25030 -30
rect 24975 -70 25030 -60
rect 25060 -30 25115 -20
rect 25060 -60 25070 -30
rect 25105 -60 25115 -30
rect 25060 -70 25115 -60
rect 25145 -30 25200 -20
rect 25145 -60 25155 -30
rect 25190 -60 25200 -30
rect 25145 -70 25200 -60
rect 25230 -30 25285 -20
rect 25230 -60 25240 -30
rect 25275 -60 25285 -30
rect 25230 -70 25285 -60
rect 25315 -30 25370 -20
rect 25315 -60 25325 -30
rect 25360 -60 25370 -30
rect 25315 -70 25370 -60
rect 25400 -30 25455 -20
rect 25400 -60 25410 -30
rect 25445 -60 25455 -30
rect 25400 -70 25455 -60
rect 25485 -30 25540 -20
rect 25485 -60 25495 -30
rect 25530 -60 25540 -30
rect 25485 -70 25540 -60
rect 25570 -30 25625 -20
rect 25570 -60 25580 -30
rect 25615 -60 25625 -30
rect 25570 -70 25625 -60
rect 25655 -30 25710 -20
rect 25655 -60 25665 -30
rect 25700 -60 25710 -30
rect 25655 -70 25710 -60
rect 25740 -30 25795 -20
rect 25740 -60 25750 -30
rect 25785 -60 25795 -30
rect 25740 -70 25795 -60
rect 25825 -30 25880 -20
rect 25825 -60 25835 -30
rect 25870 -60 25880 -30
rect 25825 -70 25880 -60
rect 25910 -30 25965 -20
rect 25910 -60 25920 -30
rect 25955 -60 25965 -30
rect 25910 -70 25965 -60
rect 25995 -30 26050 -20
rect 25995 -60 26005 -30
rect 26040 -60 26050 -30
rect 25995 -70 26050 -60
rect 26080 -30 26135 -20
rect 26080 -60 26090 -30
rect 26125 -60 26135 -30
rect 26080 -70 26135 -60
rect 26165 -30 26220 -20
rect 26165 -60 26175 -30
rect 26210 -60 26220 -30
rect 26165 -70 26220 -60
rect 26250 -30 26305 -20
rect 26250 -60 26260 -30
rect 26295 -60 26305 -30
rect 26250 -70 26305 -60
rect 26335 -30 26390 -20
rect 26335 -60 26345 -30
rect 26380 -60 26390 -30
rect 26335 -70 26390 -60
rect 26420 -30 26475 -20
rect 26420 -60 26430 -30
rect 26465 -60 26475 -30
rect 26420 -70 26475 -60
rect 26505 -30 26560 -20
rect 26505 -60 26515 -30
rect 26550 -60 26560 -30
rect 26505 -70 26560 -60
rect 26590 -30 26645 -20
rect 26590 -60 26600 -30
rect 26635 -60 26645 -30
rect 26590 -70 26645 -60
rect 26675 -30 26730 -20
rect 26675 -60 26685 -30
rect 26720 -60 26730 -30
rect 26675 -70 26730 -60
rect 26760 -30 26815 -20
rect 26760 -60 26770 -30
rect 26805 -60 26815 -30
rect 26760 -70 26815 -60
rect 26845 -30 26900 -20
rect 26845 -60 26855 -30
rect 26890 -60 26900 -30
rect 26845 -70 26900 -60
rect 26930 -30 26985 -20
rect 26930 -60 26940 -30
rect 26975 -60 26985 -30
rect 26930 -70 26985 -60
rect 27015 -30 27070 -20
rect 27015 -60 27025 -30
rect 27060 -60 27070 -30
rect 27015 -70 27070 -60
rect 27100 -30 27155 -20
rect 27100 -60 27110 -30
rect 27145 -60 27155 -30
rect 27100 -70 27155 -60
rect 27185 -30 27240 -20
rect 27185 -60 27195 -30
rect 27230 -60 27240 -30
rect 27185 -70 27240 -60
rect 27270 -30 27325 -20
rect 27270 -60 27280 -30
rect 27315 -60 27325 -30
rect 27270 -70 27325 -60
rect 27355 -30 27410 -20
rect 27355 -60 27365 -30
rect 27400 -60 27410 -30
rect 27355 -70 27410 -60
rect 27440 -30 27495 -20
rect 27440 -60 27450 -30
rect 27485 -60 27495 -30
rect 27440 -70 27495 -60
rect 27525 -30 27580 -20
rect 27525 -60 27535 -30
rect 27570 -60 27580 -30
rect 27525 -70 27580 -60
rect 27610 -30 27665 -20
rect 27610 -60 27620 -30
rect 27655 -60 27665 -30
rect 27610 -70 27665 -60
rect 27695 -30 27750 -20
rect 27695 -60 27705 -30
rect 27740 -60 27750 -30
rect 27695 -70 27750 -60
rect 27780 -30 27835 -20
rect 27780 -60 27790 -30
rect 27825 -60 27835 -30
rect 27780 -70 27835 -60
rect 27865 -30 27920 -20
rect 27865 -60 27875 -30
rect 27910 -60 27920 -30
rect 27865 -70 27920 -60
rect 27950 -30 28005 -20
rect 27950 -60 27960 -30
rect 27995 -60 28005 -30
rect 27950 -70 28005 -60
rect 28035 -30 28090 -20
rect 28035 -60 28045 -30
rect 28080 -60 28090 -30
rect 28035 -70 28090 -60
rect 28120 -30 28175 -20
rect 28120 -60 28130 -30
rect 28165 -60 28175 -30
rect 28120 -70 28175 -60
rect 28205 -30 28260 -20
rect 28205 -60 28215 -30
rect 28250 -60 28260 -30
rect 28205 -70 28260 -60
rect 28290 -30 28345 -20
rect 28290 -60 28300 -30
rect 28335 -60 28345 -30
rect 28290 -70 28345 -60
rect 28375 -30 28430 -20
rect 28375 -60 28385 -30
rect 28420 -60 28430 -30
rect 28375 -70 28430 -60
rect 28460 -30 28515 -20
rect 28460 -60 28470 -30
rect 28505 -60 28515 -30
rect 28460 -70 28515 -60
rect 28545 -30 28600 -20
rect 28545 -60 28555 -30
rect 28590 -60 28600 -30
rect 28545 -70 28600 -60
rect 28630 -30 28685 -20
rect 28630 -60 28640 -30
rect 28675 -60 28685 -30
rect 28630 -70 28685 -60
rect 28715 -30 28770 -20
rect 28715 -60 28725 -30
rect 28760 -60 28770 -30
rect 28715 -70 28770 -60
rect 28800 -30 28855 -20
rect 28800 -60 28810 -30
rect 28845 -60 28855 -30
rect 28800 -70 28855 -60
rect 28885 -30 28940 -20
rect 28885 -60 28895 -30
rect 28930 -60 28940 -30
rect 28885 -70 28940 -60
rect 28970 -30 29025 -20
rect 28970 -60 28980 -30
rect 29015 -60 29025 -30
rect 28970 -70 29025 -60
rect 29055 -30 29110 -20
rect 29055 -60 29065 -30
rect 29100 -60 29110 -30
rect 29055 -70 29110 -60
rect 29140 -30 29195 -20
rect 29140 -60 29150 -30
rect 29185 -60 29195 -30
rect 29140 -70 29195 -60
rect 29225 -30 29280 -20
rect 29225 -60 29235 -30
rect 29270 -60 29280 -30
rect 29225 -70 29280 -60
rect 29310 -30 29365 -20
rect 29310 -60 29320 -30
rect 29355 -60 29365 -30
rect 29310 -70 29365 -60
rect 29395 -30 29450 -20
rect 29395 -60 29405 -30
rect 29440 -60 29450 -30
rect 29395 -70 29450 -60
rect 29480 -30 29535 -20
rect 29480 -60 29490 -30
rect 29525 -60 29535 -30
rect 29480 -70 29535 -60
rect 29565 -30 29620 -20
rect 29565 -60 29575 -30
rect 29610 -60 29620 -30
rect 29565 -70 29620 -60
rect 105 -265 160 -255
rect 105 -295 115 -265
rect 150 -295 160 -265
rect 105 -305 160 -295
rect 190 -265 245 -255
rect 190 -295 200 -265
rect 235 -295 245 -265
rect 190 -305 245 -295
rect 275 -265 330 -255
rect 275 -295 285 -265
rect 320 -295 330 -265
rect 275 -305 330 -295
rect 360 -265 415 -255
rect 360 -295 370 -265
rect 405 -295 415 -265
rect 360 -305 415 -295
rect 445 -265 500 -255
rect 445 -295 455 -265
rect 490 -295 500 -265
rect 445 -305 500 -295
rect 530 -265 585 -255
rect 530 -295 540 -265
rect 575 -295 585 -265
rect 530 -305 585 -295
rect 615 -265 670 -255
rect 615 -295 625 -265
rect 660 -295 670 -265
rect 615 -305 670 -295
rect 700 -265 755 -255
rect 700 -295 710 -265
rect 745 -295 755 -265
rect 700 -305 755 -295
rect 785 -265 840 -255
rect 785 -295 795 -265
rect 830 -295 840 -265
rect 785 -305 840 -295
rect 870 -265 925 -255
rect 870 -295 880 -265
rect 915 -295 925 -265
rect 870 -305 925 -295
rect 955 -265 1010 -255
rect 955 -295 965 -265
rect 1000 -295 1010 -265
rect 955 -305 1010 -295
rect 1040 -265 1095 -255
rect 1040 -295 1050 -265
rect 1085 -295 1095 -265
rect 1040 -305 1095 -295
rect 1125 -265 1180 -255
rect 1125 -295 1135 -265
rect 1170 -295 1180 -265
rect 1125 -305 1180 -295
rect 1210 -265 1265 -255
rect 1210 -295 1220 -265
rect 1255 -295 1265 -265
rect 1210 -305 1265 -295
rect 1295 -265 1350 -255
rect 1295 -295 1305 -265
rect 1340 -295 1350 -265
rect 1295 -305 1350 -295
rect 1380 -265 1435 -255
rect 1380 -295 1390 -265
rect 1425 -295 1435 -265
rect 1380 -305 1435 -295
rect 1465 -265 1520 -255
rect 1465 -295 1475 -265
rect 1510 -295 1520 -265
rect 1465 -305 1520 -295
rect 1550 -265 1605 -255
rect 1550 -295 1560 -265
rect 1595 -295 1605 -265
rect 1550 -305 1605 -295
rect 1635 -265 1690 -255
rect 1635 -295 1645 -265
rect 1680 -295 1690 -265
rect 1635 -305 1690 -295
rect 1720 -265 1775 -255
rect 1720 -295 1730 -265
rect 1765 -295 1775 -265
rect 1720 -305 1775 -295
rect 1805 -265 1860 -255
rect 1805 -295 1815 -265
rect 1850 -295 1860 -265
rect 1805 -305 1860 -295
rect 1890 -265 1945 -255
rect 1890 -295 1900 -265
rect 1935 -295 1945 -265
rect 1890 -305 1945 -295
rect 1975 -265 2030 -255
rect 1975 -295 1985 -265
rect 2020 -295 2030 -265
rect 1975 -305 2030 -295
rect 2060 -265 2115 -255
rect 2060 -295 2070 -265
rect 2105 -295 2115 -265
rect 2060 -305 2115 -295
rect 2145 -265 2200 -255
rect 2145 -295 2155 -265
rect 2190 -295 2200 -265
rect 2145 -305 2200 -295
rect 2230 -265 2285 -255
rect 2230 -295 2240 -265
rect 2275 -295 2285 -265
rect 2230 -305 2285 -295
rect 2315 -265 2370 -255
rect 2315 -295 2325 -265
rect 2360 -295 2370 -265
rect 2315 -305 2370 -295
rect 2400 -265 2455 -255
rect 2400 -295 2410 -265
rect 2445 -295 2455 -265
rect 2400 -305 2455 -295
rect 2485 -265 2540 -255
rect 2485 -295 2495 -265
rect 2530 -295 2540 -265
rect 2485 -305 2540 -295
rect 2570 -265 2625 -255
rect 2570 -295 2580 -265
rect 2615 -295 2625 -265
rect 2570 -305 2625 -295
rect 2655 -265 2710 -255
rect 2655 -295 2665 -265
rect 2700 -295 2710 -265
rect 2655 -305 2710 -295
rect 2740 -265 2795 -255
rect 2740 -295 2750 -265
rect 2785 -295 2795 -265
rect 2740 -305 2795 -295
rect 2825 -265 2880 -255
rect 2825 -295 2835 -265
rect 2870 -295 2880 -265
rect 2825 -305 2880 -295
rect 2910 -265 2965 -255
rect 2910 -295 2920 -265
rect 2955 -295 2965 -265
rect 2910 -305 2965 -295
rect 2995 -265 3050 -255
rect 2995 -295 3005 -265
rect 3040 -295 3050 -265
rect 2995 -305 3050 -295
rect 3080 -265 3135 -255
rect 3080 -295 3090 -265
rect 3125 -295 3135 -265
rect 3080 -305 3135 -295
rect 3165 -265 3220 -255
rect 3165 -295 3175 -265
rect 3210 -295 3220 -265
rect 3165 -305 3220 -295
rect 3250 -265 3305 -255
rect 3250 -295 3260 -265
rect 3295 -295 3305 -265
rect 3250 -305 3305 -295
rect 3335 -265 3390 -255
rect 3335 -295 3345 -265
rect 3380 -295 3390 -265
rect 3335 -305 3390 -295
rect 3420 -265 3475 -255
rect 3420 -295 3430 -265
rect 3465 -295 3475 -265
rect 3420 -305 3475 -295
rect 3505 -265 3560 -255
rect 3505 -295 3515 -265
rect 3550 -295 3560 -265
rect 3505 -305 3560 -295
rect 3590 -265 3645 -255
rect 3590 -295 3600 -265
rect 3635 -295 3645 -265
rect 3590 -305 3645 -295
rect 3675 -265 3730 -255
rect 3675 -295 3685 -265
rect 3720 -295 3730 -265
rect 3675 -305 3730 -295
rect 3760 -265 3815 -255
rect 3760 -295 3770 -265
rect 3805 -295 3815 -265
rect 3760 -305 3815 -295
rect 3845 -265 3900 -255
rect 3845 -295 3855 -265
rect 3890 -295 3900 -265
rect 3845 -305 3900 -295
rect 3930 -265 3985 -255
rect 3930 -295 3940 -265
rect 3975 -295 3985 -265
rect 3930 -305 3985 -295
rect 4015 -265 4070 -255
rect 4015 -295 4025 -265
rect 4060 -295 4070 -265
rect 4015 -305 4070 -295
rect 4100 -265 4155 -255
rect 4100 -295 4110 -265
rect 4145 -295 4155 -265
rect 4100 -305 4155 -295
rect 4185 -265 4240 -255
rect 4185 -295 4195 -265
rect 4230 -295 4240 -265
rect 4185 -305 4240 -295
rect 4270 -265 4325 -255
rect 4270 -295 4280 -265
rect 4315 -295 4325 -265
rect 4270 -305 4325 -295
rect 4355 -265 4410 -255
rect 4355 -295 4365 -265
rect 4400 -295 4410 -265
rect 4355 -305 4410 -295
rect 4440 -265 4495 -255
rect 4440 -295 4450 -265
rect 4485 -295 4495 -265
rect 4440 -305 4495 -295
rect 4525 -265 4580 -255
rect 4525 -295 4535 -265
rect 4570 -295 4580 -265
rect 4525 -305 4580 -295
rect 4610 -265 4665 -255
rect 4610 -295 4620 -265
rect 4655 -295 4665 -265
rect 4610 -305 4665 -295
rect 4695 -265 4750 -255
rect 4695 -295 4705 -265
rect 4740 -295 4750 -265
rect 4695 -305 4750 -295
rect 4780 -265 4835 -255
rect 4780 -295 4790 -265
rect 4825 -295 4835 -265
rect 4780 -305 4835 -295
rect 4865 -265 4920 -255
rect 4865 -295 4875 -265
rect 4910 -295 4920 -265
rect 4865 -305 4920 -295
rect 4950 -265 5005 -255
rect 4950 -295 4960 -265
rect 4995 -295 5005 -265
rect 4950 -305 5005 -295
rect 5035 -265 5090 -255
rect 5035 -295 5045 -265
rect 5080 -295 5090 -265
rect 5035 -305 5090 -295
rect 5120 -265 5175 -255
rect 5120 -295 5130 -265
rect 5165 -295 5175 -265
rect 5120 -305 5175 -295
rect 5205 -265 5260 -255
rect 5205 -295 5215 -265
rect 5250 -295 5260 -265
rect 5205 -305 5260 -295
rect 5290 -265 5345 -255
rect 5290 -295 5300 -265
rect 5335 -295 5345 -265
rect 5290 -305 5345 -295
rect 5375 -265 5430 -255
rect 5375 -295 5385 -265
rect 5420 -295 5430 -265
rect 5375 -305 5430 -295
rect 5460 -265 5515 -255
rect 5460 -295 5470 -265
rect 5505 -295 5515 -265
rect 5460 -305 5515 -295
rect 5545 -265 5600 -255
rect 5545 -295 5555 -265
rect 5590 -295 5600 -265
rect 5545 -305 5600 -295
rect 5630 -265 5685 -255
rect 5630 -295 5640 -265
rect 5675 -295 5685 -265
rect 5630 -305 5685 -295
rect 5715 -265 5770 -255
rect 5715 -295 5725 -265
rect 5760 -295 5770 -265
rect 5715 -305 5770 -295
rect 5800 -265 5855 -255
rect 5800 -295 5810 -265
rect 5845 -295 5855 -265
rect 5800 -305 5855 -295
rect 5885 -265 5940 -255
rect 5885 -295 5895 -265
rect 5930 -295 5940 -265
rect 5885 -305 5940 -295
rect 5970 -265 6025 -255
rect 5970 -295 5980 -265
rect 6015 -295 6025 -265
rect 5970 -305 6025 -295
rect 6055 -265 6110 -255
rect 6055 -295 6065 -265
rect 6100 -295 6110 -265
rect 6055 -305 6110 -295
rect 6140 -265 6195 -255
rect 6140 -295 6150 -265
rect 6185 -295 6195 -265
rect 6140 -305 6195 -295
rect 6225 -265 6280 -255
rect 6225 -295 6235 -265
rect 6270 -295 6280 -265
rect 6225 -305 6280 -295
rect 6310 -265 6365 -255
rect 6310 -295 6320 -265
rect 6355 -295 6365 -265
rect 6310 -305 6365 -295
rect 6395 -265 6450 -255
rect 6395 -295 6405 -265
rect 6440 -295 6450 -265
rect 6395 -305 6450 -295
rect 6480 -265 6535 -255
rect 6480 -295 6490 -265
rect 6525 -295 6535 -265
rect 6480 -305 6535 -295
rect 6565 -265 6620 -255
rect 6565 -295 6575 -265
rect 6610 -295 6620 -265
rect 6565 -305 6620 -295
rect 6650 -265 6705 -255
rect 6650 -295 6660 -265
rect 6695 -295 6705 -265
rect 6650 -305 6705 -295
rect 6735 -265 6790 -255
rect 6735 -295 6745 -265
rect 6780 -295 6790 -265
rect 6735 -305 6790 -295
rect 6820 -265 6875 -255
rect 6820 -295 6830 -265
rect 6865 -295 6875 -265
rect 6820 -305 6875 -295
rect 6905 -265 6960 -255
rect 6905 -295 6915 -265
rect 6950 -295 6960 -265
rect 6905 -305 6960 -295
rect 6990 -265 7045 -255
rect 6990 -295 7000 -265
rect 7035 -295 7045 -265
rect 6990 -305 7045 -295
rect 7075 -265 7130 -255
rect 7075 -295 7085 -265
rect 7120 -295 7130 -265
rect 7075 -305 7130 -295
rect 7160 -265 7215 -255
rect 7160 -295 7170 -265
rect 7205 -295 7215 -265
rect 7160 -305 7215 -295
rect 7245 -265 7300 -255
rect 7245 -295 7255 -265
rect 7290 -295 7300 -265
rect 7245 -305 7300 -295
rect 7330 -265 7385 -255
rect 7330 -295 7340 -265
rect 7375 -295 7385 -265
rect 7330 -305 7385 -295
rect 7415 -265 7470 -255
rect 7415 -295 7425 -265
rect 7460 -295 7470 -265
rect 7415 -305 7470 -295
rect 7500 -265 7555 -255
rect 7500 -295 7510 -265
rect 7545 -295 7555 -265
rect 7500 -305 7555 -295
rect 7585 -265 7640 -255
rect 7585 -295 7595 -265
rect 7630 -295 7640 -265
rect 7585 -305 7640 -295
rect 7670 -265 7725 -255
rect 7670 -295 7680 -265
rect 7715 -295 7725 -265
rect 7670 -305 7725 -295
rect 7755 -265 7810 -255
rect 7755 -295 7765 -265
rect 7800 -295 7810 -265
rect 7755 -305 7810 -295
rect 7840 -265 7895 -255
rect 7840 -295 7850 -265
rect 7885 -295 7895 -265
rect 7840 -305 7895 -295
rect 7925 -265 7980 -255
rect 7925 -295 7935 -265
rect 7970 -295 7980 -265
rect 7925 -305 7980 -295
rect 8010 -265 8065 -255
rect 8010 -295 8020 -265
rect 8055 -295 8065 -265
rect 8010 -305 8065 -295
rect 8095 -265 8150 -255
rect 8095 -295 8105 -265
rect 8140 -295 8150 -265
rect 8095 -305 8150 -295
rect 8180 -265 8235 -255
rect 8180 -295 8190 -265
rect 8225 -295 8235 -265
rect 8180 -305 8235 -295
rect 8265 -265 8320 -255
rect 8265 -295 8275 -265
rect 8310 -295 8320 -265
rect 8265 -305 8320 -295
rect 8350 -265 8405 -255
rect 8350 -295 8360 -265
rect 8395 -295 8405 -265
rect 8350 -305 8405 -295
rect 8435 -265 8490 -255
rect 8435 -295 8445 -265
rect 8480 -295 8490 -265
rect 8435 -305 8490 -295
rect 8520 -265 8575 -255
rect 8520 -295 8530 -265
rect 8565 -295 8575 -265
rect 8520 -305 8575 -295
rect 8605 -265 8660 -255
rect 8605 -295 8615 -265
rect 8650 -295 8660 -265
rect 8605 -305 8660 -295
rect 8690 -265 8745 -255
rect 8690 -295 8700 -265
rect 8735 -295 8745 -265
rect 8690 -305 8745 -295
rect 8775 -265 8830 -255
rect 8775 -295 8785 -265
rect 8820 -295 8830 -265
rect 8775 -305 8830 -295
rect 8860 -265 8915 -255
rect 8860 -295 8870 -265
rect 8905 -295 8915 -265
rect 8860 -305 8915 -295
rect 8945 -265 9000 -255
rect 8945 -295 8955 -265
rect 8990 -295 9000 -265
rect 8945 -305 9000 -295
rect 9030 -265 9085 -255
rect 9030 -295 9040 -265
rect 9075 -295 9085 -265
rect 9030 -305 9085 -295
rect 9115 -265 9170 -255
rect 9115 -295 9125 -265
rect 9160 -295 9170 -265
rect 9115 -305 9170 -295
rect 9200 -265 9255 -255
rect 9200 -295 9210 -265
rect 9245 -295 9255 -265
rect 9200 -305 9255 -295
rect 9285 -265 9340 -255
rect 9285 -295 9295 -265
rect 9330 -295 9340 -265
rect 9285 -305 9340 -295
rect 9370 -265 9425 -255
rect 9370 -295 9380 -265
rect 9415 -295 9425 -265
rect 9370 -305 9425 -295
rect 9455 -265 9510 -255
rect 9455 -295 9465 -265
rect 9500 -295 9510 -265
rect 9455 -305 9510 -295
rect 9540 -265 9595 -255
rect 9540 -295 9550 -265
rect 9585 -295 9595 -265
rect 9540 -305 9595 -295
rect 9625 -265 9680 -255
rect 9625 -295 9635 -265
rect 9670 -295 9680 -265
rect 9625 -305 9680 -295
rect 9710 -265 9765 -255
rect 9710 -295 9720 -265
rect 9755 -295 9765 -265
rect 9710 -305 9765 -295
rect 9795 -265 9850 -255
rect 9795 -295 9805 -265
rect 9840 -295 9850 -265
rect 9795 -305 9850 -295
rect 9880 -265 9935 -255
rect 9880 -295 9890 -265
rect 9925 -295 9935 -265
rect 9880 -305 9935 -295
rect 9965 -265 10020 -255
rect 9965 -295 9975 -265
rect 10010 -295 10020 -265
rect 9965 -305 10020 -295
rect 10050 -265 10105 -255
rect 10050 -295 10060 -265
rect 10095 -295 10105 -265
rect 10050 -305 10105 -295
rect 10135 -265 10190 -255
rect 10135 -295 10145 -265
rect 10180 -295 10190 -265
rect 10135 -305 10190 -295
rect 10220 -265 10275 -255
rect 10220 -295 10230 -265
rect 10265 -295 10275 -265
rect 10220 -305 10275 -295
rect 10305 -265 10360 -255
rect 10305 -295 10315 -265
rect 10350 -295 10360 -265
rect 10305 -305 10360 -295
rect 10390 -265 10445 -255
rect 10390 -295 10400 -265
rect 10435 -295 10445 -265
rect 10390 -305 10445 -295
rect 10475 -265 10530 -255
rect 10475 -295 10485 -265
rect 10520 -295 10530 -265
rect 10475 -305 10530 -295
rect 10560 -265 10615 -255
rect 10560 -295 10570 -265
rect 10605 -295 10615 -265
rect 10560 -305 10615 -295
rect 10645 -265 10700 -255
rect 10645 -295 10655 -265
rect 10690 -295 10700 -265
rect 10645 -305 10700 -295
rect 10730 -265 10785 -255
rect 10730 -295 10740 -265
rect 10775 -295 10785 -265
rect 10730 -305 10785 -295
rect 10815 -265 10870 -255
rect 10815 -295 10825 -265
rect 10860 -295 10870 -265
rect 10815 -305 10870 -295
rect 10900 -265 10955 -255
rect 10900 -295 10910 -265
rect 10945 -295 10955 -265
rect 10900 -305 10955 -295
rect 10985 -265 11040 -255
rect 10985 -295 10995 -265
rect 11030 -295 11040 -265
rect 10985 -305 11040 -295
rect 11070 -265 11125 -255
rect 11070 -295 11080 -265
rect 11115 -295 11125 -265
rect 11070 -305 11125 -295
rect 11155 -265 11210 -255
rect 11155 -295 11165 -265
rect 11200 -295 11210 -265
rect 11155 -305 11210 -295
rect 11240 -265 11295 -255
rect 11240 -295 11250 -265
rect 11285 -295 11295 -265
rect 11240 -305 11295 -295
rect 11325 -265 11380 -255
rect 11325 -295 11335 -265
rect 11370 -295 11380 -265
rect 11325 -305 11380 -295
rect 11410 -265 11465 -255
rect 11410 -295 11420 -265
rect 11455 -295 11465 -265
rect 11410 -305 11465 -295
rect 11495 -265 11550 -255
rect 11495 -295 11505 -265
rect 11540 -295 11550 -265
rect 11495 -305 11550 -295
rect 11580 -265 11635 -255
rect 11580 -295 11590 -265
rect 11625 -295 11635 -265
rect 11580 -305 11635 -295
rect 11665 -265 11720 -255
rect 11665 -295 11675 -265
rect 11710 -295 11720 -265
rect 11665 -305 11720 -295
rect 11750 -265 11805 -255
rect 11750 -295 11760 -265
rect 11795 -295 11805 -265
rect 11750 -305 11805 -295
rect 11835 -265 11890 -255
rect 11835 -295 11845 -265
rect 11880 -295 11890 -265
rect 11835 -305 11890 -295
rect 11920 -265 11975 -255
rect 11920 -295 11930 -265
rect 11965 -295 11975 -265
rect 11920 -305 11975 -295
rect 12005 -265 12060 -255
rect 12005 -295 12015 -265
rect 12050 -295 12060 -265
rect 12005 -305 12060 -295
rect 12090 -265 12145 -255
rect 12090 -295 12100 -265
rect 12135 -295 12145 -265
rect 12090 -305 12145 -295
rect 12175 -265 12230 -255
rect 12175 -295 12185 -265
rect 12220 -295 12230 -265
rect 12175 -305 12230 -295
rect 12260 -265 12315 -255
rect 12260 -295 12270 -265
rect 12305 -295 12315 -265
rect 12260 -305 12315 -295
rect 12345 -265 12400 -255
rect 12345 -295 12355 -265
rect 12390 -295 12400 -265
rect 12345 -305 12400 -295
rect 12430 -265 12485 -255
rect 12430 -295 12440 -265
rect 12475 -295 12485 -265
rect 12430 -305 12485 -295
rect 12515 -265 12570 -255
rect 12515 -295 12525 -265
rect 12560 -295 12570 -265
rect 12515 -305 12570 -295
rect 12600 -265 12655 -255
rect 12600 -295 12610 -265
rect 12645 -295 12655 -265
rect 12600 -305 12655 -295
rect 12685 -265 12740 -255
rect 12685 -295 12695 -265
rect 12730 -295 12740 -265
rect 12685 -305 12740 -295
rect 12770 -265 12825 -255
rect 12770 -295 12780 -265
rect 12815 -295 12825 -265
rect 12770 -305 12825 -295
rect 12855 -265 12910 -255
rect 12855 -295 12865 -265
rect 12900 -295 12910 -265
rect 12855 -305 12910 -295
rect 12940 -265 12995 -255
rect 12940 -295 12950 -265
rect 12985 -295 12995 -265
rect 12940 -305 12995 -295
rect 13025 -265 13080 -255
rect 13025 -295 13035 -265
rect 13070 -295 13080 -265
rect 13025 -305 13080 -295
rect 13110 -265 13165 -255
rect 13110 -295 13120 -265
rect 13155 -295 13165 -265
rect 13110 -305 13165 -295
rect 13195 -265 13250 -255
rect 13195 -295 13205 -265
rect 13240 -295 13250 -265
rect 13195 -305 13250 -295
rect 13280 -265 13335 -255
rect 13280 -295 13290 -265
rect 13325 -295 13335 -265
rect 13280 -305 13335 -295
rect 13365 -265 13420 -255
rect 13365 -295 13375 -265
rect 13410 -295 13420 -265
rect 13365 -305 13420 -295
rect 13450 -265 13505 -255
rect 13450 -295 13460 -265
rect 13495 -295 13505 -265
rect 13450 -305 13505 -295
rect 13535 -265 13590 -255
rect 13535 -295 13545 -265
rect 13580 -295 13590 -265
rect 13535 -305 13590 -295
rect 13620 -265 13675 -255
rect 13620 -295 13630 -265
rect 13665 -295 13675 -265
rect 13620 -305 13675 -295
rect 13705 -265 13760 -255
rect 13705 -295 13715 -265
rect 13750 -295 13760 -265
rect 13705 -305 13760 -295
rect 13790 -265 13845 -255
rect 13790 -295 13800 -265
rect 13835 -295 13845 -265
rect 13790 -305 13845 -295
rect 13875 -265 13930 -255
rect 13875 -295 13885 -265
rect 13920 -295 13930 -265
rect 13875 -305 13930 -295
rect 13960 -265 14015 -255
rect 13960 -295 13970 -265
rect 14005 -295 14015 -265
rect 13960 -305 14015 -295
rect 14045 -265 14100 -255
rect 14045 -295 14055 -265
rect 14090 -295 14100 -265
rect 14045 -305 14100 -295
rect 14130 -265 14185 -255
rect 14130 -295 14140 -265
rect 14175 -295 14185 -265
rect 14130 -305 14185 -295
rect 14215 -265 14270 -255
rect 14215 -295 14225 -265
rect 14260 -295 14270 -265
rect 14215 -305 14270 -295
rect 14300 -265 14355 -255
rect 14300 -295 14310 -265
rect 14345 -295 14355 -265
rect 14300 -305 14355 -295
rect 14385 -265 14440 -255
rect 14385 -295 14395 -265
rect 14430 -295 14440 -265
rect 14385 -305 14440 -295
rect 14470 -265 14525 -255
rect 14470 -295 14480 -265
rect 14515 -295 14525 -265
rect 14470 -305 14525 -295
rect 14555 -265 14610 -255
rect 14555 -295 14565 -265
rect 14600 -295 14610 -265
rect 14555 -305 14610 -295
rect 14640 -265 14695 -255
rect 14640 -295 14650 -265
rect 14685 -295 14695 -265
rect 14640 -305 14695 -295
rect 14725 -265 14780 -255
rect 14725 -295 14735 -265
rect 14770 -295 14780 -265
rect 14725 -305 14780 -295
rect 14810 -265 14865 -255
rect 14810 -295 14820 -265
rect 14855 -295 14865 -265
rect 14810 -305 14865 -295
rect 14895 -265 14950 -255
rect 14895 -295 14905 -265
rect 14940 -295 14950 -265
rect 14895 -305 14950 -295
rect 14980 -265 15035 -255
rect 14980 -295 14990 -265
rect 15025 -295 15035 -265
rect 14980 -305 15035 -295
rect 15065 -265 15120 -255
rect 15065 -295 15075 -265
rect 15110 -295 15120 -265
rect 15065 -305 15120 -295
rect 15150 -265 15205 -255
rect 15150 -295 15160 -265
rect 15195 -295 15205 -265
rect 15150 -305 15205 -295
rect 15235 -265 15290 -255
rect 15235 -295 15245 -265
rect 15280 -295 15290 -265
rect 15235 -305 15290 -295
rect 15320 -265 15375 -255
rect 15320 -295 15330 -265
rect 15365 -295 15375 -265
rect 15320 -305 15375 -295
rect 15405 -265 15460 -255
rect 15405 -295 15415 -265
rect 15450 -295 15460 -265
rect 15405 -305 15460 -295
rect 15490 -265 15545 -255
rect 15490 -295 15500 -265
rect 15535 -295 15545 -265
rect 15490 -305 15545 -295
rect 15575 -265 15630 -255
rect 15575 -295 15585 -265
rect 15620 -295 15630 -265
rect 15575 -305 15630 -295
rect 15660 -265 15715 -255
rect 15660 -295 15670 -265
rect 15705 -295 15715 -265
rect 15660 -305 15715 -295
rect 15745 -265 15800 -255
rect 15745 -295 15755 -265
rect 15790 -295 15800 -265
rect 15745 -305 15800 -295
rect 15830 -265 15885 -255
rect 15830 -295 15840 -265
rect 15875 -295 15885 -265
rect 15830 -305 15885 -295
rect 15915 -265 15970 -255
rect 15915 -295 15925 -265
rect 15960 -295 15970 -265
rect 15915 -305 15970 -295
rect 16000 -265 16055 -255
rect 16000 -295 16010 -265
rect 16045 -295 16055 -265
rect 16000 -305 16055 -295
rect 16085 -265 16140 -255
rect 16085 -295 16095 -265
rect 16130 -295 16140 -265
rect 16085 -305 16140 -295
rect 16170 -265 16225 -255
rect 16170 -295 16180 -265
rect 16215 -295 16225 -265
rect 16170 -305 16225 -295
rect 16255 -265 16310 -255
rect 16255 -295 16265 -265
rect 16300 -295 16310 -265
rect 16255 -305 16310 -295
rect 16340 -265 16395 -255
rect 16340 -295 16350 -265
rect 16385 -295 16395 -265
rect 16340 -305 16395 -295
rect 16425 -265 16480 -255
rect 16425 -295 16435 -265
rect 16470 -295 16480 -265
rect 16425 -305 16480 -295
rect 16510 -265 16565 -255
rect 16510 -295 16520 -265
rect 16555 -295 16565 -265
rect 16510 -305 16565 -295
rect 16595 -265 16650 -255
rect 16595 -295 16605 -265
rect 16640 -295 16650 -265
rect 16595 -305 16650 -295
rect 16680 -265 16735 -255
rect 16680 -295 16690 -265
rect 16725 -295 16735 -265
rect 16680 -305 16735 -295
rect 16765 -265 16820 -255
rect 16765 -295 16775 -265
rect 16810 -295 16820 -265
rect 16765 -305 16820 -295
rect 16850 -265 16905 -255
rect 16850 -295 16860 -265
rect 16895 -295 16905 -265
rect 16850 -305 16905 -295
rect 16935 -265 16990 -255
rect 16935 -295 16945 -265
rect 16980 -295 16990 -265
rect 16935 -305 16990 -295
rect 17020 -265 17075 -255
rect 17020 -295 17030 -265
rect 17065 -295 17075 -265
rect 17020 -305 17075 -295
rect 17105 -265 17160 -255
rect 17105 -295 17115 -265
rect 17150 -295 17160 -265
rect 17105 -305 17160 -295
rect 17190 -265 17245 -255
rect 17190 -295 17200 -265
rect 17235 -295 17245 -265
rect 17190 -305 17245 -295
rect 17275 -265 17330 -255
rect 17275 -295 17285 -265
rect 17320 -295 17330 -265
rect 17275 -305 17330 -295
rect 17360 -265 17415 -255
rect 17360 -295 17370 -265
rect 17405 -295 17415 -265
rect 17360 -305 17415 -295
rect 17445 -265 17500 -255
rect 17445 -295 17455 -265
rect 17490 -295 17500 -265
rect 17445 -305 17500 -295
rect 17530 -265 17585 -255
rect 17530 -295 17540 -265
rect 17575 -295 17585 -265
rect 17530 -305 17585 -295
rect 17615 -265 17670 -255
rect 17615 -295 17625 -265
rect 17660 -295 17670 -265
rect 17615 -305 17670 -295
rect 17700 -265 17755 -255
rect 17700 -295 17710 -265
rect 17745 -295 17755 -265
rect 17700 -305 17755 -295
rect 17785 -265 17840 -255
rect 17785 -295 17795 -265
rect 17830 -295 17840 -265
rect 17785 -305 17840 -295
rect 17870 -265 17925 -255
rect 17870 -295 17880 -265
rect 17915 -295 17925 -265
rect 17870 -305 17925 -295
rect 17955 -265 18010 -255
rect 17955 -295 17965 -265
rect 18000 -295 18010 -265
rect 17955 -305 18010 -295
rect 18040 -265 18095 -255
rect 18040 -295 18050 -265
rect 18085 -295 18095 -265
rect 18040 -305 18095 -295
rect 18125 -265 18180 -255
rect 18125 -295 18135 -265
rect 18170 -295 18180 -265
rect 18125 -305 18180 -295
rect 18210 -265 18265 -255
rect 18210 -295 18220 -265
rect 18255 -295 18265 -265
rect 18210 -305 18265 -295
rect 18295 -265 18350 -255
rect 18295 -295 18305 -265
rect 18340 -295 18350 -265
rect 18295 -305 18350 -295
rect 18380 -265 18435 -255
rect 18380 -295 18390 -265
rect 18425 -295 18435 -265
rect 18380 -305 18435 -295
rect 18465 -265 18520 -255
rect 18465 -295 18475 -265
rect 18510 -295 18520 -265
rect 18465 -305 18520 -295
rect 18550 -265 18605 -255
rect 18550 -295 18560 -265
rect 18595 -295 18605 -265
rect 18550 -305 18605 -295
rect 18635 -265 18690 -255
rect 18635 -295 18645 -265
rect 18680 -295 18690 -265
rect 18635 -305 18690 -295
rect 18720 -265 18775 -255
rect 18720 -295 18730 -265
rect 18765 -295 18775 -265
rect 18720 -305 18775 -295
rect 18805 -265 18860 -255
rect 18805 -295 18815 -265
rect 18850 -295 18860 -265
rect 18805 -305 18860 -295
rect 18890 -265 18945 -255
rect 18890 -295 18900 -265
rect 18935 -295 18945 -265
rect 18890 -305 18945 -295
rect 18975 -265 19030 -255
rect 18975 -295 18985 -265
rect 19020 -295 19030 -265
rect 18975 -305 19030 -295
rect 19060 -265 19115 -255
rect 19060 -295 19070 -265
rect 19105 -295 19115 -265
rect 19060 -305 19115 -295
rect 19145 -265 19200 -255
rect 19145 -295 19155 -265
rect 19190 -295 19200 -265
rect 19145 -305 19200 -295
rect 19230 -265 19285 -255
rect 19230 -295 19240 -265
rect 19275 -295 19285 -265
rect 19230 -305 19285 -295
rect 19315 -265 19370 -255
rect 19315 -295 19325 -265
rect 19360 -295 19370 -265
rect 19315 -305 19370 -295
rect 19400 -265 19455 -255
rect 19400 -295 19410 -265
rect 19445 -295 19455 -265
rect 19400 -305 19455 -295
rect 19485 -265 19540 -255
rect 19485 -295 19495 -265
rect 19530 -295 19540 -265
rect 19485 -305 19540 -295
rect 19570 -265 19625 -255
rect 19570 -295 19580 -265
rect 19615 -295 19625 -265
rect 19570 -305 19625 -295
rect 19655 -265 19710 -255
rect 19655 -295 19665 -265
rect 19700 -295 19710 -265
rect 19655 -305 19710 -295
rect 19740 -265 19795 -255
rect 19740 -295 19750 -265
rect 19785 -295 19795 -265
rect 19740 -305 19795 -295
rect 19825 -265 19880 -255
rect 19825 -295 19835 -265
rect 19870 -295 19880 -265
rect 19825 -305 19880 -295
rect 19910 -265 19965 -255
rect 19910 -295 19920 -265
rect 19955 -295 19965 -265
rect 19910 -305 19965 -295
rect 19995 -265 20050 -255
rect 19995 -295 20005 -265
rect 20040 -295 20050 -265
rect 19995 -305 20050 -295
rect 20080 -265 20135 -255
rect 20080 -295 20090 -265
rect 20125 -295 20135 -265
rect 20080 -305 20135 -295
rect 20165 -265 20220 -255
rect 20165 -295 20175 -265
rect 20210 -295 20220 -265
rect 20165 -305 20220 -295
rect 20250 -265 20305 -255
rect 20250 -295 20260 -265
rect 20295 -295 20305 -265
rect 20250 -305 20305 -295
rect 20335 -265 20390 -255
rect 20335 -295 20345 -265
rect 20380 -295 20390 -265
rect 20335 -305 20390 -295
rect 20420 -265 20475 -255
rect 20420 -295 20430 -265
rect 20465 -295 20475 -265
rect 20420 -305 20475 -295
rect 20505 -265 20560 -255
rect 20505 -295 20515 -265
rect 20550 -295 20560 -265
rect 20505 -305 20560 -295
rect 20590 -265 20645 -255
rect 20590 -295 20600 -265
rect 20635 -295 20645 -265
rect 20590 -305 20645 -295
rect 20675 -265 20730 -255
rect 20675 -295 20685 -265
rect 20720 -295 20730 -265
rect 20675 -305 20730 -295
rect 20760 -265 20815 -255
rect 20760 -295 20770 -265
rect 20805 -295 20815 -265
rect 20760 -305 20815 -295
rect 20845 -265 20900 -255
rect 20845 -295 20855 -265
rect 20890 -295 20900 -265
rect 20845 -305 20900 -295
rect 20930 -265 20985 -255
rect 20930 -295 20940 -265
rect 20975 -295 20985 -265
rect 20930 -305 20985 -295
rect 21015 -265 21070 -255
rect 21015 -295 21025 -265
rect 21060 -295 21070 -265
rect 21015 -305 21070 -295
rect 21100 -265 21155 -255
rect 21100 -295 21110 -265
rect 21145 -295 21155 -265
rect 21100 -305 21155 -295
rect 21185 -265 21240 -255
rect 21185 -295 21195 -265
rect 21230 -295 21240 -265
rect 21185 -305 21240 -295
rect 21270 -265 21325 -255
rect 21270 -295 21280 -265
rect 21315 -295 21325 -265
rect 21270 -305 21325 -295
rect 21355 -265 21410 -255
rect 21355 -295 21365 -265
rect 21400 -295 21410 -265
rect 21355 -305 21410 -295
rect 21440 -265 21495 -255
rect 21440 -295 21450 -265
rect 21485 -295 21495 -265
rect 21440 -305 21495 -295
rect 21525 -265 21580 -255
rect 21525 -295 21535 -265
rect 21570 -295 21580 -265
rect 21525 -305 21580 -295
rect 21610 -265 21665 -255
rect 21610 -295 21620 -265
rect 21655 -295 21665 -265
rect 21610 -305 21665 -295
rect 21695 -265 21750 -255
rect 21695 -295 21705 -265
rect 21740 -295 21750 -265
rect 21695 -305 21750 -295
rect 21780 -265 21835 -255
rect 21780 -295 21790 -265
rect 21825 -295 21835 -265
rect 21780 -305 21835 -295
rect 21865 -265 21920 -255
rect 21865 -295 21875 -265
rect 21910 -295 21920 -265
rect 21865 -305 21920 -295
rect 21950 -265 22005 -255
rect 21950 -295 21960 -265
rect 21995 -295 22005 -265
rect 21950 -305 22005 -295
rect 22035 -265 22090 -255
rect 22035 -295 22045 -265
rect 22080 -295 22090 -265
rect 22035 -305 22090 -295
rect 22120 -265 22175 -255
rect 22120 -295 22130 -265
rect 22165 -295 22175 -265
rect 22120 -305 22175 -295
rect 22205 -265 22260 -255
rect 22205 -295 22215 -265
rect 22250 -295 22260 -265
rect 22205 -305 22260 -295
rect 22290 -265 22345 -255
rect 22290 -295 22300 -265
rect 22335 -295 22345 -265
rect 22290 -305 22345 -295
rect 22375 -265 22430 -255
rect 22375 -295 22385 -265
rect 22420 -295 22430 -265
rect 22375 -305 22430 -295
rect 22460 -265 22515 -255
rect 22460 -295 22470 -265
rect 22505 -295 22515 -265
rect 22460 -305 22515 -295
rect 22545 -265 22600 -255
rect 22545 -295 22555 -265
rect 22590 -295 22600 -265
rect 22545 -305 22600 -295
rect 22630 -265 22685 -255
rect 22630 -295 22640 -265
rect 22675 -295 22685 -265
rect 22630 -305 22685 -295
rect 22715 -265 22770 -255
rect 22715 -295 22725 -265
rect 22760 -295 22770 -265
rect 22715 -305 22770 -295
rect 22800 -265 22855 -255
rect 22800 -295 22810 -265
rect 22845 -295 22855 -265
rect 22800 -305 22855 -295
rect 22885 -265 22940 -255
rect 22885 -295 22895 -265
rect 22930 -295 22940 -265
rect 22885 -305 22940 -295
rect 22970 -265 23025 -255
rect 22970 -295 22980 -265
rect 23015 -295 23025 -265
rect 22970 -305 23025 -295
rect 23055 -265 23110 -255
rect 23055 -295 23065 -265
rect 23100 -295 23110 -265
rect 23055 -305 23110 -295
rect 23140 -265 23195 -255
rect 23140 -295 23150 -265
rect 23185 -295 23195 -265
rect 23140 -305 23195 -295
rect 23225 -265 23280 -255
rect 23225 -295 23235 -265
rect 23270 -295 23280 -265
rect 23225 -305 23280 -295
rect 23310 -265 23365 -255
rect 23310 -295 23320 -265
rect 23355 -295 23365 -265
rect 23310 -305 23365 -295
rect 23395 -265 23450 -255
rect 23395 -295 23405 -265
rect 23440 -295 23450 -265
rect 23395 -305 23450 -295
rect 23480 -265 23535 -255
rect 23480 -295 23490 -265
rect 23525 -295 23535 -265
rect 23480 -305 23535 -295
rect 23565 -265 23620 -255
rect 23565 -295 23575 -265
rect 23610 -295 23620 -265
rect 23565 -305 23620 -295
rect 23650 -265 23705 -255
rect 23650 -295 23660 -265
rect 23695 -295 23705 -265
rect 23650 -305 23705 -295
rect 23735 -265 23790 -255
rect 23735 -295 23745 -265
rect 23780 -295 23790 -265
rect 23735 -305 23790 -295
rect 23820 -265 23875 -255
rect 23820 -295 23830 -265
rect 23865 -295 23875 -265
rect 23820 -305 23875 -295
rect 23905 -265 23960 -255
rect 23905 -295 23915 -265
rect 23950 -295 23960 -265
rect 23905 -305 23960 -295
rect 23990 -265 24045 -255
rect 23990 -295 24000 -265
rect 24035 -295 24045 -265
rect 23990 -305 24045 -295
rect 24075 -265 24130 -255
rect 24075 -295 24085 -265
rect 24120 -295 24130 -265
rect 24075 -305 24130 -295
rect 24160 -265 24215 -255
rect 24160 -295 24170 -265
rect 24205 -295 24215 -265
rect 24160 -305 24215 -295
rect 24245 -265 24300 -255
rect 24245 -295 24255 -265
rect 24290 -295 24300 -265
rect 24245 -305 24300 -295
rect 24330 -265 24385 -255
rect 24330 -295 24340 -265
rect 24375 -295 24385 -265
rect 24330 -305 24385 -295
rect 24415 -265 24470 -255
rect 24415 -295 24425 -265
rect 24460 -295 24470 -265
rect 24415 -305 24470 -295
rect 24500 -265 24555 -255
rect 24500 -295 24510 -265
rect 24545 -295 24555 -265
rect 24500 -305 24555 -295
rect 24585 -265 24640 -255
rect 24585 -295 24595 -265
rect 24630 -295 24640 -265
rect 24585 -305 24640 -295
rect 24670 -265 24725 -255
rect 24670 -295 24680 -265
rect 24715 -295 24725 -265
rect 24670 -305 24725 -295
rect 24755 -265 24810 -255
rect 24755 -295 24765 -265
rect 24800 -295 24810 -265
rect 24755 -305 24810 -295
rect 24840 -265 24895 -255
rect 24840 -295 24850 -265
rect 24885 -295 24895 -265
rect 24840 -305 24895 -295
rect 24925 -265 24980 -255
rect 24925 -295 24935 -265
rect 24970 -295 24980 -265
rect 24925 -305 24980 -295
rect 25010 -265 25065 -255
rect 25010 -295 25020 -265
rect 25055 -295 25065 -265
rect 25010 -305 25065 -295
rect 25095 -265 25150 -255
rect 25095 -295 25105 -265
rect 25140 -295 25150 -265
rect 25095 -305 25150 -295
rect 25180 -265 25235 -255
rect 25180 -295 25190 -265
rect 25225 -295 25235 -265
rect 25180 -305 25235 -295
rect 25265 -265 25320 -255
rect 25265 -295 25275 -265
rect 25310 -295 25320 -265
rect 25265 -305 25320 -295
rect 25350 -265 25405 -255
rect 25350 -295 25360 -265
rect 25395 -295 25405 -265
rect 25350 -305 25405 -295
rect 25435 -265 25490 -255
rect 25435 -295 25445 -265
rect 25480 -295 25490 -265
rect 25435 -305 25490 -295
rect 25520 -265 25575 -255
rect 25520 -295 25530 -265
rect 25565 -295 25575 -265
rect 25520 -305 25575 -295
rect 25605 -265 25660 -255
rect 25605 -295 25615 -265
rect 25650 -295 25660 -265
rect 25605 -305 25660 -295
rect 25690 -265 25745 -255
rect 25690 -295 25700 -265
rect 25735 -295 25745 -265
rect 25690 -305 25745 -295
rect 25775 -265 25830 -255
rect 25775 -295 25785 -265
rect 25820 -295 25830 -265
rect 25775 -305 25830 -295
rect 25860 -265 25915 -255
rect 25860 -295 25870 -265
rect 25905 -295 25915 -265
rect 25860 -305 25915 -295
rect 25945 -265 26000 -255
rect 25945 -295 25955 -265
rect 25990 -295 26000 -265
rect 25945 -305 26000 -295
rect 26030 -265 26085 -255
rect 26030 -295 26040 -265
rect 26075 -295 26085 -265
rect 26030 -305 26085 -295
rect 26115 -265 26170 -255
rect 26115 -295 26125 -265
rect 26160 -295 26170 -265
rect 26115 -305 26170 -295
rect 26200 -265 26255 -255
rect 26200 -295 26210 -265
rect 26245 -295 26255 -265
rect 26200 -305 26255 -295
rect 26285 -265 26340 -255
rect 26285 -295 26295 -265
rect 26330 -295 26340 -265
rect 26285 -305 26340 -295
rect 26370 -265 26425 -255
rect 26370 -295 26380 -265
rect 26415 -295 26425 -265
rect 26370 -305 26425 -295
rect 26455 -265 26510 -255
rect 26455 -295 26465 -265
rect 26500 -295 26510 -265
rect 26455 -305 26510 -295
rect 26540 -265 26595 -255
rect 26540 -295 26550 -265
rect 26585 -295 26595 -265
rect 26540 -305 26595 -295
rect 26625 -265 26680 -255
rect 26625 -295 26635 -265
rect 26670 -295 26680 -265
rect 26625 -305 26680 -295
rect 26710 -265 26765 -255
rect 26710 -295 26720 -265
rect 26755 -295 26765 -265
rect 26710 -305 26765 -295
rect 26795 -265 26850 -255
rect 26795 -295 26805 -265
rect 26840 -295 26850 -265
rect 26795 -305 26850 -295
rect 26880 -265 26935 -255
rect 26880 -295 26890 -265
rect 26925 -295 26935 -265
rect 26880 -305 26935 -295
rect 26965 -265 27020 -255
rect 26965 -295 26975 -265
rect 27010 -295 27020 -265
rect 26965 -305 27020 -295
rect 27050 -265 27105 -255
rect 27050 -295 27060 -265
rect 27095 -295 27105 -265
rect 27050 -305 27105 -295
rect 27135 -265 27190 -255
rect 27135 -295 27145 -265
rect 27180 -295 27190 -265
rect 27135 -305 27190 -295
rect 27220 -265 27275 -255
rect 27220 -295 27230 -265
rect 27265 -295 27275 -265
rect 27220 -305 27275 -295
rect 27305 -265 27360 -255
rect 27305 -295 27315 -265
rect 27350 -295 27360 -265
rect 27305 -305 27360 -295
rect 27390 -265 27445 -255
rect 27390 -295 27400 -265
rect 27435 -295 27445 -265
rect 27390 -305 27445 -295
rect 27475 -265 27530 -255
rect 27475 -295 27485 -265
rect 27520 -295 27530 -265
rect 27475 -305 27530 -295
rect 27560 -265 27615 -255
rect 27560 -295 27570 -265
rect 27605 -295 27615 -265
rect 27560 -305 27615 -295
rect 27645 -265 27700 -255
rect 27645 -295 27655 -265
rect 27690 -295 27700 -265
rect 27645 -305 27700 -295
rect 27730 -265 27785 -255
rect 27730 -295 27740 -265
rect 27775 -295 27785 -265
rect 27730 -305 27785 -295
rect 27815 -265 27870 -255
rect 27815 -295 27825 -265
rect 27860 -295 27870 -265
rect 27815 -305 27870 -295
rect 27900 -265 27955 -255
rect 27900 -295 27910 -265
rect 27945 -295 27955 -265
rect 27900 -305 27955 -295
rect 27985 -265 28040 -255
rect 27985 -295 27995 -265
rect 28030 -295 28040 -265
rect 27985 -305 28040 -295
rect 28070 -265 28125 -255
rect 28070 -295 28080 -265
rect 28115 -295 28125 -265
rect 28070 -305 28125 -295
rect 28155 -265 28210 -255
rect 28155 -295 28165 -265
rect 28200 -295 28210 -265
rect 28155 -305 28210 -295
rect 28240 -265 28295 -255
rect 28240 -295 28250 -265
rect 28285 -295 28295 -265
rect 28240 -305 28295 -295
rect 28325 -265 28380 -255
rect 28325 -295 28335 -265
rect 28370 -295 28380 -265
rect 28325 -305 28380 -295
rect 28410 -265 28465 -255
rect 28410 -295 28420 -265
rect 28455 -295 28465 -265
rect 28410 -305 28465 -295
rect 28495 -265 28550 -255
rect 28495 -295 28505 -265
rect 28540 -295 28550 -265
rect 28495 -305 28550 -295
rect 28580 -265 28635 -255
rect 28580 -295 28590 -265
rect 28625 -295 28635 -265
rect 28580 -305 28635 -295
rect 28665 -265 28720 -255
rect 28665 -295 28675 -265
rect 28710 -295 28720 -265
rect 28665 -305 28720 -295
rect 28750 -265 28805 -255
rect 28750 -295 28760 -265
rect 28795 -295 28805 -265
rect 28750 -305 28805 -295
rect 28835 -265 28890 -255
rect 28835 -295 28845 -265
rect 28880 -295 28890 -265
rect 28835 -305 28890 -295
rect 28920 -265 28975 -255
rect 28920 -295 28930 -265
rect 28965 -295 28975 -265
rect 28920 -305 28975 -295
rect 29005 -265 29060 -255
rect 29005 -295 29015 -265
rect 29050 -295 29060 -265
rect 29005 -305 29060 -295
rect 29090 -265 29145 -255
rect 29090 -295 29100 -265
rect 29135 -295 29145 -265
rect 29090 -305 29145 -295
rect 29175 -265 29230 -255
rect 29175 -295 29185 -265
rect 29220 -295 29230 -265
rect 29175 -305 29230 -295
rect 29260 -265 29315 -255
rect 29260 -295 29270 -265
rect 29305 -295 29315 -265
rect 29260 -305 29315 -295
rect 29345 -265 29400 -255
rect 29345 -295 29355 -265
rect 29390 -295 29400 -265
rect 29345 -305 29400 -295
rect 29430 -265 29485 -255
rect 29430 -295 29440 -265
rect 29475 -295 29485 -265
rect 29430 -305 29485 -295
rect 29515 -265 29570 -255
rect 29515 -295 29525 -265
rect 29560 -295 29570 -265
rect 29515 -305 29570 -295
rect 29600 -265 29655 -255
rect 29600 -295 29610 -265
rect 29645 -295 29655 -265
rect 29600 -305 29655 -295
rect 29685 -265 29740 -255
rect 29685 -295 29695 -265
rect 29730 -295 29740 -265
rect 29685 -305 29740 -295
rect 29770 -265 29825 -255
rect 29770 -295 29780 -265
rect 29815 -295 29825 -265
rect 29770 -305 29825 -295
rect 29855 -265 29910 -255
rect 29855 -295 29865 -265
rect 29900 -295 29910 -265
rect 29855 -305 29910 -295
rect 29940 -265 29995 -255
rect 29940 -295 29950 -265
rect 29985 -295 29995 -265
rect 29940 -305 29995 -295
rect 30025 -265 30080 -255
rect 30025 -295 30035 -265
rect 30070 -295 30080 -265
rect 30025 -305 30080 -295
rect 30110 -265 30165 -255
rect 30110 -295 30120 -265
rect 30155 -295 30165 -265
rect 30110 -305 30165 -295
rect 30195 -265 30250 -255
rect 30195 -295 30205 -265
rect 30240 -295 30250 -265
rect 30195 -305 30250 -295
rect 30280 -265 30335 -255
rect 30280 -295 30290 -265
rect 30325 -295 30335 -265
rect 30280 -305 30335 -295
rect 30365 -265 30420 -255
rect 30365 -295 30375 -265
rect 30410 -295 30420 -265
rect 30365 -305 30420 -295
rect 30450 -265 30505 -255
rect 30450 -295 30460 -265
rect 30495 -295 30505 -265
rect 30450 -305 30505 -295
rect 30535 -265 30590 -255
rect 30535 -295 30545 -265
rect 30580 -295 30590 -265
rect 30535 -305 30590 -295
rect 30620 -265 30675 -255
rect 30620 -295 30630 -265
rect 30665 -295 30675 -265
rect 30620 -305 30675 -295
rect 30705 -265 30760 -255
rect 30705 -295 30715 -265
rect 30750 -295 30760 -265
rect 30705 -305 30760 -295
rect 30790 -265 30845 -255
rect 30790 -295 30800 -265
rect 30835 -295 30845 -265
rect 30790 -305 30845 -295
rect 30875 -265 30930 -255
rect 30875 -295 30885 -265
rect 30920 -295 30930 -265
rect 30875 -305 30930 -295
rect 30960 -265 31015 -255
rect 30960 -295 30970 -265
rect 31005 -295 31015 -265
rect 30960 -305 31015 -295
rect 31045 -265 31100 -255
rect 31045 -295 31055 -265
rect 31090 -295 31100 -265
rect 31045 -305 31100 -295
rect 31130 -265 31185 -255
rect 31130 -295 31140 -265
rect 31175 -295 31185 -265
rect 31130 -305 31185 -295
rect 31215 -265 31270 -255
rect 31215 -295 31225 -265
rect 31260 -295 31270 -265
rect 31215 -305 31270 -295
rect 31300 -265 31355 -255
rect 31300 -295 31310 -265
rect 31345 -295 31355 -265
rect 31300 -305 31355 -295
rect 31385 -265 31440 -255
rect 31385 -295 31395 -265
rect 31430 -295 31440 -265
rect 31385 -305 31440 -295
rect 31470 -265 31525 -255
rect 31470 -295 31480 -265
rect 31515 -295 31525 -265
rect 31470 -305 31525 -295
rect 31555 -265 31610 -255
rect 31555 -295 31565 -265
rect 31600 -295 31610 -265
rect 31555 -305 31610 -295
rect 31640 -265 31695 -255
rect 31640 -295 31650 -265
rect 31685 -295 31695 -265
rect 31640 -305 31695 -295
rect 31725 -265 31780 -255
rect 31725 -295 31735 -265
rect 31770 -295 31780 -265
rect 31725 -305 31780 -295
rect 31810 -265 31865 -255
rect 31810 -295 31820 -265
rect 31855 -295 31865 -265
rect 31810 -305 31865 -295
rect 31895 -265 31950 -255
rect 31895 -295 31905 -265
rect 31940 -295 31950 -265
rect 31895 -305 31950 -295
rect 31980 -265 32035 -255
rect 31980 -295 31990 -265
rect 32025 -295 32035 -265
rect 31980 -305 32035 -295
rect 32065 -265 32120 -255
rect 32065 -295 32075 -265
rect 32110 -295 32120 -265
rect 32065 -305 32120 -295
rect 32150 -265 32205 -255
rect 32150 -295 32160 -265
rect 32195 -295 32205 -265
rect 32150 -305 32205 -295
rect 32235 -265 32290 -255
rect 32235 -295 32245 -265
rect 32280 -295 32290 -265
rect 32235 -305 32290 -295
rect 32320 -265 32375 -255
rect 32320 -295 32330 -265
rect 32365 -295 32375 -265
rect 32320 -305 32375 -295
rect 32405 -265 32460 -255
rect 32405 -295 32415 -265
rect 32450 -295 32460 -265
rect 32405 -305 32460 -295
rect 32490 -265 32545 -255
rect 32490 -295 32500 -265
rect 32535 -295 32545 -265
rect 32490 -305 32545 -295
rect 32575 -265 32630 -255
rect 32575 -295 32585 -265
rect 32620 -295 32630 -265
rect 32575 -305 32630 -295
rect 32660 -265 32715 -255
rect 32660 -295 32670 -265
rect 32705 -295 32715 -265
rect 32660 -305 32715 -295
rect 32745 -265 32800 -255
rect 32745 -295 32755 -265
rect 32790 -295 32800 -265
rect 32745 -305 32800 -295
rect 32830 -265 32885 -255
rect 32830 -295 32840 -265
rect 32875 -295 32885 -265
rect 32830 -305 32885 -295
rect 32915 -265 32970 -255
rect 32915 -295 32925 -265
rect 32960 -295 32970 -265
rect 32915 -305 32970 -295
rect 33000 -265 33055 -255
rect 33000 -295 33010 -265
rect 33045 -295 33055 -265
rect 33000 -305 33055 -295
rect 33085 -265 33140 -255
rect 33085 -295 33095 -265
rect 33130 -295 33140 -265
rect 33085 -305 33140 -295
rect 33170 -265 33225 -255
rect 33170 -295 33180 -265
rect 33215 -295 33225 -265
rect 33170 -305 33225 -295
rect 33255 -265 33310 -255
rect 33255 -295 33265 -265
rect 33300 -295 33310 -265
rect 33255 -305 33310 -295
rect 33340 -265 33395 -255
rect 33340 -295 33350 -265
rect 33385 -295 33395 -265
rect 33340 -305 33395 -295
rect 33425 -265 33480 -255
rect 33425 -295 33435 -265
rect 33470 -295 33480 -265
rect 33425 -305 33480 -295
rect 33510 -265 33565 -255
rect 33510 -295 33520 -265
rect 33555 -295 33565 -265
rect 33510 -305 33565 -295
rect 33595 -265 33650 -255
rect 33595 -295 33605 -265
rect 33640 -295 33650 -265
rect 33595 -305 33650 -295
rect 33680 -265 33735 -255
rect 33680 -295 33690 -265
rect 33725 -295 33735 -265
rect 33680 -305 33735 -295
rect 33765 -265 33820 -255
rect 33765 -295 33775 -265
rect 33810 -295 33820 -265
rect 33765 -305 33820 -295
rect 33850 -265 33905 -255
rect 33850 -295 33860 -265
rect 33895 -295 33905 -265
rect 33850 -305 33905 -295
rect 33935 -265 33990 -255
rect 33935 -295 33945 -265
rect 33980 -295 33990 -265
rect 33935 -305 33990 -295
rect 34020 -265 34075 -255
rect 34020 -295 34030 -265
rect 34065 -295 34075 -265
rect 34020 -305 34075 -295
rect 34105 -265 34160 -255
rect 34105 -295 34115 -265
rect 34150 -295 34160 -265
rect 34105 -305 34160 -295
rect 34190 -265 34245 -255
rect 34190 -295 34200 -265
rect 34235 -295 34245 -265
rect 34190 -305 34245 -295
rect 34275 -265 34330 -255
rect 34275 -295 34285 -265
rect 34320 -295 34330 -265
rect 34275 -305 34330 -295
rect 34360 -265 34415 -255
rect 34360 -295 34370 -265
rect 34405 -295 34415 -265
rect 34360 -305 34415 -295
rect 34445 -265 34500 -255
rect 34445 -295 34455 -265
rect 34490 -295 34500 -265
rect 34445 -305 34500 -295
rect 34530 -265 34585 -255
rect 34530 -295 34540 -265
rect 34575 -295 34585 -265
rect 34530 -305 34585 -295
rect 34615 -265 34670 -255
rect 34615 -295 34625 -265
rect 34660 -295 34670 -265
rect 34615 -305 34670 -295
rect 34700 -265 34755 -255
rect 34700 -295 34710 -265
rect 34745 -295 34755 -265
rect 34700 -305 34755 -295
rect 34785 -265 34840 -255
rect 34785 -295 34795 -265
rect 34830 -295 34840 -265
rect 34785 -305 34840 -295
rect 34870 -265 34925 -255
rect 34870 -295 34880 -265
rect 34915 -295 34925 -265
rect 34870 -305 34925 -295
rect 34955 -265 35010 -255
rect 34955 -295 34965 -265
rect 35000 -295 35010 -265
rect 34955 -305 35010 -295
rect 35040 -265 35095 -255
rect 35040 -295 35050 -265
rect 35085 -295 35095 -265
rect 35040 -305 35095 -295
rect 35125 -265 35180 -255
rect 35125 -295 35135 -265
rect 35170 -295 35180 -265
rect 35125 -305 35180 -295
rect 35210 -265 35265 -255
rect 35210 -295 35220 -265
rect 35255 -295 35265 -265
rect 35210 -305 35265 -295
rect 35295 -265 35350 -255
rect 35295 -295 35305 -265
rect 35340 -295 35350 -265
rect 35295 -305 35350 -295
rect 35380 -265 35435 -255
rect 35380 -295 35390 -265
rect 35425 -295 35435 -265
rect 35380 -305 35435 -295
rect 35465 -265 35520 -255
rect 35465 -295 35475 -265
rect 35510 -295 35520 -265
rect 35465 -305 35520 -295
rect 35550 -265 35605 -255
rect 35550 -295 35560 -265
rect 35595 -295 35605 -265
rect 35550 -305 35605 -295
rect 35635 -265 35690 -255
rect 35635 -295 35645 -265
rect 35680 -295 35690 -265
rect 35635 -305 35690 -295
rect 35720 -265 35775 -255
rect 35720 -295 35730 -265
rect 35765 -295 35775 -265
rect 35720 -305 35775 -295
rect 35805 -265 35860 -255
rect 35805 -295 35815 -265
rect 35850 -295 35860 -265
rect 35805 -305 35860 -295
rect 35890 -265 35945 -255
rect 35890 -295 35900 -265
rect 35935 -295 35945 -265
rect 35890 -305 35945 -295
rect 35975 -265 36030 -255
rect 35975 -295 35985 -265
rect 36020 -295 36030 -265
rect 35975 -305 36030 -295
rect 36060 -265 36115 -255
rect 36060 -295 36070 -265
rect 36105 -295 36115 -265
rect 36060 -305 36115 -295
rect 36145 -265 36200 -255
rect 36145 -295 36155 -265
rect 36190 -295 36200 -265
rect 36145 -305 36200 -295
rect 36230 -265 36285 -255
rect 36230 -295 36240 -265
rect 36275 -295 36285 -265
rect 36230 -305 36285 -295
rect 36315 -265 36370 -255
rect 36315 -295 36325 -265
rect 36360 -295 36370 -265
rect 36315 -305 36370 -295
rect 36400 -265 36455 -255
rect 36400 -295 36410 -265
rect 36445 -295 36455 -265
rect 36400 -305 36455 -295
rect 36485 -265 36540 -255
rect 36485 -295 36495 -265
rect 36530 -295 36540 -265
rect 36485 -305 36540 -295
rect 36570 -265 36625 -255
rect 36570 -295 36580 -265
rect 36615 -295 36625 -265
rect 36570 -305 36625 -295
rect 36655 -265 36710 -255
rect 36655 -295 36665 -265
rect 36700 -295 36710 -265
rect 36655 -305 36710 -295
rect 36740 -265 36795 -255
rect 36740 -295 36750 -265
rect 36785 -295 36795 -265
rect 36740 -305 36795 -295
rect 36825 -265 36880 -255
rect 36825 -295 36835 -265
rect 36870 -295 36880 -265
rect 36825 -305 36880 -295
rect 36910 -265 36965 -255
rect 36910 -295 36920 -265
rect 36955 -295 36965 -265
rect 36910 -305 36965 -295
rect 36995 -265 37050 -255
rect 36995 -295 37005 -265
rect 37040 -295 37050 -265
rect 36995 -305 37050 -295
rect 37080 -265 37135 -255
rect 37080 -295 37090 -265
rect 37125 -295 37135 -265
rect 37080 -305 37135 -295
rect 37165 -265 37220 -255
rect 37165 -295 37175 -265
rect 37210 -295 37220 -265
rect 37165 -305 37220 -295
rect 37250 -265 37305 -255
rect 37250 -295 37260 -265
rect 37295 -295 37305 -265
rect 37250 -305 37305 -295
rect 37335 -265 37390 -255
rect 37335 -295 37345 -265
rect 37380 -295 37390 -265
rect 37335 -305 37390 -295
rect 37420 -265 37475 -255
rect 37420 -295 37430 -265
rect 37465 -295 37475 -265
rect 37420 -305 37475 -295
rect 37505 -265 37560 -255
rect 37505 -295 37515 -265
rect 37550 -295 37560 -265
rect 37505 -305 37560 -295
rect 37590 -265 37645 -255
rect 37590 -295 37600 -265
rect 37635 -295 37645 -265
rect 37590 -305 37645 -295
rect 37675 -265 37730 -255
rect 37675 -295 37685 -265
rect 37720 -295 37730 -265
rect 37675 -305 37730 -295
rect 37760 -265 37815 -255
rect 37760 -295 37770 -265
rect 37805 -295 37815 -265
rect 37760 -305 37815 -295
rect 37845 -265 37900 -255
rect 37845 -295 37855 -265
rect 37890 -295 37900 -265
rect 37845 -305 37900 -295
rect 37930 -265 37985 -255
rect 37930 -295 37940 -265
rect 37975 -295 37985 -265
rect 37930 -305 37985 -295
rect 38015 -265 38070 -255
rect 38015 -295 38025 -265
rect 38060 -295 38070 -265
rect 38015 -305 38070 -295
rect 38100 -265 38155 -255
rect 38100 -295 38110 -265
rect 38145 -295 38155 -265
rect 38100 -305 38155 -295
rect 38185 -265 38240 -255
rect 38185 -295 38195 -265
rect 38230 -295 38240 -265
rect 38185 -305 38240 -295
rect 38270 -265 38325 -255
rect 38270 -295 38280 -265
rect 38315 -295 38325 -265
rect 38270 -305 38325 -295
rect 38355 -265 38410 -255
rect 38355 -295 38365 -265
rect 38400 -295 38410 -265
rect 38355 -305 38410 -295
rect 38440 -265 38495 -255
rect 38440 -295 38450 -265
rect 38485 -295 38495 -265
rect 38440 -305 38495 -295
rect 38525 -265 38580 -255
rect 38525 -295 38535 -265
rect 38570 -295 38580 -265
rect 38525 -305 38580 -295
rect 38610 -265 38665 -255
rect 38610 -295 38620 -265
rect 38655 -295 38665 -265
rect 38610 -305 38665 -295
rect 38695 -265 38750 -255
rect 38695 -295 38705 -265
rect 38740 -295 38750 -265
rect 38695 -305 38750 -295
rect 38780 -265 38835 -255
rect 38780 -295 38790 -265
rect 38825 -295 38835 -265
rect 38780 -305 38835 -295
rect 38865 -265 38920 -255
rect 38865 -295 38875 -265
rect 38910 -295 38920 -265
rect 38865 -305 38920 -295
rect 38950 -265 39005 -255
rect 38950 -295 38960 -265
rect 38995 -295 39005 -265
rect 38950 -305 39005 -295
rect 39035 -265 39090 -255
rect 39035 -295 39045 -265
rect 39080 -295 39090 -265
rect 39035 -305 39090 -295
rect 39120 -265 39175 -255
rect 39120 -295 39130 -265
rect 39165 -295 39175 -265
rect 39120 -305 39175 -295
rect 39205 -265 39260 -255
rect 39205 -295 39215 -265
rect 39250 -295 39260 -265
rect 39205 -305 39260 -295
rect 39290 -265 39345 -255
rect 39290 -295 39300 -265
rect 39335 -295 39345 -265
rect 39290 -305 39345 -295
rect 39375 -265 39430 -255
rect 39375 -295 39385 -265
rect 39420 -295 39430 -265
rect 39375 -305 39430 -295
rect 39460 -265 39515 -255
rect 39460 -295 39470 -265
rect 39505 -295 39515 -265
rect 39460 -305 39515 -295
rect 39545 -265 39600 -255
rect 39545 -295 39555 -265
rect 39590 -295 39600 -265
rect 39545 -305 39600 -295
rect 39630 -265 39685 -255
rect 39630 -295 39640 -265
rect 39675 -295 39685 -265
rect 39630 -305 39685 -295
rect 39715 -265 39770 -255
rect 39715 -295 39725 -265
rect 39760 -295 39770 -265
rect 39715 -305 39770 -295
rect 39800 -265 39855 -255
rect 39800 -295 39810 -265
rect 39845 -295 39855 -265
rect 39800 -305 39855 -295
rect 39885 -265 39940 -255
rect 39885 -295 39895 -265
rect 39930 -295 39940 -265
rect 39885 -305 39940 -295
rect 39970 -265 40025 -255
rect 39970 -295 39980 -265
rect 40015 -295 40025 -265
rect 39970 -305 40025 -295
rect 40055 -265 40110 -255
rect 40055 -295 40065 -265
rect 40100 -295 40110 -265
rect 40055 -305 40110 -295
rect 40140 -265 40195 -255
rect 40140 -295 40150 -265
rect 40185 -295 40195 -265
rect 40140 -305 40195 -295
rect 40225 -265 40280 -255
rect 40225 -295 40235 -265
rect 40270 -295 40280 -265
rect 40225 -305 40280 -295
rect 40310 -265 40365 -255
rect 40310 -295 40320 -265
rect 40355 -295 40365 -265
rect 40310 -305 40365 -295
rect 40395 -265 40450 -255
rect 40395 -295 40405 -265
rect 40440 -295 40450 -265
rect 40395 -305 40450 -295
rect 40480 -265 40535 -255
rect 40480 -295 40490 -265
rect 40525 -295 40535 -265
rect 40480 -305 40535 -295
rect 40565 -265 40620 -255
rect 40565 -295 40575 -265
rect 40610 -295 40620 -265
rect 40565 -305 40620 -295
rect 40650 -265 40705 -255
rect 40650 -295 40660 -265
rect 40695 -295 40705 -265
rect 40650 -305 40705 -295
rect 40735 -265 40790 -255
rect 40735 -295 40745 -265
rect 40780 -295 40790 -265
rect 40735 -305 40790 -295
rect 40820 -265 40875 -255
rect 40820 -295 40830 -265
rect 40865 -295 40875 -265
rect 40820 -305 40875 -295
rect 40905 -265 40960 -255
rect 40905 -295 40915 -265
rect 40950 -295 40960 -265
rect 40905 -305 40960 -295
rect 40990 -265 41045 -255
rect 40990 -295 41000 -265
rect 41035 -295 41045 -265
rect 40990 -305 41045 -295
rect 41075 -265 41130 -255
rect 41075 -295 41085 -265
rect 41120 -295 41130 -265
rect 41075 -305 41130 -295
rect 41160 -265 41215 -255
rect 41160 -295 41170 -265
rect 41205 -295 41215 -265
rect 41160 -305 41215 -295
rect 41245 -265 41300 -255
rect 41245 -295 41255 -265
rect 41290 -295 41300 -265
rect 41245 -305 41300 -295
rect 41330 -265 41385 -255
rect 41330 -295 41340 -265
rect 41375 -295 41385 -265
rect 41330 -305 41385 -295
rect 41415 -265 41470 -255
rect 41415 -295 41425 -265
rect 41460 -295 41470 -265
rect 41415 -305 41470 -295
rect 41500 -265 41555 -255
rect 41500 -295 41510 -265
rect 41545 -295 41555 -265
rect 41500 -305 41555 -295
rect 41585 -265 41640 -255
rect 41585 -295 41595 -265
rect 41630 -295 41640 -265
rect 41585 -305 41640 -295
rect 41670 -265 41725 -255
rect 41670 -295 41680 -265
rect 41715 -295 41725 -265
rect 41670 -305 41725 -295
rect 41755 -265 41810 -255
rect 41755 -295 41765 -265
rect 41800 -295 41810 -265
rect 41755 -305 41810 -295
rect 41840 -265 41895 -255
rect 41840 -295 41850 -265
rect 41885 -295 41895 -265
rect 41840 -305 41895 -295
rect 41925 -265 41980 -255
rect 41925 -295 41935 -265
rect 41970 -295 41980 -265
rect 41925 -305 41980 -295
rect 42010 -265 42065 -255
rect 42010 -295 42020 -265
rect 42055 -295 42065 -265
rect 42010 -305 42065 -295
rect 42095 -265 42150 -255
rect 42095 -295 42105 -265
rect 42140 -295 42150 -265
rect 42095 -305 42150 -295
rect 42180 -265 42235 -255
rect 42180 -295 42190 -265
rect 42225 -295 42235 -265
rect 42180 -305 42235 -295
rect 42265 -265 42320 -255
rect 42265 -295 42275 -265
rect 42310 -295 42320 -265
rect 42265 -305 42320 -295
rect 42350 -265 42405 -255
rect 42350 -295 42360 -265
rect 42395 -295 42405 -265
rect 42350 -305 42405 -295
rect 42435 -265 42490 -255
rect 42435 -295 42445 -265
rect 42480 -295 42490 -265
rect 42435 -305 42490 -295
rect 42520 -265 42575 -255
rect 42520 -295 42530 -265
rect 42565 -295 42575 -265
rect 42520 -305 42575 -295
rect 42605 -265 42660 -255
rect 42605 -295 42615 -265
rect 42650 -295 42660 -265
rect 42605 -305 42660 -295
rect 42690 -265 42745 -255
rect 42690 -295 42700 -265
rect 42735 -295 42745 -265
rect 42690 -305 42745 -295
rect 42775 -265 42830 -255
rect 42775 -295 42785 -265
rect 42820 -295 42830 -265
rect 42775 -305 42830 -295
rect 42860 -265 42915 -255
rect 42860 -295 42870 -265
rect 42905 -295 42915 -265
rect 42860 -305 42915 -295
rect 42945 -265 43000 -255
rect 42945 -295 42955 -265
rect 42990 -295 43000 -265
rect 42945 -305 43000 -295
rect 43030 -265 43085 -255
rect 43030 -295 43040 -265
rect 43075 -295 43085 -265
rect 43030 -305 43085 -295
rect 43115 -265 43170 -255
rect 43115 -295 43125 -265
rect 43160 -295 43170 -265
rect 43115 -305 43170 -295
rect 43200 -265 43255 -255
rect 43200 -295 43210 -265
rect 43245 -295 43255 -265
rect 43200 -305 43255 -295
rect 43285 -265 43340 -255
rect 43285 -295 43295 -265
rect 43330 -295 43340 -265
rect 43285 -305 43340 -295
rect 43370 -265 43425 -255
rect 43370 -295 43380 -265
rect 43415 -295 43425 -265
rect 43370 -305 43425 -295
rect 43455 -265 43510 -255
rect 43455 -295 43465 -265
rect 43500 -295 43510 -265
rect 43455 -305 43510 -295
rect 43540 -265 43595 -255
rect 43540 -295 43550 -265
rect 43585 -295 43595 -265
rect 43540 -305 43595 -295
rect 65 -335 115 -325
rect 65 -365 75 -335
rect 105 -365 115 -335
rect 65 -375 115 -365
rect 235 -335 285 -325
rect 235 -365 245 -335
rect 275 -365 285 -335
rect 235 -375 285 -365
rect 405 -335 455 -325
rect 405 -365 415 -335
rect 445 -365 455 -335
rect 405 -375 455 -365
rect 575 -335 625 -325
rect 575 -365 585 -335
rect 615 -365 625 -335
rect 575 -375 625 -365
rect 745 -335 795 -325
rect 745 -365 755 -335
rect 785 -365 795 -335
rect 745 -375 795 -365
rect 915 -335 965 -325
rect 915 -365 925 -335
rect 955 -365 965 -335
rect 915 -375 965 -365
rect 1085 -335 1135 -325
rect 1085 -365 1095 -335
rect 1125 -365 1135 -335
rect 1085 -375 1135 -365
rect 1255 -335 1305 -325
rect 1255 -365 1265 -335
rect 1295 -365 1305 -335
rect 1255 -375 1305 -365
rect 1425 -335 1475 -325
rect 1425 -365 1435 -335
rect 1465 -365 1475 -335
rect 1425 -375 1475 -365
rect 1595 -335 1645 -325
rect 1595 -365 1605 -335
rect 1635 -365 1645 -335
rect 1595 -375 1645 -365
rect 1765 -335 1815 -325
rect 1765 -365 1775 -335
rect 1805 -365 1815 -335
rect 1765 -375 1815 -365
rect 1935 -335 1985 -325
rect 1935 -365 1945 -335
rect 1975 -365 1985 -335
rect 1935 -375 1985 -365
rect 2105 -335 2155 -325
rect 2105 -365 2115 -335
rect 2145 -365 2155 -335
rect 2105 -375 2155 -365
rect 2275 -335 2325 -325
rect 2275 -365 2285 -335
rect 2315 -365 2325 -335
rect 2275 -375 2325 -365
rect 2445 -335 2495 -325
rect 2445 -365 2455 -335
rect 2485 -365 2495 -335
rect 2445 -375 2495 -365
rect 2615 -335 2665 -325
rect 2615 -365 2625 -335
rect 2655 -365 2665 -335
rect 2615 -375 2665 -365
rect 2785 -335 2835 -325
rect 2785 -365 2795 -335
rect 2825 -365 2835 -335
rect 2785 -375 2835 -365
rect 2955 -335 3005 -325
rect 2955 -365 2965 -335
rect 2995 -365 3005 -335
rect 2955 -375 3005 -365
rect 3125 -335 3175 -325
rect 3125 -365 3135 -335
rect 3165 -365 3175 -335
rect 3125 -375 3175 -365
rect 3295 -335 3345 -325
rect 3295 -365 3305 -335
rect 3335 -365 3345 -335
rect 3295 -375 3345 -365
rect 3465 -335 3515 -325
rect 3465 -365 3475 -335
rect 3505 -365 3515 -335
rect 3465 -375 3515 -365
rect 3635 -335 3685 -325
rect 3635 -365 3645 -335
rect 3675 -365 3685 -335
rect 3635 -375 3685 -365
rect 3805 -335 3855 -325
rect 3805 -365 3815 -335
rect 3845 -365 3855 -335
rect 3805 -375 3855 -365
rect 3975 -335 4025 -325
rect 3975 -365 3985 -335
rect 4015 -365 4025 -335
rect 3975 -375 4025 -365
rect 4145 -335 4195 -325
rect 4145 -365 4155 -335
rect 4185 -365 4195 -335
rect 4145 -375 4195 -365
rect 4315 -335 4365 -325
rect 4315 -365 4325 -335
rect 4355 -365 4365 -335
rect 4315 -375 4365 -365
rect 4485 -335 4535 -325
rect 4485 -365 4495 -335
rect 4525 -365 4535 -335
rect 4485 -375 4535 -365
rect 4655 -335 4705 -325
rect 4655 -365 4665 -335
rect 4695 -365 4705 -335
rect 4655 -375 4705 -365
rect 4825 -335 4875 -325
rect 4825 -365 4835 -335
rect 4865 -365 4875 -335
rect 4825 -375 4875 -365
rect 4995 -335 5045 -325
rect 4995 -365 5005 -335
rect 5035 -365 5045 -335
rect 4995 -375 5045 -365
rect 5165 -335 5215 -325
rect 5165 -365 5175 -335
rect 5205 -365 5215 -335
rect 5165 -375 5215 -365
rect 5335 -335 5385 -325
rect 5335 -365 5345 -335
rect 5375 -365 5385 -335
rect 5335 -375 5385 -365
rect 5505 -335 5555 -325
rect 5505 -365 5515 -335
rect 5545 -365 5555 -335
rect 5505 -375 5555 -365
rect 5675 -335 5725 -325
rect 5675 -365 5685 -335
rect 5715 -365 5725 -335
rect 5675 -375 5725 -365
rect 5845 -335 5895 -325
rect 5845 -365 5855 -335
rect 5885 -365 5895 -335
rect 5845 -375 5895 -365
rect 6015 -335 6065 -325
rect 6015 -365 6025 -335
rect 6055 -365 6065 -335
rect 6015 -375 6065 -365
rect 6185 -335 6235 -325
rect 6185 -365 6195 -335
rect 6225 -365 6235 -335
rect 6185 -375 6235 -365
rect 6355 -335 6405 -325
rect 6355 -365 6365 -335
rect 6395 -365 6405 -335
rect 6355 -375 6405 -365
rect 6525 -335 6575 -325
rect 6525 -365 6535 -335
rect 6565 -365 6575 -335
rect 6525 -375 6575 -365
rect 6695 -335 6745 -325
rect 6695 -365 6705 -335
rect 6735 -365 6745 -335
rect 6695 -375 6745 -365
rect 6865 -335 6915 -325
rect 6865 -365 6875 -335
rect 6905 -365 6915 -335
rect 6865 -375 6915 -365
rect 7035 -335 7085 -325
rect 7035 -365 7045 -335
rect 7075 -365 7085 -335
rect 7035 -375 7085 -365
rect 7205 -335 7255 -325
rect 7205 -365 7215 -335
rect 7245 -365 7255 -335
rect 7205 -375 7255 -365
rect 7375 -335 7425 -325
rect 7375 -365 7385 -335
rect 7415 -365 7425 -335
rect 7375 -375 7425 -365
rect 7545 -335 7595 -325
rect 7545 -365 7555 -335
rect 7585 -365 7595 -335
rect 7545 -375 7595 -365
rect 7715 -335 7765 -325
rect 7715 -365 7725 -335
rect 7755 -365 7765 -335
rect 7715 -375 7765 -365
rect 7885 -335 7935 -325
rect 7885 -365 7895 -335
rect 7925 -365 7935 -335
rect 7885 -375 7935 -365
rect 8055 -335 8105 -325
rect 8055 -365 8065 -335
rect 8095 -365 8105 -335
rect 8055 -375 8105 -365
rect 8225 -335 8275 -325
rect 8225 -365 8235 -335
rect 8265 -365 8275 -335
rect 8225 -375 8275 -365
rect 8395 -335 8445 -325
rect 8395 -365 8405 -335
rect 8435 -365 8445 -335
rect 8395 -375 8445 -365
rect 8565 -335 8615 -325
rect 8565 -365 8575 -335
rect 8605 -365 8615 -335
rect 8565 -375 8615 -365
rect 8735 -335 8785 -325
rect 8735 -365 8745 -335
rect 8775 -365 8785 -335
rect 8735 -375 8785 -365
rect 8905 -335 8955 -325
rect 8905 -365 8915 -335
rect 8945 -365 8955 -335
rect 8905 -375 8955 -365
rect 9075 -335 9125 -325
rect 9075 -365 9085 -335
rect 9115 -365 9125 -335
rect 9075 -375 9125 -365
rect 9245 -335 9295 -325
rect 9245 -365 9255 -335
rect 9285 -365 9295 -335
rect 9245 -375 9295 -365
rect 9415 -335 9465 -325
rect 9415 -365 9425 -335
rect 9455 -365 9465 -335
rect 9415 -375 9465 -365
rect 9585 -335 9635 -325
rect 9585 -365 9595 -335
rect 9625 -365 9635 -335
rect 9585 -375 9635 -365
rect 9755 -335 9805 -325
rect 9755 -365 9765 -335
rect 9795 -365 9805 -335
rect 9755 -375 9805 -365
rect 9925 -335 9975 -325
rect 9925 -365 9935 -335
rect 9965 -365 9975 -335
rect 9925 -375 9975 -365
rect 10095 -335 10145 -325
rect 10095 -365 10105 -335
rect 10135 -365 10145 -335
rect 10095 -375 10145 -365
rect 10265 -335 10315 -325
rect 10265 -365 10275 -335
rect 10305 -365 10315 -335
rect 10265 -375 10315 -365
rect 10435 -335 10485 -325
rect 10435 -365 10445 -335
rect 10475 -365 10485 -335
rect 10435 -375 10485 -365
rect 10605 -335 10655 -325
rect 10605 -365 10615 -335
rect 10645 -365 10655 -335
rect 10605 -375 10655 -365
rect 10775 -335 10825 -325
rect 10775 -365 10785 -335
rect 10815 -365 10825 -335
rect 10775 -375 10825 -365
rect 10945 -335 10995 -325
rect 10945 -365 10955 -335
rect 10985 -365 10995 -335
rect 10945 -375 10995 -365
rect 11115 -335 11165 -325
rect 11115 -365 11125 -335
rect 11155 -365 11165 -335
rect 11115 -375 11165 -365
rect 11285 -335 11335 -325
rect 11285 -365 11295 -335
rect 11325 -365 11335 -335
rect 11285 -375 11335 -365
rect 11455 -335 11505 -325
rect 11455 -365 11465 -335
rect 11495 -365 11505 -335
rect 11455 -375 11505 -365
rect 11625 -335 11675 -325
rect 11625 -365 11635 -335
rect 11665 -365 11675 -335
rect 11625 -375 11675 -365
rect 11795 -335 11845 -325
rect 11795 -365 11805 -335
rect 11835 -365 11845 -335
rect 11795 -375 11845 -365
rect 11965 -335 12015 -325
rect 11965 -365 11975 -335
rect 12005 -365 12015 -335
rect 11965 -375 12015 -365
rect 12135 -335 12185 -325
rect 12135 -365 12145 -335
rect 12175 -365 12185 -335
rect 12135 -375 12185 -365
rect 12305 -335 12355 -325
rect 12305 -365 12315 -335
rect 12345 -365 12355 -335
rect 12305 -375 12355 -365
rect 12475 -335 12525 -325
rect 12475 -365 12485 -335
rect 12515 -365 12525 -335
rect 12475 -375 12525 -365
rect 12645 -335 12695 -325
rect 12645 -365 12655 -335
rect 12685 -365 12695 -335
rect 12645 -375 12695 -365
rect 12815 -335 12865 -325
rect 12815 -365 12825 -335
rect 12855 -365 12865 -335
rect 12815 -375 12865 -365
rect 12985 -335 13035 -325
rect 12985 -365 12995 -335
rect 13025 -365 13035 -335
rect 12985 -375 13035 -365
rect 13155 -335 13205 -325
rect 13155 -365 13165 -335
rect 13195 -365 13205 -335
rect 13155 -375 13205 -365
rect 13325 -335 13375 -325
rect 13325 -365 13335 -335
rect 13365 -365 13375 -335
rect 13325 -375 13375 -365
rect 13495 -335 13545 -325
rect 13495 -365 13505 -335
rect 13535 -365 13545 -335
rect 13495 -375 13545 -365
rect 13665 -335 13715 -325
rect 13665 -365 13675 -335
rect 13705 -365 13715 -335
rect 13665 -375 13715 -365
rect 13835 -335 13885 -325
rect 13835 -365 13845 -335
rect 13875 -365 13885 -335
rect 13835 -375 13885 -365
rect 14005 -335 14055 -325
rect 14005 -365 14015 -335
rect 14045 -365 14055 -335
rect 14005 -375 14055 -365
rect 14175 -335 14225 -325
rect 14175 -365 14185 -335
rect 14215 -365 14225 -335
rect 14175 -375 14225 -365
rect 14345 -335 14395 -325
rect 14345 -365 14355 -335
rect 14385 -365 14395 -335
rect 14345 -375 14395 -365
rect 14515 -335 14565 -325
rect 14515 -365 14525 -335
rect 14555 -365 14565 -335
rect 14515 -375 14565 -365
rect 14685 -335 14735 -325
rect 14685 -365 14695 -335
rect 14725 -365 14735 -335
rect 14685 -375 14735 -365
rect 14855 -335 14905 -325
rect 14855 -365 14865 -335
rect 14895 -365 14905 -335
rect 14855 -375 14905 -365
rect 15025 -335 15075 -325
rect 15025 -365 15035 -335
rect 15065 -365 15075 -335
rect 15025 -375 15075 -365
rect 15195 -335 15245 -325
rect 15195 -365 15205 -335
rect 15235 -365 15245 -335
rect 15195 -375 15245 -365
rect 15365 -335 15415 -325
rect 15365 -365 15375 -335
rect 15405 -365 15415 -335
rect 15365 -375 15415 -365
rect 15535 -335 15585 -325
rect 15535 -365 15545 -335
rect 15575 -365 15585 -335
rect 15535 -375 15585 -365
rect 15705 -335 15755 -325
rect 15705 -365 15715 -335
rect 15745 -365 15755 -335
rect 15705 -375 15755 -365
rect 15875 -335 15925 -325
rect 15875 -365 15885 -335
rect 15915 -365 15925 -335
rect 15875 -375 15925 -365
rect 16045 -335 16095 -325
rect 16045 -365 16055 -335
rect 16085 -365 16095 -335
rect 16045 -375 16095 -365
rect 16215 -335 16265 -325
rect 16215 -365 16225 -335
rect 16255 -365 16265 -335
rect 16215 -375 16265 -365
rect 16385 -335 16435 -325
rect 16385 -365 16395 -335
rect 16425 -365 16435 -335
rect 16385 -375 16435 -365
rect 16555 -335 16605 -325
rect 16555 -365 16565 -335
rect 16595 -365 16605 -335
rect 16555 -375 16605 -365
rect 16725 -335 16775 -325
rect 16725 -365 16735 -335
rect 16765 -365 16775 -335
rect 16725 -375 16775 -365
rect 16895 -335 16945 -325
rect 16895 -365 16905 -335
rect 16935 -365 16945 -335
rect 16895 -375 16945 -365
rect 17065 -335 17115 -325
rect 17065 -365 17075 -335
rect 17105 -365 17115 -335
rect 17065 -375 17115 -365
rect 17235 -335 17285 -325
rect 17235 -365 17245 -335
rect 17275 -365 17285 -335
rect 17235 -375 17285 -365
rect 17405 -335 17455 -325
rect 17405 -365 17415 -335
rect 17445 -365 17455 -335
rect 17405 -375 17455 -365
rect 17575 -335 17625 -325
rect 17575 -365 17585 -335
rect 17615 -365 17625 -335
rect 17575 -375 17625 -365
rect 17745 -335 17795 -325
rect 17745 -365 17755 -335
rect 17785 -365 17795 -335
rect 17745 -375 17795 -365
rect 17915 -335 17965 -325
rect 17915 -365 17925 -335
rect 17955 -365 17965 -335
rect 17915 -375 17965 -365
rect 18085 -335 18135 -325
rect 18085 -365 18095 -335
rect 18125 -365 18135 -335
rect 18085 -375 18135 -365
rect 18255 -335 18305 -325
rect 18255 -365 18265 -335
rect 18295 -365 18305 -335
rect 18255 -375 18305 -365
rect 18425 -335 18475 -325
rect 18425 -365 18435 -335
rect 18465 -365 18475 -335
rect 18425 -375 18475 -365
rect 18595 -335 18645 -325
rect 18595 -365 18605 -335
rect 18635 -365 18645 -335
rect 18595 -375 18645 -365
rect 18765 -335 18815 -325
rect 18765 -365 18775 -335
rect 18805 -365 18815 -335
rect 18765 -375 18815 -365
rect 18935 -335 18985 -325
rect 18935 -365 18945 -335
rect 18975 -365 18985 -335
rect 18935 -375 18985 -365
rect 19105 -335 19155 -325
rect 19105 -365 19115 -335
rect 19145 -365 19155 -335
rect 19105 -375 19155 -365
rect 19275 -335 19325 -325
rect 19275 -365 19285 -335
rect 19315 -365 19325 -335
rect 19275 -375 19325 -365
rect 19445 -335 19495 -325
rect 19445 -365 19455 -335
rect 19485 -365 19495 -335
rect 19445 -375 19495 -365
rect 19615 -335 19665 -325
rect 19615 -365 19625 -335
rect 19655 -365 19665 -335
rect 19615 -375 19665 -365
rect 19785 -335 19835 -325
rect 19785 -365 19795 -335
rect 19825 -365 19835 -335
rect 19785 -375 19835 -365
rect 19955 -335 20005 -325
rect 19955 -365 19965 -335
rect 19995 -365 20005 -335
rect 19955 -375 20005 -365
rect 20125 -335 20175 -325
rect 20125 -365 20135 -335
rect 20165 -365 20175 -335
rect 20125 -375 20175 -365
rect 20295 -335 20345 -325
rect 20295 -365 20305 -335
rect 20335 -365 20345 -335
rect 20295 -375 20345 -365
rect 20465 -335 20515 -325
rect 20465 -365 20475 -335
rect 20505 -365 20515 -335
rect 20465 -375 20515 -365
rect 20635 -335 20685 -325
rect 20635 -365 20645 -335
rect 20675 -365 20685 -335
rect 20635 -375 20685 -365
rect 20805 -335 20855 -325
rect 20805 -365 20815 -335
rect 20845 -365 20855 -335
rect 20805 -375 20855 -365
rect 20975 -335 21025 -325
rect 20975 -365 20985 -335
rect 21015 -365 21025 -335
rect 20975 -375 21025 -365
rect 21145 -335 21195 -325
rect 21145 -365 21155 -335
rect 21185 -365 21195 -335
rect 21145 -375 21195 -365
rect 21315 -335 21365 -325
rect 21315 -365 21325 -335
rect 21355 -365 21365 -335
rect 21315 -375 21365 -365
rect 21485 -335 21535 -325
rect 21485 -365 21495 -335
rect 21525 -365 21535 -335
rect 21485 -375 21535 -365
rect 21655 -335 21705 -325
rect 21655 -365 21665 -335
rect 21695 -365 21705 -335
rect 21655 -375 21705 -365
rect 21825 -335 21875 -325
rect 21825 -365 21835 -335
rect 21865 -365 21875 -335
rect 21825 -375 21875 -365
rect 21995 -335 22045 -325
rect 21995 -365 22005 -335
rect 22035 -365 22045 -335
rect 21995 -375 22045 -365
rect 22165 -335 22215 -325
rect 22165 -365 22175 -335
rect 22205 -365 22215 -335
rect 22165 -375 22215 -365
rect 22335 -335 22385 -325
rect 22335 -365 22345 -335
rect 22375 -365 22385 -335
rect 22335 -375 22385 -365
rect 22505 -335 22555 -325
rect 22505 -365 22515 -335
rect 22545 -365 22555 -335
rect 22505 -375 22555 -365
rect 22675 -335 22725 -325
rect 22675 -365 22685 -335
rect 22715 -365 22725 -335
rect 22675 -375 22725 -365
rect 22845 -335 22895 -325
rect 22845 -365 22855 -335
rect 22885 -365 22895 -335
rect 22845 -375 22895 -365
rect 23015 -335 23065 -325
rect 23015 -365 23025 -335
rect 23055 -365 23065 -335
rect 23015 -375 23065 -365
rect 23185 -335 23235 -325
rect 23185 -365 23195 -335
rect 23225 -365 23235 -335
rect 23185 -375 23235 -365
rect 23355 -335 23405 -325
rect 23355 -365 23365 -335
rect 23395 -365 23405 -335
rect 23355 -375 23405 -365
rect 23525 -335 23575 -325
rect 23525 -365 23535 -335
rect 23565 -365 23575 -335
rect 23525 -375 23575 -365
rect 23695 -335 23745 -325
rect 23695 -365 23705 -335
rect 23735 -365 23745 -335
rect 23695 -375 23745 -365
rect 23865 -335 23915 -325
rect 23865 -365 23875 -335
rect 23905 -365 23915 -335
rect 23865 -375 23915 -365
rect 24035 -335 24085 -325
rect 24035 -365 24045 -335
rect 24075 -365 24085 -335
rect 24035 -375 24085 -365
rect 24205 -335 24255 -325
rect 24205 -365 24215 -335
rect 24245 -365 24255 -335
rect 24205 -375 24255 -365
rect 24375 -335 24425 -325
rect 24375 -365 24385 -335
rect 24415 -365 24425 -335
rect 24375 -375 24425 -365
rect 24545 -335 24595 -325
rect 24545 -365 24555 -335
rect 24585 -365 24595 -335
rect 24545 -375 24595 -365
rect 24715 -335 24765 -325
rect 24715 -365 24725 -335
rect 24755 -365 24765 -335
rect 24715 -375 24765 -365
rect 24885 -335 24935 -325
rect 24885 -365 24895 -335
rect 24925 -365 24935 -335
rect 24885 -375 24935 -365
rect 25055 -335 25105 -325
rect 25055 -365 25065 -335
rect 25095 -365 25105 -335
rect 25055 -375 25105 -365
rect 25225 -335 25275 -325
rect 25225 -365 25235 -335
rect 25265 -365 25275 -335
rect 25225 -375 25275 -365
rect 25395 -335 25445 -325
rect 25395 -365 25405 -335
rect 25435 -365 25445 -335
rect 25395 -375 25445 -365
rect 25565 -335 25615 -325
rect 25565 -365 25575 -335
rect 25605 -365 25615 -335
rect 25565 -375 25615 -365
rect 25735 -335 25785 -325
rect 25735 -365 25745 -335
rect 25775 -365 25785 -335
rect 25735 -375 25785 -365
rect 25905 -335 25955 -325
rect 25905 -365 25915 -335
rect 25945 -365 25955 -335
rect 25905 -375 25955 -365
rect 26075 -335 26125 -325
rect 26075 -365 26085 -335
rect 26115 -365 26125 -335
rect 26075 -375 26125 -365
rect 26245 -335 26295 -325
rect 26245 -365 26255 -335
rect 26285 -365 26295 -335
rect 26245 -375 26295 -365
rect 26415 -335 26465 -325
rect 26415 -365 26425 -335
rect 26455 -365 26465 -335
rect 26415 -375 26465 -365
rect 26585 -335 26635 -325
rect 26585 -365 26595 -335
rect 26625 -365 26635 -335
rect 26585 -375 26635 -365
rect 26755 -335 26805 -325
rect 26755 -365 26765 -335
rect 26795 -365 26805 -335
rect 26755 -375 26805 -365
rect 26925 -335 26975 -325
rect 26925 -365 26935 -335
rect 26965 -365 26975 -335
rect 26925 -375 26975 -365
rect 27095 -335 27145 -325
rect 27095 -365 27105 -335
rect 27135 -365 27145 -335
rect 27095 -375 27145 -365
rect 27265 -335 27315 -325
rect 27265 -365 27275 -335
rect 27305 -365 27315 -335
rect 27265 -375 27315 -365
rect 27435 -335 27485 -325
rect 27435 -365 27445 -335
rect 27475 -365 27485 -335
rect 27435 -375 27485 -365
rect 27605 -335 27655 -325
rect 27605 -365 27615 -335
rect 27645 -365 27655 -335
rect 27605 -375 27655 -365
rect 27775 -335 27825 -325
rect 27775 -365 27785 -335
rect 27815 -365 27825 -335
rect 27775 -375 27825 -365
rect 27945 -335 27995 -325
rect 27945 -365 27955 -335
rect 27985 -365 27995 -335
rect 27945 -375 27995 -365
rect 28115 -335 28165 -325
rect 28115 -365 28125 -335
rect 28155 -365 28165 -335
rect 28115 -375 28165 -365
rect 28285 -335 28335 -325
rect 28285 -365 28295 -335
rect 28325 -365 28335 -335
rect 28285 -375 28335 -365
rect 28455 -335 28505 -325
rect 28455 -365 28465 -335
rect 28495 -365 28505 -335
rect 28455 -375 28505 -365
rect 28625 -335 28675 -325
rect 28625 -365 28635 -335
rect 28665 -365 28675 -335
rect 28625 -375 28675 -365
rect 28795 -335 28845 -325
rect 28795 -365 28805 -335
rect 28835 -365 28845 -335
rect 28795 -375 28845 -365
rect 28965 -335 29015 -325
rect 28965 -365 28975 -335
rect 29005 -365 29015 -335
rect 28965 -375 29015 -365
rect 29135 -335 29185 -325
rect 29135 -365 29145 -335
rect 29175 -365 29185 -335
rect 29135 -375 29185 -365
rect 29305 -335 29355 -325
rect 29305 -365 29315 -335
rect 29345 -365 29355 -335
rect 29305 -375 29355 -365
rect 29475 -335 29525 -325
rect 29475 -365 29485 -335
rect 29515 -365 29525 -335
rect 29475 -375 29525 -365
rect 29645 -335 29695 -325
rect 29645 -365 29655 -335
rect 29685 -365 29695 -335
rect 29645 -375 29695 -365
rect 29815 -335 29865 -325
rect 29815 -365 29825 -335
rect 29855 -365 29865 -335
rect 29815 -375 29865 -365
rect 29985 -335 30035 -325
rect 29985 -365 29995 -335
rect 30025 -365 30035 -335
rect 29985 -375 30035 -365
rect 30155 -335 30205 -325
rect 30155 -365 30165 -335
rect 30195 -365 30205 -335
rect 30155 -375 30205 -365
rect 30325 -335 30375 -325
rect 30325 -365 30335 -335
rect 30365 -365 30375 -335
rect 30325 -375 30375 -365
rect 30495 -335 30545 -325
rect 30495 -365 30505 -335
rect 30535 -365 30545 -335
rect 30495 -375 30545 -365
rect 30665 -335 30715 -325
rect 30665 -365 30675 -335
rect 30705 -365 30715 -335
rect 30665 -375 30715 -365
rect 30835 -335 30885 -325
rect 30835 -365 30845 -335
rect 30875 -365 30885 -335
rect 30835 -375 30885 -365
rect 31005 -335 31055 -325
rect 31005 -365 31015 -335
rect 31045 -365 31055 -335
rect 31005 -375 31055 -365
rect 31175 -335 31225 -325
rect 31175 -365 31185 -335
rect 31215 -365 31225 -335
rect 31175 -375 31225 -365
rect 31345 -335 31395 -325
rect 31345 -365 31355 -335
rect 31385 -365 31395 -335
rect 31345 -375 31395 -365
rect 31515 -335 31565 -325
rect 31515 -365 31525 -335
rect 31555 -365 31565 -335
rect 31515 -375 31565 -365
rect 31685 -335 31735 -325
rect 31685 -365 31695 -335
rect 31725 -365 31735 -335
rect 31685 -375 31735 -365
rect 31855 -335 31905 -325
rect 31855 -365 31865 -335
rect 31895 -365 31905 -335
rect 31855 -375 31905 -365
rect 32025 -335 32075 -325
rect 32025 -365 32035 -335
rect 32065 -365 32075 -335
rect 32025 -375 32075 -365
rect 32195 -335 32245 -325
rect 32195 -365 32205 -335
rect 32235 -365 32245 -335
rect 32195 -375 32245 -365
rect 32365 -335 32415 -325
rect 32365 -365 32375 -335
rect 32405 -365 32415 -335
rect 32365 -375 32415 -365
rect 32535 -335 32585 -325
rect 32535 -365 32545 -335
rect 32575 -365 32585 -335
rect 32535 -375 32585 -365
rect 32705 -335 32755 -325
rect 32705 -365 32715 -335
rect 32745 -365 32755 -335
rect 32705 -375 32755 -365
rect 32875 -335 32925 -325
rect 32875 -365 32885 -335
rect 32915 -365 32925 -335
rect 32875 -375 32925 -365
rect 33045 -335 33095 -325
rect 33045 -365 33055 -335
rect 33085 -365 33095 -335
rect 33045 -375 33095 -365
rect 33215 -335 33265 -325
rect 33215 -365 33225 -335
rect 33255 -365 33265 -335
rect 33215 -375 33265 -365
rect 33385 -335 33435 -325
rect 33385 -365 33395 -335
rect 33425 -365 33435 -335
rect 33385 -375 33435 -365
rect 33555 -335 33605 -325
rect 33555 -365 33565 -335
rect 33595 -365 33605 -335
rect 33555 -375 33605 -365
rect 33725 -335 33775 -325
rect 33725 -365 33735 -335
rect 33765 -365 33775 -335
rect 33725 -375 33775 -365
rect 33895 -335 33945 -325
rect 33895 -365 33905 -335
rect 33935 -365 33945 -335
rect 33895 -375 33945 -365
rect 34065 -335 34115 -325
rect 34065 -365 34075 -335
rect 34105 -365 34115 -335
rect 34065 -375 34115 -365
rect 34235 -335 34285 -325
rect 34235 -365 34245 -335
rect 34275 -365 34285 -335
rect 34235 -375 34285 -365
rect 34405 -335 34455 -325
rect 34405 -365 34415 -335
rect 34445 -365 34455 -335
rect 34405 -375 34455 -365
rect 34575 -335 34625 -325
rect 34575 -365 34585 -335
rect 34615 -365 34625 -335
rect 34575 -375 34625 -365
rect 34745 -335 34795 -325
rect 34745 -365 34755 -335
rect 34785 -365 34795 -335
rect 34745 -375 34795 -365
rect 34915 -335 34965 -325
rect 34915 -365 34925 -335
rect 34955 -365 34965 -335
rect 34915 -375 34965 -365
rect 35085 -335 35135 -325
rect 35085 -365 35095 -335
rect 35125 -365 35135 -335
rect 35085 -375 35135 -365
rect 35255 -335 35305 -325
rect 35255 -365 35265 -335
rect 35295 -365 35305 -335
rect 35255 -375 35305 -365
rect 35425 -335 35475 -325
rect 35425 -365 35435 -335
rect 35465 -365 35475 -335
rect 35425 -375 35475 -365
rect 35595 -335 35645 -325
rect 35595 -365 35605 -335
rect 35635 -365 35645 -335
rect 35595 -375 35645 -365
rect 35765 -335 35815 -325
rect 35765 -365 35775 -335
rect 35805 -365 35815 -335
rect 35765 -375 35815 -365
rect 35935 -335 35985 -325
rect 35935 -365 35945 -335
rect 35975 -365 35985 -335
rect 35935 -375 35985 -365
rect 36105 -335 36155 -325
rect 36105 -365 36115 -335
rect 36145 -365 36155 -335
rect 36105 -375 36155 -365
rect 36275 -335 36325 -325
rect 36275 -365 36285 -335
rect 36315 -365 36325 -335
rect 36275 -375 36325 -365
rect 36445 -335 36495 -325
rect 36445 -365 36455 -335
rect 36485 -365 36495 -335
rect 36445 -375 36495 -365
rect 36615 -335 36665 -325
rect 36615 -365 36625 -335
rect 36655 -365 36665 -335
rect 36615 -375 36665 -365
rect 36785 -335 36835 -325
rect 36785 -365 36795 -335
rect 36825 -365 36835 -335
rect 36785 -375 36835 -365
rect 36955 -335 37005 -325
rect 36955 -365 36965 -335
rect 36995 -365 37005 -335
rect 36955 -375 37005 -365
rect 37125 -335 37175 -325
rect 37125 -365 37135 -335
rect 37165 -365 37175 -335
rect 37125 -375 37175 -365
rect 37295 -335 37345 -325
rect 37295 -365 37305 -335
rect 37335 -365 37345 -335
rect 37295 -375 37345 -365
rect 37465 -335 37515 -325
rect 37465 -365 37475 -335
rect 37505 -365 37515 -335
rect 37465 -375 37515 -365
rect 37635 -335 37685 -325
rect 37635 -365 37645 -335
rect 37675 -365 37685 -335
rect 37635 -375 37685 -365
rect 37805 -335 37855 -325
rect 37805 -365 37815 -335
rect 37845 -365 37855 -335
rect 37805 -375 37855 -365
rect 37975 -335 38025 -325
rect 37975 -365 37985 -335
rect 38015 -365 38025 -335
rect 37975 -375 38025 -365
rect 38145 -335 38195 -325
rect 38145 -365 38155 -335
rect 38185 -365 38195 -335
rect 38145 -375 38195 -365
rect 38315 -335 38365 -325
rect 38315 -365 38325 -335
rect 38355 -365 38365 -335
rect 38315 -375 38365 -365
rect 38485 -335 38535 -325
rect 38485 -365 38495 -335
rect 38525 -365 38535 -335
rect 38485 -375 38535 -365
rect 38655 -335 38705 -325
rect 38655 -365 38665 -335
rect 38695 -365 38705 -335
rect 38655 -375 38705 -365
rect 38825 -335 38875 -325
rect 38825 -365 38835 -335
rect 38865 -365 38875 -335
rect 38825 -375 38875 -365
rect 38995 -335 39045 -325
rect 38995 -365 39005 -335
rect 39035 -365 39045 -335
rect 38995 -375 39045 -365
rect 39165 -335 39215 -325
rect 39165 -365 39175 -335
rect 39205 -365 39215 -335
rect 39165 -375 39215 -365
rect 39335 -335 39385 -325
rect 39335 -365 39345 -335
rect 39375 -365 39385 -335
rect 39335 -375 39385 -365
rect 39505 -335 39555 -325
rect 39505 -365 39515 -335
rect 39545 -365 39555 -335
rect 39505 -375 39555 -365
rect 39675 -335 39725 -325
rect 39675 -365 39685 -335
rect 39715 -365 39725 -335
rect 39675 -375 39725 -365
rect 39845 -335 39895 -325
rect 39845 -365 39855 -335
rect 39885 -365 39895 -335
rect 39845 -375 39895 -365
rect 40015 -335 40065 -325
rect 40015 -365 40025 -335
rect 40055 -365 40065 -335
rect 40015 -375 40065 -365
rect 40185 -335 40235 -325
rect 40185 -365 40195 -335
rect 40225 -365 40235 -335
rect 40185 -375 40235 -365
rect 40355 -335 40405 -325
rect 40355 -365 40365 -335
rect 40395 -365 40405 -335
rect 40355 -375 40405 -365
rect 40525 -335 40575 -325
rect 40525 -365 40535 -335
rect 40565 -365 40575 -335
rect 40525 -375 40575 -365
rect 40695 -335 40745 -325
rect 40695 -365 40705 -335
rect 40735 -365 40745 -335
rect 40695 -375 40745 -365
rect 40865 -335 40915 -325
rect 40865 -365 40875 -335
rect 40905 -365 40915 -335
rect 40865 -375 40915 -365
rect 41035 -335 41085 -325
rect 41035 -365 41045 -335
rect 41075 -365 41085 -335
rect 41035 -375 41085 -365
rect 41205 -335 41255 -325
rect 41205 -365 41215 -335
rect 41245 -365 41255 -335
rect 41205 -375 41255 -365
rect 41375 -335 41425 -325
rect 41375 -365 41385 -335
rect 41415 -365 41425 -335
rect 41375 -375 41425 -365
rect 41545 -335 41595 -325
rect 41545 -365 41555 -335
rect 41585 -365 41595 -335
rect 41545 -375 41595 -365
rect 41715 -335 41765 -325
rect 41715 -365 41725 -335
rect 41755 -365 41765 -335
rect 41715 -375 41765 -365
rect 41885 -335 41935 -325
rect 41885 -365 41895 -335
rect 41925 -365 41935 -335
rect 41885 -375 41935 -365
rect 42055 -335 42105 -325
rect 42055 -365 42065 -335
rect 42095 -365 42105 -335
rect 42055 -375 42105 -365
rect 42225 -335 42275 -325
rect 42225 -365 42235 -335
rect 42265 -365 42275 -335
rect 42225 -375 42275 -365
rect 42395 -335 42445 -325
rect 42395 -365 42405 -335
rect 42435 -365 42445 -335
rect 42395 -375 42445 -365
rect 42565 -335 42615 -325
rect 42565 -365 42575 -335
rect 42605 -365 42615 -335
rect 42565 -375 42615 -365
rect 42735 -335 42785 -325
rect 42735 -365 42745 -335
rect 42775 -365 42785 -335
rect 42735 -375 42785 -365
rect 42905 -335 42955 -325
rect 42905 -365 42915 -335
rect 42945 -365 42955 -335
rect 42905 -375 42955 -365
rect 43075 -335 43125 -325
rect 43075 -365 43085 -335
rect 43115 -365 43125 -335
rect 43075 -375 43125 -365
rect 43245 -335 43295 -325
rect 43245 -365 43255 -335
rect 43285 -365 43295 -335
rect 43245 -375 43295 -365
rect 43415 -335 43465 -325
rect 43415 -365 43425 -335
rect 43455 -365 43465 -335
rect 43415 -375 43465 -365
rect 43585 -335 43635 -325
rect 43585 -365 43595 -335
rect 43625 -365 43635 -335
rect 43585 -375 43635 -365
rect 150 -385 200 -375
rect 150 -415 160 -385
rect 190 -415 200 -385
rect 150 -440 200 -415
rect 150 -475 160 -440
rect 190 -475 200 -440
rect 150 -500 200 -475
rect 150 -530 160 -500
rect 190 -530 200 -500
rect 65 -550 115 -540
rect 65 -580 75 -550
rect 105 -580 115 -550
rect 65 -590 115 -580
rect 150 -600 200 -530
rect 320 -385 370 -375
rect 320 -415 330 -385
rect 360 -415 370 -385
rect 320 -440 370 -415
rect 320 -475 330 -440
rect 360 -475 370 -440
rect 320 -500 370 -475
rect 320 -530 330 -500
rect 360 -530 370 -500
rect 235 -550 285 -540
rect 235 -580 245 -550
rect 275 -580 285 -550
rect 235 -590 285 -580
rect 150 -630 160 -600
rect 190 -630 200 -600
rect 150 -635 200 -630
rect 320 -600 370 -530
rect 490 -385 540 -375
rect 490 -415 500 -385
rect 530 -415 540 -385
rect 490 -440 540 -415
rect 490 -475 500 -440
rect 530 -475 540 -440
rect 490 -500 540 -475
rect 490 -530 500 -500
rect 530 -530 540 -500
rect 405 -550 455 -540
rect 405 -580 415 -550
rect 445 -580 455 -550
rect 405 -590 455 -580
rect 320 -630 330 -600
rect 360 -630 370 -600
rect 320 -635 370 -630
rect 490 -600 540 -530
rect 660 -385 710 -375
rect 660 -415 670 -385
rect 700 -415 710 -385
rect 660 -440 710 -415
rect 660 -475 670 -440
rect 700 -475 710 -440
rect 660 -500 710 -475
rect 660 -530 670 -500
rect 700 -530 710 -500
rect 575 -550 625 -540
rect 575 -580 585 -550
rect 615 -580 625 -550
rect 575 -590 625 -580
rect 490 -630 500 -600
rect 530 -630 540 -600
rect 490 -635 540 -630
rect 660 -600 710 -530
rect 830 -385 880 -375
rect 830 -415 840 -385
rect 870 -415 880 -385
rect 830 -440 880 -415
rect 830 -475 840 -440
rect 870 -475 880 -440
rect 830 -500 880 -475
rect 830 -530 840 -500
rect 870 -530 880 -500
rect 745 -550 795 -540
rect 745 -580 755 -550
rect 785 -580 795 -550
rect 745 -590 795 -580
rect 660 -630 670 -600
rect 700 -630 710 -600
rect 660 -635 710 -630
rect 830 -600 880 -530
rect 1000 -385 1050 -375
rect 1000 -415 1010 -385
rect 1040 -415 1050 -385
rect 1000 -440 1050 -415
rect 1000 -475 1010 -440
rect 1040 -475 1050 -440
rect 1000 -500 1050 -475
rect 1000 -530 1010 -500
rect 1040 -530 1050 -500
rect 915 -550 965 -540
rect 915 -580 925 -550
rect 955 -580 965 -550
rect 915 -590 965 -580
rect 830 -630 840 -600
rect 870 -630 880 -600
rect 830 -635 880 -630
rect 1000 -600 1050 -530
rect 1170 -385 1220 -375
rect 1170 -415 1180 -385
rect 1210 -415 1220 -385
rect 1170 -440 1220 -415
rect 1170 -475 1180 -440
rect 1210 -475 1220 -440
rect 1170 -500 1220 -475
rect 1170 -530 1180 -500
rect 1210 -530 1220 -500
rect 1085 -550 1135 -540
rect 1085 -580 1095 -550
rect 1125 -580 1135 -550
rect 1085 -590 1135 -580
rect 1000 -630 1010 -600
rect 1040 -630 1050 -600
rect 1000 -635 1050 -630
rect 1170 -600 1220 -530
rect 1340 -385 1390 -375
rect 1340 -415 1350 -385
rect 1380 -415 1390 -385
rect 1340 -440 1390 -415
rect 1340 -475 1350 -440
rect 1380 -475 1390 -440
rect 1340 -500 1390 -475
rect 1340 -530 1350 -500
rect 1380 -530 1390 -500
rect 1255 -550 1305 -540
rect 1255 -580 1265 -550
rect 1295 -580 1305 -550
rect 1255 -590 1305 -580
rect 1170 -630 1180 -600
rect 1210 -630 1220 -600
rect 1170 -635 1220 -630
rect 1340 -600 1390 -530
rect 1510 -385 1560 -375
rect 1510 -415 1520 -385
rect 1550 -415 1560 -385
rect 1510 -440 1560 -415
rect 1510 -475 1520 -440
rect 1550 -475 1560 -440
rect 1510 -500 1560 -475
rect 1510 -530 1520 -500
rect 1550 -530 1560 -500
rect 1425 -550 1475 -540
rect 1425 -580 1435 -550
rect 1465 -580 1475 -550
rect 1425 -590 1475 -580
rect 1340 -630 1350 -600
rect 1380 -630 1390 -600
rect 1340 -635 1390 -630
rect 1510 -600 1560 -530
rect 1680 -385 1730 -375
rect 1680 -415 1690 -385
rect 1720 -415 1730 -385
rect 1680 -440 1730 -415
rect 1680 -475 1690 -440
rect 1720 -475 1730 -440
rect 1680 -500 1730 -475
rect 1680 -530 1690 -500
rect 1720 -530 1730 -500
rect 1595 -550 1645 -540
rect 1595 -580 1605 -550
rect 1635 -580 1645 -550
rect 1595 -590 1645 -580
rect 1510 -630 1520 -600
rect 1550 -630 1560 -600
rect 1510 -635 1560 -630
rect 1680 -600 1730 -530
rect 1850 -385 1900 -375
rect 1850 -415 1860 -385
rect 1890 -415 1900 -385
rect 1850 -440 1900 -415
rect 1850 -475 1860 -440
rect 1890 -475 1900 -440
rect 1850 -500 1900 -475
rect 1850 -530 1860 -500
rect 1890 -530 1900 -500
rect 1765 -550 1815 -540
rect 1765 -580 1775 -550
rect 1805 -580 1815 -550
rect 1765 -590 1815 -580
rect 1680 -630 1690 -600
rect 1720 -630 1730 -600
rect 1680 -635 1730 -630
rect 1850 -600 1900 -530
rect 2020 -385 2070 -375
rect 2020 -415 2030 -385
rect 2060 -415 2070 -385
rect 2020 -440 2070 -415
rect 2020 -475 2030 -440
rect 2060 -475 2070 -440
rect 2020 -500 2070 -475
rect 2020 -530 2030 -500
rect 2060 -530 2070 -500
rect 1935 -550 1985 -540
rect 1935 -580 1945 -550
rect 1975 -580 1985 -550
rect 1935 -590 1985 -580
rect 1850 -630 1860 -600
rect 1890 -630 1900 -600
rect 1850 -635 1900 -630
rect 2020 -600 2070 -530
rect 2190 -385 2240 -375
rect 2190 -415 2200 -385
rect 2230 -415 2240 -385
rect 2190 -440 2240 -415
rect 2190 -475 2200 -440
rect 2230 -475 2240 -440
rect 2190 -500 2240 -475
rect 2190 -530 2200 -500
rect 2230 -530 2240 -500
rect 2105 -550 2155 -540
rect 2105 -580 2115 -550
rect 2145 -580 2155 -550
rect 2105 -590 2155 -580
rect 2020 -630 2030 -600
rect 2060 -630 2070 -600
rect 2020 -635 2070 -630
rect 2190 -600 2240 -530
rect 2360 -385 2410 -375
rect 2360 -415 2370 -385
rect 2400 -415 2410 -385
rect 2360 -440 2410 -415
rect 2360 -475 2370 -440
rect 2400 -475 2410 -440
rect 2360 -500 2410 -475
rect 2360 -530 2370 -500
rect 2400 -530 2410 -500
rect 2275 -550 2325 -540
rect 2275 -580 2285 -550
rect 2315 -580 2325 -550
rect 2275 -590 2325 -580
rect 2190 -630 2200 -600
rect 2230 -630 2240 -600
rect 2190 -635 2240 -630
rect 2360 -600 2410 -530
rect 2530 -385 2580 -375
rect 2530 -415 2540 -385
rect 2570 -415 2580 -385
rect 2530 -440 2580 -415
rect 2530 -475 2540 -440
rect 2570 -475 2580 -440
rect 2530 -500 2580 -475
rect 2530 -530 2540 -500
rect 2570 -530 2580 -500
rect 2445 -550 2495 -540
rect 2445 -580 2455 -550
rect 2485 -580 2495 -550
rect 2445 -590 2495 -580
rect 2360 -630 2370 -600
rect 2400 -630 2410 -600
rect 2360 -635 2410 -630
rect 2530 -600 2580 -530
rect 2700 -385 2750 -375
rect 2700 -415 2710 -385
rect 2740 -415 2750 -385
rect 2700 -440 2750 -415
rect 2700 -475 2710 -440
rect 2740 -475 2750 -440
rect 2700 -500 2750 -475
rect 2700 -530 2710 -500
rect 2740 -530 2750 -500
rect 2615 -550 2665 -540
rect 2615 -580 2625 -550
rect 2655 -580 2665 -550
rect 2615 -590 2665 -580
rect 2530 -630 2540 -600
rect 2570 -630 2580 -600
rect 2530 -635 2580 -630
rect 2700 -600 2750 -530
rect 2870 -385 2920 -375
rect 2870 -415 2880 -385
rect 2910 -415 2920 -385
rect 2870 -440 2920 -415
rect 2870 -475 2880 -440
rect 2910 -475 2920 -440
rect 2870 -500 2920 -475
rect 2870 -530 2880 -500
rect 2910 -530 2920 -500
rect 2785 -550 2835 -540
rect 2785 -580 2795 -550
rect 2825 -580 2835 -550
rect 2785 -590 2835 -580
rect 2700 -630 2710 -600
rect 2740 -630 2750 -600
rect 2700 -635 2750 -630
rect 2870 -600 2920 -530
rect 3040 -385 3090 -375
rect 3040 -415 3050 -385
rect 3080 -415 3090 -385
rect 3040 -440 3090 -415
rect 3040 -475 3050 -440
rect 3080 -475 3090 -440
rect 3040 -500 3090 -475
rect 3040 -530 3050 -500
rect 3080 -530 3090 -500
rect 2955 -550 3005 -540
rect 2955 -580 2965 -550
rect 2995 -580 3005 -550
rect 2955 -590 3005 -580
rect 2870 -630 2880 -600
rect 2910 -630 2920 -600
rect 2870 -635 2920 -630
rect 3040 -600 3090 -530
rect 3210 -385 3260 -375
rect 3210 -415 3220 -385
rect 3250 -415 3260 -385
rect 3210 -440 3260 -415
rect 3210 -475 3220 -440
rect 3250 -475 3260 -440
rect 3210 -500 3260 -475
rect 3210 -530 3220 -500
rect 3250 -530 3260 -500
rect 3125 -550 3175 -540
rect 3125 -580 3135 -550
rect 3165 -580 3175 -550
rect 3125 -590 3175 -580
rect 3040 -630 3050 -600
rect 3080 -630 3090 -600
rect 3040 -635 3090 -630
rect 3210 -600 3260 -530
rect 3380 -385 3430 -375
rect 3380 -415 3390 -385
rect 3420 -415 3430 -385
rect 3380 -440 3430 -415
rect 3380 -475 3390 -440
rect 3420 -475 3430 -440
rect 3380 -500 3430 -475
rect 3380 -530 3390 -500
rect 3420 -530 3430 -500
rect 3295 -550 3345 -540
rect 3295 -580 3305 -550
rect 3335 -580 3345 -550
rect 3295 -590 3345 -580
rect 3210 -630 3220 -600
rect 3250 -630 3260 -600
rect 3210 -635 3260 -630
rect 3380 -600 3430 -530
rect 3550 -385 3600 -375
rect 3550 -415 3560 -385
rect 3590 -415 3600 -385
rect 3550 -440 3600 -415
rect 3550 -475 3560 -440
rect 3590 -475 3600 -440
rect 3550 -500 3600 -475
rect 3550 -530 3560 -500
rect 3590 -530 3600 -500
rect 3465 -550 3515 -540
rect 3465 -580 3475 -550
rect 3505 -580 3515 -550
rect 3465 -590 3515 -580
rect 3380 -630 3390 -600
rect 3420 -630 3430 -600
rect 3380 -635 3430 -630
rect 3550 -600 3600 -530
rect 3720 -385 3770 -375
rect 3720 -415 3730 -385
rect 3760 -415 3770 -385
rect 3720 -440 3770 -415
rect 3720 -475 3730 -440
rect 3760 -475 3770 -440
rect 3720 -500 3770 -475
rect 3720 -530 3730 -500
rect 3760 -530 3770 -500
rect 3635 -550 3685 -540
rect 3635 -580 3645 -550
rect 3675 -580 3685 -550
rect 3635 -590 3685 -580
rect 3550 -630 3560 -600
rect 3590 -630 3600 -600
rect 3550 -635 3600 -630
rect 3720 -600 3770 -530
rect 3890 -385 3940 -375
rect 3890 -415 3900 -385
rect 3930 -415 3940 -385
rect 3890 -440 3940 -415
rect 3890 -475 3900 -440
rect 3930 -475 3940 -440
rect 3890 -500 3940 -475
rect 3890 -530 3900 -500
rect 3930 -530 3940 -500
rect 3805 -550 3855 -540
rect 3805 -580 3815 -550
rect 3845 -580 3855 -550
rect 3805 -590 3855 -580
rect 3720 -630 3730 -600
rect 3760 -630 3770 -600
rect 3720 -635 3770 -630
rect 3890 -600 3940 -530
rect 4060 -385 4110 -375
rect 4060 -415 4070 -385
rect 4100 -415 4110 -385
rect 4060 -440 4110 -415
rect 4060 -475 4070 -440
rect 4100 -475 4110 -440
rect 4060 -500 4110 -475
rect 4060 -530 4070 -500
rect 4100 -530 4110 -500
rect 3975 -550 4025 -540
rect 3975 -580 3985 -550
rect 4015 -580 4025 -550
rect 3975 -590 4025 -580
rect 3890 -630 3900 -600
rect 3930 -630 3940 -600
rect 3890 -635 3940 -630
rect 4060 -600 4110 -530
rect 4230 -385 4280 -375
rect 4230 -415 4240 -385
rect 4270 -415 4280 -385
rect 4230 -440 4280 -415
rect 4230 -475 4240 -440
rect 4270 -475 4280 -440
rect 4230 -500 4280 -475
rect 4230 -530 4240 -500
rect 4270 -530 4280 -500
rect 4145 -550 4195 -540
rect 4145 -580 4155 -550
rect 4185 -580 4195 -550
rect 4145 -590 4195 -580
rect 4060 -630 4070 -600
rect 4100 -630 4110 -600
rect 4060 -635 4110 -630
rect 4230 -600 4280 -530
rect 4400 -385 4450 -375
rect 4400 -415 4410 -385
rect 4440 -415 4450 -385
rect 4400 -440 4450 -415
rect 4400 -475 4410 -440
rect 4440 -475 4450 -440
rect 4400 -500 4450 -475
rect 4400 -530 4410 -500
rect 4440 -530 4450 -500
rect 4315 -550 4365 -540
rect 4315 -580 4325 -550
rect 4355 -580 4365 -550
rect 4315 -590 4365 -580
rect 4230 -630 4240 -600
rect 4270 -630 4280 -600
rect 4230 -635 4280 -630
rect 4400 -600 4450 -530
rect 4570 -385 4620 -375
rect 4570 -415 4580 -385
rect 4610 -415 4620 -385
rect 4570 -440 4620 -415
rect 4570 -475 4580 -440
rect 4610 -475 4620 -440
rect 4570 -500 4620 -475
rect 4570 -530 4580 -500
rect 4610 -530 4620 -500
rect 4485 -550 4535 -540
rect 4485 -580 4495 -550
rect 4525 -580 4535 -550
rect 4485 -590 4535 -580
rect 4400 -630 4410 -600
rect 4440 -630 4450 -600
rect 4400 -635 4450 -630
rect 4570 -600 4620 -530
rect 4740 -385 4790 -375
rect 4740 -415 4750 -385
rect 4780 -415 4790 -385
rect 4740 -440 4790 -415
rect 4740 -475 4750 -440
rect 4780 -475 4790 -440
rect 4740 -500 4790 -475
rect 4740 -530 4750 -500
rect 4780 -530 4790 -500
rect 4655 -550 4705 -540
rect 4655 -580 4665 -550
rect 4695 -580 4705 -550
rect 4655 -590 4705 -580
rect 4570 -630 4580 -600
rect 4610 -630 4620 -600
rect 4570 -635 4620 -630
rect 4740 -600 4790 -530
rect 4910 -385 4960 -375
rect 4910 -415 4920 -385
rect 4950 -415 4960 -385
rect 4910 -440 4960 -415
rect 4910 -475 4920 -440
rect 4950 -475 4960 -440
rect 4910 -500 4960 -475
rect 4910 -530 4920 -500
rect 4950 -530 4960 -500
rect 4825 -550 4875 -540
rect 4825 -580 4835 -550
rect 4865 -580 4875 -550
rect 4825 -590 4875 -580
rect 4740 -630 4750 -600
rect 4780 -630 4790 -600
rect 4740 -635 4790 -630
rect 4910 -600 4960 -530
rect 5080 -385 5130 -375
rect 5080 -415 5090 -385
rect 5120 -415 5130 -385
rect 5080 -440 5130 -415
rect 5080 -475 5090 -440
rect 5120 -475 5130 -440
rect 5080 -500 5130 -475
rect 5080 -530 5090 -500
rect 5120 -530 5130 -500
rect 4995 -550 5045 -540
rect 4995 -580 5005 -550
rect 5035 -580 5045 -550
rect 4995 -590 5045 -580
rect 4910 -630 4920 -600
rect 4950 -630 4960 -600
rect 4910 -635 4960 -630
rect 5080 -600 5130 -530
rect 5250 -385 5300 -375
rect 5250 -415 5260 -385
rect 5290 -415 5300 -385
rect 5250 -440 5300 -415
rect 5250 -475 5260 -440
rect 5290 -475 5300 -440
rect 5250 -500 5300 -475
rect 5250 -530 5260 -500
rect 5290 -530 5300 -500
rect 5165 -550 5215 -540
rect 5165 -580 5175 -550
rect 5205 -580 5215 -550
rect 5165 -590 5215 -580
rect 5080 -630 5090 -600
rect 5120 -630 5130 -600
rect 5080 -635 5130 -630
rect 5250 -600 5300 -530
rect 5420 -385 5470 -375
rect 5420 -415 5430 -385
rect 5460 -415 5470 -385
rect 5420 -440 5470 -415
rect 5420 -475 5430 -440
rect 5460 -475 5470 -440
rect 5420 -500 5470 -475
rect 5420 -530 5430 -500
rect 5460 -530 5470 -500
rect 5335 -550 5385 -540
rect 5335 -580 5345 -550
rect 5375 -580 5385 -550
rect 5335 -590 5385 -580
rect 5250 -630 5260 -600
rect 5290 -630 5300 -600
rect 5250 -635 5300 -630
rect 5420 -600 5470 -530
rect 5590 -385 5640 -375
rect 5590 -415 5600 -385
rect 5630 -415 5640 -385
rect 5590 -440 5640 -415
rect 5590 -475 5600 -440
rect 5630 -475 5640 -440
rect 5590 -500 5640 -475
rect 5590 -530 5600 -500
rect 5630 -530 5640 -500
rect 5505 -550 5555 -540
rect 5505 -580 5515 -550
rect 5545 -580 5555 -550
rect 5505 -590 5555 -580
rect 5420 -630 5430 -600
rect 5460 -630 5470 -600
rect 5420 -635 5470 -630
rect 5590 -600 5640 -530
rect 5760 -385 5810 -375
rect 5760 -415 5770 -385
rect 5800 -415 5810 -385
rect 5760 -440 5810 -415
rect 5760 -475 5770 -440
rect 5800 -475 5810 -440
rect 5760 -500 5810 -475
rect 5760 -530 5770 -500
rect 5800 -530 5810 -500
rect 5675 -550 5725 -540
rect 5675 -580 5685 -550
rect 5715 -580 5725 -550
rect 5675 -590 5725 -580
rect 5590 -630 5600 -600
rect 5630 -630 5640 -600
rect 5590 -635 5640 -630
rect 5760 -600 5810 -530
rect 5930 -385 5980 -375
rect 5930 -415 5940 -385
rect 5970 -415 5980 -385
rect 5930 -440 5980 -415
rect 5930 -475 5940 -440
rect 5970 -475 5980 -440
rect 5930 -500 5980 -475
rect 5930 -530 5940 -500
rect 5970 -530 5980 -500
rect 5845 -550 5895 -540
rect 5845 -580 5855 -550
rect 5885 -580 5895 -550
rect 5845 -590 5895 -580
rect 5760 -630 5770 -600
rect 5800 -630 5810 -600
rect 5760 -635 5810 -630
rect 5930 -600 5980 -530
rect 6100 -385 6150 -375
rect 6100 -415 6110 -385
rect 6140 -415 6150 -385
rect 6100 -440 6150 -415
rect 6100 -475 6110 -440
rect 6140 -475 6150 -440
rect 6100 -500 6150 -475
rect 6100 -530 6110 -500
rect 6140 -530 6150 -500
rect 6015 -550 6065 -540
rect 6015 -580 6025 -550
rect 6055 -580 6065 -550
rect 6015 -590 6065 -580
rect 5930 -630 5940 -600
rect 5970 -630 5980 -600
rect 5930 -635 5980 -630
rect 6100 -600 6150 -530
rect 6270 -385 6320 -375
rect 6270 -415 6280 -385
rect 6310 -415 6320 -385
rect 6270 -440 6320 -415
rect 6270 -475 6280 -440
rect 6310 -475 6320 -440
rect 6270 -500 6320 -475
rect 6270 -530 6280 -500
rect 6310 -530 6320 -500
rect 6185 -550 6235 -540
rect 6185 -580 6195 -550
rect 6225 -580 6235 -550
rect 6185 -590 6235 -580
rect 6100 -630 6110 -600
rect 6140 -630 6150 -600
rect 6100 -635 6150 -630
rect 6270 -600 6320 -530
rect 6440 -385 6490 -375
rect 6440 -415 6450 -385
rect 6480 -415 6490 -385
rect 6440 -440 6490 -415
rect 6440 -475 6450 -440
rect 6480 -475 6490 -440
rect 6440 -500 6490 -475
rect 6440 -530 6450 -500
rect 6480 -530 6490 -500
rect 6355 -550 6405 -540
rect 6355 -580 6365 -550
rect 6395 -580 6405 -550
rect 6355 -590 6405 -580
rect 6270 -630 6280 -600
rect 6310 -630 6320 -600
rect 6270 -635 6320 -630
rect 6440 -600 6490 -530
rect 6610 -385 6660 -375
rect 6610 -415 6620 -385
rect 6650 -415 6660 -385
rect 6610 -440 6660 -415
rect 6610 -475 6620 -440
rect 6650 -475 6660 -440
rect 6610 -500 6660 -475
rect 6610 -530 6620 -500
rect 6650 -530 6660 -500
rect 6525 -550 6575 -540
rect 6525 -580 6535 -550
rect 6565 -580 6575 -550
rect 6525 -590 6575 -580
rect 6440 -630 6450 -600
rect 6480 -630 6490 -600
rect 6440 -635 6490 -630
rect 6610 -600 6660 -530
rect 6780 -385 6830 -375
rect 6780 -415 6790 -385
rect 6820 -415 6830 -385
rect 6780 -440 6830 -415
rect 6780 -475 6790 -440
rect 6820 -475 6830 -440
rect 6780 -500 6830 -475
rect 6780 -530 6790 -500
rect 6820 -530 6830 -500
rect 6695 -550 6745 -540
rect 6695 -580 6705 -550
rect 6735 -580 6745 -550
rect 6695 -590 6745 -580
rect 6610 -630 6620 -600
rect 6650 -630 6660 -600
rect 6610 -635 6660 -630
rect 6780 -600 6830 -530
rect 6950 -385 7000 -375
rect 6950 -415 6960 -385
rect 6990 -415 7000 -385
rect 6950 -440 7000 -415
rect 6950 -475 6960 -440
rect 6990 -475 7000 -440
rect 6950 -500 7000 -475
rect 6950 -530 6960 -500
rect 6990 -530 7000 -500
rect 6865 -550 6915 -540
rect 6865 -580 6875 -550
rect 6905 -580 6915 -550
rect 6865 -590 6915 -580
rect 6780 -630 6790 -600
rect 6820 -630 6830 -600
rect 6780 -635 6830 -630
rect 6950 -600 7000 -530
rect 7120 -385 7170 -375
rect 7120 -415 7130 -385
rect 7160 -415 7170 -385
rect 7120 -440 7170 -415
rect 7120 -475 7130 -440
rect 7160 -475 7170 -440
rect 7120 -500 7170 -475
rect 7120 -530 7130 -500
rect 7160 -530 7170 -500
rect 7035 -550 7085 -540
rect 7035 -580 7045 -550
rect 7075 -580 7085 -550
rect 7035 -590 7085 -580
rect 6950 -630 6960 -600
rect 6990 -630 7000 -600
rect 6950 -635 7000 -630
rect 7120 -600 7170 -530
rect 7290 -385 7340 -375
rect 7290 -415 7300 -385
rect 7330 -415 7340 -385
rect 7290 -440 7340 -415
rect 7290 -475 7300 -440
rect 7330 -475 7340 -440
rect 7290 -500 7340 -475
rect 7290 -530 7300 -500
rect 7330 -530 7340 -500
rect 7205 -550 7255 -540
rect 7205 -580 7215 -550
rect 7245 -580 7255 -550
rect 7205 -590 7255 -580
rect 7120 -630 7130 -600
rect 7160 -630 7170 -600
rect 7120 -635 7170 -630
rect 7290 -600 7340 -530
rect 7460 -385 7510 -375
rect 7460 -415 7470 -385
rect 7500 -415 7510 -385
rect 7460 -440 7510 -415
rect 7460 -475 7470 -440
rect 7500 -475 7510 -440
rect 7460 -500 7510 -475
rect 7460 -530 7470 -500
rect 7500 -530 7510 -500
rect 7375 -550 7425 -540
rect 7375 -580 7385 -550
rect 7415 -580 7425 -550
rect 7375 -590 7425 -580
rect 7290 -630 7300 -600
rect 7330 -630 7340 -600
rect 7290 -635 7340 -630
rect 7460 -600 7510 -530
rect 7630 -385 7680 -375
rect 7630 -415 7640 -385
rect 7670 -415 7680 -385
rect 7630 -440 7680 -415
rect 7630 -475 7640 -440
rect 7670 -475 7680 -440
rect 7630 -500 7680 -475
rect 7630 -530 7640 -500
rect 7670 -530 7680 -500
rect 7545 -550 7595 -540
rect 7545 -580 7555 -550
rect 7585 -580 7595 -550
rect 7545 -590 7595 -580
rect 7460 -630 7470 -600
rect 7500 -630 7510 -600
rect 7460 -635 7510 -630
rect 7630 -600 7680 -530
rect 7800 -385 7850 -375
rect 7800 -415 7810 -385
rect 7840 -415 7850 -385
rect 7800 -440 7850 -415
rect 7800 -475 7810 -440
rect 7840 -475 7850 -440
rect 7800 -500 7850 -475
rect 7800 -530 7810 -500
rect 7840 -530 7850 -500
rect 7715 -550 7765 -540
rect 7715 -580 7725 -550
rect 7755 -580 7765 -550
rect 7715 -590 7765 -580
rect 7630 -630 7640 -600
rect 7670 -630 7680 -600
rect 7630 -635 7680 -630
rect 7800 -600 7850 -530
rect 7970 -385 8020 -375
rect 7970 -415 7980 -385
rect 8010 -415 8020 -385
rect 7970 -440 8020 -415
rect 7970 -475 7980 -440
rect 8010 -475 8020 -440
rect 7970 -500 8020 -475
rect 7970 -530 7980 -500
rect 8010 -530 8020 -500
rect 7885 -550 7935 -540
rect 7885 -580 7895 -550
rect 7925 -580 7935 -550
rect 7885 -590 7935 -580
rect 7800 -630 7810 -600
rect 7840 -630 7850 -600
rect 7800 -635 7850 -630
rect 7970 -600 8020 -530
rect 8140 -385 8190 -375
rect 8140 -415 8150 -385
rect 8180 -415 8190 -385
rect 8140 -440 8190 -415
rect 8140 -475 8150 -440
rect 8180 -475 8190 -440
rect 8140 -500 8190 -475
rect 8140 -530 8150 -500
rect 8180 -530 8190 -500
rect 8055 -550 8105 -540
rect 8055 -580 8065 -550
rect 8095 -580 8105 -550
rect 8055 -590 8105 -580
rect 7970 -630 7980 -600
rect 8010 -630 8020 -600
rect 7970 -635 8020 -630
rect 8140 -600 8190 -530
rect 8310 -385 8360 -375
rect 8310 -415 8320 -385
rect 8350 -415 8360 -385
rect 8310 -440 8360 -415
rect 8310 -475 8320 -440
rect 8350 -475 8360 -440
rect 8310 -500 8360 -475
rect 8310 -530 8320 -500
rect 8350 -530 8360 -500
rect 8225 -550 8275 -540
rect 8225 -580 8235 -550
rect 8265 -580 8275 -550
rect 8225 -590 8275 -580
rect 8140 -630 8150 -600
rect 8180 -630 8190 -600
rect 8140 -635 8190 -630
rect 8310 -600 8360 -530
rect 8480 -385 8530 -375
rect 8480 -415 8490 -385
rect 8520 -415 8530 -385
rect 8480 -440 8530 -415
rect 8480 -475 8490 -440
rect 8520 -475 8530 -440
rect 8480 -500 8530 -475
rect 8480 -530 8490 -500
rect 8520 -530 8530 -500
rect 8395 -550 8445 -540
rect 8395 -580 8405 -550
rect 8435 -580 8445 -550
rect 8395 -590 8445 -580
rect 8310 -630 8320 -600
rect 8350 -630 8360 -600
rect 8310 -635 8360 -630
rect 8480 -600 8530 -530
rect 8650 -385 8700 -375
rect 8650 -415 8660 -385
rect 8690 -415 8700 -385
rect 8650 -440 8700 -415
rect 8650 -475 8660 -440
rect 8690 -475 8700 -440
rect 8650 -500 8700 -475
rect 8650 -530 8660 -500
rect 8690 -530 8700 -500
rect 8565 -550 8615 -540
rect 8565 -580 8575 -550
rect 8605 -580 8615 -550
rect 8565 -590 8615 -580
rect 8480 -630 8490 -600
rect 8520 -630 8530 -600
rect 8480 -635 8530 -630
rect 8650 -600 8700 -530
rect 8820 -385 8870 -375
rect 8820 -415 8830 -385
rect 8860 -415 8870 -385
rect 8820 -440 8870 -415
rect 8820 -475 8830 -440
rect 8860 -475 8870 -440
rect 8820 -500 8870 -475
rect 8820 -530 8830 -500
rect 8860 -530 8870 -500
rect 8735 -550 8785 -540
rect 8735 -580 8745 -550
rect 8775 -580 8785 -550
rect 8735 -590 8785 -580
rect 8650 -630 8660 -600
rect 8690 -630 8700 -600
rect 8650 -635 8700 -630
rect 8820 -600 8870 -530
rect 8990 -385 9040 -375
rect 8990 -415 9000 -385
rect 9030 -415 9040 -385
rect 8990 -440 9040 -415
rect 8990 -475 9000 -440
rect 9030 -475 9040 -440
rect 8990 -500 9040 -475
rect 8990 -530 9000 -500
rect 9030 -530 9040 -500
rect 8905 -550 8955 -540
rect 8905 -580 8915 -550
rect 8945 -580 8955 -550
rect 8905 -590 8955 -580
rect 8820 -630 8830 -600
rect 8860 -630 8870 -600
rect 8820 -635 8870 -630
rect 8990 -600 9040 -530
rect 9160 -385 9210 -375
rect 9160 -415 9170 -385
rect 9200 -415 9210 -385
rect 9160 -440 9210 -415
rect 9160 -475 9170 -440
rect 9200 -475 9210 -440
rect 9160 -500 9210 -475
rect 9160 -530 9170 -500
rect 9200 -530 9210 -500
rect 9075 -550 9125 -540
rect 9075 -580 9085 -550
rect 9115 -580 9125 -550
rect 9075 -590 9125 -580
rect 8990 -630 9000 -600
rect 9030 -630 9040 -600
rect 8990 -635 9040 -630
rect 9160 -600 9210 -530
rect 9330 -385 9380 -375
rect 9330 -415 9340 -385
rect 9370 -415 9380 -385
rect 9330 -440 9380 -415
rect 9330 -475 9340 -440
rect 9370 -475 9380 -440
rect 9330 -500 9380 -475
rect 9330 -530 9340 -500
rect 9370 -530 9380 -500
rect 9245 -550 9295 -540
rect 9245 -580 9255 -550
rect 9285 -580 9295 -550
rect 9245 -590 9295 -580
rect 9160 -630 9170 -600
rect 9200 -630 9210 -600
rect 9160 -635 9210 -630
rect 9330 -600 9380 -530
rect 9500 -385 9550 -375
rect 9500 -415 9510 -385
rect 9540 -415 9550 -385
rect 9500 -440 9550 -415
rect 9500 -475 9510 -440
rect 9540 -475 9550 -440
rect 9500 -500 9550 -475
rect 9500 -530 9510 -500
rect 9540 -530 9550 -500
rect 9415 -550 9465 -540
rect 9415 -580 9425 -550
rect 9455 -580 9465 -550
rect 9415 -590 9465 -580
rect 9330 -630 9340 -600
rect 9370 -630 9380 -600
rect 9330 -635 9380 -630
rect 9500 -600 9550 -530
rect 9670 -385 9720 -375
rect 9670 -415 9680 -385
rect 9710 -415 9720 -385
rect 9670 -440 9720 -415
rect 9670 -475 9680 -440
rect 9710 -475 9720 -440
rect 9670 -500 9720 -475
rect 9670 -530 9680 -500
rect 9710 -530 9720 -500
rect 9585 -550 9635 -540
rect 9585 -580 9595 -550
rect 9625 -580 9635 -550
rect 9585 -590 9635 -580
rect 9500 -630 9510 -600
rect 9540 -630 9550 -600
rect 9500 -635 9550 -630
rect 9670 -600 9720 -530
rect 9840 -385 9890 -375
rect 9840 -415 9850 -385
rect 9880 -415 9890 -385
rect 9840 -440 9890 -415
rect 9840 -475 9850 -440
rect 9880 -475 9890 -440
rect 9840 -500 9890 -475
rect 9840 -530 9850 -500
rect 9880 -530 9890 -500
rect 9755 -550 9805 -540
rect 9755 -580 9765 -550
rect 9795 -580 9805 -550
rect 9755 -590 9805 -580
rect 9670 -630 9680 -600
rect 9710 -630 9720 -600
rect 9670 -635 9720 -630
rect 9840 -600 9890 -530
rect 10010 -385 10060 -375
rect 10010 -415 10020 -385
rect 10050 -415 10060 -385
rect 10010 -440 10060 -415
rect 10010 -475 10020 -440
rect 10050 -475 10060 -440
rect 10010 -500 10060 -475
rect 10010 -530 10020 -500
rect 10050 -530 10060 -500
rect 9925 -550 9975 -540
rect 9925 -580 9935 -550
rect 9965 -580 9975 -550
rect 9925 -590 9975 -580
rect 9840 -630 9850 -600
rect 9880 -630 9890 -600
rect 9840 -635 9890 -630
rect 10010 -600 10060 -530
rect 10180 -385 10230 -375
rect 10180 -415 10190 -385
rect 10220 -415 10230 -385
rect 10180 -440 10230 -415
rect 10180 -475 10190 -440
rect 10220 -475 10230 -440
rect 10180 -500 10230 -475
rect 10180 -530 10190 -500
rect 10220 -530 10230 -500
rect 10095 -550 10145 -540
rect 10095 -580 10105 -550
rect 10135 -580 10145 -550
rect 10095 -590 10145 -580
rect 10010 -630 10020 -600
rect 10050 -630 10060 -600
rect 10010 -635 10060 -630
rect 10180 -600 10230 -530
rect 10350 -385 10400 -375
rect 10350 -415 10360 -385
rect 10390 -415 10400 -385
rect 10350 -440 10400 -415
rect 10350 -475 10360 -440
rect 10390 -475 10400 -440
rect 10350 -500 10400 -475
rect 10350 -530 10360 -500
rect 10390 -530 10400 -500
rect 10265 -550 10315 -540
rect 10265 -580 10275 -550
rect 10305 -580 10315 -550
rect 10265 -590 10315 -580
rect 10180 -630 10190 -600
rect 10220 -630 10230 -600
rect 10180 -635 10230 -630
rect 10350 -600 10400 -530
rect 10520 -385 10570 -375
rect 10520 -415 10530 -385
rect 10560 -415 10570 -385
rect 10520 -440 10570 -415
rect 10520 -475 10530 -440
rect 10560 -475 10570 -440
rect 10520 -500 10570 -475
rect 10520 -530 10530 -500
rect 10560 -530 10570 -500
rect 10435 -550 10485 -540
rect 10435 -580 10445 -550
rect 10475 -580 10485 -550
rect 10435 -590 10485 -580
rect 10350 -630 10360 -600
rect 10390 -630 10400 -600
rect 10350 -635 10400 -630
rect 10520 -600 10570 -530
rect 10690 -385 10740 -375
rect 10690 -415 10700 -385
rect 10730 -415 10740 -385
rect 10690 -440 10740 -415
rect 10690 -475 10700 -440
rect 10730 -475 10740 -440
rect 10690 -500 10740 -475
rect 10690 -530 10700 -500
rect 10730 -530 10740 -500
rect 10605 -550 10655 -540
rect 10605 -580 10615 -550
rect 10645 -580 10655 -550
rect 10605 -590 10655 -580
rect 10520 -630 10530 -600
rect 10560 -630 10570 -600
rect 10520 -635 10570 -630
rect 10690 -600 10740 -530
rect 10860 -385 10910 -375
rect 10860 -415 10870 -385
rect 10900 -415 10910 -385
rect 10860 -440 10910 -415
rect 10860 -475 10870 -440
rect 10900 -475 10910 -440
rect 10860 -500 10910 -475
rect 10860 -530 10870 -500
rect 10900 -530 10910 -500
rect 10775 -550 10825 -540
rect 10775 -580 10785 -550
rect 10815 -580 10825 -550
rect 10775 -590 10825 -580
rect 10690 -630 10700 -600
rect 10730 -630 10740 -600
rect 10690 -635 10740 -630
rect 10860 -600 10910 -530
rect 11030 -385 11080 -375
rect 11030 -415 11040 -385
rect 11070 -415 11080 -385
rect 11030 -440 11080 -415
rect 11030 -475 11040 -440
rect 11070 -475 11080 -440
rect 11030 -500 11080 -475
rect 11030 -530 11040 -500
rect 11070 -530 11080 -500
rect 10945 -550 10995 -540
rect 10945 -580 10955 -550
rect 10985 -580 10995 -550
rect 10945 -590 10995 -580
rect 10860 -630 10870 -600
rect 10900 -630 10910 -600
rect 10860 -635 10910 -630
rect 11030 -600 11080 -530
rect 11200 -385 11250 -375
rect 11200 -415 11210 -385
rect 11240 -415 11250 -385
rect 11200 -440 11250 -415
rect 11200 -475 11210 -440
rect 11240 -475 11250 -440
rect 11200 -500 11250 -475
rect 11200 -530 11210 -500
rect 11240 -530 11250 -500
rect 11115 -550 11165 -540
rect 11115 -580 11125 -550
rect 11155 -580 11165 -550
rect 11115 -590 11165 -580
rect 11030 -630 11040 -600
rect 11070 -630 11080 -600
rect 11030 -635 11080 -630
rect 11200 -600 11250 -530
rect 11370 -385 11420 -375
rect 11370 -415 11380 -385
rect 11410 -415 11420 -385
rect 11370 -440 11420 -415
rect 11370 -475 11380 -440
rect 11410 -475 11420 -440
rect 11370 -500 11420 -475
rect 11370 -530 11380 -500
rect 11410 -530 11420 -500
rect 11285 -550 11335 -540
rect 11285 -580 11295 -550
rect 11325 -580 11335 -550
rect 11285 -590 11335 -580
rect 11200 -630 11210 -600
rect 11240 -630 11250 -600
rect 11200 -635 11250 -630
rect 11370 -600 11420 -530
rect 11540 -385 11590 -375
rect 11540 -415 11550 -385
rect 11580 -415 11590 -385
rect 11540 -440 11590 -415
rect 11540 -475 11550 -440
rect 11580 -475 11590 -440
rect 11540 -500 11590 -475
rect 11540 -530 11550 -500
rect 11580 -530 11590 -500
rect 11455 -550 11505 -540
rect 11455 -580 11465 -550
rect 11495 -580 11505 -550
rect 11455 -590 11505 -580
rect 11370 -630 11380 -600
rect 11410 -630 11420 -600
rect 11370 -635 11420 -630
rect 11540 -600 11590 -530
rect 11710 -385 11760 -375
rect 11710 -415 11720 -385
rect 11750 -415 11760 -385
rect 11710 -440 11760 -415
rect 11710 -475 11720 -440
rect 11750 -475 11760 -440
rect 11710 -500 11760 -475
rect 11710 -530 11720 -500
rect 11750 -530 11760 -500
rect 11625 -550 11675 -540
rect 11625 -580 11635 -550
rect 11665 -580 11675 -550
rect 11625 -590 11675 -580
rect 11540 -630 11550 -600
rect 11580 -630 11590 -600
rect 11540 -635 11590 -630
rect 11710 -600 11760 -530
rect 11880 -385 11930 -375
rect 11880 -415 11890 -385
rect 11920 -415 11930 -385
rect 11880 -440 11930 -415
rect 11880 -475 11890 -440
rect 11920 -475 11930 -440
rect 11880 -500 11930 -475
rect 11880 -530 11890 -500
rect 11920 -530 11930 -500
rect 11795 -550 11845 -540
rect 11795 -580 11805 -550
rect 11835 -580 11845 -550
rect 11795 -590 11845 -580
rect 11710 -630 11720 -600
rect 11750 -630 11760 -600
rect 11710 -635 11760 -630
rect 11880 -600 11930 -530
rect 12050 -385 12100 -375
rect 12050 -415 12060 -385
rect 12090 -415 12100 -385
rect 12050 -440 12100 -415
rect 12050 -475 12060 -440
rect 12090 -475 12100 -440
rect 12050 -500 12100 -475
rect 12050 -530 12060 -500
rect 12090 -530 12100 -500
rect 11965 -550 12015 -540
rect 11965 -580 11975 -550
rect 12005 -580 12015 -550
rect 11965 -590 12015 -580
rect 11880 -630 11890 -600
rect 11920 -630 11930 -600
rect 11880 -635 11930 -630
rect 12050 -600 12100 -530
rect 12220 -385 12270 -375
rect 12220 -415 12230 -385
rect 12260 -415 12270 -385
rect 12220 -440 12270 -415
rect 12220 -475 12230 -440
rect 12260 -475 12270 -440
rect 12220 -500 12270 -475
rect 12220 -530 12230 -500
rect 12260 -530 12270 -500
rect 12135 -550 12185 -540
rect 12135 -580 12145 -550
rect 12175 -580 12185 -550
rect 12135 -590 12185 -580
rect 12050 -630 12060 -600
rect 12090 -630 12100 -600
rect 12050 -635 12100 -630
rect 12220 -600 12270 -530
rect 12390 -385 12440 -375
rect 12390 -415 12400 -385
rect 12430 -415 12440 -385
rect 12390 -440 12440 -415
rect 12390 -475 12400 -440
rect 12430 -475 12440 -440
rect 12390 -500 12440 -475
rect 12390 -530 12400 -500
rect 12430 -530 12440 -500
rect 12305 -550 12355 -540
rect 12305 -580 12315 -550
rect 12345 -580 12355 -550
rect 12305 -590 12355 -580
rect 12220 -630 12230 -600
rect 12260 -630 12270 -600
rect 12220 -635 12270 -630
rect 12390 -600 12440 -530
rect 12560 -385 12610 -375
rect 12560 -415 12570 -385
rect 12600 -415 12610 -385
rect 12560 -440 12610 -415
rect 12560 -475 12570 -440
rect 12600 -475 12610 -440
rect 12560 -500 12610 -475
rect 12560 -530 12570 -500
rect 12600 -530 12610 -500
rect 12475 -550 12525 -540
rect 12475 -580 12485 -550
rect 12515 -580 12525 -550
rect 12475 -590 12525 -580
rect 12390 -630 12400 -600
rect 12430 -630 12440 -600
rect 12390 -635 12440 -630
rect 12560 -600 12610 -530
rect 12730 -385 12780 -375
rect 12730 -415 12740 -385
rect 12770 -415 12780 -385
rect 12730 -440 12780 -415
rect 12730 -475 12740 -440
rect 12770 -475 12780 -440
rect 12730 -500 12780 -475
rect 12730 -530 12740 -500
rect 12770 -530 12780 -500
rect 12645 -550 12695 -540
rect 12645 -580 12655 -550
rect 12685 -580 12695 -550
rect 12645 -590 12695 -580
rect 12560 -630 12570 -600
rect 12600 -630 12610 -600
rect 12560 -635 12610 -630
rect 12730 -600 12780 -530
rect 12900 -385 12950 -375
rect 12900 -415 12910 -385
rect 12940 -415 12950 -385
rect 12900 -440 12950 -415
rect 12900 -475 12910 -440
rect 12940 -475 12950 -440
rect 12900 -500 12950 -475
rect 12900 -530 12910 -500
rect 12940 -530 12950 -500
rect 12815 -550 12865 -540
rect 12815 -580 12825 -550
rect 12855 -580 12865 -550
rect 12815 -590 12865 -580
rect 12730 -630 12740 -600
rect 12770 -630 12780 -600
rect 12730 -635 12780 -630
rect 12900 -600 12950 -530
rect 13070 -385 13120 -375
rect 13070 -415 13080 -385
rect 13110 -415 13120 -385
rect 13070 -440 13120 -415
rect 13070 -475 13080 -440
rect 13110 -475 13120 -440
rect 13070 -500 13120 -475
rect 13070 -530 13080 -500
rect 13110 -530 13120 -500
rect 12985 -550 13035 -540
rect 12985 -580 12995 -550
rect 13025 -580 13035 -550
rect 12985 -590 13035 -580
rect 12900 -630 12910 -600
rect 12940 -630 12950 -600
rect 12900 -635 12950 -630
rect 13070 -600 13120 -530
rect 13240 -385 13290 -375
rect 13240 -415 13250 -385
rect 13280 -415 13290 -385
rect 13240 -440 13290 -415
rect 13240 -475 13250 -440
rect 13280 -475 13290 -440
rect 13240 -500 13290 -475
rect 13240 -530 13250 -500
rect 13280 -530 13290 -500
rect 13155 -550 13205 -540
rect 13155 -580 13165 -550
rect 13195 -580 13205 -550
rect 13155 -590 13205 -580
rect 13070 -630 13080 -600
rect 13110 -630 13120 -600
rect 13070 -635 13120 -630
rect 13240 -600 13290 -530
rect 13410 -385 13460 -375
rect 13410 -415 13420 -385
rect 13450 -415 13460 -385
rect 13410 -440 13460 -415
rect 13410 -475 13420 -440
rect 13450 -475 13460 -440
rect 13410 -500 13460 -475
rect 13410 -530 13420 -500
rect 13450 -530 13460 -500
rect 13325 -550 13375 -540
rect 13325 -580 13335 -550
rect 13365 -580 13375 -550
rect 13325 -590 13375 -580
rect 13240 -630 13250 -600
rect 13280 -630 13290 -600
rect 13240 -635 13290 -630
rect 13410 -600 13460 -530
rect 13580 -385 13630 -375
rect 13580 -415 13590 -385
rect 13620 -415 13630 -385
rect 13580 -440 13630 -415
rect 13580 -475 13590 -440
rect 13620 -475 13630 -440
rect 13580 -500 13630 -475
rect 13580 -530 13590 -500
rect 13620 -530 13630 -500
rect 13495 -550 13545 -540
rect 13495 -580 13505 -550
rect 13535 -580 13545 -550
rect 13495 -590 13545 -580
rect 13410 -630 13420 -600
rect 13450 -630 13460 -600
rect 13410 -635 13460 -630
rect 13580 -600 13630 -530
rect 13750 -385 13800 -375
rect 13750 -415 13760 -385
rect 13790 -415 13800 -385
rect 13750 -440 13800 -415
rect 13750 -475 13760 -440
rect 13790 -475 13800 -440
rect 13750 -500 13800 -475
rect 13750 -530 13760 -500
rect 13790 -530 13800 -500
rect 13665 -550 13715 -540
rect 13665 -580 13675 -550
rect 13705 -580 13715 -550
rect 13665 -590 13715 -580
rect 13580 -630 13590 -600
rect 13620 -630 13630 -600
rect 13580 -635 13630 -630
rect 13750 -600 13800 -530
rect 13920 -385 13970 -375
rect 13920 -415 13930 -385
rect 13960 -415 13970 -385
rect 13920 -440 13970 -415
rect 13920 -475 13930 -440
rect 13960 -475 13970 -440
rect 13920 -500 13970 -475
rect 13920 -530 13930 -500
rect 13960 -530 13970 -500
rect 13835 -550 13885 -540
rect 13835 -580 13845 -550
rect 13875 -580 13885 -550
rect 13835 -590 13885 -580
rect 13750 -630 13760 -600
rect 13790 -630 13800 -600
rect 13750 -635 13800 -630
rect 13920 -600 13970 -530
rect 14090 -385 14140 -375
rect 14090 -415 14100 -385
rect 14130 -415 14140 -385
rect 14090 -440 14140 -415
rect 14090 -475 14100 -440
rect 14130 -475 14140 -440
rect 14090 -500 14140 -475
rect 14090 -530 14100 -500
rect 14130 -530 14140 -500
rect 14005 -550 14055 -540
rect 14005 -580 14015 -550
rect 14045 -580 14055 -550
rect 14005 -590 14055 -580
rect 13920 -630 13930 -600
rect 13960 -630 13970 -600
rect 13920 -635 13970 -630
rect 14090 -600 14140 -530
rect 14260 -385 14310 -375
rect 14260 -415 14270 -385
rect 14300 -415 14310 -385
rect 14260 -440 14310 -415
rect 14260 -475 14270 -440
rect 14300 -475 14310 -440
rect 14260 -500 14310 -475
rect 14260 -530 14270 -500
rect 14300 -530 14310 -500
rect 14175 -550 14225 -540
rect 14175 -580 14185 -550
rect 14215 -580 14225 -550
rect 14175 -590 14225 -580
rect 14090 -630 14100 -600
rect 14130 -630 14140 -600
rect 14090 -635 14140 -630
rect 14260 -600 14310 -530
rect 14430 -385 14480 -375
rect 14430 -415 14440 -385
rect 14470 -415 14480 -385
rect 14430 -440 14480 -415
rect 14430 -475 14440 -440
rect 14470 -475 14480 -440
rect 14430 -500 14480 -475
rect 14430 -530 14440 -500
rect 14470 -530 14480 -500
rect 14345 -550 14395 -540
rect 14345 -580 14355 -550
rect 14385 -580 14395 -550
rect 14345 -590 14395 -580
rect 14260 -630 14270 -600
rect 14300 -630 14310 -600
rect 14260 -635 14310 -630
rect 14430 -600 14480 -530
rect 14600 -385 14650 -375
rect 14600 -415 14610 -385
rect 14640 -415 14650 -385
rect 14600 -440 14650 -415
rect 14600 -475 14610 -440
rect 14640 -475 14650 -440
rect 14600 -500 14650 -475
rect 14600 -530 14610 -500
rect 14640 -530 14650 -500
rect 14515 -550 14565 -540
rect 14515 -580 14525 -550
rect 14555 -580 14565 -550
rect 14515 -590 14565 -580
rect 14430 -630 14440 -600
rect 14470 -630 14480 -600
rect 14430 -635 14480 -630
rect 14600 -600 14650 -530
rect 14770 -385 14820 -375
rect 14770 -415 14780 -385
rect 14810 -415 14820 -385
rect 14770 -440 14820 -415
rect 14770 -475 14780 -440
rect 14810 -475 14820 -440
rect 14770 -500 14820 -475
rect 14770 -530 14780 -500
rect 14810 -530 14820 -500
rect 14685 -550 14735 -540
rect 14685 -580 14695 -550
rect 14725 -580 14735 -550
rect 14685 -590 14735 -580
rect 14600 -630 14610 -600
rect 14640 -630 14650 -600
rect 14600 -635 14650 -630
rect 14770 -600 14820 -530
rect 14940 -385 14990 -375
rect 14940 -415 14950 -385
rect 14980 -415 14990 -385
rect 14940 -440 14990 -415
rect 14940 -475 14950 -440
rect 14980 -475 14990 -440
rect 14940 -500 14990 -475
rect 14940 -530 14950 -500
rect 14980 -530 14990 -500
rect 14855 -550 14905 -540
rect 14855 -580 14865 -550
rect 14895 -580 14905 -550
rect 14855 -590 14905 -580
rect 14770 -630 14780 -600
rect 14810 -630 14820 -600
rect 14770 -635 14820 -630
rect 14940 -600 14990 -530
rect 15110 -385 15160 -375
rect 15110 -415 15120 -385
rect 15150 -415 15160 -385
rect 15110 -440 15160 -415
rect 15110 -475 15120 -440
rect 15150 -475 15160 -440
rect 15110 -500 15160 -475
rect 15110 -530 15120 -500
rect 15150 -530 15160 -500
rect 15025 -550 15075 -540
rect 15025 -580 15035 -550
rect 15065 -580 15075 -550
rect 15025 -590 15075 -580
rect 14940 -630 14950 -600
rect 14980 -630 14990 -600
rect 14940 -635 14990 -630
rect 15110 -600 15160 -530
rect 15280 -385 15330 -375
rect 15280 -415 15290 -385
rect 15320 -415 15330 -385
rect 15280 -440 15330 -415
rect 15280 -475 15290 -440
rect 15320 -475 15330 -440
rect 15280 -500 15330 -475
rect 15280 -530 15290 -500
rect 15320 -530 15330 -500
rect 15195 -550 15245 -540
rect 15195 -580 15205 -550
rect 15235 -580 15245 -550
rect 15195 -590 15245 -580
rect 15110 -630 15120 -600
rect 15150 -630 15160 -600
rect 15110 -635 15160 -630
rect 15280 -600 15330 -530
rect 15450 -385 15500 -375
rect 15450 -415 15460 -385
rect 15490 -415 15500 -385
rect 15450 -440 15500 -415
rect 15450 -475 15460 -440
rect 15490 -475 15500 -440
rect 15450 -500 15500 -475
rect 15450 -530 15460 -500
rect 15490 -530 15500 -500
rect 15365 -550 15415 -540
rect 15365 -580 15375 -550
rect 15405 -580 15415 -550
rect 15365 -590 15415 -580
rect 15280 -630 15290 -600
rect 15320 -630 15330 -600
rect 15280 -635 15330 -630
rect 15450 -600 15500 -530
rect 15620 -385 15670 -375
rect 15620 -415 15630 -385
rect 15660 -415 15670 -385
rect 15620 -440 15670 -415
rect 15620 -475 15630 -440
rect 15660 -475 15670 -440
rect 15620 -500 15670 -475
rect 15620 -530 15630 -500
rect 15660 -530 15670 -500
rect 15535 -550 15585 -540
rect 15535 -580 15545 -550
rect 15575 -580 15585 -550
rect 15535 -590 15585 -580
rect 15450 -630 15460 -600
rect 15490 -630 15500 -600
rect 15450 -635 15500 -630
rect 15620 -600 15670 -530
rect 15790 -385 15840 -375
rect 15790 -415 15800 -385
rect 15830 -415 15840 -385
rect 15790 -440 15840 -415
rect 15790 -475 15800 -440
rect 15830 -475 15840 -440
rect 15790 -500 15840 -475
rect 15790 -530 15800 -500
rect 15830 -530 15840 -500
rect 15705 -550 15755 -540
rect 15705 -580 15715 -550
rect 15745 -580 15755 -550
rect 15705 -590 15755 -580
rect 15620 -630 15630 -600
rect 15660 -630 15670 -600
rect 15620 -635 15670 -630
rect 15790 -600 15840 -530
rect 15960 -385 16010 -375
rect 15960 -415 15970 -385
rect 16000 -415 16010 -385
rect 15960 -440 16010 -415
rect 15960 -475 15970 -440
rect 16000 -475 16010 -440
rect 15960 -500 16010 -475
rect 15960 -530 15970 -500
rect 16000 -530 16010 -500
rect 15875 -550 15925 -540
rect 15875 -580 15885 -550
rect 15915 -580 15925 -550
rect 15875 -590 15925 -580
rect 15790 -630 15800 -600
rect 15830 -630 15840 -600
rect 15790 -635 15840 -630
rect 15960 -600 16010 -530
rect 16130 -385 16180 -375
rect 16130 -415 16140 -385
rect 16170 -415 16180 -385
rect 16130 -440 16180 -415
rect 16130 -475 16140 -440
rect 16170 -475 16180 -440
rect 16130 -500 16180 -475
rect 16130 -530 16140 -500
rect 16170 -530 16180 -500
rect 16045 -550 16095 -540
rect 16045 -580 16055 -550
rect 16085 -580 16095 -550
rect 16045 -590 16095 -580
rect 15960 -630 15970 -600
rect 16000 -630 16010 -600
rect 15960 -635 16010 -630
rect 16130 -600 16180 -530
rect 16300 -385 16350 -375
rect 16300 -415 16310 -385
rect 16340 -415 16350 -385
rect 16300 -440 16350 -415
rect 16300 -475 16310 -440
rect 16340 -475 16350 -440
rect 16300 -500 16350 -475
rect 16300 -530 16310 -500
rect 16340 -530 16350 -500
rect 16215 -550 16265 -540
rect 16215 -580 16225 -550
rect 16255 -580 16265 -550
rect 16215 -590 16265 -580
rect 16130 -630 16140 -600
rect 16170 -630 16180 -600
rect 16130 -635 16180 -630
rect 16300 -600 16350 -530
rect 16470 -385 16520 -375
rect 16470 -415 16480 -385
rect 16510 -415 16520 -385
rect 16470 -440 16520 -415
rect 16470 -475 16480 -440
rect 16510 -475 16520 -440
rect 16470 -500 16520 -475
rect 16470 -530 16480 -500
rect 16510 -530 16520 -500
rect 16385 -550 16435 -540
rect 16385 -580 16395 -550
rect 16425 -580 16435 -550
rect 16385 -590 16435 -580
rect 16300 -630 16310 -600
rect 16340 -630 16350 -600
rect 16300 -635 16350 -630
rect 16470 -600 16520 -530
rect 16640 -385 16690 -375
rect 16640 -415 16650 -385
rect 16680 -415 16690 -385
rect 16640 -440 16690 -415
rect 16640 -475 16650 -440
rect 16680 -475 16690 -440
rect 16640 -500 16690 -475
rect 16640 -530 16650 -500
rect 16680 -530 16690 -500
rect 16555 -550 16605 -540
rect 16555 -580 16565 -550
rect 16595 -580 16605 -550
rect 16555 -590 16605 -580
rect 16470 -630 16480 -600
rect 16510 -630 16520 -600
rect 16470 -635 16520 -630
rect 16640 -600 16690 -530
rect 16810 -385 16860 -375
rect 16810 -415 16820 -385
rect 16850 -415 16860 -385
rect 16810 -440 16860 -415
rect 16810 -475 16820 -440
rect 16850 -475 16860 -440
rect 16810 -500 16860 -475
rect 16810 -530 16820 -500
rect 16850 -530 16860 -500
rect 16725 -550 16775 -540
rect 16725 -580 16735 -550
rect 16765 -580 16775 -550
rect 16725 -590 16775 -580
rect 16640 -630 16650 -600
rect 16680 -630 16690 -600
rect 16640 -635 16690 -630
rect 16810 -600 16860 -530
rect 16980 -385 17030 -375
rect 16980 -415 16990 -385
rect 17020 -415 17030 -385
rect 16980 -440 17030 -415
rect 16980 -475 16990 -440
rect 17020 -475 17030 -440
rect 16980 -500 17030 -475
rect 16980 -530 16990 -500
rect 17020 -530 17030 -500
rect 16895 -550 16945 -540
rect 16895 -580 16905 -550
rect 16935 -580 16945 -550
rect 16895 -590 16945 -580
rect 16810 -630 16820 -600
rect 16850 -630 16860 -600
rect 16810 -635 16860 -630
rect 16980 -600 17030 -530
rect 17150 -385 17200 -375
rect 17150 -415 17160 -385
rect 17190 -415 17200 -385
rect 17150 -440 17200 -415
rect 17150 -475 17160 -440
rect 17190 -475 17200 -440
rect 17150 -500 17200 -475
rect 17150 -530 17160 -500
rect 17190 -530 17200 -500
rect 17065 -550 17115 -540
rect 17065 -580 17075 -550
rect 17105 -580 17115 -550
rect 17065 -590 17115 -580
rect 16980 -630 16990 -600
rect 17020 -630 17030 -600
rect 16980 -635 17030 -630
rect 17150 -600 17200 -530
rect 17320 -385 17370 -375
rect 17320 -415 17330 -385
rect 17360 -415 17370 -385
rect 17320 -440 17370 -415
rect 17320 -475 17330 -440
rect 17360 -475 17370 -440
rect 17320 -500 17370 -475
rect 17320 -530 17330 -500
rect 17360 -530 17370 -500
rect 17235 -550 17285 -540
rect 17235 -580 17245 -550
rect 17275 -580 17285 -550
rect 17235 -590 17285 -580
rect 17150 -630 17160 -600
rect 17190 -630 17200 -600
rect 17150 -635 17200 -630
rect 17320 -600 17370 -530
rect 17490 -385 17540 -375
rect 17490 -415 17500 -385
rect 17530 -415 17540 -385
rect 17490 -440 17540 -415
rect 17490 -475 17500 -440
rect 17530 -475 17540 -440
rect 17490 -500 17540 -475
rect 17490 -530 17500 -500
rect 17530 -530 17540 -500
rect 17405 -550 17455 -540
rect 17405 -580 17415 -550
rect 17445 -580 17455 -550
rect 17405 -590 17455 -580
rect 17320 -630 17330 -600
rect 17360 -630 17370 -600
rect 17320 -635 17370 -630
rect 17490 -600 17540 -530
rect 17660 -385 17710 -375
rect 17660 -415 17670 -385
rect 17700 -415 17710 -385
rect 17660 -440 17710 -415
rect 17660 -475 17670 -440
rect 17700 -475 17710 -440
rect 17660 -500 17710 -475
rect 17660 -530 17670 -500
rect 17700 -530 17710 -500
rect 17575 -550 17625 -540
rect 17575 -580 17585 -550
rect 17615 -580 17625 -550
rect 17575 -590 17625 -580
rect 17490 -630 17500 -600
rect 17530 -630 17540 -600
rect 17490 -635 17540 -630
rect 17660 -600 17710 -530
rect 17830 -385 17880 -375
rect 17830 -415 17840 -385
rect 17870 -415 17880 -385
rect 17830 -440 17880 -415
rect 17830 -475 17840 -440
rect 17870 -475 17880 -440
rect 17830 -500 17880 -475
rect 17830 -530 17840 -500
rect 17870 -530 17880 -500
rect 17745 -550 17795 -540
rect 17745 -580 17755 -550
rect 17785 -580 17795 -550
rect 17745 -590 17795 -580
rect 17660 -630 17670 -600
rect 17700 -630 17710 -600
rect 17660 -635 17710 -630
rect 17830 -600 17880 -530
rect 18000 -385 18050 -375
rect 18000 -415 18010 -385
rect 18040 -415 18050 -385
rect 18000 -440 18050 -415
rect 18000 -475 18010 -440
rect 18040 -475 18050 -440
rect 18000 -500 18050 -475
rect 18000 -530 18010 -500
rect 18040 -530 18050 -500
rect 17915 -550 17965 -540
rect 17915 -580 17925 -550
rect 17955 -580 17965 -550
rect 17915 -590 17965 -580
rect 17830 -630 17840 -600
rect 17870 -630 17880 -600
rect 17830 -635 17880 -630
rect 18000 -600 18050 -530
rect 18170 -385 18220 -375
rect 18170 -415 18180 -385
rect 18210 -415 18220 -385
rect 18170 -440 18220 -415
rect 18170 -475 18180 -440
rect 18210 -475 18220 -440
rect 18170 -500 18220 -475
rect 18170 -530 18180 -500
rect 18210 -530 18220 -500
rect 18085 -550 18135 -540
rect 18085 -580 18095 -550
rect 18125 -580 18135 -550
rect 18085 -590 18135 -580
rect 18000 -630 18010 -600
rect 18040 -630 18050 -600
rect 18000 -635 18050 -630
rect 18170 -600 18220 -530
rect 18340 -385 18390 -375
rect 18340 -415 18350 -385
rect 18380 -415 18390 -385
rect 18340 -440 18390 -415
rect 18340 -475 18350 -440
rect 18380 -475 18390 -440
rect 18340 -500 18390 -475
rect 18340 -530 18350 -500
rect 18380 -530 18390 -500
rect 18255 -550 18305 -540
rect 18255 -580 18265 -550
rect 18295 -580 18305 -550
rect 18255 -590 18305 -580
rect 18170 -630 18180 -600
rect 18210 -630 18220 -600
rect 18170 -635 18220 -630
rect 18340 -600 18390 -530
rect 18510 -385 18560 -375
rect 18510 -415 18520 -385
rect 18550 -415 18560 -385
rect 18510 -440 18560 -415
rect 18510 -475 18520 -440
rect 18550 -475 18560 -440
rect 18510 -500 18560 -475
rect 18510 -530 18520 -500
rect 18550 -530 18560 -500
rect 18425 -550 18475 -540
rect 18425 -580 18435 -550
rect 18465 -580 18475 -550
rect 18425 -590 18475 -580
rect 18340 -630 18350 -600
rect 18380 -630 18390 -600
rect 18340 -635 18390 -630
rect 18510 -600 18560 -530
rect 18680 -385 18730 -375
rect 18680 -415 18690 -385
rect 18720 -415 18730 -385
rect 18680 -440 18730 -415
rect 18680 -475 18690 -440
rect 18720 -475 18730 -440
rect 18680 -500 18730 -475
rect 18680 -530 18690 -500
rect 18720 -530 18730 -500
rect 18595 -550 18645 -540
rect 18595 -580 18605 -550
rect 18635 -580 18645 -550
rect 18595 -590 18645 -580
rect 18510 -630 18520 -600
rect 18550 -630 18560 -600
rect 18510 -635 18560 -630
rect 18680 -600 18730 -530
rect 18850 -385 18900 -375
rect 18850 -415 18860 -385
rect 18890 -415 18900 -385
rect 18850 -440 18900 -415
rect 18850 -475 18860 -440
rect 18890 -475 18900 -440
rect 18850 -500 18900 -475
rect 18850 -530 18860 -500
rect 18890 -530 18900 -500
rect 18765 -550 18815 -540
rect 18765 -580 18775 -550
rect 18805 -580 18815 -550
rect 18765 -590 18815 -580
rect 18680 -630 18690 -600
rect 18720 -630 18730 -600
rect 18680 -635 18730 -630
rect 18850 -600 18900 -530
rect 19020 -385 19070 -375
rect 19020 -415 19030 -385
rect 19060 -415 19070 -385
rect 19020 -440 19070 -415
rect 19020 -475 19030 -440
rect 19060 -475 19070 -440
rect 19020 -500 19070 -475
rect 19020 -530 19030 -500
rect 19060 -530 19070 -500
rect 18935 -550 18985 -540
rect 18935 -580 18945 -550
rect 18975 -580 18985 -550
rect 18935 -590 18985 -580
rect 18850 -630 18860 -600
rect 18890 -630 18900 -600
rect 18850 -635 18900 -630
rect 19020 -600 19070 -530
rect 19190 -385 19240 -375
rect 19190 -415 19200 -385
rect 19230 -415 19240 -385
rect 19190 -440 19240 -415
rect 19190 -475 19200 -440
rect 19230 -475 19240 -440
rect 19190 -500 19240 -475
rect 19190 -530 19200 -500
rect 19230 -530 19240 -500
rect 19105 -550 19155 -540
rect 19105 -580 19115 -550
rect 19145 -580 19155 -550
rect 19105 -590 19155 -580
rect 19020 -630 19030 -600
rect 19060 -630 19070 -600
rect 19020 -635 19070 -630
rect 19190 -600 19240 -530
rect 19360 -385 19410 -375
rect 19360 -415 19370 -385
rect 19400 -415 19410 -385
rect 19360 -440 19410 -415
rect 19360 -475 19370 -440
rect 19400 -475 19410 -440
rect 19360 -500 19410 -475
rect 19360 -530 19370 -500
rect 19400 -530 19410 -500
rect 19275 -550 19325 -540
rect 19275 -580 19285 -550
rect 19315 -580 19325 -550
rect 19275 -590 19325 -580
rect 19190 -630 19200 -600
rect 19230 -630 19240 -600
rect 19190 -635 19240 -630
rect 19360 -600 19410 -530
rect 19530 -385 19580 -375
rect 19530 -415 19540 -385
rect 19570 -415 19580 -385
rect 19530 -440 19580 -415
rect 19530 -475 19540 -440
rect 19570 -475 19580 -440
rect 19530 -500 19580 -475
rect 19530 -530 19540 -500
rect 19570 -530 19580 -500
rect 19445 -550 19495 -540
rect 19445 -580 19455 -550
rect 19485 -580 19495 -550
rect 19445 -590 19495 -580
rect 19360 -630 19370 -600
rect 19400 -630 19410 -600
rect 19360 -635 19410 -630
rect 19530 -600 19580 -530
rect 19700 -385 19750 -375
rect 19700 -415 19710 -385
rect 19740 -415 19750 -385
rect 19700 -440 19750 -415
rect 19700 -475 19710 -440
rect 19740 -475 19750 -440
rect 19700 -500 19750 -475
rect 19700 -530 19710 -500
rect 19740 -530 19750 -500
rect 19615 -550 19665 -540
rect 19615 -580 19625 -550
rect 19655 -580 19665 -550
rect 19615 -590 19665 -580
rect 19530 -630 19540 -600
rect 19570 -630 19580 -600
rect 19530 -635 19580 -630
rect 19700 -600 19750 -530
rect 19870 -385 19920 -375
rect 19870 -415 19880 -385
rect 19910 -415 19920 -385
rect 19870 -440 19920 -415
rect 19870 -475 19880 -440
rect 19910 -475 19920 -440
rect 19870 -500 19920 -475
rect 19870 -530 19880 -500
rect 19910 -530 19920 -500
rect 19785 -550 19835 -540
rect 19785 -580 19795 -550
rect 19825 -580 19835 -550
rect 19785 -590 19835 -580
rect 19700 -630 19710 -600
rect 19740 -630 19750 -600
rect 19700 -635 19750 -630
rect 19870 -600 19920 -530
rect 20040 -385 20090 -375
rect 20040 -415 20050 -385
rect 20080 -415 20090 -385
rect 20040 -440 20090 -415
rect 20040 -475 20050 -440
rect 20080 -475 20090 -440
rect 20040 -500 20090 -475
rect 20040 -530 20050 -500
rect 20080 -530 20090 -500
rect 19955 -550 20005 -540
rect 19955 -580 19965 -550
rect 19995 -580 20005 -550
rect 19955 -590 20005 -580
rect 19870 -630 19880 -600
rect 19910 -630 19920 -600
rect 19870 -635 19920 -630
rect 20040 -600 20090 -530
rect 20210 -385 20260 -375
rect 20210 -415 20220 -385
rect 20250 -415 20260 -385
rect 20210 -440 20260 -415
rect 20210 -475 20220 -440
rect 20250 -475 20260 -440
rect 20210 -500 20260 -475
rect 20210 -530 20220 -500
rect 20250 -530 20260 -500
rect 20125 -550 20175 -540
rect 20125 -580 20135 -550
rect 20165 -580 20175 -550
rect 20125 -590 20175 -580
rect 20040 -630 20050 -600
rect 20080 -630 20090 -600
rect 20040 -635 20090 -630
rect 20210 -600 20260 -530
rect 20380 -385 20430 -375
rect 20380 -415 20390 -385
rect 20420 -415 20430 -385
rect 20380 -440 20430 -415
rect 20380 -475 20390 -440
rect 20420 -475 20430 -440
rect 20380 -500 20430 -475
rect 20380 -530 20390 -500
rect 20420 -530 20430 -500
rect 20295 -550 20345 -540
rect 20295 -580 20305 -550
rect 20335 -580 20345 -550
rect 20295 -590 20345 -580
rect 20210 -630 20220 -600
rect 20250 -630 20260 -600
rect 20210 -635 20260 -630
rect 20380 -600 20430 -530
rect 20550 -385 20600 -375
rect 20550 -415 20560 -385
rect 20590 -415 20600 -385
rect 20550 -440 20600 -415
rect 20550 -475 20560 -440
rect 20590 -475 20600 -440
rect 20550 -500 20600 -475
rect 20550 -530 20560 -500
rect 20590 -530 20600 -500
rect 20465 -550 20515 -540
rect 20465 -580 20475 -550
rect 20505 -580 20515 -550
rect 20465 -590 20515 -580
rect 20380 -630 20390 -600
rect 20420 -630 20430 -600
rect 20380 -635 20430 -630
rect 20550 -600 20600 -530
rect 20720 -385 20770 -375
rect 20720 -415 20730 -385
rect 20760 -415 20770 -385
rect 20720 -440 20770 -415
rect 20720 -475 20730 -440
rect 20760 -475 20770 -440
rect 20720 -500 20770 -475
rect 20720 -530 20730 -500
rect 20760 -530 20770 -500
rect 20635 -550 20685 -540
rect 20635 -580 20645 -550
rect 20675 -580 20685 -550
rect 20635 -590 20685 -580
rect 20550 -630 20560 -600
rect 20590 -630 20600 -600
rect 20550 -635 20600 -630
rect 20720 -600 20770 -530
rect 20890 -385 20940 -375
rect 20890 -415 20900 -385
rect 20930 -415 20940 -385
rect 20890 -440 20940 -415
rect 20890 -475 20900 -440
rect 20930 -475 20940 -440
rect 20890 -500 20940 -475
rect 20890 -530 20900 -500
rect 20930 -530 20940 -500
rect 20805 -550 20855 -540
rect 20805 -580 20815 -550
rect 20845 -580 20855 -550
rect 20805 -590 20855 -580
rect 20720 -630 20730 -600
rect 20760 -630 20770 -600
rect 20720 -635 20770 -630
rect 20890 -600 20940 -530
rect 21060 -385 21110 -375
rect 21060 -415 21070 -385
rect 21100 -415 21110 -385
rect 21060 -440 21110 -415
rect 21060 -475 21070 -440
rect 21100 -475 21110 -440
rect 21060 -500 21110 -475
rect 21060 -530 21070 -500
rect 21100 -530 21110 -500
rect 20975 -550 21025 -540
rect 20975 -580 20985 -550
rect 21015 -580 21025 -550
rect 20975 -590 21025 -580
rect 20890 -630 20900 -600
rect 20930 -630 20940 -600
rect 20890 -635 20940 -630
rect 21060 -600 21110 -530
rect 21230 -385 21280 -375
rect 21230 -415 21240 -385
rect 21270 -415 21280 -385
rect 21230 -440 21280 -415
rect 21230 -475 21240 -440
rect 21270 -475 21280 -440
rect 21230 -500 21280 -475
rect 21230 -530 21240 -500
rect 21270 -530 21280 -500
rect 21145 -550 21195 -540
rect 21145 -580 21155 -550
rect 21185 -580 21195 -550
rect 21145 -590 21195 -580
rect 21060 -630 21070 -600
rect 21100 -630 21110 -600
rect 21060 -635 21110 -630
rect 21230 -600 21280 -530
rect 21400 -385 21450 -375
rect 21400 -415 21410 -385
rect 21440 -415 21450 -385
rect 21400 -440 21450 -415
rect 21400 -475 21410 -440
rect 21440 -475 21450 -440
rect 21400 -500 21450 -475
rect 21400 -530 21410 -500
rect 21440 -530 21450 -500
rect 21315 -550 21365 -540
rect 21315 -580 21325 -550
rect 21355 -580 21365 -550
rect 21315 -590 21365 -580
rect 21230 -630 21240 -600
rect 21270 -630 21280 -600
rect 21230 -635 21280 -630
rect 21400 -600 21450 -530
rect 21570 -385 21620 -375
rect 21570 -415 21580 -385
rect 21610 -415 21620 -385
rect 21570 -440 21620 -415
rect 21570 -475 21580 -440
rect 21610 -475 21620 -440
rect 21570 -500 21620 -475
rect 21570 -530 21580 -500
rect 21610 -530 21620 -500
rect 21485 -550 21535 -540
rect 21485 -580 21495 -550
rect 21525 -580 21535 -550
rect 21485 -590 21535 -580
rect 21400 -630 21410 -600
rect 21440 -630 21450 -600
rect 21400 -635 21450 -630
rect 21570 -600 21620 -530
rect 21740 -385 21790 -375
rect 21740 -415 21750 -385
rect 21780 -415 21790 -385
rect 21740 -440 21790 -415
rect 21740 -475 21750 -440
rect 21780 -475 21790 -440
rect 21740 -500 21790 -475
rect 21740 -530 21750 -500
rect 21780 -530 21790 -500
rect 21655 -550 21705 -540
rect 21655 -580 21665 -550
rect 21695 -580 21705 -550
rect 21655 -590 21705 -580
rect 21570 -630 21580 -600
rect 21610 -630 21620 -600
rect 21570 -635 21620 -630
rect 21740 -600 21790 -530
rect 21910 -385 21960 -375
rect 21910 -415 21920 -385
rect 21950 -415 21960 -385
rect 21910 -440 21960 -415
rect 21910 -475 21920 -440
rect 21950 -475 21960 -440
rect 21910 -500 21960 -475
rect 21910 -530 21920 -500
rect 21950 -530 21960 -500
rect 21825 -550 21875 -540
rect 21825 -580 21835 -550
rect 21865 -580 21875 -550
rect 21825 -590 21875 -580
rect 21740 -630 21750 -600
rect 21780 -630 21790 -600
rect 21740 -635 21790 -630
rect 21910 -600 21960 -530
rect 22080 -385 22130 -375
rect 22080 -415 22090 -385
rect 22120 -415 22130 -385
rect 22080 -440 22130 -415
rect 22080 -475 22090 -440
rect 22120 -475 22130 -440
rect 22080 -500 22130 -475
rect 22080 -530 22090 -500
rect 22120 -530 22130 -500
rect 21995 -550 22045 -540
rect 21995 -580 22005 -550
rect 22035 -580 22045 -550
rect 21995 -590 22045 -580
rect 21910 -630 21920 -600
rect 21950 -630 21960 -600
rect 21910 -635 21960 -630
rect 22080 -600 22130 -530
rect 22250 -385 22300 -375
rect 22250 -415 22260 -385
rect 22290 -415 22300 -385
rect 22250 -440 22300 -415
rect 22250 -475 22260 -440
rect 22290 -475 22300 -440
rect 22250 -500 22300 -475
rect 22250 -530 22260 -500
rect 22290 -530 22300 -500
rect 22165 -550 22215 -540
rect 22165 -580 22175 -550
rect 22205 -580 22215 -550
rect 22165 -590 22215 -580
rect 22080 -630 22090 -600
rect 22120 -630 22130 -600
rect 22080 -635 22130 -630
rect 22250 -600 22300 -530
rect 22420 -385 22470 -375
rect 22420 -415 22430 -385
rect 22460 -415 22470 -385
rect 22420 -440 22470 -415
rect 22420 -475 22430 -440
rect 22460 -475 22470 -440
rect 22420 -500 22470 -475
rect 22420 -530 22430 -500
rect 22460 -530 22470 -500
rect 22335 -550 22385 -540
rect 22335 -580 22345 -550
rect 22375 -580 22385 -550
rect 22335 -590 22385 -580
rect 22250 -630 22260 -600
rect 22290 -630 22300 -600
rect 22250 -635 22300 -630
rect 22420 -600 22470 -530
rect 22590 -385 22640 -375
rect 22590 -415 22600 -385
rect 22630 -415 22640 -385
rect 22590 -440 22640 -415
rect 22590 -475 22600 -440
rect 22630 -475 22640 -440
rect 22590 -500 22640 -475
rect 22590 -530 22600 -500
rect 22630 -530 22640 -500
rect 22505 -550 22555 -540
rect 22505 -580 22515 -550
rect 22545 -580 22555 -550
rect 22505 -590 22555 -580
rect 22420 -630 22430 -600
rect 22460 -630 22470 -600
rect 22420 -635 22470 -630
rect 22590 -600 22640 -530
rect 22760 -385 22810 -375
rect 22760 -415 22770 -385
rect 22800 -415 22810 -385
rect 22760 -440 22810 -415
rect 22760 -475 22770 -440
rect 22800 -475 22810 -440
rect 22760 -500 22810 -475
rect 22760 -530 22770 -500
rect 22800 -530 22810 -500
rect 22675 -550 22725 -540
rect 22675 -580 22685 -550
rect 22715 -580 22725 -550
rect 22675 -590 22725 -580
rect 22590 -630 22600 -600
rect 22630 -630 22640 -600
rect 22590 -635 22640 -630
rect 22760 -600 22810 -530
rect 22930 -385 22980 -375
rect 22930 -415 22940 -385
rect 22970 -415 22980 -385
rect 22930 -440 22980 -415
rect 22930 -475 22940 -440
rect 22970 -475 22980 -440
rect 22930 -500 22980 -475
rect 22930 -530 22940 -500
rect 22970 -530 22980 -500
rect 22845 -550 22895 -540
rect 22845 -580 22855 -550
rect 22885 -580 22895 -550
rect 22845 -590 22895 -580
rect 22760 -630 22770 -600
rect 22800 -630 22810 -600
rect 22760 -635 22810 -630
rect 22930 -600 22980 -530
rect 23100 -385 23150 -375
rect 23100 -415 23110 -385
rect 23140 -415 23150 -385
rect 23100 -440 23150 -415
rect 23100 -475 23110 -440
rect 23140 -475 23150 -440
rect 23100 -500 23150 -475
rect 23100 -530 23110 -500
rect 23140 -530 23150 -500
rect 23015 -550 23065 -540
rect 23015 -580 23025 -550
rect 23055 -580 23065 -550
rect 23015 -590 23065 -580
rect 22930 -630 22940 -600
rect 22970 -630 22980 -600
rect 22930 -635 22980 -630
rect 23100 -600 23150 -530
rect 23270 -385 23320 -375
rect 23270 -415 23280 -385
rect 23310 -415 23320 -385
rect 23270 -440 23320 -415
rect 23270 -475 23280 -440
rect 23310 -475 23320 -440
rect 23270 -500 23320 -475
rect 23270 -530 23280 -500
rect 23310 -530 23320 -500
rect 23185 -550 23235 -540
rect 23185 -580 23195 -550
rect 23225 -580 23235 -550
rect 23185 -590 23235 -580
rect 23100 -630 23110 -600
rect 23140 -630 23150 -600
rect 23100 -635 23150 -630
rect 23270 -600 23320 -530
rect 23440 -385 23490 -375
rect 23440 -415 23450 -385
rect 23480 -415 23490 -385
rect 23440 -440 23490 -415
rect 23440 -475 23450 -440
rect 23480 -475 23490 -440
rect 23440 -500 23490 -475
rect 23440 -530 23450 -500
rect 23480 -530 23490 -500
rect 23355 -550 23405 -540
rect 23355 -580 23365 -550
rect 23395 -580 23405 -550
rect 23355 -590 23405 -580
rect 23270 -630 23280 -600
rect 23310 -630 23320 -600
rect 23270 -635 23320 -630
rect 23440 -600 23490 -530
rect 23610 -385 23660 -375
rect 23610 -415 23620 -385
rect 23650 -415 23660 -385
rect 23610 -440 23660 -415
rect 23610 -475 23620 -440
rect 23650 -475 23660 -440
rect 23610 -500 23660 -475
rect 23610 -530 23620 -500
rect 23650 -530 23660 -500
rect 23525 -550 23575 -540
rect 23525 -580 23535 -550
rect 23565 -580 23575 -550
rect 23525 -590 23575 -580
rect 23440 -630 23450 -600
rect 23480 -630 23490 -600
rect 23440 -635 23490 -630
rect 23610 -600 23660 -530
rect 23780 -385 23830 -375
rect 23780 -415 23790 -385
rect 23820 -415 23830 -385
rect 23780 -440 23830 -415
rect 23780 -475 23790 -440
rect 23820 -475 23830 -440
rect 23780 -500 23830 -475
rect 23780 -530 23790 -500
rect 23820 -530 23830 -500
rect 23695 -550 23745 -540
rect 23695 -580 23705 -550
rect 23735 -580 23745 -550
rect 23695 -590 23745 -580
rect 23610 -630 23620 -600
rect 23650 -630 23660 -600
rect 23610 -635 23660 -630
rect 23780 -600 23830 -530
rect 23950 -385 24000 -375
rect 23950 -415 23960 -385
rect 23990 -415 24000 -385
rect 23950 -440 24000 -415
rect 23950 -475 23960 -440
rect 23990 -475 24000 -440
rect 23950 -500 24000 -475
rect 23950 -530 23960 -500
rect 23990 -530 24000 -500
rect 23865 -550 23915 -540
rect 23865 -580 23875 -550
rect 23905 -580 23915 -550
rect 23865 -590 23915 -580
rect 23780 -630 23790 -600
rect 23820 -630 23830 -600
rect 23780 -635 23830 -630
rect 23950 -600 24000 -530
rect 24120 -385 24170 -375
rect 24120 -415 24130 -385
rect 24160 -415 24170 -385
rect 24120 -440 24170 -415
rect 24120 -475 24130 -440
rect 24160 -475 24170 -440
rect 24120 -500 24170 -475
rect 24120 -530 24130 -500
rect 24160 -530 24170 -500
rect 24035 -550 24085 -540
rect 24035 -580 24045 -550
rect 24075 -580 24085 -550
rect 24035 -590 24085 -580
rect 23950 -630 23960 -600
rect 23990 -630 24000 -600
rect 23950 -635 24000 -630
rect 24120 -600 24170 -530
rect 24290 -385 24340 -375
rect 24290 -415 24300 -385
rect 24330 -415 24340 -385
rect 24290 -440 24340 -415
rect 24290 -475 24300 -440
rect 24330 -475 24340 -440
rect 24290 -500 24340 -475
rect 24290 -530 24300 -500
rect 24330 -530 24340 -500
rect 24205 -550 24255 -540
rect 24205 -580 24215 -550
rect 24245 -580 24255 -550
rect 24205 -590 24255 -580
rect 24120 -630 24130 -600
rect 24160 -630 24170 -600
rect 24120 -635 24170 -630
rect 24290 -600 24340 -530
rect 24460 -385 24510 -375
rect 24460 -415 24470 -385
rect 24500 -415 24510 -385
rect 24460 -440 24510 -415
rect 24460 -475 24470 -440
rect 24500 -475 24510 -440
rect 24460 -500 24510 -475
rect 24460 -530 24470 -500
rect 24500 -530 24510 -500
rect 24375 -550 24425 -540
rect 24375 -580 24385 -550
rect 24415 -580 24425 -550
rect 24375 -590 24425 -580
rect 24290 -630 24300 -600
rect 24330 -630 24340 -600
rect 24290 -635 24340 -630
rect 24460 -600 24510 -530
rect 24630 -385 24680 -375
rect 24630 -415 24640 -385
rect 24670 -415 24680 -385
rect 24630 -440 24680 -415
rect 24630 -475 24640 -440
rect 24670 -475 24680 -440
rect 24630 -500 24680 -475
rect 24630 -530 24640 -500
rect 24670 -530 24680 -500
rect 24545 -550 24595 -540
rect 24545 -580 24555 -550
rect 24585 -580 24595 -550
rect 24545 -590 24595 -580
rect 24460 -630 24470 -600
rect 24500 -630 24510 -600
rect 24460 -635 24510 -630
rect 24630 -600 24680 -530
rect 24800 -385 24850 -375
rect 24800 -415 24810 -385
rect 24840 -415 24850 -385
rect 24800 -440 24850 -415
rect 24800 -475 24810 -440
rect 24840 -475 24850 -440
rect 24800 -500 24850 -475
rect 24800 -530 24810 -500
rect 24840 -530 24850 -500
rect 24715 -550 24765 -540
rect 24715 -580 24725 -550
rect 24755 -580 24765 -550
rect 24715 -590 24765 -580
rect 24630 -630 24640 -600
rect 24670 -630 24680 -600
rect 24630 -635 24680 -630
rect 24800 -600 24850 -530
rect 24970 -385 25020 -375
rect 24970 -415 24980 -385
rect 25010 -415 25020 -385
rect 24970 -440 25020 -415
rect 24970 -475 24980 -440
rect 25010 -475 25020 -440
rect 24970 -500 25020 -475
rect 24970 -530 24980 -500
rect 25010 -530 25020 -500
rect 24885 -550 24935 -540
rect 24885 -580 24895 -550
rect 24925 -580 24935 -550
rect 24885 -590 24935 -580
rect 24800 -630 24810 -600
rect 24840 -630 24850 -600
rect 24800 -635 24850 -630
rect 24970 -600 25020 -530
rect 25140 -385 25190 -375
rect 25140 -415 25150 -385
rect 25180 -415 25190 -385
rect 25140 -440 25190 -415
rect 25140 -475 25150 -440
rect 25180 -475 25190 -440
rect 25140 -500 25190 -475
rect 25140 -530 25150 -500
rect 25180 -530 25190 -500
rect 25055 -550 25105 -540
rect 25055 -580 25065 -550
rect 25095 -580 25105 -550
rect 25055 -590 25105 -580
rect 24970 -630 24980 -600
rect 25010 -630 25020 -600
rect 24970 -635 25020 -630
rect 25140 -600 25190 -530
rect 25310 -385 25360 -375
rect 25310 -415 25320 -385
rect 25350 -415 25360 -385
rect 25310 -440 25360 -415
rect 25310 -475 25320 -440
rect 25350 -475 25360 -440
rect 25310 -500 25360 -475
rect 25310 -530 25320 -500
rect 25350 -530 25360 -500
rect 25225 -550 25275 -540
rect 25225 -580 25235 -550
rect 25265 -580 25275 -550
rect 25225 -590 25275 -580
rect 25140 -630 25150 -600
rect 25180 -630 25190 -600
rect 25140 -635 25190 -630
rect 25310 -600 25360 -530
rect 25480 -385 25530 -375
rect 25480 -415 25490 -385
rect 25520 -415 25530 -385
rect 25480 -440 25530 -415
rect 25480 -475 25490 -440
rect 25520 -475 25530 -440
rect 25480 -500 25530 -475
rect 25480 -530 25490 -500
rect 25520 -530 25530 -500
rect 25395 -550 25445 -540
rect 25395 -580 25405 -550
rect 25435 -580 25445 -550
rect 25395 -590 25445 -580
rect 25310 -630 25320 -600
rect 25350 -630 25360 -600
rect 25310 -635 25360 -630
rect 25480 -600 25530 -530
rect 25650 -385 25700 -375
rect 25650 -415 25660 -385
rect 25690 -415 25700 -385
rect 25650 -440 25700 -415
rect 25650 -475 25660 -440
rect 25690 -475 25700 -440
rect 25650 -500 25700 -475
rect 25650 -530 25660 -500
rect 25690 -530 25700 -500
rect 25565 -550 25615 -540
rect 25565 -580 25575 -550
rect 25605 -580 25615 -550
rect 25565 -590 25615 -580
rect 25480 -630 25490 -600
rect 25520 -630 25530 -600
rect 25480 -635 25530 -630
rect 25650 -600 25700 -530
rect 25820 -385 25870 -375
rect 25820 -415 25830 -385
rect 25860 -415 25870 -385
rect 25820 -440 25870 -415
rect 25820 -475 25830 -440
rect 25860 -475 25870 -440
rect 25820 -500 25870 -475
rect 25820 -530 25830 -500
rect 25860 -530 25870 -500
rect 25735 -550 25785 -540
rect 25735 -580 25745 -550
rect 25775 -580 25785 -550
rect 25735 -590 25785 -580
rect 25650 -630 25660 -600
rect 25690 -630 25700 -600
rect 25650 -635 25700 -630
rect 25820 -600 25870 -530
rect 25990 -385 26040 -375
rect 25990 -415 26000 -385
rect 26030 -415 26040 -385
rect 25990 -440 26040 -415
rect 25990 -475 26000 -440
rect 26030 -475 26040 -440
rect 25990 -500 26040 -475
rect 25990 -530 26000 -500
rect 26030 -530 26040 -500
rect 25905 -550 25955 -540
rect 25905 -580 25915 -550
rect 25945 -580 25955 -550
rect 25905 -590 25955 -580
rect 25820 -630 25830 -600
rect 25860 -630 25870 -600
rect 25820 -635 25870 -630
rect 25990 -600 26040 -530
rect 26160 -385 26210 -375
rect 26160 -415 26170 -385
rect 26200 -415 26210 -385
rect 26160 -440 26210 -415
rect 26160 -475 26170 -440
rect 26200 -475 26210 -440
rect 26160 -500 26210 -475
rect 26160 -530 26170 -500
rect 26200 -530 26210 -500
rect 26075 -550 26125 -540
rect 26075 -580 26085 -550
rect 26115 -580 26125 -550
rect 26075 -590 26125 -580
rect 25990 -630 26000 -600
rect 26030 -630 26040 -600
rect 25990 -635 26040 -630
rect 26160 -600 26210 -530
rect 26330 -385 26380 -375
rect 26330 -415 26340 -385
rect 26370 -415 26380 -385
rect 26330 -440 26380 -415
rect 26330 -475 26340 -440
rect 26370 -475 26380 -440
rect 26330 -500 26380 -475
rect 26330 -530 26340 -500
rect 26370 -530 26380 -500
rect 26245 -550 26295 -540
rect 26245 -580 26255 -550
rect 26285 -580 26295 -550
rect 26245 -590 26295 -580
rect 26160 -630 26170 -600
rect 26200 -630 26210 -600
rect 26160 -635 26210 -630
rect 26330 -600 26380 -530
rect 26500 -385 26550 -375
rect 26500 -415 26510 -385
rect 26540 -415 26550 -385
rect 26500 -440 26550 -415
rect 26500 -475 26510 -440
rect 26540 -475 26550 -440
rect 26500 -500 26550 -475
rect 26500 -530 26510 -500
rect 26540 -530 26550 -500
rect 26415 -550 26465 -540
rect 26415 -580 26425 -550
rect 26455 -580 26465 -550
rect 26415 -590 26465 -580
rect 26330 -630 26340 -600
rect 26370 -630 26380 -600
rect 26330 -635 26380 -630
rect 26500 -600 26550 -530
rect 26670 -385 26720 -375
rect 26670 -415 26680 -385
rect 26710 -415 26720 -385
rect 26670 -440 26720 -415
rect 26670 -475 26680 -440
rect 26710 -475 26720 -440
rect 26670 -500 26720 -475
rect 26670 -530 26680 -500
rect 26710 -530 26720 -500
rect 26585 -550 26635 -540
rect 26585 -580 26595 -550
rect 26625 -580 26635 -550
rect 26585 -590 26635 -580
rect 26500 -630 26510 -600
rect 26540 -630 26550 -600
rect 26500 -635 26550 -630
rect 26670 -600 26720 -530
rect 26840 -385 26890 -375
rect 26840 -415 26850 -385
rect 26880 -415 26890 -385
rect 26840 -440 26890 -415
rect 26840 -475 26850 -440
rect 26880 -475 26890 -440
rect 26840 -500 26890 -475
rect 26840 -530 26850 -500
rect 26880 -530 26890 -500
rect 26755 -550 26805 -540
rect 26755 -580 26765 -550
rect 26795 -580 26805 -550
rect 26755 -590 26805 -580
rect 26670 -630 26680 -600
rect 26710 -630 26720 -600
rect 26670 -635 26720 -630
rect 26840 -600 26890 -530
rect 27010 -385 27060 -375
rect 27010 -415 27020 -385
rect 27050 -415 27060 -385
rect 27010 -440 27060 -415
rect 27010 -475 27020 -440
rect 27050 -475 27060 -440
rect 27010 -500 27060 -475
rect 27010 -530 27020 -500
rect 27050 -530 27060 -500
rect 26925 -550 26975 -540
rect 26925 -580 26935 -550
rect 26965 -580 26975 -550
rect 26925 -590 26975 -580
rect 26840 -630 26850 -600
rect 26880 -630 26890 -600
rect 26840 -635 26890 -630
rect 27010 -600 27060 -530
rect 27180 -385 27230 -375
rect 27180 -415 27190 -385
rect 27220 -415 27230 -385
rect 27180 -440 27230 -415
rect 27180 -475 27190 -440
rect 27220 -475 27230 -440
rect 27180 -500 27230 -475
rect 27180 -530 27190 -500
rect 27220 -530 27230 -500
rect 27095 -550 27145 -540
rect 27095 -580 27105 -550
rect 27135 -580 27145 -550
rect 27095 -590 27145 -580
rect 27010 -630 27020 -600
rect 27050 -630 27060 -600
rect 27010 -635 27060 -630
rect 27180 -600 27230 -530
rect 27350 -385 27400 -375
rect 27350 -415 27360 -385
rect 27390 -415 27400 -385
rect 27350 -440 27400 -415
rect 27350 -475 27360 -440
rect 27390 -475 27400 -440
rect 27350 -500 27400 -475
rect 27350 -530 27360 -500
rect 27390 -530 27400 -500
rect 27265 -550 27315 -540
rect 27265 -580 27275 -550
rect 27305 -580 27315 -550
rect 27265 -590 27315 -580
rect 27180 -630 27190 -600
rect 27220 -630 27230 -600
rect 27180 -635 27230 -630
rect 27350 -600 27400 -530
rect 27520 -385 27570 -375
rect 27520 -415 27530 -385
rect 27560 -415 27570 -385
rect 27520 -440 27570 -415
rect 27520 -475 27530 -440
rect 27560 -475 27570 -440
rect 27520 -500 27570 -475
rect 27520 -530 27530 -500
rect 27560 -530 27570 -500
rect 27435 -550 27485 -540
rect 27435 -580 27445 -550
rect 27475 -580 27485 -550
rect 27435 -590 27485 -580
rect 27350 -630 27360 -600
rect 27390 -630 27400 -600
rect 27350 -635 27400 -630
rect 27520 -600 27570 -530
rect 27690 -385 27740 -375
rect 27690 -415 27700 -385
rect 27730 -415 27740 -385
rect 27690 -440 27740 -415
rect 27690 -475 27700 -440
rect 27730 -475 27740 -440
rect 27690 -500 27740 -475
rect 27690 -530 27700 -500
rect 27730 -530 27740 -500
rect 27605 -550 27655 -540
rect 27605 -580 27615 -550
rect 27645 -580 27655 -550
rect 27605 -590 27655 -580
rect 27520 -630 27530 -600
rect 27560 -630 27570 -600
rect 27520 -635 27570 -630
rect 27690 -600 27740 -530
rect 27860 -385 27910 -375
rect 27860 -415 27870 -385
rect 27900 -415 27910 -385
rect 27860 -440 27910 -415
rect 27860 -475 27870 -440
rect 27900 -475 27910 -440
rect 27860 -500 27910 -475
rect 27860 -530 27870 -500
rect 27900 -530 27910 -500
rect 27775 -550 27825 -540
rect 27775 -580 27785 -550
rect 27815 -580 27825 -550
rect 27775 -590 27825 -580
rect 27690 -630 27700 -600
rect 27730 -630 27740 -600
rect 27690 -635 27740 -630
rect 27860 -600 27910 -530
rect 28030 -385 28080 -375
rect 28030 -415 28040 -385
rect 28070 -415 28080 -385
rect 28030 -440 28080 -415
rect 28030 -475 28040 -440
rect 28070 -475 28080 -440
rect 28030 -500 28080 -475
rect 28030 -530 28040 -500
rect 28070 -530 28080 -500
rect 27945 -550 27995 -540
rect 27945 -580 27955 -550
rect 27985 -580 27995 -550
rect 27945 -590 27995 -580
rect 27860 -630 27870 -600
rect 27900 -630 27910 -600
rect 27860 -635 27910 -630
rect 28030 -600 28080 -530
rect 28200 -385 28250 -375
rect 28200 -415 28210 -385
rect 28240 -415 28250 -385
rect 28200 -440 28250 -415
rect 28200 -475 28210 -440
rect 28240 -475 28250 -440
rect 28200 -500 28250 -475
rect 28200 -530 28210 -500
rect 28240 -530 28250 -500
rect 28115 -550 28165 -540
rect 28115 -580 28125 -550
rect 28155 -580 28165 -550
rect 28115 -590 28165 -580
rect 28030 -630 28040 -600
rect 28070 -630 28080 -600
rect 28030 -635 28080 -630
rect 28200 -600 28250 -530
rect 28370 -385 28420 -375
rect 28370 -415 28380 -385
rect 28410 -415 28420 -385
rect 28370 -440 28420 -415
rect 28370 -475 28380 -440
rect 28410 -475 28420 -440
rect 28370 -500 28420 -475
rect 28370 -530 28380 -500
rect 28410 -530 28420 -500
rect 28285 -550 28335 -540
rect 28285 -580 28295 -550
rect 28325 -580 28335 -550
rect 28285 -590 28335 -580
rect 28200 -630 28210 -600
rect 28240 -630 28250 -600
rect 28200 -635 28250 -630
rect 28370 -600 28420 -530
rect 28540 -385 28590 -375
rect 28540 -415 28550 -385
rect 28580 -415 28590 -385
rect 28540 -440 28590 -415
rect 28540 -475 28550 -440
rect 28580 -475 28590 -440
rect 28540 -500 28590 -475
rect 28540 -530 28550 -500
rect 28580 -530 28590 -500
rect 28455 -550 28505 -540
rect 28455 -580 28465 -550
rect 28495 -580 28505 -550
rect 28455 -590 28505 -580
rect 28370 -630 28380 -600
rect 28410 -630 28420 -600
rect 28370 -635 28420 -630
rect 28540 -600 28590 -530
rect 28710 -385 28760 -375
rect 28710 -415 28720 -385
rect 28750 -415 28760 -385
rect 28710 -440 28760 -415
rect 28710 -475 28720 -440
rect 28750 -475 28760 -440
rect 28710 -500 28760 -475
rect 28710 -530 28720 -500
rect 28750 -530 28760 -500
rect 28625 -550 28675 -540
rect 28625 -580 28635 -550
rect 28665 -580 28675 -550
rect 28625 -590 28675 -580
rect 28540 -630 28550 -600
rect 28580 -630 28590 -600
rect 28540 -635 28590 -630
rect 28710 -600 28760 -530
rect 28880 -385 28930 -375
rect 28880 -415 28890 -385
rect 28920 -415 28930 -385
rect 28880 -440 28930 -415
rect 28880 -475 28890 -440
rect 28920 -475 28930 -440
rect 28880 -500 28930 -475
rect 28880 -530 28890 -500
rect 28920 -530 28930 -500
rect 28795 -550 28845 -540
rect 28795 -580 28805 -550
rect 28835 -580 28845 -550
rect 28795 -590 28845 -580
rect 28710 -630 28720 -600
rect 28750 -630 28760 -600
rect 28710 -635 28760 -630
rect 28880 -600 28930 -530
rect 29050 -385 29100 -375
rect 29050 -415 29060 -385
rect 29090 -415 29100 -385
rect 29050 -440 29100 -415
rect 29050 -475 29060 -440
rect 29090 -475 29100 -440
rect 29050 -500 29100 -475
rect 29050 -530 29060 -500
rect 29090 -530 29100 -500
rect 28965 -550 29015 -540
rect 28965 -580 28975 -550
rect 29005 -580 29015 -550
rect 28965 -590 29015 -580
rect 28880 -630 28890 -600
rect 28920 -630 28930 -600
rect 28880 -635 28930 -630
rect 29050 -600 29100 -530
rect 29220 -385 29270 -375
rect 29220 -415 29230 -385
rect 29260 -415 29270 -385
rect 29220 -440 29270 -415
rect 29220 -475 29230 -440
rect 29260 -475 29270 -440
rect 29220 -500 29270 -475
rect 29220 -530 29230 -500
rect 29260 -530 29270 -500
rect 29135 -550 29185 -540
rect 29135 -580 29145 -550
rect 29175 -580 29185 -550
rect 29135 -590 29185 -580
rect 29050 -630 29060 -600
rect 29090 -630 29100 -600
rect 29050 -635 29100 -630
rect 29220 -600 29270 -530
rect 29390 -385 29440 -375
rect 29390 -415 29400 -385
rect 29430 -415 29440 -385
rect 29390 -440 29440 -415
rect 29390 -475 29400 -440
rect 29430 -475 29440 -440
rect 29390 -500 29440 -475
rect 29390 -530 29400 -500
rect 29430 -530 29440 -500
rect 29305 -550 29355 -540
rect 29305 -580 29315 -550
rect 29345 -580 29355 -550
rect 29305 -590 29355 -580
rect 29220 -630 29230 -600
rect 29260 -630 29270 -600
rect 29220 -635 29270 -630
rect 29390 -600 29440 -530
rect 29560 -385 29610 -375
rect 29560 -415 29570 -385
rect 29600 -415 29610 -385
rect 29560 -440 29610 -415
rect 29560 -475 29570 -440
rect 29600 -475 29610 -440
rect 29560 -500 29610 -475
rect 29560 -530 29570 -500
rect 29600 -530 29610 -500
rect 29475 -550 29525 -540
rect 29475 -580 29485 -550
rect 29515 -580 29525 -550
rect 29475 -590 29525 -580
rect 29390 -630 29400 -600
rect 29430 -630 29440 -600
rect 29390 -635 29440 -630
rect 29560 -600 29610 -530
rect 29730 -385 29780 -375
rect 29730 -415 29740 -385
rect 29770 -415 29780 -385
rect 29730 -440 29780 -415
rect 29730 -475 29740 -440
rect 29770 -475 29780 -440
rect 29730 -500 29780 -475
rect 29730 -530 29740 -500
rect 29770 -530 29780 -500
rect 29645 -550 29695 -540
rect 29645 -580 29655 -550
rect 29685 -580 29695 -550
rect 29645 -590 29695 -580
rect 29560 -630 29570 -600
rect 29600 -630 29610 -600
rect 29560 -635 29610 -630
rect 29730 -600 29780 -530
rect 29900 -385 29950 -375
rect 29900 -415 29910 -385
rect 29940 -415 29950 -385
rect 29900 -440 29950 -415
rect 29900 -475 29910 -440
rect 29940 -475 29950 -440
rect 29900 -500 29950 -475
rect 29900 -530 29910 -500
rect 29940 -530 29950 -500
rect 29815 -550 29865 -540
rect 29815 -580 29825 -550
rect 29855 -580 29865 -550
rect 29815 -590 29865 -580
rect 29730 -630 29740 -600
rect 29770 -630 29780 -600
rect 29730 -635 29780 -630
rect 29900 -600 29950 -530
rect 30070 -385 30120 -375
rect 30070 -415 30080 -385
rect 30110 -415 30120 -385
rect 30070 -440 30120 -415
rect 30070 -475 30080 -440
rect 30110 -475 30120 -440
rect 30070 -500 30120 -475
rect 30070 -530 30080 -500
rect 30110 -530 30120 -500
rect 29985 -550 30035 -540
rect 29985 -580 29995 -550
rect 30025 -580 30035 -550
rect 29985 -590 30035 -580
rect 29900 -630 29910 -600
rect 29940 -630 29950 -600
rect 29900 -635 29950 -630
rect 30070 -600 30120 -530
rect 30240 -385 30290 -375
rect 30240 -415 30250 -385
rect 30280 -415 30290 -385
rect 30240 -440 30290 -415
rect 30240 -475 30250 -440
rect 30280 -475 30290 -440
rect 30240 -500 30290 -475
rect 30240 -530 30250 -500
rect 30280 -530 30290 -500
rect 30155 -550 30205 -540
rect 30155 -580 30165 -550
rect 30195 -580 30205 -550
rect 30155 -590 30205 -580
rect 30070 -630 30080 -600
rect 30110 -630 30120 -600
rect 30070 -635 30120 -630
rect 30240 -600 30290 -530
rect 30410 -385 30460 -375
rect 30410 -415 30420 -385
rect 30450 -415 30460 -385
rect 30410 -440 30460 -415
rect 30410 -475 30420 -440
rect 30450 -475 30460 -440
rect 30410 -500 30460 -475
rect 30410 -530 30420 -500
rect 30450 -530 30460 -500
rect 30325 -550 30375 -540
rect 30325 -580 30335 -550
rect 30365 -580 30375 -550
rect 30325 -590 30375 -580
rect 30240 -630 30250 -600
rect 30280 -630 30290 -600
rect 30240 -635 30290 -630
rect 30410 -600 30460 -530
rect 30580 -385 30630 -375
rect 30580 -415 30590 -385
rect 30620 -415 30630 -385
rect 30580 -440 30630 -415
rect 30580 -475 30590 -440
rect 30620 -475 30630 -440
rect 30580 -500 30630 -475
rect 30580 -530 30590 -500
rect 30620 -530 30630 -500
rect 30495 -550 30545 -540
rect 30495 -580 30505 -550
rect 30535 -580 30545 -550
rect 30495 -590 30545 -580
rect 30410 -630 30420 -600
rect 30450 -630 30460 -600
rect 30410 -635 30460 -630
rect 30580 -600 30630 -530
rect 30750 -385 30800 -375
rect 30750 -415 30760 -385
rect 30790 -415 30800 -385
rect 30750 -440 30800 -415
rect 30750 -475 30760 -440
rect 30790 -475 30800 -440
rect 30750 -500 30800 -475
rect 30750 -530 30760 -500
rect 30790 -530 30800 -500
rect 30665 -550 30715 -540
rect 30665 -580 30675 -550
rect 30705 -580 30715 -550
rect 30665 -590 30715 -580
rect 30580 -630 30590 -600
rect 30620 -630 30630 -600
rect 30580 -635 30630 -630
rect 30750 -600 30800 -530
rect 30920 -385 30970 -375
rect 30920 -415 30930 -385
rect 30960 -415 30970 -385
rect 30920 -440 30970 -415
rect 30920 -475 30930 -440
rect 30960 -475 30970 -440
rect 30920 -500 30970 -475
rect 30920 -530 30930 -500
rect 30960 -530 30970 -500
rect 30835 -550 30885 -540
rect 30835 -580 30845 -550
rect 30875 -580 30885 -550
rect 30835 -590 30885 -580
rect 30750 -630 30760 -600
rect 30790 -630 30800 -600
rect 30750 -635 30800 -630
rect 30920 -600 30970 -530
rect 31090 -385 31140 -375
rect 31090 -415 31100 -385
rect 31130 -415 31140 -385
rect 31090 -440 31140 -415
rect 31090 -475 31100 -440
rect 31130 -475 31140 -440
rect 31090 -500 31140 -475
rect 31090 -530 31100 -500
rect 31130 -530 31140 -500
rect 31005 -550 31055 -540
rect 31005 -580 31015 -550
rect 31045 -580 31055 -550
rect 31005 -590 31055 -580
rect 30920 -630 30930 -600
rect 30960 -630 30970 -600
rect 30920 -635 30970 -630
rect 31090 -600 31140 -530
rect 31260 -385 31310 -375
rect 31260 -415 31270 -385
rect 31300 -415 31310 -385
rect 31260 -440 31310 -415
rect 31260 -475 31270 -440
rect 31300 -475 31310 -440
rect 31260 -500 31310 -475
rect 31260 -530 31270 -500
rect 31300 -530 31310 -500
rect 31175 -550 31225 -540
rect 31175 -580 31185 -550
rect 31215 -580 31225 -550
rect 31175 -590 31225 -580
rect 31090 -630 31100 -600
rect 31130 -630 31140 -600
rect 31090 -635 31140 -630
rect 31260 -600 31310 -530
rect 31430 -385 31480 -375
rect 31430 -415 31440 -385
rect 31470 -415 31480 -385
rect 31430 -440 31480 -415
rect 31430 -475 31440 -440
rect 31470 -475 31480 -440
rect 31430 -500 31480 -475
rect 31430 -530 31440 -500
rect 31470 -530 31480 -500
rect 31345 -550 31395 -540
rect 31345 -580 31355 -550
rect 31385 -580 31395 -550
rect 31345 -590 31395 -580
rect 31260 -630 31270 -600
rect 31300 -630 31310 -600
rect 31260 -635 31310 -630
rect 31430 -600 31480 -530
rect 31600 -385 31650 -375
rect 31600 -415 31610 -385
rect 31640 -415 31650 -385
rect 31600 -440 31650 -415
rect 31600 -475 31610 -440
rect 31640 -475 31650 -440
rect 31600 -500 31650 -475
rect 31600 -530 31610 -500
rect 31640 -530 31650 -500
rect 31515 -550 31565 -540
rect 31515 -580 31525 -550
rect 31555 -580 31565 -550
rect 31515 -590 31565 -580
rect 31430 -630 31440 -600
rect 31470 -630 31480 -600
rect 31430 -635 31480 -630
rect 31600 -600 31650 -530
rect 31770 -385 31820 -375
rect 31770 -415 31780 -385
rect 31810 -415 31820 -385
rect 31770 -440 31820 -415
rect 31770 -475 31780 -440
rect 31810 -475 31820 -440
rect 31770 -500 31820 -475
rect 31770 -530 31780 -500
rect 31810 -530 31820 -500
rect 31685 -550 31735 -540
rect 31685 -580 31695 -550
rect 31725 -580 31735 -550
rect 31685 -590 31735 -580
rect 31600 -630 31610 -600
rect 31640 -630 31650 -600
rect 31600 -635 31650 -630
rect 31770 -600 31820 -530
rect 31940 -385 31990 -375
rect 31940 -415 31950 -385
rect 31980 -415 31990 -385
rect 31940 -440 31990 -415
rect 31940 -475 31950 -440
rect 31980 -475 31990 -440
rect 31940 -500 31990 -475
rect 31940 -530 31950 -500
rect 31980 -530 31990 -500
rect 31855 -550 31905 -540
rect 31855 -580 31865 -550
rect 31895 -580 31905 -550
rect 31855 -590 31905 -580
rect 31770 -630 31780 -600
rect 31810 -630 31820 -600
rect 31770 -635 31820 -630
rect 31940 -600 31990 -530
rect 32110 -385 32160 -375
rect 32110 -415 32120 -385
rect 32150 -415 32160 -385
rect 32110 -440 32160 -415
rect 32110 -475 32120 -440
rect 32150 -475 32160 -440
rect 32110 -500 32160 -475
rect 32110 -530 32120 -500
rect 32150 -530 32160 -500
rect 32025 -550 32075 -540
rect 32025 -580 32035 -550
rect 32065 -580 32075 -550
rect 32025 -590 32075 -580
rect 31940 -630 31950 -600
rect 31980 -630 31990 -600
rect 31940 -635 31990 -630
rect 32110 -600 32160 -530
rect 32280 -385 32330 -375
rect 32280 -415 32290 -385
rect 32320 -415 32330 -385
rect 32280 -440 32330 -415
rect 32280 -475 32290 -440
rect 32320 -475 32330 -440
rect 32280 -500 32330 -475
rect 32280 -530 32290 -500
rect 32320 -530 32330 -500
rect 32195 -550 32245 -540
rect 32195 -580 32205 -550
rect 32235 -580 32245 -550
rect 32195 -590 32245 -580
rect 32110 -630 32120 -600
rect 32150 -630 32160 -600
rect 32110 -635 32160 -630
rect 32280 -600 32330 -530
rect 32450 -385 32500 -375
rect 32450 -415 32460 -385
rect 32490 -415 32500 -385
rect 32450 -440 32500 -415
rect 32450 -475 32460 -440
rect 32490 -475 32500 -440
rect 32450 -500 32500 -475
rect 32450 -530 32460 -500
rect 32490 -530 32500 -500
rect 32365 -550 32415 -540
rect 32365 -580 32375 -550
rect 32405 -580 32415 -550
rect 32365 -590 32415 -580
rect 32280 -630 32290 -600
rect 32320 -630 32330 -600
rect 32280 -635 32330 -630
rect 32450 -600 32500 -530
rect 32620 -385 32670 -375
rect 32620 -415 32630 -385
rect 32660 -415 32670 -385
rect 32620 -440 32670 -415
rect 32620 -475 32630 -440
rect 32660 -475 32670 -440
rect 32620 -500 32670 -475
rect 32620 -530 32630 -500
rect 32660 -530 32670 -500
rect 32535 -550 32585 -540
rect 32535 -580 32545 -550
rect 32575 -580 32585 -550
rect 32535 -590 32585 -580
rect 32450 -630 32460 -600
rect 32490 -630 32500 -600
rect 32450 -635 32500 -630
rect 32620 -600 32670 -530
rect 32790 -385 32840 -375
rect 32790 -415 32800 -385
rect 32830 -415 32840 -385
rect 32790 -440 32840 -415
rect 32790 -475 32800 -440
rect 32830 -475 32840 -440
rect 32790 -500 32840 -475
rect 32790 -530 32800 -500
rect 32830 -530 32840 -500
rect 32705 -550 32755 -540
rect 32705 -580 32715 -550
rect 32745 -580 32755 -550
rect 32705 -590 32755 -580
rect 32620 -630 32630 -600
rect 32660 -630 32670 -600
rect 32620 -635 32670 -630
rect 32790 -600 32840 -530
rect 32960 -385 33010 -375
rect 32960 -415 32970 -385
rect 33000 -415 33010 -385
rect 32960 -440 33010 -415
rect 32960 -475 32970 -440
rect 33000 -475 33010 -440
rect 32960 -500 33010 -475
rect 32960 -530 32970 -500
rect 33000 -530 33010 -500
rect 32875 -550 32925 -540
rect 32875 -580 32885 -550
rect 32915 -580 32925 -550
rect 32875 -590 32925 -580
rect 32790 -630 32800 -600
rect 32830 -630 32840 -600
rect 32790 -635 32840 -630
rect 32960 -600 33010 -530
rect 33130 -385 33180 -375
rect 33130 -415 33140 -385
rect 33170 -415 33180 -385
rect 33130 -440 33180 -415
rect 33130 -475 33140 -440
rect 33170 -475 33180 -440
rect 33130 -500 33180 -475
rect 33130 -530 33140 -500
rect 33170 -530 33180 -500
rect 33045 -550 33095 -540
rect 33045 -580 33055 -550
rect 33085 -580 33095 -550
rect 33045 -590 33095 -580
rect 32960 -630 32970 -600
rect 33000 -630 33010 -600
rect 32960 -635 33010 -630
rect 33130 -600 33180 -530
rect 33300 -385 33350 -375
rect 33300 -415 33310 -385
rect 33340 -415 33350 -385
rect 33300 -440 33350 -415
rect 33300 -475 33310 -440
rect 33340 -475 33350 -440
rect 33300 -500 33350 -475
rect 33300 -530 33310 -500
rect 33340 -530 33350 -500
rect 33215 -550 33265 -540
rect 33215 -580 33225 -550
rect 33255 -580 33265 -550
rect 33215 -590 33265 -580
rect 33130 -630 33140 -600
rect 33170 -630 33180 -600
rect 33130 -635 33180 -630
rect 33300 -600 33350 -530
rect 33470 -385 33520 -375
rect 33470 -415 33480 -385
rect 33510 -415 33520 -385
rect 33470 -440 33520 -415
rect 33470 -475 33480 -440
rect 33510 -475 33520 -440
rect 33470 -500 33520 -475
rect 33470 -530 33480 -500
rect 33510 -530 33520 -500
rect 33385 -550 33435 -540
rect 33385 -580 33395 -550
rect 33425 -580 33435 -550
rect 33385 -590 33435 -580
rect 33300 -630 33310 -600
rect 33340 -630 33350 -600
rect 33300 -635 33350 -630
rect 33470 -600 33520 -530
rect 33640 -385 33690 -375
rect 33640 -415 33650 -385
rect 33680 -415 33690 -385
rect 33640 -440 33690 -415
rect 33640 -475 33650 -440
rect 33680 -475 33690 -440
rect 33640 -500 33690 -475
rect 33640 -530 33650 -500
rect 33680 -530 33690 -500
rect 33555 -550 33605 -540
rect 33555 -580 33565 -550
rect 33595 -580 33605 -550
rect 33555 -590 33605 -580
rect 33470 -630 33480 -600
rect 33510 -630 33520 -600
rect 33470 -635 33520 -630
rect 33640 -600 33690 -530
rect 33810 -385 33860 -375
rect 33810 -415 33820 -385
rect 33850 -415 33860 -385
rect 33810 -440 33860 -415
rect 33810 -475 33820 -440
rect 33850 -475 33860 -440
rect 33810 -500 33860 -475
rect 33810 -530 33820 -500
rect 33850 -530 33860 -500
rect 33725 -550 33775 -540
rect 33725 -580 33735 -550
rect 33765 -580 33775 -550
rect 33725 -590 33775 -580
rect 33640 -630 33650 -600
rect 33680 -630 33690 -600
rect 33640 -635 33690 -630
rect 33810 -600 33860 -530
rect 33980 -385 34030 -375
rect 33980 -415 33990 -385
rect 34020 -415 34030 -385
rect 33980 -440 34030 -415
rect 33980 -475 33990 -440
rect 34020 -475 34030 -440
rect 33980 -500 34030 -475
rect 33980 -530 33990 -500
rect 34020 -530 34030 -500
rect 33895 -550 33945 -540
rect 33895 -580 33905 -550
rect 33935 -580 33945 -550
rect 33895 -590 33945 -580
rect 33810 -630 33820 -600
rect 33850 -630 33860 -600
rect 33810 -635 33860 -630
rect 33980 -600 34030 -530
rect 34150 -385 34200 -375
rect 34150 -415 34160 -385
rect 34190 -415 34200 -385
rect 34150 -440 34200 -415
rect 34150 -475 34160 -440
rect 34190 -475 34200 -440
rect 34150 -500 34200 -475
rect 34150 -530 34160 -500
rect 34190 -530 34200 -500
rect 34065 -550 34115 -540
rect 34065 -580 34075 -550
rect 34105 -580 34115 -550
rect 34065 -590 34115 -580
rect 33980 -630 33990 -600
rect 34020 -630 34030 -600
rect 33980 -635 34030 -630
rect 34150 -600 34200 -530
rect 34320 -385 34370 -375
rect 34320 -415 34330 -385
rect 34360 -415 34370 -385
rect 34320 -440 34370 -415
rect 34320 -475 34330 -440
rect 34360 -475 34370 -440
rect 34320 -500 34370 -475
rect 34320 -530 34330 -500
rect 34360 -530 34370 -500
rect 34235 -550 34285 -540
rect 34235 -580 34245 -550
rect 34275 -580 34285 -550
rect 34235 -590 34285 -580
rect 34150 -630 34160 -600
rect 34190 -630 34200 -600
rect 34150 -635 34200 -630
rect 34320 -600 34370 -530
rect 34490 -385 34540 -375
rect 34490 -415 34500 -385
rect 34530 -415 34540 -385
rect 34490 -440 34540 -415
rect 34490 -475 34500 -440
rect 34530 -475 34540 -440
rect 34490 -500 34540 -475
rect 34490 -530 34500 -500
rect 34530 -530 34540 -500
rect 34405 -550 34455 -540
rect 34405 -580 34415 -550
rect 34445 -580 34455 -550
rect 34405 -590 34455 -580
rect 34320 -630 34330 -600
rect 34360 -630 34370 -600
rect 34320 -635 34370 -630
rect 34490 -600 34540 -530
rect 34660 -385 34710 -375
rect 34660 -415 34670 -385
rect 34700 -415 34710 -385
rect 34660 -440 34710 -415
rect 34660 -475 34670 -440
rect 34700 -475 34710 -440
rect 34660 -500 34710 -475
rect 34660 -530 34670 -500
rect 34700 -530 34710 -500
rect 34575 -550 34625 -540
rect 34575 -580 34585 -550
rect 34615 -580 34625 -550
rect 34575 -590 34625 -580
rect 34490 -630 34500 -600
rect 34530 -630 34540 -600
rect 34490 -635 34540 -630
rect 34660 -600 34710 -530
rect 34830 -385 34880 -375
rect 34830 -415 34840 -385
rect 34870 -415 34880 -385
rect 34830 -440 34880 -415
rect 34830 -475 34840 -440
rect 34870 -475 34880 -440
rect 34830 -500 34880 -475
rect 34830 -530 34840 -500
rect 34870 -530 34880 -500
rect 34745 -550 34795 -540
rect 34745 -580 34755 -550
rect 34785 -580 34795 -550
rect 34745 -590 34795 -580
rect 34660 -630 34670 -600
rect 34700 -630 34710 -600
rect 34660 -635 34710 -630
rect 34830 -600 34880 -530
rect 35000 -385 35050 -375
rect 35000 -415 35010 -385
rect 35040 -415 35050 -385
rect 35000 -440 35050 -415
rect 35000 -475 35010 -440
rect 35040 -475 35050 -440
rect 35000 -500 35050 -475
rect 35000 -530 35010 -500
rect 35040 -530 35050 -500
rect 34915 -550 34965 -540
rect 34915 -580 34925 -550
rect 34955 -580 34965 -550
rect 34915 -590 34965 -580
rect 34830 -630 34840 -600
rect 34870 -630 34880 -600
rect 34830 -635 34880 -630
rect 35000 -600 35050 -530
rect 35170 -385 35220 -375
rect 35170 -415 35180 -385
rect 35210 -415 35220 -385
rect 35170 -440 35220 -415
rect 35170 -475 35180 -440
rect 35210 -475 35220 -440
rect 35170 -500 35220 -475
rect 35170 -530 35180 -500
rect 35210 -530 35220 -500
rect 35085 -550 35135 -540
rect 35085 -580 35095 -550
rect 35125 -580 35135 -550
rect 35085 -590 35135 -580
rect 35000 -630 35010 -600
rect 35040 -630 35050 -600
rect 35000 -635 35050 -630
rect 35170 -600 35220 -530
rect 35340 -385 35390 -375
rect 35340 -415 35350 -385
rect 35380 -415 35390 -385
rect 35340 -440 35390 -415
rect 35340 -475 35350 -440
rect 35380 -475 35390 -440
rect 35340 -500 35390 -475
rect 35340 -530 35350 -500
rect 35380 -530 35390 -500
rect 35255 -550 35305 -540
rect 35255 -580 35265 -550
rect 35295 -580 35305 -550
rect 35255 -590 35305 -580
rect 35170 -630 35180 -600
rect 35210 -630 35220 -600
rect 35170 -635 35220 -630
rect 35340 -600 35390 -530
rect 35510 -385 35560 -375
rect 35510 -415 35520 -385
rect 35550 -415 35560 -385
rect 35510 -440 35560 -415
rect 35510 -475 35520 -440
rect 35550 -475 35560 -440
rect 35510 -500 35560 -475
rect 35510 -530 35520 -500
rect 35550 -530 35560 -500
rect 35425 -550 35475 -540
rect 35425 -580 35435 -550
rect 35465 -580 35475 -550
rect 35425 -590 35475 -580
rect 35340 -630 35350 -600
rect 35380 -630 35390 -600
rect 35340 -635 35390 -630
rect 35510 -600 35560 -530
rect 35680 -385 35730 -375
rect 35680 -415 35690 -385
rect 35720 -415 35730 -385
rect 35680 -440 35730 -415
rect 35680 -475 35690 -440
rect 35720 -475 35730 -440
rect 35680 -500 35730 -475
rect 35680 -530 35690 -500
rect 35720 -530 35730 -500
rect 35595 -550 35645 -540
rect 35595 -580 35605 -550
rect 35635 -580 35645 -550
rect 35595 -590 35645 -580
rect 35510 -630 35520 -600
rect 35550 -630 35560 -600
rect 35510 -635 35560 -630
rect 35680 -600 35730 -530
rect 35850 -385 35900 -375
rect 35850 -415 35860 -385
rect 35890 -415 35900 -385
rect 35850 -440 35900 -415
rect 35850 -475 35860 -440
rect 35890 -475 35900 -440
rect 35850 -500 35900 -475
rect 35850 -530 35860 -500
rect 35890 -530 35900 -500
rect 35765 -550 35815 -540
rect 35765 -580 35775 -550
rect 35805 -580 35815 -550
rect 35765 -590 35815 -580
rect 35680 -630 35690 -600
rect 35720 -630 35730 -600
rect 35680 -635 35730 -630
rect 35850 -600 35900 -530
rect 36020 -385 36070 -375
rect 36020 -415 36030 -385
rect 36060 -415 36070 -385
rect 36020 -440 36070 -415
rect 36020 -475 36030 -440
rect 36060 -475 36070 -440
rect 36020 -500 36070 -475
rect 36020 -530 36030 -500
rect 36060 -530 36070 -500
rect 35935 -550 35985 -540
rect 35935 -580 35945 -550
rect 35975 -580 35985 -550
rect 35935 -590 35985 -580
rect 35850 -630 35860 -600
rect 35890 -630 35900 -600
rect 35850 -635 35900 -630
rect 36020 -600 36070 -530
rect 36190 -385 36240 -375
rect 36190 -415 36200 -385
rect 36230 -415 36240 -385
rect 36190 -440 36240 -415
rect 36190 -475 36200 -440
rect 36230 -475 36240 -440
rect 36190 -500 36240 -475
rect 36190 -530 36200 -500
rect 36230 -530 36240 -500
rect 36105 -550 36155 -540
rect 36105 -580 36115 -550
rect 36145 -580 36155 -550
rect 36105 -590 36155 -580
rect 36020 -630 36030 -600
rect 36060 -630 36070 -600
rect 36020 -635 36070 -630
rect 36190 -600 36240 -530
rect 36360 -385 36410 -375
rect 36360 -415 36370 -385
rect 36400 -415 36410 -385
rect 36360 -440 36410 -415
rect 36360 -475 36370 -440
rect 36400 -475 36410 -440
rect 36360 -500 36410 -475
rect 36360 -530 36370 -500
rect 36400 -530 36410 -500
rect 36275 -550 36325 -540
rect 36275 -580 36285 -550
rect 36315 -580 36325 -550
rect 36275 -590 36325 -580
rect 36190 -630 36200 -600
rect 36230 -630 36240 -600
rect 36190 -635 36240 -630
rect 36360 -600 36410 -530
rect 36530 -385 36580 -375
rect 36530 -415 36540 -385
rect 36570 -415 36580 -385
rect 36530 -440 36580 -415
rect 36530 -475 36540 -440
rect 36570 -475 36580 -440
rect 36530 -500 36580 -475
rect 36530 -530 36540 -500
rect 36570 -530 36580 -500
rect 36445 -550 36495 -540
rect 36445 -580 36455 -550
rect 36485 -580 36495 -550
rect 36445 -590 36495 -580
rect 36360 -630 36370 -600
rect 36400 -630 36410 -600
rect 36360 -635 36410 -630
rect 36530 -600 36580 -530
rect 36700 -385 36750 -375
rect 36700 -415 36710 -385
rect 36740 -415 36750 -385
rect 36700 -440 36750 -415
rect 36700 -475 36710 -440
rect 36740 -475 36750 -440
rect 36700 -500 36750 -475
rect 36700 -530 36710 -500
rect 36740 -530 36750 -500
rect 36615 -550 36665 -540
rect 36615 -580 36625 -550
rect 36655 -580 36665 -550
rect 36615 -590 36665 -580
rect 36530 -630 36540 -600
rect 36570 -630 36580 -600
rect 36530 -635 36580 -630
rect 36700 -600 36750 -530
rect 36870 -385 36920 -375
rect 36870 -415 36880 -385
rect 36910 -415 36920 -385
rect 36870 -440 36920 -415
rect 36870 -475 36880 -440
rect 36910 -475 36920 -440
rect 36870 -500 36920 -475
rect 36870 -530 36880 -500
rect 36910 -530 36920 -500
rect 36785 -550 36835 -540
rect 36785 -580 36795 -550
rect 36825 -580 36835 -550
rect 36785 -590 36835 -580
rect 36700 -630 36710 -600
rect 36740 -630 36750 -600
rect 36700 -635 36750 -630
rect 36870 -600 36920 -530
rect 37040 -385 37090 -375
rect 37040 -415 37050 -385
rect 37080 -415 37090 -385
rect 37040 -440 37090 -415
rect 37040 -475 37050 -440
rect 37080 -475 37090 -440
rect 37040 -500 37090 -475
rect 37040 -530 37050 -500
rect 37080 -530 37090 -500
rect 36955 -550 37005 -540
rect 36955 -580 36965 -550
rect 36995 -580 37005 -550
rect 36955 -590 37005 -580
rect 36870 -630 36880 -600
rect 36910 -630 36920 -600
rect 36870 -635 36920 -630
rect 37040 -600 37090 -530
rect 37210 -385 37260 -375
rect 37210 -415 37220 -385
rect 37250 -415 37260 -385
rect 37210 -440 37260 -415
rect 37210 -475 37220 -440
rect 37250 -475 37260 -440
rect 37210 -500 37260 -475
rect 37210 -530 37220 -500
rect 37250 -530 37260 -500
rect 37125 -550 37175 -540
rect 37125 -580 37135 -550
rect 37165 -580 37175 -550
rect 37125 -590 37175 -580
rect 37040 -630 37050 -600
rect 37080 -630 37090 -600
rect 37040 -635 37090 -630
rect 37210 -600 37260 -530
rect 37380 -385 37430 -375
rect 37380 -415 37390 -385
rect 37420 -415 37430 -385
rect 37380 -440 37430 -415
rect 37380 -475 37390 -440
rect 37420 -475 37430 -440
rect 37380 -500 37430 -475
rect 37380 -530 37390 -500
rect 37420 -530 37430 -500
rect 37295 -550 37345 -540
rect 37295 -580 37305 -550
rect 37335 -580 37345 -550
rect 37295 -590 37345 -580
rect 37210 -630 37220 -600
rect 37250 -630 37260 -600
rect 37210 -635 37260 -630
rect 37380 -600 37430 -530
rect 37550 -385 37600 -375
rect 37550 -415 37560 -385
rect 37590 -415 37600 -385
rect 37550 -440 37600 -415
rect 37550 -475 37560 -440
rect 37590 -475 37600 -440
rect 37550 -500 37600 -475
rect 37550 -530 37560 -500
rect 37590 -530 37600 -500
rect 37465 -550 37515 -540
rect 37465 -580 37475 -550
rect 37505 -580 37515 -550
rect 37465 -590 37515 -580
rect 37380 -630 37390 -600
rect 37420 -630 37430 -600
rect 37380 -635 37430 -630
rect 37550 -600 37600 -530
rect 37720 -385 37770 -375
rect 37720 -415 37730 -385
rect 37760 -415 37770 -385
rect 37720 -440 37770 -415
rect 37720 -475 37730 -440
rect 37760 -475 37770 -440
rect 37720 -500 37770 -475
rect 37720 -530 37730 -500
rect 37760 -530 37770 -500
rect 37635 -550 37685 -540
rect 37635 -580 37645 -550
rect 37675 -580 37685 -550
rect 37635 -590 37685 -580
rect 37550 -630 37560 -600
rect 37590 -630 37600 -600
rect 37550 -635 37600 -630
rect 37720 -600 37770 -530
rect 37890 -385 37940 -375
rect 37890 -415 37900 -385
rect 37930 -415 37940 -385
rect 37890 -440 37940 -415
rect 37890 -475 37900 -440
rect 37930 -475 37940 -440
rect 37890 -500 37940 -475
rect 37890 -530 37900 -500
rect 37930 -530 37940 -500
rect 37805 -550 37855 -540
rect 37805 -580 37815 -550
rect 37845 -580 37855 -550
rect 37805 -590 37855 -580
rect 37720 -630 37730 -600
rect 37760 -630 37770 -600
rect 37720 -635 37770 -630
rect 37890 -600 37940 -530
rect 38060 -385 38110 -375
rect 38060 -415 38070 -385
rect 38100 -415 38110 -385
rect 38060 -440 38110 -415
rect 38060 -475 38070 -440
rect 38100 -475 38110 -440
rect 38060 -500 38110 -475
rect 38060 -530 38070 -500
rect 38100 -530 38110 -500
rect 37975 -550 38025 -540
rect 37975 -580 37985 -550
rect 38015 -580 38025 -550
rect 37975 -590 38025 -580
rect 37890 -630 37900 -600
rect 37930 -630 37940 -600
rect 37890 -635 37940 -630
rect 38060 -600 38110 -530
rect 38230 -385 38280 -375
rect 38230 -415 38240 -385
rect 38270 -415 38280 -385
rect 38230 -440 38280 -415
rect 38230 -475 38240 -440
rect 38270 -475 38280 -440
rect 38230 -500 38280 -475
rect 38230 -530 38240 -500
rect 38270 -530 38280 -500
rect 38145 -550 38195 -540
rect 38145 -580 38155 -550
rect 38185 -580 38195 -550
rect 38145 -590 38195 -580
rect 38060 -630 38070 -600
rect 38100 -630 38110 -600
rect 38060 -635 38110 -630
rect 38230 -600 38280 -530
rect 38400 -385 38450 -375
rect 38400 -415 38410 -385
rect 38440 -415 38450 -385
rect 38400 -440 38450 -415
rect 38400 -475 38410 -440
rect 38440 -475 38450 -440
rect 38400 -500 38450 -475
rect 38400 -530 38410 -500
rect 38440 -530 38450 -500
rect 38315 -550 38365 -540
rect 38315 -580 38325 -550
rect 38355 -580 38365 -550
rect 38315 -590 38365 -580
rect 38230 -630 38240 -600
rect 38270 -630 38280 -600
rect 38230 -635 38280 -630
rect 38400 -600 38450 -530
rect 38570 -385 38620 -375
rect 38570 -415 38580 -385
rect 38610 -415 38620 -385
rect 38570 -440 38620 -415
rect 38570 -475 38580 -440
rect 38610 -475 38620 -440
rect 38570 -500 38620 -475
rect 38570 -530 38580 -500
rect 38610 -530 38620 -500
rect 38485 -550 38535 -540
rect 38485 -580 38495 -550
rect 38525 -580 38535 -550
rect 38485 -590 38535 -580
rect 38400 -630 38410 -600
rect 38440 -630 38450 -600
rect 38400 -635 38450 -630
rect 38570 -600 38620 -530
rect 38740 -385 38790 -375
rect 38740 -415 38750 -385
rect 38780 -415 38790 -385
rect 38740 -440 38790 -415
rect 38740 -475 38750 -440
rect 38780 -475 38790 -440
rect 38740 -500 38790 -475
rect 38740 -530 38750 -500
rect 38780 -530 38790 -500
rect 38655 -550 38705 -540
rect 38655 -580 38665 -550
rect 38695 -580 38705 -550
rect 38655 -590 38705 -580
rect 38570 -630 38580 -600
rect 38610 -630 38620 -600
rect 38570 -635 38620 -630
rect 38740 -600 38790 -530
rect 38910 -385 38960 -375
rect 38910 -415 38920 -385
rect 38950 -415 38960 -385
rect 38910 -440 38960 -415
rect 38910 -475 38920 -440
rect 38950 -475 38960 -440
rect 38910 -500 38960 -475
rect 38910 -530 38920 -500
rect 38950 -530 38960 -500
rect 38825 -550 38875 -540
rect 38825 -580 38835 -550
rect 38865 -580 38875 -550
rect 38825 -590 38875 -580
rect 38740 -630 38750 -600
rect 38780 -630 38790 -600
rect 38740 -635 38790 -630
rect 38910 -600 38960 -530
rect 39080 -385 39130 -375
rect 39080 -415 39090 -385
rect 39120 -415 39130 -385
rect 39080 -440 39130 -415
rect 39080 -475 39090 -440
rect 39120 -475 39130 -440
rect 39080 -500 39130 -475
rect 39080 -530 39090 -500
rect 39120 -530 39130 -500
rect 38995 -550 39045 -540
rect 38995 -580 39005 -550
rect 39035 -580 39045 -550
rect 38995 -590 39045 -580
rect 38910 -630 38920 -600
rect 38950 -630 38960 -600
rect 38910 -635 38960 -630
rect 39080 -600 39130 -530
rect 39250 -385 39300 -375
rect 39250 -415 39260 -385
rect 39290 -415 39300 -385
rect 39250 -440 39300 -415
rect 39250 -475 39260 -440
rect 39290 -475 39300 -440
rect 39250 -500 39300 -475
rect 39250 -530 39260 -500
rect 39290 -530 39300 -500
rect 39165 -550 39215 -540
rect 39165 -580 39175 -550
rect 39205 -580 39215 -550
rect 39165 -590 39215 -580
rect 39080 -630 39090 -600
rect 39120 -630 39130 -600
rect 39080 -635 39130 -630
rect 39250 -600 39300 -530
rect 39420 -385 39470 -375
rect 39420 -415 39430 -385
rect 39460 -415 39470 -385
rect 39420 -440 39470 -415
rect 39420 -475 39430 -440
rect 39460 -475 39470 -440
rect 39420 -500 39470 -475
rect 39420 -530 39430 -500
rect 39460 -530 39470 -500
rect 39335 -550 39385 -540
rect 39335 -580 39345 -550
rect 39375 -580 39385 -550
rect 39335 -590 39385 -580
rect 39250 -630 39260 -600
rect 39290 -630 39300 -600
rect 39250 -635 39300 -630
rect 39420 -600 39470 -530
rect 39590 -385 39640 -375
rect 39590 -415 39600 -385
rect 39630 -415 39640 -385
rect 39590 -440 39640 -415
rect 39590 -475 39600 -440
rect 39630 -475 39640 -440
rect 39590 -500 39640 -475
rect 39590 -530 39600 -500
rect 39630 -530 39640 -500
rect 39505 -550 39555 -540
rect 39505 -580 39515 -550
rect 39545 -580 39555 -550
rect 39505 -590 39555 -580
rect 39420 -630 39430 -600
rect 39460 -630 39470 -600
rect 39420 -635 39470 -630
rect 39590 -600 39640 -530
rect 39760 -385 39810 -375
rect 39760 -415 39770 -385
rect 39800 -415 39810 -385
rect 39760 -440 39810 -415
rect 39760 -475 39770 -440
rect 39800 -475 39810 -440
rect 39760 -500 39810 -475
rect 39760 -530 39770 -500
rect 39800 -530 39810 -500
rect 39675 -550 39725 -540
rect 39675 -580 39685 -550
rect 39715 -580 39725 -550
rect 39675 -590 39725 -580
rect 39590 -630 39600 -600
rect 39630 -630 39640 -600
rect 39590 -635 39640 -630
rect 39760 -600 39810 -530
rect 39930 -385 39980 -375
rect 39930 -415 39940 -385
rect 39970 -415 39980 -385
rect 39930 -440 39980 -415
rect 39930 -475 39940 -440
rect 39970 -475 39980 -440
rect 39930 -500 39980 -475
rect 39930 -530 39940 -500
rect 39970 -530 39980 -500
rect 39845 -550 39895 -540
rect 39845 -580 39855 -550
rect 39885 -580 39895 -550
rect 39845 -590 39895 -580
rect 39760 -630 39770 -600
rect 39800 -630 39810 -600
rect 39760 -635 39810 -630
rect 39930 -600 39980 -530
rect 40100 -385 40150 -375
rect 40100 -415 40110 -385
rect 40140 -415 40150 -385
rect 40100 -440 40150 -415
rect 40100 -475 40110 -440
rect 40140 -475 40150 -440
rect 40100 -500 40150 -475
rect 40100 -530 40110 -500
rect 40140 -530 40150 -500
rect 40015 -550 40065 -540
rect 40015 -580 40025 -550
rect 40055 -580 40065 -550
rect 40015 -590 40065 -580
rect 39930 -630 39940 -600
rect 39970 -630 39980 -600
rect 39930 -635 39980 -630
rect 40100 -600 40150 -530
rect 40270 -385 40320 -375
rect 40270 -415 40280 -385
rect 40310 -415 40320 -385
rect 40270 -440 40320 -415
rect 40270 -475 40280 -440
rect 40310 -475 40320 -440
rect 40270 -500 40320 -475
rect 40270 -530 40280 -500
rect 40310 -530 40320 -500
rect 40185 -550 40235 -540
rect 40185 -580 40195 -550
rect 40225 -580 40235 -550
rect 40185 -590 40235 -580
rect 40100 -630 40110 -600
rect 40140 -630 40150 -600
rect 40100 -635 40150 -630
rect 40270 -600 40320 -530
rect 40440 -385 40490 -375
rect 40440 -415 40450 -385
rect 40480 -415 40490 -385
rect 40440 -440 40490 -415
rect 40440 -475 40450 -440
rect 40480 -475 40490 -440
rect 40440 -500 40490 -475
rect 40440 -530 40450 -500
rect 40480 -530 40490 -500
rect 40355 -550 40405 -540
rect 40355 -580 40365 -550
rect 40395 -580 40405 -550
rect 40355 -590 40405 -580
rect 40270 -630 40280 -600
rect 40310 -630 40320 -600
rect 40270 -635 40320 -630
rect 40440 -600 40490 -530
rect 40610 -385 40660 -375
rect 40610 -415 40620 -385
rect 40650 -415 40660 -385
rect 40610 -440 40660 -415
rect 40610 -475 40620 -440
rect 40650 -475 40660 -440
rect 40610 -500 40660 -475
rect 40610 -530 40620 -500
rect 40650 -530 40660 -500
rect 40525 -550 40575 -540
rect 40525 -580 40535 -550
rect 40565 -580 40575 -550
rect 40525 -590 40575 -580
rect 40440 -630 40450 -600
rect 40480 -630 40490 -600
rect 40440 -635 40490 -630
rect 40610 -600 40660 -530
rect 40780 -385 40830 -375
rect 40780 -415 40790 -385
rect 40820 -415 40830 -385
rect 40780 -440 40830 -415
rect 40780 -475 40790 -440
rect 40820 -475 40830 -440
rect 40780 -500 40830 -475
rect 40780 -530 40790 -500
rect 40820 -530 40830 -500
rect 40695 -550 40745 -540
rect 40695 -580 40705 -550
rect 40735 -580 40745 -550
rect 40695 -590 40745 -580
rect 40610 -630 40620 -600
rect 40650 -630 40660 -600
rect 40610 -635 40660 -630
rect 40780 -600 40830 -530
rect 40950 -385 41000 -375
rect 40950 -415 40960 -385
rect 40990 -415 41000 -385
rect 40950 -440 41000 -415
rect 40950 -475 40960 -440
rect 40990 -475 41000 -440
rect 40950 -500 41000 -475
rect 40950 -530 40960 -500
rect 40990 -530 41000 -500
rect 40865 -550 40915 -540
rect 40865 -580 40875 -550
rect 40905 -580 40915 -550
rect 40865 -590 40915 -580
rect 40780 -630 40790 -600
rect 40820 -630 40830 -600
rect 40780 -635 40830 -630
rect 40950 -600 41000 -530
rect 41120 -385 41170 -375
rect 41120 -415 41130 -385
rect 41160 -415 41170 -385
rect 41120 -440 41170 -415
rect 41120 -475 41130 -440
rect 41160 -475 41170 -440
rect 41120 -500 41170 -475
rect 41120 -530 41130 -500
rect 41160 -530 41170 -500
rect 41035 -550 41085 -540
rect 41035 -580 41045 -550
rect 41075 -580 41085 -550
rect 41035 -590 41085 -580
rect 40950 -630 40960 -600
rect 40990 -630 41000 -600
rect 40950 -635 41000 -630
rect 41120 -600 41170 -530
rect 41290 -385 41340 -375
rect 41290 -415 41300 -385
rect 41330 -415 41340 -385
rect 41290 -440 41340 -415
rect 41290 -475 41300 -440
rect 41330 -475 41340 -440
rect 41290 -500 41340 -475
rect 41290 -530 41300 -500
rect 41330 -530 41340 -500
rect 41205 -550 41255 -540
rect 41205 -580 41215 -550
rect 41245 -580 41255 -550
rect 41205 -590 41255 -580
rect 41120 -630 41130 -600
rect 41160 -630 41170 -600
rect 41120 -635 41170 -630
rect 41290 -600 41340 -530
rect 41460 -385 41510 -375
rect 41460 -415 41470 -385
rect 41500 -415 41510 -385
rect 41460 -440 41510 -415
rect 41460 -475 41470 -440
rect 41500 -475 41510 -440
rect 41460 -500 41510 -475
rect 41460 -530 41470 -500
rect 41500 -530 41510 -500
rect 41375 -550 41425 -540
rect 41375 -580 41385 -550
rect 41415 -580 41425 -550
rect 41375 -590 41425 -580
rect 41290 -630 41300 -600
rect 41330 -630 41340 -600
rect 41290 -635 41340 -630
rect 41460 -600 41510 -530
rect 41630 -385 41680 -375
rect 41630 -415 41640 -385
rect 41670 -415 41680 -385
rect 41630 -440 41680 -415
rect 41630 -475 41640 -440
rect 41670 -475 41680 -440
rect 41630 -500 41680 -475
rect 41630 -530 41640 -500
rect 41670 -530 41680 -500
rect 41545 -550 41595 -540
rect 41545 -580 41555 -550
rect 41585 -580 41595 -550
rect 41545 -590 41595 -580
rect 41460 -630 41470 -600
rect 41500 -630 41510 -600
rect 41460 -635 41510 -630
rect 41630 -600 41680 -530
rect 41800 -385 41850 -375
rect 41800 -415 41810 -385
rect 41840 -415 41850 -385
rect 41800 -440 41850 -415
rect 41800 -475 41810 -440
rect 41840 -475 41850 -440
rect 41800 -500 41850 -475
rect 41800 -530 41810 -500
rect 41840 -530 41850 -500
rect 41715 -550 41765 -540
rect 41715 -580 41725 -550
rect 41755 -580 41765 -550
rect 41715 -590 41765 -580
rect 41630 -630 41640 -600
rect 41670 -630 41680 -600
rect 41630 -635 41680 -630
rect 41800 -600 41850 -530
rect 41970 -385 42020 -375
rect 41970 -415 41980 -385
rect 42010 -415 42020 -385
rect 41970 -440 42020 -415
rect 41970 -475 41980 -440
rect 42010 -475 42020 -440
rect 41970 -500 42020 -475
rect 41970 -530 41980 -500
rect 42010 -530 42020 -500
rect 41885 -550 41935 -540
rect 41885 -580 41895 -550
rect 41925 -580 41935 -550
rect 41885 -590 41935 -580
rect 41800 -630 41810 -600
rect 41840 -630 41850 -600
rect 41800 -635 41850 -630
rect 41970 -600 42020 -530
rect 42140 -385 42190 -375
rect 42140 -415 42150 -385
rect 42180 -415 42190 -385
rect 42140 -440 42190 -415
rect 42140 -475 42150 -440
rect 42180 -475 42190 -440
rect 42140 -500 42190 -475
rect 42140 -530 42150 -500
rect 42180 -530 42190 -500
rect 42055 -550 42105 -540
rect 42055 -580 42065 -550
rect 42095 -580 42105 -550
rect 42055 -590 42105 -580
rect 41970 -630 41980 -600
rect 42010 -630 42020 -600
rect 41970 -635 42020 -630
rect 42140 -600 42190 -530
rect 42310 -385 42360 -375
rect 42310 -415 42320 -385
rect 42350 -415 42360 -385
rect 42310 -440 42360 -415
rect 42310 -475 42320 -440
rect 42350 -475 42360 -440
rect 42310 -500 42360 -475
rect 42310 -530 42320 -500
rect 42350 -530 42360 -500
rect 42225 -550 42275 -540
rect 42225 -580 42235 -550
rect 42265 -580 42275 -550
rect 42225 -590 42275 -580
rect 42140 -630 42150 -600
rect 42180 -630 42190 -600
rect 42140 -635 42190 -630
rect 42310 -600 42360 -530
rect 42480 -385 42530 -375
rect 42480 -415 42490 -385
rect 42520 -415 42530 -385
rect 42480 -440 42530 -415
rect 42480 -475 42490 -440
rect 42520 -475 42530 -440
rect 42480 -500 42530 -475
rect 42480 -530 42490 -500
rect 42520 -530 42530 -500
rect 42395 -550 42445 -540
rect 42395 -580 42405 -550
rect 42435 -580 42445 -550
rect 42395 -590 42445 -580
rect 42310 -630 42320 -600
rect 42350 -630 42360 -600
rect 42310 -635 42360 -630
rect 42480 -600 42530 -530
rect 42650 -385 42700 -375
rect 42650 -415 42660 -385
rect 42690 -415 42700 -385
rect 42650 -440 42700 -415
rect 42650 -475 42660 -440
rect 42690 -475 42700 -440
rect 42650 -500 42700 -475
rect 42650 -530 42660 -500
rect 42690 -530 42700 -500
rect 42565 -550 42615 -540
rect 42565 -580 42575 -550
rect 42605 -580 42615 -550
rect 42565 -590 42615 -580
rect 42480 -630 42490 -600
rect 42520 -630 42530 -600
rect 42480 -635 42530 -630
rect 42650 -600 42700 -530
rect 42820 -385 42870 -375
rect 42820 -415 42830 -385
rect 42860 -415 42870 -385
rect 42820 -440 42870 -415
rect 42820 -475 42830 -440
rect 42860 -475 42870 -440
rect 42820 -500 42870 -475
rect 42820 -530 42830 -500
rect 42860 -530 42870 -500
rect 42735 -550 42785 -540
rect 42735 -580 42745 -550
rect 42775 -580 42785 -550
rect 42735 -590 42785 -580
rect 42650 -630 42660 -600
rect 42690 -630 42700 -600
rect 42650 -635 42700 -630
rect 42820 -600 42870 -530
rect 42990 -385 43040 -375
rect 42990 -415 43000 -385
rect 43030 -415 43040 -385
rect 42990 -440 43040 -415
rect 42990 -475 43000 -440
rect 43030 -475 43040 -440
rect 42990 -500 43040 -475
rect 42990 -530 43000 -500
rect 43030 -530 43040 -500
rect 42905 -550 42955 -540
rect 42905 -580 42915 -550
rect 42945 -580 42955 -550
rect 42905 -590 42955 -580
rect 42820 -630 42830 -600
rect 42860 -630 42870 -600
rect 42820 -635 42870 -630
rect 42990 -600 43040 -530
rect 43160 -385 43210 -375
rect 43160 -415 43170 -385
rect 43200 -415 43210 -385
rect 43160 -440 43210 -415
rect 43160 -475 43170 -440
rect 43200 -475 43210 -440
rect 43160 -500 43210 -475
rect 43160 -530 43170 -500
rect 43200 -530 43210 -500
rect 43075 -550 43125 -540
rect 43075 -580 43085 -550
rect 43115 -580 43125 -550
rect 43075 -590 43125 -580
rect 42990 -630 43000 -600
rect 43030 -630 43040 -600
rect 42990 -635 43040 -630
rect 43160 -600 43210 -530
rect 43330 -385 43380 -375
rect 43330 -415 43340 -385
rect 43370 -415 43380 -385
rect 43330 -440 43380 -415
rect 43330 -475 43340 -440
rect 43370 -475 43380 -440
rect 43330 -500 43380 -475
rect 43330 -530 43340 -500
rect 43370 -530 43380 -500
rect 43245 -550 43295 -540
rect 43245 -580 43255 -550
rect 43285 -580 43295 -550
rect 43245 -590 43295 -580
rect 43160 -630 43170 -600
rect 43200 -630 43210 -600
rect 43160 -635 43210 -630
rect 43330 -600 43380 -530
rect 43500 -385 43550 -375
rect 43500 -415 43510 -385
rect 43540 -415 43550 -385
rect 43500 -440 43550 -415
rect 43500 -475 43510 -440
rect 43540 -475 43550 -440
rect 43500 -500 43550 -475
rect 43500 -530 43510 -500
rect 43540 -530 43550 -500
rect 43415 -550 43465 -540
rect 43415 -580 43425 -550
rect 43455 -580 43465 -550
rect 43415 -590 43465 -580
rect 43330 -630 43340 -600
rect 43370 -630 43380 -600
rect 43330 -635 43380 -630
rect 43500 -600 43550 -530
rect 43585 -550 43635 -540
rect 43585 -580 43595 -550
rect 43625 -580 43635 -550
rect 43585 -590 43635 -580
rect 43500 -630 43510 -600
rect 43540 -630 43550 -600
rect 43500 -635 43550 -630
rect 65 -650 115 -640
rect 65 -680 75 -650
rect 105 -680 115 -650
rect 65 -690 115 -680
rect 235 -650 285 -640
rect 235 -680 245 -650
rect 275 -680 285 -650
rect 235 -690 285 -680
rect 405 -650 455 -640
rect 405 -680 415 -650
rect 445 -680 455 -650
rect 405 -690 455 -680
rect 575 -650 625 -640
rect 575 -680 585 -650
rect 615 -680 625 -650
rect 575 -690 625 -680
rect 745 -650 795 -640
rect 745 -680 755 -650
rect 785 -680 795 -650
rect 745 -690 795 -680
rect 915 -650 965 -640
rect 915 -680 925 -650
rect 955 -680 965 -650
rect 915 -690 965 -680
rect 1085 -650 1135 -640
rect 1085 -680 1095 -650
rect 1125 -680 1135 -650
rect 1085 -690 1135 -680
rect 1255 -650 1305 -640
rect 1255 -680 1265 -650
rect 1295 -680 1305 -650
rect 1255 -690 1305 -680
rect 1425 -650 1475 -640
rect 1425 -680 1435 -650
rect 1465 -680 1475 -650
rect 1425 -690 1475 -680
rect 1595 -650 1645 -640
rect 1595 -680 1605 -650
rect 1635 -680 1645 -650
rect 1595 -690 1645 -680
rect 1765 -650 1815 -640
rect 1765 -680 1775 -650
rect 1805 -680 1815 -650
rect 1765 -690 1815 -680
rect 1935 -650 1985 -640
rect 1935 -680 1945 -650
rect 1975 -680 1985 -650
rect 1935 -690 1985 -680
rect 2105 -650 2155 -640
rect 2105 -680 2115 -650
rect 2145 -680 2155 -650
rect 2105 -690 2155 -680
rect 2275 -650 2325 -640
rect 2275 -680 2285 -650
rect 2315 -680 2325 -650
rect 2275 -690 2325 -680
rect 2445 -650 2495 -640
rect 2445 -680 2455 -650
rect 2485 -680 2495 -650
rect 2445 -690 2495 -680
rect 2615 -650 2665 -640
rect 2615 -680 2625 -650
rect 2655 -680 2665 -650
rect 2615 -690 2665 -680
rect 2785 -650 2835 -640
rect 2785 -680 2795 -650
rect 2825 -680 2835 -650
rect 2785 -690 2835 -680
rect 2955 -650 3005 -640
rect 2955 -680 2965 -650
rect 2995 -680 3005 -650
rect 2955 -690 3005 -680
rect 3125 -650 3175 -640
rect 3125 -680 3135 -650
rect 3165 -680 3175 -650
rect 3125 -690 3175 -680
rect 3295 -650 3345 -640
rect 3295 -680 3305 -650
rect 3335 -680 3345 -650
rect 3295 -690 3345 -680
rect 3465 -650 3515 -640
rect 3465 -680 3475 -650
rect 3505 -680 3515 -650
rect 3465 -690 3515 -680
rect 3635 -650 3685 -640
rect 3635 -680 3645 -650
rect 3675 -680 3685 -650
rect 3635 -690 3685 -680
rect 3805 -650 3855 -640
rect 3805 -680 3815 -650
rect 3845 -680 3855 -650
rect 3805 -690 3855 -680
rect 3975 -650 4025 -640
rect 3975 -680 3985 -650
rect 4015 -680 4025 -650
rect 3975 -690 4025 -680
rect 4145 -650 4195 -640
rect 4145 -680 4155 -650
rect 4185 -680 4195 -650
rect 4145 -690 4195 -680
rect 4315 -650 4365 -640
rect 4315 -680 4325 -650
rect 4355 -680 4365 -650
rect 4315 -690 4365 -680
rect 4485 -650 4535 -640
rect 4485 -680 4495 -650
rect 4525 -680 4535 -650
rect 4485 -690 4535 -680
rect 4655 -650 4705 -640
rect 4655 -680 4665 -650
rect 4695 -680 4705 -650
rect 4655 -690 4705 -680
rect 4825 -650 4875 -640
rect 4825 -680 4835 -650
rect 4865 -680 4875 -650
rect 4825 -690 4875 -680
rect 4995 -650 5045 -640
rect 4995 -680 5005 -650
rect 5035 -680 5045 -650
rect 4995 -690 5045 -680
rect 5165 -650 5215 -640
rect 5165 -680 5175 -650
rect 5205 -680 5215 -650
rect 5165 -690 5215 -680
rect 5335 -650 5385 -640
rect 5335 -680 5345 -650
rect 5375 -680 5385 -650
rect 5335 -690 5385 -680
rect 5505 -650 5555 -640
rect 5505 -680 5515 -650
rect 5545 -680 5555 -650
rect 5505 -690 5555 -680
rect 5675 -650 5725 -640
rect 5675 -680 5685 -650
rect 5715 -680 5725 -650
rect 5675 -690 5725 -680
rect 5845 -650 5895 -640
rect 5845 -680 5855 -650
rect 5885 -680 5895 -650
rect 5845 -690 5895 -680
rect 6015 -650 6065 -640
rect 6015 -680 6025 -650
rect 6055 -680 6065 -650
rect 6015 -690 6065 -680
rect 6185 -650 6235 -640
rect 6185 -680 6195 -650
rect 6225 -680 6235 -650
rect 6185 -690 6235 -680
rect 6355 -650 6405 -640
rect 6355 -680 6365 -650
rect 6395 -680 6405 -650
rect 6355 -690 6405 -680
rect 6525 -650 6575 -640
rect 6525 -680 6535 -650
rect 6565 -680 6575 -650
rect 6525 -690 6575 -680
rect 6695 -650 6745 -640
rect 6695 -680 6705 -650
rect 6735 -680 6745 -650
rect 6695 -690 6745 -680
rect 6865 -650 6915 -640
rect 6865 -680 6875 -650
rect 6905 -680 6915 -650
rect 6865 -690 6915 -680
rect 7035 -650 7085 -640
rect 7035 -680 7045 -650
rect 7075 -680 7085 -650
rect 7035 -690 7085 -680
rect 7205 -650 7255 -640
rect 7205 -680 7215 -650
rect 7245 -680 7255 -650
rect 7205 -690 7255 -680
rect 7375 -650 7425 -640
rect 7375 -680 7385 -650
rect 7415 -680 7425 -650
rect 7375 -690 7425 -680
rect 7545 -650 7595 -640
rect 7545 -680 7555 -650
rect 7585 -680 7595 -650
rect 7545 -690 7595 -680
rect 7715 -650 7765 -640
rect 7715 -680 7725 -650
rect 7755 -680 7765 -650
rect 7715 -690 7765 -680
rect 7885 -650 7935 -640
rect 7885 -680 7895 -650
rect 7925 -680 7935 -650
rect 7885 -690 7935 -680
rect 8055 -650 8105 -640
rect 8055 -680 8065 -650
rect 8095 -680 8105 -650
rect 8055 -690 8105 -680
rect 8225 -650 8275 -640
rect 8225 -680 8235 -650
rect 8265 -680 8275 -650
rect 8225 -690 8275 -680
rect 8395 -650 8445 -640
rect 8395 -680 8405 -650
rect 8435 -680 8445 -650
rect 8395 -690 8445 -680
rect 8565 -650 8615 -640
rect 8565 -680 8575 -650
rect 8605 -680 8615 -650
rect 8565 -690 8615 -680
rect 8735 -650 8785 -640
rect 8735 -680 8745 -650
rect 8775 -680 8785 -650
rect 8735 -690 8785 -680
rect 8905 -650 8955 -640
rect 8905 -680 8915 -650
rect 8945 -680 8955 -650
rect 8905 -690 8955 -680
rect 9075 -650 9125 -640
rect 9075 -680 9085 -650
rect 9115 -680 9125 -650
rect 9075 -690 9125 -680
rect 9245 -650 9295 -640
rect 9245 -680 9255 -650
rect 9285 -680 9295 -650
rect 9245 -690 9295 -680
rect 9415 -650 9465 -640
rect 9415 -680 9425 -650
rect 9455 -680 9465 -650
rect 9415 -690 9465 -680
rect 9585 -650 9635 -640
rect 9585 -680 9595 -650
rect 9625 -680 9635 -650
rect 9585 -690 9635 -680
rect 9755 -650 9805 -640
rect 9755 -680 9765 -650
rect 9795 -680 9805 -650
rect 9755 -690 9805 -680
rect 9925 -650 9975 -640
rect 9925 -680 9935 -650
rect 9965 -680 9975 -650
rect 9925 -690 9975 -680
rect 10095 -650 10145 -640
rect 10095 -680 10105 -650
rect 10135 -680 10145 -650
rect 10095 -690 10145 -680
rect 10265 -650 10315 -640
rect 10265 -680 10275 -650
rect 10305 -680 10315 -650
rect 10265 -690 10315 -680
rect 10435 -650 10485 -640
rect 10435 -680 10445 -650
rect 10475 -680 10485 -650
rect 10435 -690 10485 -680
rect 10605 -650 10655 -640
rect 10605 -680 10615 -650
rect 10645 -680 10655 -650
rect 10605 -690 10655 -680
rect 10775 -650 10825 -640
rect 10775 -680 10785 -650
rect 10815 -680 10825 -650
rect 10775 -690 10825 -680
rect 10945 -650 10995 -640
rect 10945 -680 10955 -650
rect 10985 -680 10995 -650
rect 10945 -690 10995 -680
rect 11115 -650 11165 -640
rect 11115 -680 11125 -650
rect 11155 -680 11165 -650
rect 11115 -690 11165 -680
rect 11285 -650 11335 -640
rect 11285 -680 11295 -650
rect 11325 -680 11335 -650
rect 11285 -690 11335 -680
rect 11455 -650 11505 -640
rect 11455 -680 11465 -650
rect 11495 -680 11505 -650
rect 11455 -690 11505 -680
rect 11625 -650 11675 -640
rect 11625 -680 11635 -650
rect 11665 -680 11675 -650
rect 11625 -690 11675 -680
rect 11795 -650 11845 -640
rect 11795 -680 11805 -650
rect 11835 -680 11845 -650
rect 11795 -690 11845 -680
rect 11965 -650 12015 -640
rect 11965 -680 11975 -650
rect 12005 -680 12015 -650
rect 11965 -690 12015 -680
rect 12135 -650 12185 -640
rect 12135 -680 12145 -650
rect 12175 -680 12185 -650
rect 12135 -690 12185 -680
rect 12305 -650 12355 -640
rect 12305 -680 12315 -650
rect 12345 -680 12355 -650
rect 12305 -690 12355 -680
rect 12475 -650 12525 -640
rect 12475 -680 12485 -650
rect 12515 -680 12525 -650
rect 12475 -690 12525 -680
rect 12645 -650 12695 -640
rect 12645 -680 12655 -650
rect 12685 -680 12695 -650
rect 12645 -690 12695 -680
rect 12815 -650 12865 -640
rect 12815 -680 12825 -650
rect 12855 -680 12865 -650
rect 12815 -690 12865 -680
rect 12985 -650 13035 -640
rect 12985 -680 12995 -650
rect 13025 -680 13035 -650
rect 12985 -690 13035 -680
rect 13155 -650 13205 -640
rect 13155 -680 13165 -650
rect 13195 -680 13205 -650
rect 13155 -690 13205 -680
rect 13325 -650 13375 -640
rect 13325 -680 13335 -650
rect 13365 -680 13375 -650
rect 13325 -690 13375 -680
rect 13495 -650 13545 -640
rect 13495 -680 13505 -650
rect 13535 -680 13545 -650
rect 13495 -690 13545 -680
rect 13665 -650 13715 -640
rect 13665 -680 13675 -650
rect 13705 -680 13715 -650
rect 13665 -690 13715 -680
rect 13835 -650 13885 -640
rect 13835 -680 13845 -650
rect 13875 -680 13885 -650
rect 13835 -690 13885 -680
rect 14005 -650 14055 -640
rect 14005 -680 14015 -650
rect 14045 -680 14055 -650
rect 14005 -690 14055 -680
rect 14175 -650 14225 -640
rect 14175 -680 14185 -650
rect 14215 -680 14225 -650
rect 14175 -690 14225 -680
rect 14345 -650 14395 -640
rect 14345 -680 14355 -650
rect 14385 -680 14395 -650
rect 14345 -690 14395 -680
rect 14515 -650 14565 -640
rect 14515 -680 14525 -650
rect 14555 -680 14565 -650
rect 14515 -690 14565 -680
rect 14685 -650 14735 -640
rect 14685 -680 14695 -650
rect 14725 -680 14735 -650
rect 14685 -690 14735 -680
rect 14855 -650 14905 -640
rect 14855 -680 14865 -650
rect 14895 -680 14905 -650
rect 14855 -690 14905 -680
rect 15025 -650 15075 -640
rect 15025 -680 15035 -650
rect 15065 -680 15075 -650
rect 15025 -690 15075 -680
rect 15195 -650 15245 -640
rect 15195 -680 15205 -650
rect 15235 -680 15245 -650
rect 15195 -690 15245 -680
rect 15365 -650 15415 -640
rect 15365 -680 15375 -650
rect 15405 -680 15415 -650
rect 15365 -690 15415 -680
rect 15535 -650 15585 -640
rect 15535 -680 15545 -650
rect 15575 -680 15585 -650
rect 15535 -690 15585 -680
rect 15705 -650 15755 -640
rect 15705 -680 15715 -650
rect 15745 -680 15755 -650
rect 15705 -690 15755 -680
rect 15875 -650 15925 -640
rect 15875 -680 15885 -650
rect 15915 -680 15925 -650
rect 15875 -690 15925 -680
rect 16045 -650 16095 -640
rect 16045 -680 16055 -650
rect 16085 -680 16095 -650
rect 16045 -690 16095 -680
rect 16215 -650 16265 -640
rect 16215 -680 16225 -650
rect 16255 -680 16265 -650
rect 16215 -690 16265 -680
rect 16385 -650 16435 -640
rect 16385 -680 16395 -650
rect 16425 -680 16435 -650
rect 16385 -690 16435 -680
rect 16555 -650 16605 -640
rect 16555 -680 16565 -650
rect 16595 -680 16605 -650
rect 16555 -690 16605 -680
rect 16725 -650 16775 -640
rect 16725 -680 16735 -650
rect 16765 -680 16775 -650
rect 16725 -690 16775 -680
rect 16895 -650 16945 -640
rect 16895 -680 16905 -650
rect 16935 -680 16945 -650
rect 16895 -690 16945 -680
rect 17065 -650 17115 -640
rect 17065 -680 17075 -650
rect 17105 -680 17115 -650
rect 17065 -690 17115 -680
rect 17235 -650 17285 -640
rect 17235 -680 17245 -650
rect 17275 -680 17285 -650
rect 17235 -690 17285 -680
rect 17405 -650 17455 -640
rect 17405 -680 17415 -650
rect 17445 -680 17455 -650
rect 17405 -690 17455 -680
rect 17575 -650 17625 -640
rect 17575 -680 17585 -650
rect 17615 -680 17625 -650
rect 17575 -690 17625 -680
rect 17745 -650 17795 -640
rect 17745 -680 17755 -650
rect 17785 -680 17795 -650
rect 17745 -690 17795 -680
rect 17915 -650 17965 -640
rect 17915 -680 17925 -650
rect 17955 -680 17965 -650
rect 17915 -690 17965 -680
rect 18085 -650 18135 -640
rect 18085 -680 18095 -650
rect 18125 -680 18135 -650
rect 18085 -690 18135 -680
rect 18255 -650 18305 -640
rect 18255 -680 18265 -650
rect 18295 -680 18305 -650
rect 18255 -690 18305 -680
rect 18425 -650 18475 -640
rect 18425 -680 18435 -650
rect 18465 -680 18475 -650
rect 18425 -690 18475 -680
rect 18595 -650 18645 -640
rect 18595 -680 18605 -650
rect 18635 -680 18645 -650
rect 18595 -690 18645 -680
rect 18765 -650 18815 -640
rect 18765 -680 18775 -650
rect 18805 -680 18815 -650
rect 18765 -690 18815 -680
rect 18935 -650 18985 -640
rect 18935 -680 18945 -650
rect 18975 -680 18985 -650
rect 18935 -690 18985 -680
rect 19105 -650 19155 -640
rect 19105 -680 19115 -650
rect 19145 -680 19155 -650
rect 19105 -690 19155 -680
rect 19275 -650 19325 -640
rect 19275 -680 19285 -650
rect 19315 -680 19325 -650
rect 19275 -690 19325 -680
rect 19445 -650 19495 -640
rect 19445 -680 19455 -650
rect 19485 -680 19495 -650
rect 19445 -690 19495 -680
rect 19615 -650 19665 -640
rect 19615 -680 19625 -650
rect 19655 -680 19665 -650
rect 19615 -690 19665 -680
rect 19785 -650 19835 -640
rect 19785 -680 19795 -650
rect 19825 -680 19835 -650
rect 19785 -690 19835 -680
rect 19955 -650 20005 -640
rect 19955 -680 19965 -650
rect 19995 -680 20005 -650
rect 19955 -690 20005 -680
rect 20125 -650 20175 -640
rect 20125 -680 20135 -650
rect 20165 -680 20175 -650
rect 20125 -690 20175 -680
rect 20295 -650 20345 -640
rect 20295 -680 20305 -650
rect 20335 -680 20345 -650
rect 20295 -690 20345 -680
rect 20465 -650 20515 -640
rect 20465 -680 20475 -650
rect 20505 -680 20515 -650
rect 20465 -690 20515 -680
rect 20635 -650 20685 -640
rect 20635 -680 20645 -650
rect 20675 -680 20685 -650
rect 20635 -690 20685 -680
rect 20805 -650 20855 -640
rect 20805 -680 20815 -650
rect 20845 -680 20855 -650
rect 20805 -690 20855 -680
rect 20975 -650 21025 -640
rect 20975 -680 20985 -650
rect 21015 -680 21025 -650
rect 20975 -690 21025 -680
rect 21145 -650 21195 -640
rect 21145 -680 21155 -650
rect 21185 -680 21195 -650
rect 21145 -690 21195 -680
rect 21315 -650 21365 -640
rect 21315 -680 21325 -650
rect 21355 -680 21365 -650
rect 21315 -690 21365 -680
rect 21485 -650 21535 -640
rect 21485 -680 21495 -650
rect 21525 -680 21535 -650
rect 21485 -690 21535 -680
rect 21655 -650 21705 -640
rect 21655 -680 21665 -650
rect 21695 -680 21705 -650
rect 21655 -690 21705 -680
rect 21825 -650 21875 -640
rect 21825 -680 21835 -650
rect 21865 -680 21875 -650
rect 21825 -690 21875 -680
rect 21995 -650 22045 -640
rect 21995 -680 22005 -650
rect 22035 -680 22045 -650
rect 21995 -690 22045 -680
rect 22165 -650 22215 -640
rect 22165 -680 22175 -650
rect 22205 -680 22215 -650
rect 22165 -690 22215 -680
rect 22335 -650 22385 -640
rect 22335 -680 22345 -650
rect 22375 -680 22385 -650
rect 22335 -690 22385 -680
rect 22505 -650 22555 -640
rect 22505 -680 22515 -650
rect 22545 -680 22555 -650
rect 22505 -690 22555 -680
rect 22675 -650 22725 -640
rect 22675 -680 22685 -650
rect 22715 -680 22725 -650
rect 22675 -690 22725 -680
rect 22845 -650 22895 -640
rect 22845 -680 22855 -650
rect 22885 -680 22895 -650
rect 22845 -690 22895 -680
rect 23015 -650 23065 -640
rect 23015 -680 23025 -650
rect 23055 -680 23065 -650
rect 23015 -690 23065 -680
rect 23185 -650 23235 -640
rect 23185 -680 23195 -650
rect 23225 -680 23235 -650
rect 23185 -690 23235 -680
rect 23355 -650 23405 -640
rect 23355 -680 23365 -650
rect 23395 -680 23405 -650
rect 23355 -690 23405 -680
rect 23525 -650 23575 -640
rect 23525 -680 23535 -650
rect 23565 -680 23575 -650
rect 23525 -690 23575 -680
rect 23695 -650 23745 -640
rect 23695 -680 23705 -650
rect 23735 -680 23745 -650
rect 23695 -690 23745 -680
rect 23865 -650 23915 -640
rect 23865 -680 23875 -650
rect 23905 -680 23915 -650
rect 23865 -690 23915 -680
rect 24035 -650 24085 -640
rect 24035 -680 24045 -650
rect 24075 -680 24085 -650
rect 24035 -690 24085 -680
rect 24205 -650 24255 -640
rect 24205 -680 24215 -650
rect 24245 -680 24255 -650
rect 24205 -690 24255 -680
rect 24375 -650 24425 -640
rect 24375 -680 24385 -650
rect 24415 -680 24425 -650
rect 24375 -690 24425 -680
rect 24545 -650 24595 -640
rect 24545 -680 24555 -650
rect 24585 -680 24595 -650
rect 24545 -690 24595 -680
rect 24715 -650 24765 -640
rect 24715 -680 24725 -650
rect 24755 -680 24765 -650
rect 24715 -690 24765 -680
rect 24885 -650 24935 -640
rect 24885 -680 24895 -650
rect 24925 -680 24935 -650
rect 24885 -690 24935 -680
rect 25055 -650 25105 -640
rect 25055 -680 25065 -650
rect 25095 -680 25105 -650
rect 25055 -690 25105 -680
rect 25225 -650 25275 -640
rect 25225 -680 25235 -650
rect 25265 -680 25275 -650
rect 25225 -690 25275 -680
rect 25395 -650 25445 -640
rect 25395 -680 25405 -650
rect 25435 -680 25445 -650
rect 25395 -690 25445 -680
rect 25565 -650 25615 -640
rect 25565 -680 25575 -650
rect 25605 -680 25615 -650
rect 25565 -690 25615 -680
rect 25735 -650 25785 -640
rect 25735 -680 25745 -650
rect 25775 -680 25785 -650
rect 25735 -690 25785 -680
rect 25905 -650 25955 -640
rect 25905 -680 25915 -650
rect 25945 -680 25955 -650
rect 25905 -690 25955 -680
rect 26075 -650 26125 -640
rect 26075 -680 26085 -650
rect 26115 -680 26125 -650
rect 26075 -690 26125 -680
rect 26245 -650 26295 -640
rect 26245 -680 26255 -650
rect 26285 -680 26295 -650
rect 26245 -690 26295 -680
rect 26415 -650 26465 -640
rect 26415 -680 26425 -650
rect 26455 -680 26465 -650
rect 26415 -690 26465 -680
rect 26585 -650 26635 -640
rect 26585 -680 26595 -650
rect 26625 -680 26635 -650
rect 26585 -690 26635 -680
rect 26755 -650 26805 -640
rect 26755 -680 26765 -650
rect 26795 -680 26805 -650
rect 26755 -690 26805 -680
rect 26925 -650 26975 -640
rect 26925 -680 26935 -650
rect 26965 -680 26975 -650
rect 26925 -690 26975 -680
rect 27095 -650 27145 -640
rect 27095 -680 27105 -650
rect 27135 -680 27145 -650
rect 27095 -690 27145 -680
rect 27265 -650 27315 -640
rect 27265 -680 27275 -650
rect 27305 -680 27315 -650
rect 27265 -690 27315 -680
rect 27435 -650 27485 -640
rect 27435 -680 27445 -650
rect 27475 -680 27485 -650
rect 27435 -690 27485 -680
rect 27605 -650 27655 -640
rect 27605 -680 27615 -650
rect 27645 -680 27655 -650
rect 27605 -690 27655 -680
rect 27775 -650 27825 -640
rect 27775 -680 27785 -650
rect 27815 -680 27825 -650
rect 27775 -690 27825 -680
rect 27945 -650 27995 -640
rect 27945 -680 27955 -650
rect 27985 -680 27995 -650
rect 27945 -690 27995 -680
rect 28115 -650 28165 -640
rect 28115 -680 28125 -650
rect 28155 -680 28165 -650
rect 28115 -690 28165 -680
rect 28285 -650 28335 -640
rect 28285 -680 28295 -650
rect 28325 -680 28335 -650
rect 28285 -690 28335 -680
rect 28455 -650 28505 -640
rect 28455 -680 28465 -650
rect 28495 -680 28505 -650
rect 28455 -690 28505 -680
rect 28625 -650 28675 -640
rect 28625 -680 28635 -650
rect 28665 -680 28675 -650
rect 28625 -690 28675 -680
rect 28795 -650 28845 -640
rect 28795 -680 28805 -650
rect 28835 -680 28845 -650
rect 28795 -690 28845 -680
rect 28965 -650 29015 -640
rect 28965 -680 28975 -650
rect 29005 -680 29015 -650
rect 28965 -690 29015 -680
rect 29135 -650 29185 -640
rect 29135 -680 29145 -650
rect 29175 -680 29185 -650
rect 29135 -690 29185 -680
rect 29305 -650 29355 -640
rect 29305 -680 29315 -650
rect 29345 -680 29355 -650
rect 29305 -690 29355 -680
rect 29475 -650 29525 -640
rect 29475 -680 29485 -650
rect 29515 -680 29525 -650
rect 29475 -690 29525 -680
rect 29645 -650 29695 -640
rect 29645 -680 29655 -650
rect 29685 -680 29695 -650
rect 29645 -690 29695 -680
rect 29815 -650 29865 -640
rect 29815 -680 29825 -650
rect 29855 -680 29865 -650
rect 29815 -690 29865 -680
rect 29985 -650 30035 -640
rect 29985 -680 29995 -650
rect 30025 -680 30035 -650
rect 29985 -690 30035 -680
rect 30155 -650 30205 -640
rect 30155 -680 30165 -650
rect 30195 -680 30205 -650
rect 30155 -690 30205 -680
rect 30325 -650 30375 -640
rect 30325 -680 30335 -650
rect 30365 -680 30375 -650
rect 30325 -690 30375 -680
rect 30495 -650 30545 -640
rect 30495 -680 30505 -650
rect 30535 -680 30545 -650
rect 30495 -690 30545 -680
rect 30665 -650 30715 -640
rect 30665 -680 30675 -650
rect 30705 -680 30715 -650
rect 30665 -690 30715 -680
rect 30835 -650 30885 -640
rect 30835 -680 30845 -650
rect 30875 -680 30885 -650
rect 30835 -690 30885 -680
rect 31005 -650 31055 -640
rect 31005 -680 31015 -650
rect 31045 -680 31055 -650
rect 31005 -690 31055 -680
rect 31175 -650 31225 -640
rect 31175 -680 31185 -650
rect 31215 -680 31225 -650
rect 31175 -690 31225 -680
rect 31345 -650 31395 -640
rect 31345 -680 31355 -650
rect 31385 -680 31395 -650
rect 31345 -690 31395 -680
rect 31515 -650 31565 -640
rect 31515 -680 31525 -650
rect 31555 -680 31565 -650
rect 31515 -690 31565 -680
rect 31685 -650 31735 -640
rect 31685 -680 31695 -650
rect 31725 -680 31735 -650
rect 31685 -690 31735 -680
rect 31855 -650 31905 -640
rect 31855 -680 31865 -650
rect 31895 -680 31905 -650
rect 31855 -690 31905 -680
rect 32025 -650 32075 -640
rect 32025 -680 32035 -650
rect 32065 -680 32075 -650
rect 32025 -690 32075 -680
rect 32195 -650 32245 -640
rect 32195 -680 32205 -650
rect 32235 -680 32245 -650
rect 32195 -690 32245 -680
rect 32365 -650 32415 -640
rect 32365 -680 32375 -650
rect 32405 -680 32415 -650
rect 32365 -690 32415 -680
rect 32535 -650 32585 -640
rect 32535 -680 32545 -650
rect 32575 -680 32585 -650
rect 32535 -690 32585 -680
rect 32705 -650 32755 -640
rect 32705 -680 32715 -650
rect 32745 -680 32755 -650
rect 32705 -690 32755 -680
rect 32875 -650 32925 -640
rect 32875 -680 32885 -650
rect 32915 -680 32925 -650
rect 32875 -690 32925 -680
rect 33045 -650 33095 -640
rect 33045 -680 33055 -650
rect 33085 -680 33095 -650
rect 33045 -690 33095 -680
rect 33215 -650 33265 -640
rect 33215 -680 33225 -650
rect 33255 -680 33265 -650
rect 33215 -690 33265 -680
rect 33385 -650 33435 -640
rect 33385 -680 33395 -650
rect 33425 -680 33435 -650
rect 33385 -690 33435 -680
rect 33555 -650 33605 -640
rect 33555 -680 33565 -650
rect 33595 -680 33605 -650
rect 33555 -690 33605 -680
rect 33725 -650 33775 -640
rect 33725 -680 33735 -650
rect 33765 -680 33775 -650
rect 33725 -690 33775 -680
rect 33895 -650 33945 -640
rect 33895 -680 33905 -650
rect 33935 -680 33945 -650
rect 33895 -690 33945 -680
rect 34065 -650 34115 -640
rect 34065 -680 34075 -650
rect 34105 -680 34115 -650
rect 34065 -690 34115 -680
rect 34235 -650 34285 -640
rect 34235 -680 34245 -650
rect 34275 -680 34285 -650
rect 34235 -690 34285 -680
rect 34405 -650 34455 -640
rect 34405 -680 34415 -650
rect 34445 -680 34455 -650
rect 34405 -690 34455 -680
rect 34575 -650 34625 -640
rect 34575 -680 34585 -650
rect 34615 -680 34625 -650
rect 34575 -690 34625 -680
rect 34745 -650 34795 -640
rect 34745 -680 34755 -650
rect 34785 -680 34795 -650
rect 34745 -690 34795 -680
rect 34915 -650 34965 -640
rect 34915 -680 34925 -650
rect 34955 -680 34965 -650
rect 34915 -690 34965 -680
rect 35085 -650 35135 -640
rect 35085 -680 35095 -650
rect 35125 -680 35135 -650
rect 35085 -690 35135 -680
rect 35255 -650 35305 -640
rect 35255 -680 35265 -650
rect 35295 -680 35305 -650
rect 35255 -690 35305 -680
rect 35425 -650 35475 -640
rect 35425 -680 35435 -650
rect 35465 -680 35475 -650
rect 35425 -690 35475 -680
rect 35595 -650 35645 -640
rect 35595 -680 35605 -650
rect 35635 -680 35645 -650
rect 35595 -690 35645 -680
rect 35765 -650 35815 -640
rect 35765 -680 35775 -650
rect 35805 -680 35815 -650
rect 35765 -690 35815 -680
rect 35935 -650 35985 -640
rect 35935 -680 35945 -650
rect 35975 -680 35985 -650
rect 35935 -690 35985 -680
rect 36105 -650 36155 -640
rect 36105 -680 36115 -650
rect 36145 -680 36155 -650
rect 36105 -690 36155 -680
rect 36275 -650 36325 -640
rect 36275 -680 36285 -650
rect 36315 -680 36325 -650
rect 36275 -690 36325 -680
rect 36445 -650 36495 -640
rect 36445 -680 36455 -650
rect 36485 -680 36495 -650
rect 36445 -690 36495 -680
rect 36615 -650 36665 -640
rect 36615 -680 36625 -650
rect 36655 -680 36665 -650
rect 36615 -690 36665 -680
rect 36785 -650 36835 -640
rect 36785 -680 36795 -650
rect 36825 -680 36835 -650
rect 36785 -690 36835 -680
rect 36955 -650 37005 -640
rect 36955 -680 36965 -650
rect 36995 -680 37005 -650
rect 36955 -690 37005 -680
rect 37125 -650 37175 -640
rect 37125 -680 37135 -650
rect 37165 -680 37175 -650
rect 37125 -690 37175 -680
rect 37295 -650 37345 -640
rect 37295 -680 37305 -650
rect 37335 -680 37345 -650
rect 37295 -690 37345 -680
rect 37465 -650 37515 -640
rect 37465 -680 37475 -650
rect 37505 -680 37515 -650
rect 37465 -690 37515 -680
rect 37635 -650 37685 -640
rect 37635 -680 37645 -650
rect 37675 -680 37685 -650
rect 37635 -690 37685 -680
rect 37805 -650 37855 -640
rect 37805 -680 37815 -650
rect 37845 -680 37855 -650
rect 37805 -690 37855 -680
rect 37975 -650 38025 -640
rect 37975 -680 37985 -650
rect 38015 -680 38025 -650
rect 37975 -690 38025 -680
rect 38145 -650 38195 -640
rect 38145 -680 38155 -650
rect 38185 -680 38195 -650
rect 38145 -690 38195 -680
rect 38315 -650 38365 -640
rect 38315 -680 38325 -650
rect 38355 -680 38365 -650
rect 38315 -690 38365 -680
rect 38485 -650 38535 -640
rect 38485 -680 38495 -650
rect 38525 -680 38535 -650
rect 38485 -690 38535 -680
rect 38655 -650 38705 -640
rect 38655 -680 38665 -650
rect 38695 -680 38705 -650
rect 38655 -690 38705 -680
rect 38825 -650 38875 -640
rect 38825 -680 38835 -650
rect 38865 -680 38875 -650
rect 38825 -690 38875 -680
rect 38995 -650 39045 -640
rect 38995 -680 39005 -650
rect 39035 -680 39045 -650
rect 38995 -690 39045 -680
rect 39165 -650 39215 -640
rect 39165 -680 39175 -650
rect 39205 -680 39215 -650
rect 39165 -690 39215 -680
rect 39335 -650 39385 -640
rect 39335 -680 39345 -650
rect 39375 -680 39385 -650
rect 39335 -690 39385 -680
rect 39505 -650 39555 -640
rect 39505 -680 39515 -650
rect 39545 -680 39555 -650
rect 39505 -690 39555 -680
rect 39675 -650 39725 -640
rect 39675 -680 39685 -650
rect 39715 -680 39725 -650
rect 39675 -690 39725 -680
rect 39845 -650 39895 -640
rect 39845 -680 39855 -650
rect 39885 -680 39895 -650
rect 39845 -690 39895 -680
rect 40015 -650 40065 -640
rect 40015 -680 40025 -650
rect 40055 -680 40065 -650
rect 40015 -690 40065 -680
rect 40185 -650 40235 -640
rect 40185 -680 40195 -650
rect 40225 -680 40235 -650
rect 40185 -690 40235 -680
rect 40355 -650 40405 -640
rect 40355 -680 40365 -650
rect 40395 -680 40405 -650
rect 40355 -690 40405 -680
rect 40525 -650 40575 -640
rect 40525 -680 40535 -650
rect 40565 -680 40575 -650
rect 40525 -690 40575 -680
rect 40695 -650 40745 -640
rect 40695 -680 40705 -650
rect 40735 -680 40745 -650
rect 40695 -690 40745 -680
rect 40865 -650 40915 -640
rect 40865 -680 40875 -650
rect 40905 -680 40915 -650
rect 40865 -690 40915 -680
rect 41035 -650 41085 -640
rect 41035 -680 41045 -650
rect 41075 -680 41085 -650
rect 41035 -690 41085 -680
rect 41205 -650 41255 -640
rect 41205 -680 41215 -650
rect 41245 -680 41255 -650
rect 41205 -690 41255 -680
rect 41375 -650 41425 -640
rect 41375 -680 41385 -650
rect 41415 -680 41425 -650
rect 41375 -690 41425 -680
rect 41545 -650 41595 -640
rect 41545 -680 41555 -650
rect 41585 -680 41595 -650
rect 41545 -690 41595 -680
rect 41715 -650 41765 -640
rect 41715 -680 41725 -650
rect 41755 -680 41765 -650
rect 41715 -690 41765 -680
rect 41885 -650 41935 -640
rect 41885 -680 41895 -650
rect 41925 -680 41935 -650
rect 41885 -690 41935 -680
rect 42055 -650 42105 -640
rect 42055 -680 42065 -650
rect 42095 -680 42105 -650
rect 42055 -690 42105 -680
rect 42225 -650 42275 -640
rect 42225 -680 42235 -650
rect 42265 -680 42275 -650
rect 42225 -690 42275 -680
rect 42395 -650 42445 -640
rect 42395 -680 42405 -650
rect 42435 -680 42445 -650
rect 42395 -690 42445 -680
rect 42565 -650 42615 -640
rect 42565 -680 42575 -650
rect 42605 -680 42615 -650
rect 42565 -690 42615 -680
rect 42735 -650 42785 -640
rect 42735 -680 42745 -650
rect 42775 -680 42785 -650
rect 42735 -690 42785 -680
rect 42905 -650 42955 -640
rect 42905 -680 42915 -650
rect 42945 -680 42955 -650
rect 42905 -690 42955 -680
rect 43075 -650 43125 -640
rect 43075 -680 43085 -650
rect 43115 -680 43125 -650
rect 43075 -690 43125 -680
rect 43245 -650 43295 -640
rect 43245 -680 43255 -650
rect 43285 -680 43295 -650
rect 43245 -690 43295 -680
rect 43415 -650 43465 -640
rect 43415 -680 43425 -650
rect 43455 -680 43465 -650
rect 43415 -690 43465 -680
rect 43585 -650 43635 -640
rect 43585 -680 43595 -650
rect 43625 -680 43635 -650
rect 43585 -690 43635 -680
<< via1 >>
rect 35 15 65 55
rect 225 175 255 205
rect 395 175 425 205
rect 565 175 595 205
rect 760 175 790 205
rect 930 175 960 205
rect 1100 175 1130 205
rect 1270 175 1300 205
rect 1440 175 1470 205
rect 1610 175 1640 205
rect 1780 175 1810 205
rect 1950 175 1980 205
rect 2120 175 2150 205
rect 2270 175 2300 205
rect 2440 175 2470 205
rect 2610 175 2640 205
rect 2780 175 2810 205
rect 2950 175 2980 205
rect 3120 175 3150 205
rect 3290 175 3320 205
rect 3460 175 3490 205
rect 3630 175 3660 205
rect 3800 175 3830 205
rect 3970 175 4000 205
rect 4140 175 4170 205
rect 4310 175 4340 205
rect 4480 175 4510 205
rect 4650 175 4680 205
rect 4820 175 4850 205
rect 4990 175 5020 205
rect 5160 175 5190 205
rect 5330 175 5360 205
rect 5500 175 5530 205
rect 5670 175 5700 205
rect 5840 175 5870 205
rect 6010 175 6040 205
rect 6180 175 6210 205
rect 6350 175 6380 205
rect 6520 175 6550 205
rect 6690 175 6720 205
rect 6860 175 6890 205
rect 7030 175 7060 205
rect 7200 175 7230 205
rect 7370 175 7400 205
rect 7540 175 7570 205
rect 7710 175 7740 205
rect 7860 175 7890 205
rect 8030 175 8060 205
rect 8200 175 8230 205
rect 8370 175 8400 205
rect 8540 175 8570 205
rect 8710 175 8740 205
rect 8880 175 8910 205
rect 9050 175 9080 205
rect 9220 175 9250 205
rect 9390 175 9420 205
rect 9560 175 9590 205
rect 9730 175 9760 205
rect 9900 175 9930 205
rect 10070 175 10100 205
rect 10240 175 10270 205
rect 10410 175 10440 205
rect 10580 175 10610 205
rect 10750 175 10780 205
rect 10920 175 10950 205
rect 11090 175 11120 205
rect 11260 175 11290 205
rect 11430 175 11460 205
rect 11600 175 11630 205
rect 11770 175 11800 205
rect 11940 175 11970 205
rect 12110 175 12140 205
rect 12280 175 12310 205
rect 12450 175 12480 205
rect 12620 175 12650 205
rect 12790 175 12820 205
rect 12960 175 12990 205
rect 13130 175 13160 205
rect 13300 175 13330 205
rect 13470 175 13500 205
rect 13640 175 13670 205
rect 13810 175 13840 205
rect 13980 175 14010 205
rect 14150 175 14180 205
rect 14320 175 14350 205
rect 14490 175 14520 205
rect 14660 175 14690 205
rect 14830 175 14860 205
rect 15000 175 15030 205
rect 15170 175 15200 205
rect 15340 175 15370 205
rect 15510 175 15540 205
rect 15680 175 15710 205
rect 15850 175 15880 205
rect 16020 175 16050 205
rect 16190 175 16220 205
rect 16360 175 16390 205
rect 16530 175 16560 205
rect 16700 175 16730 205
rect 16870 175 16900 205
rect 17040 175 17070 205
rect 17210 175 17240 205
rect 17380 175 17410 205
rect 17550 175 17580 205
rect 17720 175 17750 205
rect 17890 175 17920 205
rect 18060 175 18090 205
rect 18230 175 18260 205
rect 18400 175 18430 205
rect 18570 175 18600 205
rect 18740 175 18770 205
rect 18910 175 18940 205
rect 19080 175 19110 205
rect 19250 175 19280 205
rect 19420 175 19450 205
rect 19590 175 19620 205
rect 19760 175 19790 205
rect 19930 175 19960 205
rect 20100 175 20130 205
rect 20270 175 20300 205
rect 20440 175 20470 205
rect 20610 175 20640 205
rect 20780 175 20810 205
rect 20950 175 20980 205
rect 21120 175 21150 205
rect 21290 175 21320 205
rect 21460 175 21490 205
rect 21630 175 21660 205
rect 21800 175 21830 205
rect 21970 175 22000 205
rect 22140 175 22170 205
rect 22310 175 22340 205
rect 22480 175 22510 205
rect 22650 175 22680 205
rect 22820 175 22850 205
rect 22990 175 23020 205
rect 23160 175 23190 205
rect 23330 175 23360 205
rect 23500 175 23530 205
rect 23670 175 23700 205
rect 23840 175 23870 205
rect 24010 175 24040 205
rect 24180 175 24210 205
rect 24350 175 24380 205
rect 24520 175 24550 205
rect 24690 175 24720 205
rect 24860 175 24890 205
rect 25030 175 25060 205
rect 25200 175 25230 205
rect 25370 175 25400 205
rect 25540 175 25570 205
rect 25710 175 25740 205
rect 25880 175 25910 205
rect 26050 175 26080 205
rect 26220 175 26250 205
rect 26390 175 26420 205
rect 26560 175 26590 205
rect 26730 175 26760 205
rect 26900 175 26930 205
rect 27070 175 27100 205
rect 27240 175 27270 205
rect 27410 175 27440 205
rect 27580 175 27610 205
rect 27750 175 27780 205
rect 27920 175 27950 205
rect 28090 175 28120 205
rect 28260 175 28290 205
rect 28430 175 28460 205
rect 28600 175 28630 205
rect 28770 175 28800 205
rect 28940 175 28970 205
rect 29110 175 29140 205
rect 29280 175 29310 205
rect 29450 175 29480 205
rect 29620 175 29650 205
rect 310 65 340 100
rect 225 10 255 40
rect 480 65 510 100
rect 395 10 425 40
rect 845 65 875 100
rect 565 10 595 40
rect 760 10 790 40
rect 1015 65 1045 100
rect 930 10 960 40
rect 1185 65 1215 100
rect 1100 10 1130 40
rect 1355 65 1385 100
rect 1270 10 1300 40
rect 1525 65 1555 100
rect 1440 10 1470 40
rect 1695 65 1725 100
rect 1610 10 1640 40
rect 1865 65 1895 100
rect 1780 10 1810 40
rect 2035 65 2065 100
rect 1950 10 1980 40
rect 2355 65 2385 100
rect 2120 10 2150 40
rect 2270 10 2300 40
rect 2525 65 2555 100
rect 2440 10 2470 40
rect 2695 65 2725 100
rect 2610 10 2640 40
rect 2865 65 2895 100
rect 2780 10 2810 40
rect 3035 65 3065 100
rect 2950 10 2980 40
rect 3205 65 3235 100
rect 3120 10 3150 40
rect 3375 65 3405 100
rect 3290 10 3320 40
rect 3545 65 3575 100
rect 3460 10 3490 40
rect 3715 65 3745 100
rect 3630 10 3660 40
rect 3885 65 3915 100
rect 3800 10 3830 40
rect 4055 65 4085 100
rect 3970 10 4000 40
rect 4225 65 4255 100
rect 4140 10 4170 40
rect 4395 65 4425 100
rect 4310 10 4340 40
rect 4565 65 4595 100
rect 4480 10 4510 40
rect 4735 65 4765 100
rect 4650 10 4680 40
rect 4905 65 4935 100
rect 4820 10 4850 40
rect 5075 65 5105 100
rect 4990 10 5020 40
rect 5245 65 5275 100
rect 5160 10 5190 40
rect 5415 65 5445 100
rect 5330 10 5360 40
rect 5585 65 5615 100
rect 5500 10 5530 40
rect 5755 65 5785 100
rect 5670 10 5700 40
rect 5925 65 5955 100
rect 5840 10 5870 40
rect 6095 65 6125 100
rect 6010 10 6040 40
rect 6265 65 6295 100
rect 6180 10 6210 40
rect 6435 65 6465 100
rect 6350 10 6380 40
rect 6605 65 6635 100
rect 6520 10 6550 40
rect 6775 65 6805 100
rect 6690 10 6720 40
rect 6945 65 6975 100
rect 6860 10 6890 40
rect 7115 65 7145 100
rect 7030 10 7060 40
rect 7285 65 7315 100
rect 7200 10 7230 40
rect 7455 65 7485 100
rect 7370 10 7400 40
rect 7625 65 7655 100
rect 7540 10 7570 40
rect 7945 65 7975 100
rect 7710 10 7740 40
rect 7860 10 7890 40
rect 8115 65 8145 100
rect 8030 10 8060 40
rect 8285 65 8315 100
rect 8200 10 8230 40
rect 8455 65 8485 100
rect 8370 10 8400 40
rect 8625 65 8655 100
rect 8540 10 8570 40
rect 8795 65 8825 100
rect 8710 10 8740 40
rect 8965 65 8995 100
rect 8880 10 8910 40
rect 9135 65 9165 100
rect 9050 10 9080 40
rect 9305 65 9335 100
rect 9220 10 9250 40
rect 9475 65 9505 100
rect 9390 10 9420 40
rect 9645 65 9675 100
rect 9560 10 9590 40
rect 9815 65 9845 100
rect 9730 10 9760 40
rect 9985 65 10015 100
rect 9900 10 9930 40
rect 10155 65 10185 100
rect 10070 10 10100 40
rect 10325 65 10355 100
rect 10240 10 10270 40
rect 10495 65 10525 100
rect 10410 10 10440 40
rect 10665 65 10695 100
rect 10580 10 10610 40
rect 10835 65 10865 100
rect 10750 10 10780 40
rect 11005 65 11035 100
rect 10920 10 10950 40
rect 11175 65 11205 100
rect 11090 10 11120 40
rect 11345 65 11375 100
rect 11260 10 11290 40
rect 11515 65 11545 100
rect 11430 10 11460 40
rect 11685 65 11715 100
rect 11600 10 11630 40
rect 11855 65 11885 100
rect 11770 10 11800 40
rect 12025 65 12055 100
rect 11940 10 11970 40
rect 12195 65 12225 100
rect 12110 10 12140 40
rect 12365 65 12395 100
rect 12280 10 12310 40
rect 12535 65 12565 100
rect 12450 10 12480 40
rect 12705 65 12735 100
rect 12620 10 12650 40
rect 12875 65 12905 100
rect 12790 10 12820 40
rect 13045 65 13075 100
rect 12960 10 12990 40
rect 13215 65 13245 100
rect 13130 10 13160 40
rect 13385 65 13415 100
rect 13300 10 13330 40
rect 13555 65 13585 100
rect 13470 10 13500 40
rect 13725 65 13755 100
rect 13640 10 13670 40
rect 13895 65 13925 100
rect 13810 10 13840 40
rect 14065 65 14095 100
rect 13980 10 14010 40
rect 14235 65 14265 100
rect 14150 10 14180 40
rect 14405 65 14435 100
rect 14320 10 14350 40
rect 14575 65 14605 100
rect 14490 10 14520 40
rect 14745 65 14775 100
rect 14660 10 14690 40
rect 14915 65 14945 100
rect 14830 10 14860 40
rect 15085 65 15115 100
rect 15000 10 15030 40
rect 15255 65 15285 100
rect 15170 10 15200 40
rect 15425 65 15455 100
rect 15340 10 15370 40
rect 15595 65 15625 100
rect 15510 10 15540 40
rect 15765 65 15795 100
rect 15680 10 15710 40
rect 15935 65 15965 100
rect 15850 10 15880 40
rect 16105 65 16135 100
rect 16020 10 16050 40
rect 16275 65 16305 100
rect 16190 10 16220 40
rect 16445 65 16475 100
rect 16360 10 16390 40
rect 16615 65 16645 100
rect 16530 10 16560 40
rect 16785 65 16815 100
rect 16700 10 16730 40
rect 16955 65 16985 100
rect 16870 10 16900 40
rect 17125 65 17155 100
rect 17040 10 17070 40
rect 17295 65 17325 100
rect 17210 10 17240 40
rect 17465 65 17495 100
rect 17380 10 17410 40
rect 17635 65 17665 100
rect 17550 10 17580 40
rect 17805 65 17835 100
rect 17720 10 17750 40
rect 17975 65 18005 100
rect 17890 10 17920 40
rect 18145 65 18175 100
rect 18060 10 18090 40
rect 18315 65 18345 100
rect 18230 10 18260 40
rect 18485 65 18515 100
rect 18400 10 18430 40
rect 18655 65 18685 100
rect 18570 10 18600 40
rect 18825 65 18855 100
rect 18740 10 18770 40
rect 18995 65 19025 100
rect 18910 10 18940 40
rect 19165 65 19195 100
rect 19080 10 19110 40
rect 19335 65 19365 100
rect 19250 10 19280 40
rect 19505 65 19535 100
rect 19420 10 19450 40
rect 19675 65 19705 100
rect 19590 10 19620 40
rect 19845 65 19875 100
rect 19760 10 19790 40
rect 20015 65 20045 100
rect 19930 10 19960 40
rect 20185 65 20215 100
rect 20100 10 20130 40
rect 20355 65 20385 100
rect 20270 10 20300 40
rect 20525 65 20555 100
rect 20440 10 20470 40
rect 20695 65 20725 100
rect 20610 10 20640 40
rect 20865 65 20895 100
rect 20780 10 20810 40
rect 21035 65 21065 100
rect 20950 10 20980 40
rect 21205 65 21235 100
rect 21120 10 21150 40
rect 21375 65 21405 100
rect 21290 10 21320 40
rect 21545 65 21575 100
rect 21460 10 21490 40
rect 21715 65 21745 100
rect 21630 10 21660 40
rect 21885 65 21915 100
rect 21800 10 21830 40
rect 22055 65 22085 100
rect 21970 10 22000 40
rect 22225 65 22255 100
rect 22140 10 22170 40
rect 22395 65 22425 100
rect 22310 10 22340 40
rect 22565 65 22595 100
rect 22480 10 22510 40
rect 22735 65 22765 100
rect 22650 10 22680 40
rect 22905 65 22935 100
rect 22820 10 22850 40
rect 23075 65 23105 100
rect 22990 10 23020 40
rect 23245 65 23275 100
rect 23160 10 23190 40
rect 23415 65 23445 100
rect 23330 10 23360 40
rect 23585 65 23615 100
rect 23500 10 23530 40
rect 23755 65 23785 100
rect 23670 10 23700 40
rect 23925 65 23955 100
rect 23840 10 23870 40
rect 24095 65 24125 100
rect 24010 10 24040 40
rect 24265 65 24295 100
rect 24180 10 24210 40
rect 24435 65 24465 100
rect 24350 10 24380 40
rect 24605 65 24635 100
rect 24520 10 24550 40
rect 24775 65 24805 100
rect 24690 10 24720 40
rect 24945 65 24975 100
rect 24860 10 24890 40
rect 25115 65 25145 100
rect 25030 10 25060 40
rect 25285 65 25315 100
rect 25200 10 25230 40
rect 25455 65 25485 100
rect 25370 10 25400 40
rect 25625 65 25655 100
rect 25540 10 25570 40
rect 25795 65 25825 100
rect 25710 10 25740 40
rect 25965 65 25995 100
rect 25880 10 25910 40
rect 26135 65 26165 100
rect 26050 10 26080 40
rect 26305 65 26335 100
rect 26220 10 26250 40
rect 26475 65 26505 100
rect 26390 10 26420 40
rect 26645 65 26675 100
rect 26560 10 26590 40
rect 26815 65 26845 100
rect 26730 10 26760 40
rect 26985 65 27015 100
rect 26900 10 26930 40
rect 27155 65 27185 100
rect 27070 10 27100 40
rect 27325 65 27355 100
rect 27240 10 27270 40
rect 27495 65 27525 100
rect 27410 10 27440 40
rect 27665 65 27695 100
rect 27580 10 27610 40
rect 27835 65 27865 100
rect 27750 10 27780 40
rect 28005 65 28035 100
rect 27920 10 27950 40
rect 28175 65 28205 100
rect 28090 10 28120 40
rect 28345 65 28375 100
rect 28260 10 28290 40
rect 28515 65 28545 100
rect 28430 10 28460 40
rect 28685 65 28715 100
rect 28600 10 28630 40
rect 28855 65 28885 100
rect 28770 10 28800 40
rect 29025 65 29055 100
rect 28940 10 28970 40
rect 29195 65 29225 100
rect 29110 10 29140 40
rect 29365 65 29395 100
rect 29280 10 29310 40
rect 29535 65 29565 100
rect 29450 10 29480 40
rect 29620 10 29650 40
rect 100 -60 130 -30
rect 265 -60 300 -30
rect 350 -60 385 -30
rect 435 -60 470 -30
rect 520 -60 555 -30
rect 800 -60 835 -30
rect 885 -60 920 -30
rect 970 -60 1005 -30
rect 1055 -60 1090 -30
rect 1140 -60 1175 -30
rect 1225 -60 1260 -30
rect 1310 -60 1345 -30
rect 1395 -60 1430 -30
rect 1480 -60 1515 -30
rect 1565 -60 1600 -30
rect 1650 -60 1685 -30
rect 1735 -60 1770 -30
rect 1820 -60 1855 -30
rect 1905 -60 1940 -30
rect 1990 -60 2025 -30
rect 2075 -60 2110 -30
rect 2310 -60 2345 -30
rect 2395 -60 2430 -30
rect 2480 -60 2515 -30
rect 2565 -60 2600 -30
rect 2650 -60 2685 -30
rect 2735 -60 2770 -30
rect 2820 -60 2855 -30
rect 2905 -60 2940 -30
rect 2990 -60 3025 -30
rect 3075 -60 3110 -30
rect 3160 -60 3195 -30
rect 3245 -60 3280 -30
rect 3330 -60 3365 -30
rect 3415 -60 3450 -30
rect 3500 -60 3535 -30
rect 3585 -60 3620 -30
rect 3670 -60 3705 -30
rect 3755 -60 3790 -30
rect 3840 -60 3875 -30
rect 3925 -60 3960 -30
rect 4010 -60 4045 -30
rect 4095 -60 4130 -30
rect 4180 -60 4215 -30
rect 4265 -60 4300 -30
rect 4350 -60 4385 -30
rect 4435 -60 4470 -30
rect 4520 -60 4555 -30
rect 4605 -60 4640 -30
rect 4690 -60 4725 -30
rect 4775 -60 4810 -30
rect 4860 -60 4895 -30
rect 4945 -60 4980 -30
rect 5030 -60 5065 -30
rect 5115 -60 5150 -30
rect 5200 -60 5235 -30
rect 5285 -60 5320 -30
rect 5370 -60 5405 -30
rect 5455 -60 5490 -30
rect 5540 -60 5575 -30
rect 5625 -60 5660 -30
rect 5710 -60 5745 -30
rect 5795 -60 5830 -30
rect 5880 -60 5915 -30
rect 5965 -60 6000 -30
rect 6050 -60 6085 -30
rect 6135 -60 6170 -30
rect 6220 -60 6255 -30
rect 6305 -60 6340 -30
rect 6390 -60 6425 -30
rect 6475 -60 6510 -30
rect 6560 -60 6595 -30
rect 6645 -60 6680 -30
rect 6730 -60 6765 -30
rect 6815 -60 6850 -30
rect 6900 -60 6935 -30
rect 6985 -60 7020 -30
rect 7070 -60 7105 -30
rect 7155 -60 7190 -30
rect 7240 -60 7275 -30
rect 7325 -60 7360 -30
rect 7410 -60 7445 -30
rect 7495 -60 7530 -30
rect 7580 -60 7615 -30
rect 7665 -60 7700 -30
rect 7900 -60 7935 -30
rect 7985 -60 8020 -30
rect 8070 -60 8105 -30
rect 8155 -60 8190 -30
rect 8240 -60 8275 -30
rect 8325 -60 8360 -30
rect 8410 -60 8445 -30
rect 8495 -60 8530 -30
rect 8580 -60 8615 -30
rect 8665 -60 8700 -30
rect 8750 -60 8785 -30
rect 8835 -60 8870 -30
rect 8920 -60 8955 -30
rect 9005 -60 9040 -30
rect 9090 -60 9125 -30
rect 9175 -60 9210 -30
rect 9260 -60 9295 -30
rect 9345 -60 9380 -30
rect 9430 -60 9465 -30
rect 9515 -60 9550 -30
rect 9600 -60 9635 -30
rect 9685 -60 9720 -30
rect 9770 -60 9805 -30
rect 9855 -60 9890 -30
rect 9940 -60 9975 -30
rect 10025 -60 10060 -30
rect 10110 -60 10145 -30
rect 10195 -60 10230 -30
rect 10280 -60 10315 -30
rect 10365 -60 10400 -30
rect 10450 -60 10485 -30
rect 10535 -60 10570 -30
rect 10620 -60 10655 -30
rect 10705 -60 10740 -30
rect 10790 -60 10825 -30
rect 10875 -60 10910 -30
rect 10960 -60 10995 -30
rect 11045 -60 11080 -30
rect 11130 -60 11165 -30
rect 11215 -60 11250 -30
rect 11300 -60 11335 -30
rect 11385 -60 11420 -30
rect 11470 -60 11505 -30
rect 11555 -60 11590 -30
rect 11640 -60 11675 -30
rect 11725 -60 11760 -30
rect 11810 -60 11845 -30
rect 11895 -60 11930 -30
rect 11980 -60 12015 -30
rect 12065 -60 12100 -30
rect 12150 -60 12185 -30
rect 12235 -60 12270 -30
rect 12320 -60 12355 -30
rect 12405 -60 12440 -30
rect 12490 -60 12525 -30
rect 12575 -60 12610 -30
rect 12660 -60 12695 -30
rect 12745 -60 12780 -30
rect 12830 -60 12865 -30
rect 12915 -60 12950 -30
rect 13000 -60 13035 -30
rect 13085 -60 13120 -30
rect 13170 -60 13205 -30
rect 13255 -60 13290 -30
rect 13340 -60 13375 -30
rect 13425 -60 13460 -30
rect 13510 -60 13545 -30
rect 13595 -60 13630 -30
rect 13680 -60 13715 -30
rect 13765 -60 13800 -30
rect 13850 -60 13885 -30
rect 13935 -60 13970 -30
rect 14020 -60 14055 -30
rect 14105 -60 14140 -30
rect 14190 -60 14225 -30
rect 14275 -60 14310 -30
rect 14360 -60 14395 -30
rect 14445 -60 14480 -30
rect 14530 -60 14565 -30
rect 14615 -60 14650 -30
rect 14700 -60 14735 -30
rect 14785 -60 14820 -30
rect 14870 -60 14905 -30
rect 14955 -60 14990 -30
rect 15040 -60 15075 -30
rect 15125 -60 15160 -30
rect 15210 -60 15245 -30
rect 15295 -60 15330 -30
rect 15380 -60 15415 -30
rect 15465 -60 15500 -30
rect 15550 -60 15585 -30
rect 15635 -60 15670 -30
rect 15720 -60 15755 -30
rect 15805 -60 15840 -30
rect 15890 -60 15925 -30
rect 15975 -60 16010 -30
rect 16060 -60 16095 -30
rect 16145 -60 16180 -30
rect 16230 -60 16265 -30
rect 16315 -60 16350 -30
rect 16400 -60 16435 -30
rect 16485 -60 16520 -30
rect 16570 -60 16605 -30
rect 16655 -60 16690 -30
rect 16740 -60 16775 -30
rect 16825 -60 16860 -30
rect 16910 -60 16945 -30
rect 16995 -60 17030 -30
rect 17080 -60 17115 -30
rect 17165 -60 17200 -30
rect 17250 -60 17285 -30
rect 17335 -60 17370 -30
rect 17420 -60 17455 -30
rect 17505 -60 17540 -30
rect 17590 -60 17625 -30
rect 17675 -60 17710 -30
rect 17760 -60 17795 -30
rect 17845 -60 17880 -30
rect 17930 -60 17965 -30
rect 18015 -60 18050 -30
rect 18100 -60 18135 -30
rect 18185 -60 18220 -30
rect 18270 -60 18305 -30
rect 18355 -60 18390 -30
rect 18440 -60 18475 -30
rect 18525 -60 18560 -30
rect 18610 -60 18645 -30
rect 18695 -60 18730 -30
rect 18780 -60 18815 -30
rect 18865 -60 18900 -30
rect 18950 -60 18985 -30
rect 19035 -60 19070 -30
rect 19120 -60 19155 -30
rect 19205 -60 19240 -30
rect 19290 -60 19325 -30
rect 19375 -60 19410 -30
rect 19460 -60 19495 -30
rect 19545 -60 19580 -30
rect 19630 -60 19665 -30
rect 19715 -60 19750 -30
rect 19800 -60 19835 -30
rect 19885 -60 19920 -30
rect 19970 -60 20005 -30
rect 20055 -60 20090 -30
rect 20140 -60 20175 -30
rect 20225 -60 20260 -30
rect 20310 -60 20345 -30
rect 20395 -60 20430 -30
rect 20480 -60 20515 -30
rect 20565 -60 20600 -30
rect 20650 -60 20685 -30
rect 20735 -60 20770 -30
rect 20820 -60 20855 -30
rect 20905 -60 20940 -30
rect 20990 -60 21025 -30
rect 21075 -60 21110 -30
rect 21160 -60 21195 -30
rect 21245 -60 21280 -30
rect 21330 -60 21365 -30
rect 21415 -60 21450 -30
rect 21500 -60 21535 -30
rect 21585 -60 21620 -30
rect 21670 -60 21705 -30
rect 21755 -60 21790 -30
rect 21840 -60 21875 -30
rect 21925 -60 21960 -30
rect 22010 -60 22045 -30
rect 22095 -60 22130 -30
rect 22180 -60 22215 -30
rect 22265 -60 22300 -30
rect 22350 -60 22385 -30
rect 22435 -60 22470 -30
rect 22520 -60 22555 -30
rect 22605 -60 22640 -30
rect 22690 -60 22725 -30
rect 22775 -60 22810 -30
rect 22860 -60 22895 -30
rect 22945 -60 22980 -30
rect 23030 -60 23065 -30
rect 23115 -60 23150 -30
rect 23200 -60 23235 -30
rect 23285 -60 23320 -30
rect 23370 -60 23405 -30
rect 23455 -60 23490 -30
rect 23540 -60 23575 -30
rect 23625 -60 23660 -30
rect 23710 -60 23745 -30
rect 23795 -60 23830 -30
rect 23880 -60 23915 -30
rect 23965 -60 24000 -30
rect 24050 -60 24085 -30
rect 24135 -60 24170 -30
rect 24220 -60 24255 -30
rect 24305 -60 24340 -30
rect 24390 -60 24425 -30
rect 24475 -60 24510 -30
rect 24560 -60 24595 -30
rect 24645 -60 24680 -30
rect 24730 -60 24765 -30
rect 24815 -60 24850 -30
rect 24900 -60 24935 -30
rect 24985 -60 25020 -30
rect 25070 -60 25105 -30
rect 25155 -60 25190 -30
rect 25240 -60 25275 -30
rect 25325 -60 25360 -30
rect 25410 -60 25445 -30
rect 25495 -60 25530 -30
rect 25580 -60 25615 -30
rect 25665 -60 25700 -30
rect 25750 -60 25785 -30
rect 25835 -60 25870 -30
rect 25920 -60 25955 -30
rect 26005 -60 26040 -30
rect 26090 -60 26125 -30
rect 26175 -60 26210 -30
rect 26260 -60 26295 -30
rect 26345 -60 26380 -30
rect 26430 -60 26465 -30
rect 26515 -60 26550 -30
rect 26600 -60 26635 -30
rect 26685 -60 26720 -30
rect 26770 -60 26805 -30
rect 26855 -60 26890 -30
rect 26940 -60 26975 -30
rect 27025 -60 27060 -30
rect 27110 -60 27145 -30
rect 27195 -60 27230 -30
rect 27280 -60 27315 -30
rect 27365 -60 27400 -30
rect 27450 -60 27485 -30
rect 27535 -60 27570 -30
rect 27620 -60 27655 -30
rect 27705 -60 27740 -30
rect 27790 -60 27825 -30
rect 27875 -60 27910 -30
rect 27960 -60 27995 -30
rect 28045 -60 28080 -30
rect 28130 -60 28165 -30
rect 28215 -60 28250 -30
rect 28300 -60 28335 -30
rect 28385 -60 28420 -30
rect 28470 -60 28505 -30
rect 28555 -60 28590 -30
rect 28640 -60 28675 -30
rect 28725 -60 28760 -30
rect 28810 -60 28845 -30
rect 28895 -60 28930 -30
rect 28980 -60 29015 -30
rect 29065 -60 29100 -30
rect 29150 -60 29185 -30
rect 29235 -60 29270 -30
rect 29320 -60 29355 -30
rect 29405 -60 29440 -30
rect 29490 -60 29525 -30
rect 29575 -60 29610 -30
rect 115 -295 150 -265
rect 200 -295 235 -265
rect 285 -295 320 -265
rect 370 -295 405 -265
rect 455 -295 490 -265
rect 540 -295 575 -265
rect 625 -295 660 -265
rect 710 -295 745 -265
rect 795 -295 830 -265
rect 880 -295 915 -265
rect 965 -295 1000 -265
rect 1050 -295 1085 -265
rect 1135 -295 1170 -265
rect 1220 -295 1255 -265
rect 1305 -295 1340 -265
rect 1390 -295 1425 -265
rect 1475 -295 1510 -265
rect 1560 -295 1595 -265
rect 1645 -295 1680 -265
rect 1730 -295 1765 -265
rect 1815 -295 1850 -265
rect 1900 -295 1935 -265
rect 1985 -295 2020 -265
rect 2070 -295 2105 -265
rect 2155 -295 2190 -265
rect 2240 -295 2275 -265
rect 2325 -295 2360 -265
rect 2410 -295 2445 -265
rect 2495 -295 2530 -265
rect 2580 -295 2615 -265
rect 2665 -295 2700 -265
rect 2750 -295 2785 -265
rect 2835 -295 2870 -265
rect 2920 -295 2955 -265
rect 3005 -295 3040 -265
rect 3090 -295 3125 -265
rect 3175 -295 3210 -265
rect 3260 -295 3295 -265
rect 3345 -295 3380 -265
rect 3430 -295 3465 -265
rect 3515 -295 3550 -265
rect 3600 -295 3635 -265
rect 3685 -295 3720 -265
rect 3770 -295 3805 -265
rect 3855 -295 3890 -265
rect 3940 -295 3975 -265
rect 4025 -295 4060 -265
rect 4110 -295 4145 -265
rect 4195 -295 4230 -265
rect 4280 -295 4315 -265
rect 4365 -295 4400 -265
rect 4450 -295 4485 -265
rect 4535 -295 4570 -265
rect 4620 -295 4655 -265
rect 4705 -295 4740 -265
rect 4790 -295 4825 -265
rect 4875 -295 4910 -265
rect 4960 -295 4995 -265
rect 5045 -295 5080 -265
rect 5130 -295 5165 -265
rect 5215 -295 5250 -265
rect 5300 -295 5335 -265
rect 5385 -295 5420 -265
rect 5470 -295 5505 -265
rect 5555 -295 5590 -265
rect 5640 -295 5675 -265
rect 5725 -295 5760 -265
rect 5810 -295 5845 -265
rect 5895 -295 5930 -265
rect 5980 -295 6015 -265
rect 6065 -295 6100 -265
rect 6150 -295 6185 -265
rect 6235 -295 6270 -265
rect 6320 -295 6355 -265
rect 6405 -295 6440 -265
rect 6490 -295 6525 -265
rect 6575 -295 6610 -265
rect 6660 -295 6695 -265
rect 6745 -295 6780 -265
rect 6830 -295 6865 -265
rect 6915 -295 6950 -265
rect 7000 -295 7035 -265
rect 7085 -295 7120 -265
rect 7170 -295 7205 -265
rect 7255 -295 7290 -265
rect 7340 -295 7375 -265
rect 7425 -295 7460 -265
rect 7510 -295 7545 -265
rect 7595 -295 7630 -265
rect 7680 -295 7715 -265
rect 7765 -295 7800 -265
rect 7850 -295 7885 -265
rect 7935 -295 7970 -265
rect 8020 -295 8055 -265
rect 8105 -295 8140 -265
rect 8190 -295 8225 -265
rect 8275 -295 8310 -265
rect 8360 -295 8395 -265
rect 8445 -295 8480 -265
rect 8530 -295 8565 -265
rect 8615 -295 8650 -265
rect 8700 -295 8735 -265
rect 8785 -295 8820 -265
rect 8870 -295 8905 -265
rect 8955 -295 8990 -265
rect 9040 -295 9075 -265
rect 9125 -295 9160 -265
rect 9210 -295 9245 -265
rect 9295 -295 9330 -265
rect 9380 -295 9415 -265
rect 9465 -295 9500 -265
rect 9550 -295 9585 -265
rect 9635 -295 9670 -265
rect 9720 -295 9755 -265
rect 9805 -295 9840 -265
rect 9890 -295 9925 -265
rect 9975 -295 10010 -265
rect 10060 -295 10095 -265
rect 10145 -295 10180 -265
rect 10230 -295 10265 -265
rect 10315 -295 10350 -265
rect 10400 -295 10435 -265
rect 10485 -295 10520 -265
rect 10570 -295 10605 -265
rect 10655 -295 10690 -265
rect 10740 -295 10775 -265
rect 10825 -295 10860 -265
rect 10910 -295 10945 -265
rect 10995 -295 11030 -265
rect 11080 -295 11115 -265
rect 11165 -295 11200 -265
rect 11250 -295 11285 -265
rect 11335 -295 11370 -265
rect 11420 -295 11455 -265
rect 11505 -295 11540 -265
rect 11590 -295 11625 -265
rect 11675 -295 11710 -265
rect 11760 -295 11795 -265
rect 11845 -295 11880 -265
rect 11930 -295 11965 -265
rect 12015 -295 12050 -265
rect 12100 -295 12135 -265
rect 12185 -295 12220 -265
rect 12270 -295 12305 -265
rect 12355 -295 12390 -265
rect 12440 -295 12475 -265
rect 12525 -295 12560 -265
rect 12610 -295 12645 -265
rect 12695 -295 12730 -265
rect 12780 -295 12815 -265
rect 12865 -295 12900 -265
rect 12950 -295 12985 -265
rect 13035 -295 13070 -265
rect 13120 -295 13155 -265
rect 13205 -295 13240 -265
rect 13290 -295 13325 -265
rect 13375 -295 13410 -265
rect 13460 -295 13495 -265
rect 13545 -295 13580 -265
rect 13630 -295 13665 -265
rect 13715 -295 13750 -265
rect 13800 -295 13835 -265
rect 13885 -295 13920 -265
rect 13970 -295 14005 -265
rect 14055 -295 14090 -265
rect 14140 -295 14175 -265
rect 14225 -295 14260 -265
rect 14310 -295 14345 -265
rect 14395 -295 14430 -265
rect 14480 -295 14515 -265
rect 14565 -295 14600 -265
rect 14650 -295 14685 -265
rect 14735 -295 14770 -265
rect 14820 -295 14855 -265
rect 14905 -295 14940 -265
rect 14990 -295 15025 -265
rect 15075 -295 15110 -265
rect 15160 -295 15195 -265
rect 15245 -295 15280 -265
rect 15330 -295 15365 -265
rect 15415 -295 15450 -265
rect 15500 -295 15535 -265
rect 15585 -295 15620 -265
rect 15670 -295 15705 -265
rect 15755 -295 15790 -265
rect 15840 -295 15875 -265
rect 15925 -295 15960 -265
rect 16010 -295 16045 -265
rect 16095 -295 16130 -265
rect 16180 -295 16215 -265
rect 16265 -295 16300 -265
rect 16350 -295 16385 -265
rect 16435 -295 16470 -265
rect 16520 -295 16555 -265
rect 16605 -295 16640 -265
rect 16690 -295 16725 -265
rect 16775 -295 16810 -265
rect 16860 -295 16895 -265
rect 16945 -295 16980 -265
rect 17030 -295 17065 -265
rect 17115 -295 17150 -265
rect 17200 -295 17235 -265
rect 17285 -295 17320 -265
rect 17370 -295 17405 -265
rect 17455 -295 17490 -265
rect 17540 -295 17575 -265
rect 17625 -295 17660 -265
rect 17710 -295 17745 -265
rect 17795 -295 17830 -265
rect 17880 -295 17915 -265
rect 17965 -295 18000 -265
rect 18050 -295 18085 -265
rect 18135 -295 18170 -265
rect 18220 -295 18255 -265
rect 18305 -295 18340 -265
rect 18390 -295 18425 -265
rect 18475 -295 18510 -265
rect 18560 -295 18595 -265
rect 18645 -295 18680 -265
rect 18730 -295 18765 -265
rect 18815 -295 18850 -265
rect 18900 -295 18935 -265
rect 18985 -295 19020 -265
rect 19070 -295 19105 -265
rect 19155 -295 19190 -265
rect 19240 -295 19275 -265
rect 19325 -295 19360 -265
rect 19410 -295 19445 -265
rect 19495 -295 19530 -265
rect 19580 -295 19615 -265
rect 19665 -295 19700 -265
rect 19750 -295 19785 -265
rect 19835 -295 19870 -265
rect 19920 -295 19955 -265
rect 20005 -295 20040 -265
rect 20090 -295 20125 -265
rect 20175 -295 20210 -265
rect 20260 -295 20295 -265
rect 20345 -295 20380 -265
rect 20430 -295 20465 -265
rect 20515 -295 20550 -265
rect 20600 -295 20635 -265
rect 20685 -295 20720 -265
rect 20770 -295 20805 -265
rect 20855 -295 20890 -265
rect 20940 -295 20975 -265
rect 21025 -295 21060 -265
rect 21110 -295 21145 -265
rect 21195 -295 21230 -265
rect 21280 -295 21315 -265
rect 21365 -295 21400 -265
rect 21450 -295 21485 -265
rect 21535 -295 21570 -265
rect 21620 -295 21655 -265
rect 21705 -295 21740 -265
rect 21790 -295 21825 -265
rect 21875 -295 21910 -265
rect 21960 -295 21995 -265
rect 22045 -295 22080 -265
rect 22130 -295 22165 -265
rect 22215 -295 22250 -265
rect 22300 -295 22335 -265
rect 22385 -295 22420 -265
rect 22470 -295 22505 -265
rect 22555 -295 22590 -265
rect 22640 -295 22675 -265
rect 22725 -295 22760 -265
rect 22810 -295 22845 -265
rect 22895 -295 22930 -265
rect 22980 -295 23015 -265
rect 23065 -295 23100 -265
rect 23150 -295 23185 -265
rect 23235 -295 23270 -265
rect 23320 -295 23355 -265
rect 23405 -295 23440 -265
rect 23490 -295 23525 -265
rect 23575 -295 23610 -265
rect 23660 -295 23695 -265
rect 23745 -295 23780 -265
rect 23830 -295 23865 -265
rect 23915 -295 23950 -265
rect 24000 -295 24035 -265
rect 24085 -295 24120 -265
rect 24170 -295 24205 -265
rect 24255 -295 24290 -265
rect 24340 -295 24375 -265
rect 24425 -295 24460 -265
rect 24510 -295 24545 -265
rect 24595 -295 24630 -265
rect 24680 -295 24715 -265
rect 24765 -295 24800 -265
rect 24850 -295 24885 -265
rect 24935 -295 24970 -265
rect 25020 -295 25055 -265
rect 25105 -295 25140 -265
rect 25190 -295 25225 -265
rect 25275 -295 25310 -265
rect 25360 -295 25395 -265
rect 25445 -295 25480 -265
rect 25530 -295 25565 -265
rect 25615 -295 25650 -265
rect 25700 -295 25735 -265
rect 25785 -295 25820 -265
rect 25870 -295 25905 -265
rect 25955 -295 25990 -265
rect 26040 -295 26075 -265
rect 26125 -295 26160 -265
rect 26210 -295 26245 -265
rect 26295 -295 26330 -265
rect 26380 -295 26415 -265
rect 26465 -295 26500 -265
rect 26550 -295 26585 -265
rect 26635 -295 26670 -265
rect 26720 -295 26755 -265
rect 26805 -295 26840 -265
rect 26890 -295 26925 -265
rect 26975 -295 27010 -265
rect 27060 -295 27095 -265
rect 27145 -295 27180 -265
rect 27230 -295 27265 -265
rect 27315 -295 27350 -265
rect 27400 -295 27435 -265
rect 27485 -295 27520 -265
rect 27570 -295 27605 -265
rect 27655 -295 27690 -265
rect 27740 -295 27775 -265
rect 27825 -295 27860 -265
rect 27910 -295 27945 -265
rect 27995 -295 28030 -265
rect 28080 -295 28115 -265
rect 28165 -295 28200 -265
rect 28250 -295 28285 -265
rect 28335 -295 28370 -265
rect 28420 -295 28455 -265
rect 28505 -295 28540 -265
rect 28590 -295 28625 -265
rect 28675 -295 28710 -265
rect 28760 -295 28795 -265
rect 28845 -295 28880 -265
rect 28930 -295 28965 -265
rect 29015 -295 29050 -265
rect 29100 -295 29135 -265
rect 29185 -295 29220 -265
rect 29270 -295 29305 -265
rect 29355 -295 29390 -265
rect 29440 -295 29475 -265
rect 29525 -295 29560 -265
rect 29610 -295 29645 -265
rect 29695 -295 29730 -265
rect 29780 -295 29815 -265
rect 29865 -295 29900 -265
rect 29950 -295 29985 -265
rect 30035 -295 30070 -265
rect 30120 -295 30155 -265
rect 30205 -295 30240 -265
rect 30290 -295 30325 -265
rect 30375 -295 30410 -265
rect 30460 -295 30495 -265
rect 30545 -295 30580 -265
rect 30630 -295 30665 -265
rect 30715 -295 30750 -265
rect 30800 -295 30835 -265
rect 30885 -295 30920 -265
rect 30970 -295 31005 -265
rect 31055 -295 31090 -265
rect 31140 -295 31175 -265
rect 31225 -295 31260 -265
rect 31310 -295 31345 -265
rect 31395 -295 31430 -265
rect 31480 -295 31515 -265
rect 31565 -295 31600 -265
rect 31650 -295 31685 -265
rect 31735 -295 31770 -265
rect 31820 -295 31855 -265
rect 31905 -295 31940 -265
rect 31990 -295 32025 -265
rect 32075 -295 32110 -265
rect 32160 -295 32195 -265
rect 32245 -295 32280 -265
rect 32330 -295 32365 -265
rect 32415 -295 32450 -265
rect 32500 -295 32535 -265
rect 32585 -295 32620 -265
rect 32670 -295 32705 -265
rect 32755 -295 32790 -265
rect 32840 -295 32875 -265
rect 32925 -295 32960 -265
rect 33010 -295 33045 -265
rect 33095 -295 33130 -265
rect 33180 -295 33215 -265
rect 33265 -295 33300 -265
rect 33350 -295 33385 -265
rect 33435 -295 33470 -265
rect 33520 -295 33555 -265
rect 33605 -295 33640 -265
rect 33690 -295 33725 -265
rect 33775 -295 33810 -265
rect 33860 -295 33895 -265
rect 33945 -295 33980 -265
rect 34030 -295 34065 -265
rect 34115 -295 34150 -265
rect 34200 -295 34235 -265
rect 34285 -295 34320 -265
rect 34370 -295 34405 -265
rect 34455 -295 34490 -265
rect 34540 -295 34575 -265
rect 34625 -295 34660 -265
rect 34710 -295 34745 -265
rect 34795 -295 34830 -265
rect 34880 -295 34915 -265
rect 34965 -295 35000 -265
rect 35050 -295 35085 -265
rect 35135 -295 35170 -265
rect 35220 -295 35255 -265
rect 35305 -295 35340 -265
rect 35390 -295 35425 -265
rect 35475 -295 35510 -265
rect 35560 -295 35595 -265
rect 35645 -295 35680 -265
rect 35730 -295 35765 -265
rect 35815 -295 35850 -265
rect 35900 -295 35935 -265
rect 35985 -295 36020 -265
rect 36070 -295 36105 -265
rect 36155 -295 36190 -265
rect 36240 -295 36275 -265
rect 36325 -295 36360 -265
rect 36410 -295 36445 -265
rect 36495 -295 36530 -265
rect 36580 -295 36615 -265
rect 36665 -295 36700 -265
rect 36750 -295 36785 -265
rect 36835 -295 36870 -265
rect 36920 -295 36955 -265
rect 37005 -295 37040 -265
rect 37090 -295 37125 -265
rect 37175 -295 37210 -265
rect 37260 -295 37295 -265
rect 37345 -295 37380 -265
rect 37430 -295 37465 -265
rect 37515 -295 37550 -265
rect 37600 -295 37635 -265
rect 37685 -295 37720 -265
rect 37770 -295 37805 -265
rect 37855 -295 37890 -265
rect 37940 -295 37975 -265
rect 38025 -295 38060 -265
rect 38110 -295 38145 -265
rect 38195 -295 38230 -265
rect 38280 -295 38315 -265
rect 38365 -295 38400 -265
rect 38450 -295 38485 -265
rect 38535 -295 38570 -265
rect 38620 -295 38655 -265
rect 38705 -295 38740 -265
rect 38790 -295 38825 -265
rect 38875 -295 38910 -265
rect 38960 -295 38995 -265
rect 39045 -295 39080 -265
rect 39130 -295 39165 -265
rect 39215 -295 39250 -265
rect 39300 -295 39335 -265
rect 39385 -295 39420 -265
rect 39470 -295 39505 -265
rect 39555 -295 39590 -265
rect 39640 -295 39675 -265
rect 39725 -295 39760 -265
rect 39810 -295 39845 -265
rect 39895 -295 39930 -265
rect 39980 -295 40015 -265
rect 40065 -295 40100 -265
rect 40150 -295 40185 -265
rect 40235 -295 40270 -265
rect 40320 -295 40355 -265
rect 40405 -295 40440 -265
rect 40490 -295 40525 -265
rect 40575 -295 40610 -265
rect 40660 -295 40695 -265
rect 40745 -295 40780 -265
rect 40830 -295 40865 -265
rect 40915 -295 40950 -265
rect 41000 -295 41035 -265
rect 41085 -295 41120 -265
rect 41170 -295 41205 -265
rect 41255 -295 41290 -265
rect 41340 -295 41375 -265
rect 41425 -295 41460 -265
rect 41510 -295 41545 -265
rect 41595 -295 41630 -265
rect 41680 -295 41715 -265
rect 41765 -295 41800 -265
rect 41850 -295 41885 -265
rect 41935 -295 41970 -265
rect 42020 -295 42055 -265
rect 42105 -295 42140 -265
rect 42190 -295 42225 -265
rect 42275 -295 42310 -265
rect 42360 -295 42395 -265
rect 42445 -295 42480 -265
rect 42530 -295 42565 -265
rect 42615 -295 42650 -265
rect 42700 -295 42735 -265
rect 42785 -295 42820 -265
rect 42870 -295 42905 -265
rect 42955 -295 42990 -265
rect 43040 -295 43075 -265
rect 43125 -295 43160 -265
rect 43210 -295 43245 -265
rect 43295 -295 43330 -265
rect 43380 -295 43415 -265
rect 43465 -295 43500 -265
rect 43550 -295 43585 -265
rect 75 -365 105 -335
rect 245 -365 275 -335
rect 415 -365 445 -335
rect 585 -365 615 -335
rect 755 -365 785 -335
rect 925 -365 955 -335
rect 1095 -365 1125 -335
rect 1265 -365 1295 -335
rect 1435 -365 1465 -335
rect 1605 -365 1635 -335
rect 1775 -365 1805 -335
rect 1945 -365 1975 -335
rect 2115 -365 2145 -335
rect 2285 -365 2315 -335
rect 2455 -365 2485 -335
rect 2625 -365 2655 -335
rect 2795 -365 2825 -335
rect 2965 -365 2995 -335
rect 3135 -365 3165 -335
rect 3305 -365 3335 -335
rect 3475 -365 3505 -335
rect 3645 -365 3675 -335
rect 3815 -365 3845 -335
rect 3985 -365 4015 -335
rect 4155 -365 4185 -335
rect 4325 -365 4355 -335
rect 4495 -365 4525 -335
rect 4665 -365 4695 -335
rect 4835 -365 4865 -335
rect 5005 -365 5035 -335
rect 5175 -365 5205 -335
rect 5345 -365 5375 -335
rect 5515 -365 5545 -335
rect 5685 -365 5715 -335
rect 5855 -365 5885 -335
rect 6025 -365 6055 -335
rect 6195 -365 6225 -335
rect 6365 -365 6395 -335
rect 6535 -365 6565 -335
rect 6705 -365 6735 -335
rect 6875 -365 6905 -335
rect 7045 -365 7075 -335
rect 7215 -365 7245 -335
rect 7385 -365 7415 -335
rect 7555 -365 7585 -335
rect 7725 -365 7755 -335
rect 7895 -365 7925 -335
rect 8065 -365 8095 -335
rect 8235 -365 8265 -335
rect 8405 -365 8435 -335
rect 8575 -365 8605 -335
rect 8745 -365 8775 -335
rect 8915 -365 8945 -335
rect 9085 -365 9115 -335
rect 9255 -365 9285 -335
rect 9425 -365 9455 -335
rect 9595 -365 9625 -335
rect 9765 -365 9795 -335
rect 9935 -365 9965 -335
rect 10105 -365 10135 -335
rect 10275 -365 10305 -335
rect 10445 -365 10475 -335
rect 10615 -365 10645 -335
rect 10785 -365 10815 -335
rect 10955 -365 10985 -335
rect 11125 -365 11155 -335
rect 11295 -365 11325 -335
rect 11465 -365 11495 -335
rect 11635 -365 11665 -335
rect 11805 -365 11835 -335
rect 11975 -365 12005 -335
rect 12145 -365 12175 -335
rect 12315 -365 12345 -335
rect 12485 -365 12515 -335
rect 12655 -365 12685 -335
rect 12825 -365 12855 -335
rect 12995 -365 13025 -335
rect 13165 -365 13195 -335
rect 13335 -365 13365 -335
rect 13505 -365 13535 -335
rect 13675 -365 13705 -335
rect 13845 -365 13875 -335
rect 14015 -365 14045 -335
rect 14185 -365 14215 -335
rect 14355 -365 14385 -335
rect 14525 -365 14555 -335
rect 14695 -365 14725 -335
rect 14865 -365 14895 -335
rect 15035 -365 15065 -335
rect 15205 -365 15235 -335
rect 15375 -365 15405 -335
rect 15545 -365 15575 -335
rect 15715 -365 15745 -335
rect 15885 -365 15915 -335
rect 16055 -365 16085 -335
rect 16225 -365 16255 -335
rect 16395 -365 16425 -335
rect 16565 -365 16595 -335
rect 16735 -365 16765 -335
rect 16905 -365 16935 -335
rect 17075 -365 17105 -335
rect 17245 -365 17275 -335
rect 17415 -365 17445 -335
rect 17585 -365 17615 -335
rect 17755 -365 17785 -335
rect 17925 -365 17955 -335
rect 18095 -365 18125 -335
rect 18265 -365 18295 -335
rect 18435 -365 18465 -335
rect 18605 -365 18635 -335
rect 18775 -365 18805 -335
rect 18945 -365 18975 -335
rect 19115 -365 19145 -335
rect 19285 -365 19315 -335
rect 19455 -365 19485 -335
rect 19625 -365 19655 -335
rect 19795 -365 19825 -335
rect 19965 -365 19995 -335
rect 20135 -365 20165 -335
rect 20305 -365 20335 -335
rect 20475 -365 20505 -335
rect 20645 -365 20675 -335
rect 20815 -365 20845 -335
rect 20985 -365 21015 -335
rect 21155 -365 21185 -335
rect 21325 -365 21355 -335
rect 21495 -365 21525 -335
rect 21665 -365 21695 -335
rect 21835 -365 21865 -335
rect 22005 -365 22035 -335
rect 22175 -365 22205 -335
rect 22345 -365 22375 -335
rect 22515 -365 22545 -335
rect 22685 -365 22715 -335
rect 22855 -365 22885 -335
rect 23025 -365 23055 -335
rect 23195 -365 23225 -335
rect 23365 -365 23395 -335
rect 23535 -365 23565 -335
rect 23705 -365 23735 -335
rect 23875 -365 23905 -335
rect 24045 -365 24075 -335
rect 24215 -365 24245 -335
rect 24385 -365 24415 -335
rect 24555 -365 24585 -335
rect 24725 -365 24755 -335
rect 24895 -365 24925 -335
rect 25065 -365 25095 -335
rect 25235 -365 25265 -335
rect 25405 -365 25435 -335
rect 25575 -365 25605 -335
rect 25745 -365 25775 -335
rect 25915 -365 25945 -335
rect 26085 -365 26115 -335
rect 26255 -365 26285 -335
rect 26425 -365 26455 -335
rect 26595 -365 26625 -335
rect 26765 -365 26795 -335
rect 26935 -365 26965 -335
rect 27105 -365 27135 -335
rect 27275 -365 27305 -335
rect 27445 -365 27475 -335
rect 27615 -365 27645 -335
rect 27785 -365 27815 -335
rect 27955 -365 27985 -335
rect 28125 -365 28155 -335
rect 28295 -365 28325 -335
rect 28465 -365 28495 -335
rect 28635 -365 28665 -335
rect 28805 -365 28835 -335
rect 28975 -365 29005 -335
rect 29145 -365 29175 -335
rect 29315 -365 29345 -335
rect 29485 -365 29515 -335
rect 29655 -365 29685 -335
rect 29825 -365 29855 -335
rect 29995 -365 30025 -335
rect 30165 -365 30195 -335
rect 30335 -365 30365 -335
rect 30505 -365 30535 -335
rect 30675 -365 30705 -335
rect 30845 -365 30875 -335
rect 31015 -365 31045 -335
rect 31185 -365 31215 -335
rect 31355 -365 31385 -335
rect 31525 -365 31555 -335
rect 31695 -365 31725 -335
rect 31865 -365 31895 -335
rect 32035 -365 32065 -335
rect 32205 -365 32235 -335
rect 32375 -365 32405 -335
rect 32545 -365 32575 -335
rect 32715 -365 32745 -335
rect 32885 -365 32915 -335
rect 33055 -365 33085 -335
rect 33225 -365 33255 -335
rect 33395 -365 33425 -335
rect 33565 -365 33595 -335
rect 33735 -365 33765 -335
rect 33905 -365 33935 -335
rect 34075 -365 34105 -335
rect 34245 -365 34275 -335
rect 34415 -365 34445 -335
rect 34585 -365 34615 -335
rect 34755 -365 34785 -335
rect 34925 -365 34955 -335
rect 35095 -365 35125 -335
rect 35265 -365 35295 -335
rect 35435 -365 35465 -335
rect 35605 -365 35635 -335
rect 35775 -365 35805 -335
rect 35945 -365 35975 -335
rect 36115 -365 36145 -335
rect 36285 -365 36315 -335
rect 36455 -365 36485 -335
rect 36625 -365 36655 -335
rect 36795 -365 36825 -335
rect 36965 -365 36995 -335
rect 37135 -365 37165 -335
rect 37305 -365 37335 -335
rect 37475 -365 37505 -335
rect 37645 -365 37675 -335
rect 37815 -365 37845 -335
rect 37985 -365 38015 -335
rect 38155 -365 38185 -335
rect 38325 -365 38355 -335
rect 38495 -365 38525 -335
rect 38665 -365 38695 -335
rect 38835 -365 38865 -335
rect 39005 -365 39035 -335
rect 39175 -365 39205 -335
rect 39345 -365 39375 -335
rect 39515 -365 39545 -335
rect 39685 -365 39715 -335
rect 39855 -365 39885 -335
rect 40025 -365 40055 -335
rect 40195 -365 40225 -335
rect 40365 -365 40395 -335
rect 40535 -365 40565 -335
rect 40705 -365 40735 -335
rect 40875 -365 40905 -335
rect 41045 -365 41075 -335
rect 41215 -365 41245 -335
rect 41385 -365 41415 -335
rect 41555 -365 41585 -335
rect 41725 -365 41755 -335
rect 41895 -365 41925 -335
rect 42065 -365 42095 -335
rect 42235 -365 42265 -335
rect 42405 -365 42435 -335
rect 42575 -365 42605 -335
rect 42745 -365 42775 -335
rect 42915 -365 42945 -335
rect 43085 -365 43115 -335
rect 43255 -365 43285 -335
rect 43425 -365 43455 -335
rect 43595 -365 43625 -335
rect 160 -475 190 -440
rect 75 -580 105 -550
rect 330 -475 360 -440
rect 245 -580 275 -550
rect 500 -475 530 -440
rect 415 -580 445 -550
rect 670 -475 700 -440
rect 585 -580 615 -550
rect 840 -475 870 -440
rect 755 -580 785 -550
rect 1010 -475 1040 -440
rect 925 -580 955 -550
rect 1180 -475 1210 -440
rect 1095 -580 1125 -550
rect 1350 -475 1380 -440
rect 1265 -580 1295 -550
rect 1520 -475 1550 -440
rect 1435 -580 1465 -550
rect 1690 -475 1720 -440
rect 1605 -580 1635 -550
rect 1860 -475 1890 -440
rect 1775 -580 1805 -550
rect 2030 -475 2060 -440
rect 1945 -580 1975 -550
rect 2200 -475 2230 -440
rect 2115 -580 2145 -550
rect 2370 -475 2400 -440
rect 2285 -580 2315 -550
rect 2540 -475 2570 -440
rect 2455 -580 2485 -550
rect 2710 -475 2740 -440
rect 2625 -580 2655 -550
rect 2880 -475 2910 -440
rect 2795 -580 2825 -550
rect 3050 -475 3080 -440
rect 2965 -580 2995 -550
rect 3220 -475 3250 -440
rect 3135 -580 3165 -550
rect 3390 -475 3420 -440
rect 3305 -580 3335 -550
rect 3560 -475 3590 -440
rect 3475 -580 3505 -550
rect 3730 -475 3760 -440
rect 3645 -580 3675 -550
rect 3900 -475 3930 -440
rect 3815 -580 3845 -550
rect 4070 -475 4100 -440
rect 3985 -580 4015 -550
rect 4240 -475 4270 -440
rect 4155 -580 4185 -550
rect 4410 -475 4440 -440
rect 4325 -580 4355 -550
rect 4580 -475 4610 -440
rect 4495 -580 4525 -550
rect 4750 -475 4780 -440
rect 4665 -580 4695 -550
rect 4920 -475 4950 -440
rect 4835 -580 4865 -550
rect 5090 -475 5120 -440
rect 5005 -580 5035 -550
rect 5260 -475 5290 -440
rect 5175 -580 5205 -550
rect 5430 -475 5460 -440
rect 5345 -580 5375 -550
rect 5600 -475 5630 -440
rect 5515 -580 5545 -550
rect 5770 -475 5800 -440
rect 5685 -580 5715 -550
rect 5940 -475 5970 -440
rect 5855 -580 5885 -550
rect 6110 -475 6140 -440
rect 6025 -580 6055 -550
rect 6280 -475 6310 -440
rect 6195 -580 6225 -550
rect 6450 -475 6480 -440
rect 6365 -580 6395 -550
rect 6620 -475 6650 -440
rect 6535 -580 6565 -550
rect 6790 -475 6820 -440
rect 6705 -580 6735 -550
rect 6960 -475 6990 -440
rect 6875 -580 6905 -550
rect 7130 -475 7160 -440
rect 7045 -580 7075 -550
rect 7300 -475 7330 -440
rect 7215 -580 7245 -550
rect 7470 -475 7500 -440
rect 7385 -580 7415 -550
rect 7640 -475 7670 -440
rect 7555 -580 7585 -550
rect 7810 -475 7840 -440
rect 7725 -580 7755 -550
rect 7980 -475 8010 -440
rect 7895 -580 7925 -550
rect 8150 -475 8180 -440
rect 8065 -580 8095 -550
rect 8320 -475 8350 -440
rect 8235 -580 8265 -550
rect 8490 -475 8520 -440
rect 8405 -580 8435 -550
rect 8660 -475 8690 -440
rect 8575 -580 8605 -550
rect 8830 -475 8860 -440
rect 8745 -580 8775 -550
rect 9000 -475 9030 -440
rect 8915 -580 8945 -550
rect 9170 -475 9200 -440
rect 9085 -580 9115 -550
rect 9340 -475 9370 -440
rect 9255 -580 9285 -550
rect 9510 -475 9540 -440
rect 9425 -580 9455 -550
rect 9680 -475 9710 -440
rect 9595 -580 9625 -550
rect 9850 -475 9880 -440
rect 9765 -580 9795 -550
rect 10020 -475 10050 -440
rect 9935 -580 9965 -550
rect 10190 -475 10220 -440
rect 10105 -580 10135 -550
rect 10360 -475 10390 -440
rect 10275 -580 10305 -550
rect 10530 -475 10560 -440
rect 10445 -580 10475 -550
rect 10700 -475 10730 -440
rect 10615 -580 10645 -550
rect 10870 -475 10900 -440
rect 10785 -580 10815 -550
rect 11040 -475 11070 -440
rect 10955 -580 10985 -550
rect 11210 -475 11240 -440
rect 11125 -580 11155 -550
rect 11380 -475 11410 -440
rect 11295 -580 11325 -550
rect 11550 -475 11580 -440
rect 11465 -580 11495 -550
rect 11720 -475 11750 -440
rect 11635 -580 11665 -550
rect 11890 -475 11920 -440
rect 11805 -580 11835 -550
rect 12060 -475 12090 -440
rect 11975 -580 12005 -550
rect 12230 -475 12260 -440
rect 12145 -580 12175 -550
rect 12400 -475 12430 -440
rect 12315 -580 12345 -550
rect 12570 -475 12600 -440
rect 12485 -580 12515 -550
rect 12740 -475 12770 -440
rect 12655 -580 12685 -550
rect 12910 -475 12940 -440
rect 12825 -580 12855 -550
rect 13080 -475 13110 -440
rect 12995 -580 13025 -550
rect 13250 -475 13280 -440
rect 13165 -580 13195 -550
rect 13420 -475 13450 -440
rect 13335 -580 13365 -550
rect 13590 -475 13620 -440
rect 13505 -580 13535 -550
rect 13760 -475 13790 -440
rect 13675 -580 13705 -550
rect 13930 -475 13960 -440
rect 13845 -580 13875 -550
rect 14100 -475 14130 -440
rect 14015 -580 14045 -550
rect 14270 -475 14300 -440
rect 14185 -580 14215 -550
rect 14440 -475 14470 -440
rect 14355 -580 14385 -550
rect 14610 -475 14640 -440
rect 14525 -580 14555 -550
rect 14780 -475 14810 -440
rect 14695 -580 14725 -550
rect 14950 -475 14980 -440
rect 14865 -580 14895 -550
rect 15120 -475 15150 -440
rect 15035 -580 15065 -550
rect 15290 -475 15320 -440
rect 15205 -580 15235 -550
rect 15460 -475 15490 -440
rect 15375 -580 15405 -550
rect 15630 -475 15660 -440
rect 15545 -580 15575 -550
rect 15800 -475 15830 -440
rect 15715 -580 15745 -550
rect 15970 -475 16000 -440
rect 15885 -580 15915 -550
rect 16140 -475 16170 -440
rect 16055 -580 16085 -550
rect 16310 -475 16340 -440
rect 16225 -580 16255 -550
rect 16480 -475 16510 -440
rect 16395 -580 16425 -550
rect 16650 -475 16680 -440
rect 16565 -580 16595 -550
rect 16820 -475 16850 -440
rect 16735 -580 16765 -550
rect 16990 -475 17020 -440
rect 16905 -580 16935 -550
rect 17160 -475 17190 -440
rect 17075 -580 17105 -550
rect 17330 -475 17360 -440
rect 17245 -580 17275 -550
rect 17500 -475 17530 -440
rect 17415 -580 17445 -550
rect 17670 -475 17700 -440
rect 17585 -580 17615 -550
rect 17840 -475 17870 -440
rect 17755 -580 17785 -550
rect 18010 -475 18040 -440
rect 17925 -580 17955 -550
rect 18180 -475 18210 -440
rect 18095 -580 18125 -550
rect 18350 -475 18380 -440
rect 18265 -580 18295 -550
rect 18520 -475 18550 -440
rect 18435 -580 18465 -550
rect 18690 -475 18720 -440
rect 18605 -580 18635 -550
rect 18860 -475 18890 -440
rect 18775 -580 18805 -550
rect 19030 -475 19060 -440
rect 18945 -580 18975 -550
rect 19200 -475 19230 -440
rect 19115 -580 19145 -550
rect 19370 -475 19400 -440
rect 19285 -580 19315 -550
rect 19540 -475 19570 -440
rect 19455 -580 19485 -550
rect 19710 -475 19740 -440
rect 19625 -580 19655 -550
rect 19880 -475 19910 -440
rect 19795 -580 19825 -550
rect 20050 -475 20080 -440
rect 19965 -580 19995 -550
rect 20220 -475 20250 -440
rect 20135 -580 20165 -550
rect 20390 -475 20420 -440
rect 20305 -580 20335 -550
rect 20560 -475 20590 -440
rect 20475 -580 20505 -550
rect 20730 -475 20760 -440
rect 20645 -580 20675 -550
rect 20900 -475 20930 -440
rect 20815 -580 20845 -550
rect 21070 -475 21100 -440
rect 20985 -580 21015 -550
rect 21240 -475 21270 -440
rect 21155 -580 21185 -550
rect 21410 -475 21440 -440
rect 21325 -580 21355 -550
rect 21580 -475 21610 -440
rect 21495 -580 21525 -550
rect 21750 -475 21780 -440
rect 21665 -580 21695 -550
rect 21920 -475 21950 -440
rect 21835 -580 21865 -550
rect 22090 -475 22120 -440
rect 22005 -580 22035 -550
rect 22260 -475 22290 -440
rect 22175 -580 22205 -550
rect 22430 -475 22460 -440
rect 22345 -580 22375 -550
rect 22600 -475 22630 -440
rect 22515 -580 22545 -550
rect 22770 -475 22800 -440
rect 22685 -580 22715 -550
rect 22940 -475 22970 -440
rect 22855 -580 22885 -550
rect 23110 -475 23140 -440
rect 23025 -580 23055 -550
rect 23280 -475 23310 -440
rect 23195 -580 23225 -550
rect 23450 -475 23480 -440
rect 23365 -580 23395 -550
rect 23620 -475 23650 -440
rect 23535 -580 23565 -550
rect 23790 -475 23820 -440
rect 23705 -580 23735 -550
rect 23960 -475 23990 -440
rect 23875 -580 23905 -550
rect 24130 -475 24160 -440
rect 24045 -580 24075 -550
rect 24300 -475 24330 -440
rect 24215 -580 24245 -550
rect 24470 -475 24500 -440
rect 24385 -580 24415 -550
rect 24640 -475 24670 -440
rect 24555 -580 24585 -550
rect 24810 -475 24840 -440
rect 24725 -580 24755 -550
rect 24980 -475 25010 -440
rect 24895 -580 24925 -550
rect 25150 -475 25180 -440
rect 25065 -580 25095 -550
rect 25320 -475 25350 -440
rect 25235 -580 25265 -550
rect 25490 -475 25520 -440
rect 25405 -580 25435 -550
rect 25660 -475 25690 -440
rect 25575 -580 25605 -550
rect 25830 -475 25860 -440
rect 25745 -580 25775 -550
rect 26000 -475 26030 -440
rect 25915 -580 25945 -550
rect 26170 -475 26200 -440
rect 26085 -580 26115 -550
rect 26340 -475 26370 -440
rect 26255 -580 26285 -550
rect 26510 -475 26540 -440
rect 26425 -580 26455 -550
rect 26680 -475 26710 -440
rect 26595 -580 26625 -550
rect 26850 -475 26880 -440
rect 26765 -580 26795 -550
rect 27020 -475 27050 -440
rect 26935 -580 26965 -550
rect 27190 -475 27220 -440
rect 27105 -580 27135 -550
rect 27360 -475 27390 -440
rect 27275 -580 27305 -550
rect 27530 -475 27560 -440
rect 27445 -580 27475 -550
rect 27700 -475 27730 -440
rect 27615 -580 27645 -550
rect 27870 -475 27900 -440
rect 27785 -580 27815 -550
rect 28040 -475 28070 -440
rect 27955 -580 27985 -550
rect 28210 -475 28240 -440
rect 28125 -580 28155 -550
rect 28380 -475 28410 -440
rect 28295 -580 28325 -550
rect 28550 -475 28580 -440
rect 28465 -580 28495 -550
rect 28720 -475 28750 -440
rect 28635 -580 28665 -550
rect 28890 -475 28920 -440
rect 28805 -580 28835 -550
rect 29060 -475 29090 -440
rect 28975 -580 29005 -550
rect 29230 -475 29260 -440
rect 29145 -580 29175 -550
rect 29400 -475 29430 -440
rect 29315 -580 29345 -550
rect 29570 -475 29600 -440
rect 29485 -580 29515 -550
rect 29740 -475 29770 -440
rect 29655 -580 29685 -550
rect 29910 -475 29940 -440
rect 29825 -580 29855 -550
rect 30080 -475 30110 -440
rect 29995 -580 30025 -550
rect 30250 -475 30280 -440
rect 30165 -580 30195 -550
rect 30420 -475 30450 -440
rect 30335 -580 30365 -550
rect 30590 -475 30620 -440
rect 30505 -580 30535 -550
rect 30760 -475 30790 -440
rect 30675 -580 30705 -550
rect 30930 -475 30960 -440
rect 30845 -580 30875 -550
rect 31100 -475 31130 -440
rect 31015 -580 31045 -550
rect 31270 -475 31300 -440
rect 31185 -580 31215 -550
rect 31440 -475 31470 -440
rect 31355 -580 31385 -550
rect 31610 -475 31640 -440
rect 31525 -580 31555 -550
rect 31780 -475 31810 -440
rect 31695 -580 31725 -550
rect 31950 -475 31980 -440
rect 31865 -580 31895 -550
rect 32120 -475 32150 -440
rect 32035 -580 32065 -550
rect 32290 -475 32320 -440
rect 32205 -580 32235 -550
rect 32460 -475 32490 -440
rect 32375 -580 32405 -550
rect 32630 -475 32660 -440
rect 32545 -580 32575 -550
rect 32800 -475 32830 -440
rect 32715 -580 32745 -550
rect 32970 -475 33000 -440
rect 32885 -580 32915 -550
rect 33140 -475 33170 -440
rect 33055 -580 33085 -550
rect 33310 -475 33340 -440
rect 33225 -580 33255 -550
rect 33480 -475 33510 -440
rect 33395 -580 33425 -550
rect 33650 -475 33680 -440
rect 33565 -580 33595 -550
rect 33820 -475 33850 -440
rect 33735 -580 33765 -550
rect 33990 -475 34020 -440
rect 33905 -580 33935 -550
rect 34160 -475 34190 -440
rect 34075 -580 34105 -550
rect 34330 -475 34360 -440
rect 34245 -580 34275 -550
rect 34500 -475 34530 -440
rect 34415 -580 34445 -550
rect 34670 -475 34700 -440
rect 34585 -580 34615 -550
rect 34840 -475 34870 -440
rect 34755 -580 34785 -550
rect 35010 -475 35040 -440
rect 34925 -580 34955 -550
rect 35180 -475 35210 -440
rect 35095 -580 35125 -550
rect 35350 -475 35380 -440
rect 35265 -580 35295 -550
rect 35520 -475 35550 -440
rect 35435 -580 35465 -550
rect 35690 -475 35720 -440
rect 35605 -580 35635 -550
rect 35860 -475 35890 -440
rect 35775 -580 35805 -550
rect 36030 -475 36060 -440
rect 35945 -580 35975 -550
rect 36200 -475 36230 -440
rect 36115 -580 36145 -550
rect 36370 -475 36400 -440
rect 36285 -580 36315 -550
rect 36540 -475 36570 -440
rect 36455 -580 36485 -550
rect 36710 -475 36740 -440
rect 36625 -580 36655 -550
rect 36880 -475 36910 -440
rect 36795 -580 36825 -550
rect 37050 -475 37080 -440
rect 36965 -580 36995 -550
rect 37220 -475 37250 -440
rect 37135 -580 37165 -550
rect 37390 -475 37420 -440
rect 37305 -580 37335 -550
rect 37560 -475 37590 -440
rect 37475 -580 37505 -550
rect 37730 -475 37760 -440
rect 37645 -580 37675 -550
rect 37900 -475 37930 -440
rect 37815 -580 37845 -550
rect 38070 -475 38100 -440
rect 37985 -580 38015 -550
rect 38240 -475 38270 -440
rect 38155 -580 38185 -550
rect 38410 -475 38440 -440
rect 38325 -580 38355 -550
rect 38580 -475 38610 -440
rect 38495 -580 38525 -550
rect 38750 -475 38780 -440
rect 38665 -580 38695 -550
rect 38920 -475 38950 -440
rect 38835 -580 38865 -550
rect 39090 -475 39120 -440
rect 39005 -580 39035 -550
rect 39260 -475 39290 -440
rect 39175 -580 39205 -550
rect 39430 -475 39460 -440
rect 39345 -580 39375 -550
rect 39600 -475 39630 -440
rect 39515 -580 39545 -550
rect 39770 -475 39800 -440
rect 39685 -580 39715 -550
rect 39940 -475 39970 -440
rect 39855 -580 39885 -550
rect 40110 -475 40140 -440
rect 40025 -580 40055 -550
rect 40280 -475 40310 -440
rect 40195 -580 40225 -550
rect 40450 -475 40480 -440
rect 40365 -580 40395 -550
rect 40620 -475 40650 -440
rect 40535 -580 40565 -550
rect 40790 -475 40820 -440
rect 40705 -580 40735 -550
rect 40960 -475 40990 -440
rect 40875 -580 40905 -550
rect 41130 -475 41160 -440
rect 41045 -580 41075 -550
rect 41300 -475 41330 -440
rect 41215 -580 41245 -550
rect 41470 -475 41500 -440
rect 41385 -580 41415 -550
rect 41640 -475 41670 -440
rect 41555 -580 41585 -550
rect 41810 -475 41840 -440
rect 41725 -580 41755 -550
rect 41980 -475 42010 -440
rect 41895 -580 41925 -550
rect 42150 -475 42180 -440
rect 42065 -580 42095 -550
rect 42320 -475 42350 -440
rect 42235 -580 42265 -550
rect 42490 -475 42520 -440
rect 42405 -580 42435 -550
rect 42660 -475 42690 -440
rect 42575 -580 42605 -550
rect 42830 -475 42860 -440
rect 42745 -580 42775 -550
rect 43000 -475 43030 -440
rect 42915 -580 42945 -550
rect 43170 -475 43200 -440
rect 43085 -580 43115 -550
rect 43340 -475 43370 -440
rect 43255 -580 43285 -550
rect 43510 -475 43540 -440
rect 43425 -580 43455 -550
rect 43595 -580 43625 -550
rect 75 -680 105 -650
rect 245 -680 275 -650
rect 415 -680 445 -650
rect 585 -680 615 -650
rect 755 -680 785 -650
rect 925 -680 955 -650
rect 1095 -680 1125 -650
rect 1265 -680 1295 -650
rect 1435 -680 1465 -650
rect 1605 -680 1635 -650
rect 1775 -680 1805 -650
rect 1945 -680 1975 -650
rect 2115 -680 2145 -650
rect 2285 -680 2315 -650
rect 2455 -680 2485 -650
rect 2625 -680 2655 -650
rect 2795 -680 2825 -650
rect 2965 -680 2995 -650
rect 3135 -680 3165 -650
rect 3305 -680 3335 -650
rect 3475 -680 3505 -650
rect 3645 -680 3675 -650
rect 3815 -680 3845 -650
rect 3985 -680 4015 -650
rect 4155 -680 4185 -650
rect 4325 -680 4355 -650
rect 4495 -680 4525 -650
rect 4665 -680 4695 -650
rect 4835 -680 4865 -650
rect 5005 -680 5035 -650
rect 5175 -680 5205 -650
rect 5345 -680 5375 -650
rect 5515 -680 5545 -650
rect 5685 -680 5715 -650
rect 5855 -680 5885 -650
rect 6025 -680 6055 -650
rect 6195 -680 6225 -650
rect 6365 -680 6395 -650
rect 6535 -680 6565 -650
rect 6705 -680 6735 -650
rect 6875 -680 6905 -650
rect 7045 -680 7075 -650
rect 7215 -680 7245 -650
rect 7385 -680 7415 -650
rect 7555 -680 7585 -650
rect 7725 -680 7755 -650
rect 7895 -680 7925 -650
rect 8065 -680 8095 -650
rect 8235 -680 8265 -650
rect 8405 -680 8435 -650
rect 8575 -680 8605 -650
rect 8745 -680 8775 -650
rect 8915 -680 8945 -650
rect 9085 -680 9115 -650
rect 9255 -680 9285 -650
rect 9425 -680 9455 -650
rect 9595 -680 9625 -650
rect 9765 -680 9795 -650
rect 9935 -680 9965 -650
rect 10105 -680 10135 -650
rect 10275 -680 10305 -650
rect 10445 -680 10475 -650
rect 10615 -680 10645 -650
rect 10785 -680 10815 -650
rect 10955 -680 10985 -650
rect 11125 -680 11155 -650
rect 11295 -680 11325 -650
rect 11465 -680 11495 -650
rect 11635 -680 11665 -650
rect 11805 -680 11835 -650
rect 11975 -680 12005 -650
rect 12145 -680 12175 -650
rect 12315 -680 12345 -650
rect 12485 -680 12515 -650
rect 12655 -680 12685 -650
rect 12825 -680 12855 -650
rect 12995 -680 13025 -650
rect 13165 -680 13195 -650
rect 13335 -680 13365 -650
rect 13505 -680 13535 -650
rect 13675 -680 13705 -650
rect 13845 -680 13875 -650
rect 14015 -680 14045 -650
rect 14185 -680 14215 -650
rect 14355 -680 14385 -650
rect 14525 -680 14555 -650
rect 14695 -680 14725 -650
rect 14865 -680 14895 -650
rect 15035 -680 15065 -650
rect 15205 -680 15235 -650
rect 15375 -680 15405 -650
rect 15545 -680 15575 -650
rect 15715 -680 15745 -650
rect 15885 -680 15915 -650
rect 16055 -680 16085 -650
rect 16225 -680 16255 -650
rect 16395 -680 16425 -650
rect 16565 -680 16595 -650
rect 16735 -680 16765 -650
rect 16905 -680 16935 -650
rect 17075 -680 17105 -650
rect 17245 -680 17275 -650
rect 17415 -680 17445 -650
rect 17585 -680 17615 -650
rect 17755 -680 17785 -650
rect 17925 -680 17955 -650
rect 18095 -680 18125 -650
rect 18265 -680 18295 -650
rect 18435 -680 18465 -650
rect 18605 -680 18635 -650
rect 18775 -680 18805 -650
rect 18945 -680 18975 -650
rect 19115 -680 19145 -650
rect 19285 -680 19315 -650
rect 19455 -680 19485 -650
rect 19625 -680 19655 -650
rect 19795 -680 19825 -650
rect 19965 -680 19995 -650
rect 20135 -680 20165 -650
rect 20305 -680 20335 -650
rect 20475 -680 20505 -650
rect 20645 -680 20675 -650
rect 20815 -680 20845 -650
rect 20985 -680 21015 -650
rect 21155 -680 21185 -650
rect 21325 -680 21355 -650
rect 21495 -680 21525 -650
rect 21665 -680 21695 -650
rect 21835 -680 21865 -650
rect 22005 -680 22035 -650
rect 22175 -680 22205 -650
rect 22345 -680 22375 -650
rect 22515 -680 22545 -650
rect 22685 -680 22715 -650
rect 22855 -680 22885 -650
rect 23025 -680 23055 -650
rect 23195 -680 23225 -650
rect 23365 -680 23395 -650
rect 23535 -680 23565 -650
rect 23705 -680 23735 -650
rect 23875 -680 23905 -650
rect 24045 -680 24075 -650
rect 24215 -680 24245 -650
rect 24385 -680 24415 -650
rect 24555 -680 24585 -650
rect 24725 -680 24755 -650
rect 24895 -680 24925 -650
rect 25065 -680 25095 -650
rect 25235 -680 25265 -650
rect 25405 -680 25435 -650
rect 25575 -680 25605 -650
rect 25745 -680 25775 -650
rect 25915 -680 25945 -650
rect 26085 -680 26115 -650
rect 26255 -680 26285 -650
rect 26425 -680 26455 -650
rect 26595 -680 26625 -650
rect 26765 -680 26795 -650
rect 26935 -680 26965 -650
rect 27105 -680 27135 -650
rect 27275 -680 27305 -650
rect 27445 -680 27475 -650
rect 27615 -680 27645 -650
rect 27785 -680 27815 -650
rect 27955 -680 27985 -650
rect 28125 -680 28155 -650
rect 28295 -680 28325 -650
rect 28465 -680 28495 -650
rect 28635 -680 28665 -650
rect 28805 -680 28835 -650
rect 28975 -680 29005 -650
rect 29145 -680 29175 -650
rect 29315 -680 29345 -650
rect 29485 -680 29515 -650
rect 29655 -680 29685 -650
rect 29825 -680 29855 -650
rect 29995 -680 30025 -650
rect 30165 -680 30195 -650
rect 30335 -680 30365 -650
rect 30505 -680 30535 -650
rect 30675 -680 30705 -650
rect 30845 -680 30875 -650
rect 31015 -680 31045 -650
rect 31185 -680 31215 -650
rect 31355 -680 31385 -650
rect 31525 -680 31555 -650
rect 31695 -680 31725 -650
rect 31865 -680 31895 -650
rect 32035 -680 32065 -650
rect 32205 -680 32235 -650
rect 32375 -680 32405 -650
rect 32545 -680 32575 -650
rect 32715 -680 32745 -650
rect 32885 -680 32915 -650
rect 33055 -680 33085 -650
rect 33225 -680 33255 -650
rect 33395 -680 33425 -650
rect 33565 -680 33595 -650
rect 33735 -680 33765 -650
rect 33905 -680 33935 -650
rect 34075 -680 34105 -650
rect 34245 -680 34275 -650
rect 34415 -680 34445 -650
rect 34585 -680 34615 -650
rect 34755 -680 34785 -650
rect 34925 -680 34955 -650
rect 35095 -680 35125 -650
rect 35265 -680 35295 -650
rect 35435 -680 35465 -650
rect 35605 -680 35635 -650
rect 35775 -680 35805 -650
rect 35945 -680 35975 -650
rect 36115 -680 36145 -650
rect 36285 -680 36315 -650
rect 36455 -680 36485 -650
rect 36625 -680 36655 -650
rect 36795 -680 36825 -650
rect 36965 -680 36995 -650
rect 37135 -680 37165 -650
rect 37305 -680 37335 -650
rect 37475 -680 37505 -650
rect 37645 -680 37675 -650
rect 37815 -680 37845 -650
rect 37985 -680 38015 -650
rect 38155 -680 38185 -650
rect 38325 -680 38355 -650
rect 38495 -680 38525 -650
rect 38665 -680 38695 -650
rect 38835 -680 38865 -650
rect 39005 -680 39035 -650
rect 39175 -680 39205 -650
rect 39345 -680 39375 -650
rect 39515 -680 39545 -650
rect 39685 -680 39715 -650
rect 39855 -680 39885 -650
rect 40025 -680 40055 -650
rect 40195 -680 40225 -650
rect 40365 -680 40395 -650
rect 40535 -680 40565 -650
rect 40705 -680 40735 -650
rect 40875 -680 40905 -650
rect 41045 -680 41075 -650
rect 41215 -680 41245 -650
rect 41385 -680 41415 -650
rect 41555 -680 41585 -650
rect 41725 -680 41755 -650
rect 41895 -680 41925 -650
rect 42065 -680 42095 -650
rect 42235 -680 42265 -650
rect 42405 -680 42435 -650
rect 42575 -680 42605 -650
rect 42745 -680 42775 -650
rect 42915 -680 42945 -650
rect 43085 -680 43115 -650
rect 43255 -680 43285 -650
rect 43425 -680 43455 -650
rect 43595 -680 43625 -650
<< metal2 >>
rect 215 205 265 215
rect 385 205 435 215
rect 555 205 605 215
rect 750 205 800 215
rect 920 205 970 215
rect 1090 205 1140 215
rect 1260 205 1310 215
rect 1430 205 1480 215
rect 1600 205 1650 215
rect 1770 205 1820 215
rect 1940 205 1990 215
rect 2110 205 2160 215
rect 2260 205 2310 215
rect 2430 205 2480 215
rect 2600 205 2650 215
rect 2770 205 2820 215
rect 2940 205 2990 215
rect 3110 205 3160 215
rect 3280 205 3330 215
rect 3450 205 3500 215
rect 3620 205 3670 215
rect 3790 205 3840 215
rect 3960 205 4010 215
rect 4130 205 4180 215
rect 4300 205 4350 215
rect 4470 205 4520 215
rect 4640 205 4690 215
rect 4810 205 4860 215
rect 4980 205 5030 215
rect 5150 205 5200 215
rect 5320 205 5370 215
rect 5490 205 5540 215
rect 5660 205 5710 215
rect 5830 205 5880 215
rect 6000 205 6050 215
rect 6170 205 6220 215
rect 6340 205 6390 215
rect 6510 205 6560 215
rect 6680 205 6730 215
rect 6850 205 6900 215
rect 7020 205 7070 215
rect 7190 205 7240 215
rect 7360 205 7410 215
rect 7530 205 7580 215
rect 7700 205 7750 215
rect 7850 205 7900 215
rect 8020 205 8070 215
rect 8190 205 8240 215
rect 8360 205 8410 215
rect 8530 205 8580 215
rect 8700 205 8750 215
rect 8870 205 8920 215
rect 9040 205 9090 215
rect 9210 205 9260 215
rect 9380 205 9430 215
rect 9550 205 9600 215
rect 9720 205 9770 215
rect 9890 205 9940 215
rect 10060 205 10110 215
rect 10230 205 10280 215
rect 10400 205 10450 215
rect 10570 205 10620 215
rect 10740 205 10790 215
rect 10910 205 10960 215
rect 11080 205 11130 215
rect 11250 205 11300 215
rect 11420 205 11470 215
rect 11590 205 11640 215
rect 11760 205 11810 215
rect 11930 205 11980 215
rect 12100 205 12150 215
rect 12270 205 12320 215
rect 12440 205 12490 215
rect 12610 205 12660 215
rect 12780 205 12830 215
rect 12950 205 13000 215
rect 13120 205 13170 215
rect 13290 205 13340 215
rect 13460 205 13510 215
rect 13630 205 13680 215
rect 13800 205 13850 215
rect 13970 205 14020 215
rect 14140 205 14190 215
rect 14310 205 14360 215
rect 14480 205 14530 215
rect 14650 205 14700 215
rect 14820 205 14870 215
rect 14990 205 15040 215
rect 15160 205 15210 215
rect 15330 205 15380 215
rect 15500 205 15550 215
rect 15670 205 15720 215
rect 15840 205 15890 215
rect 16010 205 16060 215
rect 16180 205 16230 215
rect 16350 205 16400 215
rect 16520 205 16570 215
rect 16690 205 16740 215
rect 16860 205 16910 215
rect 17030 205 17080 215
rect 17200 205 17250 215
rect 17370 205 17420 215
rect 17540 205 17590 215
rect 17710 205 17760 215
rect 17880 205 17930 215
rect 18050 205 18100 215
rect 18220 205 18270 215
rect 18390 205 18440 215
rect 18560 205 18610 215
rect 18730 205 18780 215
rect 18900 205 18950 215
rect 19070 205 19120 215
rect 19240 205 19290 215
rect 19410 205 19460 215
rect 19580 205 19630 215
rect 19750 205 19800 215
rect 19920 205 19970 215
rect 20090 205 20140 215
rect 20260 205 20310 215
rect 20430 205 20480 215
rect 20600 205 20650 215
rect 20770 205 20820 215
rect 20940 205 20990 215
rect 21110 205 21160 215
rect 21280 205 21330 215
rect 21450 205 21500 215
rect 21620 205 21670 215
rect 21790 205 21840 215
rect 21960 205 22010 215
rect 22130 205 22180 215
rect 22300 205 22350 215
rect 22470 205 22520 215
rect 22640 205 22690 215
rect 22810 205 22860 215
rect 22980 205 23030 215
rect 23150 205 23200 215
rect 23320 205 23370 215
rect 23490 205 23540 215
rect 23660 205 23710 215
rect 23830 205 23880 215
rect 24000 205 24050 215
rect 24170 205 24220 215
rect 24340 205 24390 215
rect 24510 205 24560 215
rect 24680 205 24730 215
rect 24850 205 24900 215
rect 25020 205 25070 215
rect 25190 205 25240 215
rect 25360 205 25410 215
rect 25530 205 25580 215
rect 25700 205 25750 215
rect 25870 205 25920 215
rect 26040 205 26090 215
rect 26210 205 26260 215
rect 26380 205 26430 215
rect 26550 205 26600 215
rect 26720 205 26770 215
rect 26890 205 26940 215
rect 27060 205 27110 215
rect 27230 205 27280 215
rect 27400 205 27450 215
rect 27570 205 27620 215
rect 27740 205 27790 215
rect 27910 205 27960 215
rect 28080 205 28130 215
rect 28250 205 28300 215
rect 28420 205 28470 215
rect 28590 205 28640 215
rect 28760 205 28810 215
rect 28930 205 28980 215
rect 29100 205 29150 215
rect 29270 205 29320 215
rect 29440 205 29490 215
rect 29610 205 29660 215
rect 215 175 225 205
rect 255 175 395 205
rect 425 175 565 205
rect 595 175 615 205
rect 750 175 760 205
rect 790 175 930 205
rect 960 175 1100 205
rect 1130 175 1270 205
rect 1300 175 1440 205
rect 1470 175 1610 205
rect 1640 175 1780 205
rect 1810 175 1950 205
rect 1980 175 2120 205
rect 2150 175 2170 205
rect 2260 175 2270 205
rect 2300 175 2440 205
rect 2470 175 2610 205
rect 2640 175 2780 205
rect 2810 175 2950 205
rect 2980 175 3120 205
rect 3150 175 3290 205
rect 3320 175 3460 205
rect 3490 175 3630 205
rect 3660 175 3800 205
rect 3830 175 3970 205
rect 4000 175 4140 205
rect 4170 175 4310 205
rect 4340 175 4480 205
rect 4510 175 4650 205
rect 4680 175 4820 205
rect 4850 175 4990 205
rect 5020 175 5160 205
rect 5190 175 5330 205
rect 5360 175 5500 205
rect 5530 175 5670 205
rect 5700 175 5840 205
rect 5870 175 6010 205
rect 6040 175 6180 205
rect 6210 175 6350 205
rect 6380 175 6520 205
rect 6550 175 6690 205
rect 6720 175 6860 205
rect 6890 175 7030 205
rect 7060 175 7200 205
rect 7230 175 7370 205
rect 7400 175 7540 205
rect 7570 175 7710 205
rect 7740 175 7760 205
rect 7850 175 7860 205
rect 7890 175 8030 205
rect 8060 175 8200 205
rect 8230 175 8370 205
rect 8400 175 8540 205
rect 8570 175 8710 205
rect 8740 175 8880 205
rect 8910 175 9050 205
rect 9080 175 9220 205
rect 9250 175 9390 205
rect 9420 175 9560 205
rect 9590 175 9730 205
rect 9760 175 9900 205
rect 9930 175 10070 205
rect 10100 175 10240 205
rect 10270 175 10410 205
rect 10440 175 10580 205
rect 10610 175 10750 205
rect 10780 175 10920 205
rect 10950 175 11090 205
rect 11120 175 11260 205
rect 11290 175 11430 205
rect 11460 175 11600 205
rect 11630 175 11770 205
rect 11800 175 11940 205
rect 11970 175 12110 205
rect 12140 175 12280 205
rect 12310 175 12450 205
rect 12480 175 12620 205
rect 12650 175 12790 205
rect 12820 175 12960 205
rect 12990 175 13130 205
rect 13160 175 13300 205
rect 13330 175 13470 205
rect 13500 175 13640 205
rect 13670 175 13810 205
rect 13840 175 13980 205
rect 14010 175 14150 205
rect 14180 175 14320 205
rect 14350 175 14490 205
rect 14520 175 14660 205
rect 14690 175 14830 205
rect 14860 175 15000 205
rect 15030 175 15170 205
rect 15200 175 15340 205
rect 15370 175 15510 205
rect 15540 175 15680 205
rect 15710 175 15850 205
rect 15880 175 16020 205
rect 16050 175 16190 205
rect 16220 175 16360 205
rect 16390 175 16530 205
rect 16560 175 16700 205
rect 16730 175 16870 205
rect 16900 175 17040 205
rect 17070 175 17210 205
rect 17240 175 17380 205
rect 17410 175 17550 205
rect 17580 175 17720 205
rect 17750 175 17890 205
rect 17920 175 18060 205
rect 18090 175 18230 205
rect 18260 175 18400 205
rect 18430 175 18570 205
rect 18600 175 18740 205
rect 18770 175 18910 205
rect 18940 175 19080 205
rect 19110 175 19250 205
rect 19280 175 19420 205
rect 19450 175 19590 205
rect 19620 175 19760 205
rect 19790 175 19930 205
rect 19960 175 20100 205
rect 20130 175 20270 205
rect 20300 175 20440 205
rect 20470 175 20610 205
rect 20640 175 20780 205
rect 20810 175 20950 205
rect 20980 175 21120 205
rect 21150 175 21290 205
rect 21320 175 21460 205
rect 21490 175 21630 205
rect 21660 175 21800 205
rect 21830 175 21970 205
rect 22000 175 22140 205
rect 22170 175 22310 205
rect 22340 175 22480 205
rect 22510 175 22650 205
rect 22680 175 22820 205
rect 22850 175 22990 205
rect 23020 175 23160 205
rect 23190 175 23330 205
rect 23360 175 23500 205
rect 23530 175 23670 205
rect 23700 175 23840 205
rect 23870 175 24010 205
rect 24040 175 24180 205
rect 24210 175 24350 205
rect 24380 175 24520 205
rect 24550 175 24690 205
rect 24720 175 24860 205
rect 24890 175 25030 205
rect 25060 175 25200 205
rect 25230 175 25370 205
rect 25400 175 25540 205
rect 25570 175 25710 205
rect 25740 175 25880 205
rect 25910 175 26050 205
rect 26080 175 26220 205
rect 26250 175 26390 205
rect 26420 175 26560 205
rect 26590 175 26730 205
rect 26760 175 26900 205
rect 26930 175 27070 205
rect 27100 175 27240 205
rect 27270 175 27410 205
rect 27440 175 27580 205
rect 27610 175 27750 205
rect 27780 175 27920 205
rect 27950 175 28090 205
rect 28120 175 28260 205
rect 28290 175 28430 205
rect 28460 175 28600 205
rect 28630 175 28770 205
rect 28800 175 28940 205
rect 28970 175 29110 205
rect 29140 175 29280 205
rect 29310 175 29450 205
rect 29480 175 29620 205
rect 29650 175 29660 205
rect 215 165 265 175
rect 385 165 435 175
rect 555 165 605 175
rect 750 165 800 175
rect 920 165 970 175
rect 1090 165 1140 175
rect 1260 165 1310 175
rect 1430 165 1480 175
rect 1600 165 1650 175
rect 1770 165 1820 175
rect 1940 165 1990 175
rect 2110 165 2160 175
rect 2260 165 2310 175
rect 2430 165 2480 175
rect 2600 165 2650 175
rect 2770 165 2820 175
rect 2940 165 2990 175
rect 3110 165 3160 175
rect 3280 165 3330 175
rect 3450 165 3500 175
rect 3620 165 3670 175
rect 3790 165 3840 175
rect 3960 165 4010 175
rect 4130 165 4180 175
rect 4300 165 4350 175
rect 4470 165 4520 175
rect 4640 165 4690 175
rect 4810 165 4860 175
rect 4980 165 5030 175
rect 5150 165 5200 175
rect 5320 165 5370 175
rect 5490 165 5540 175
rect 5660 165 5710 175
rect 5830 165 5880 175
rect 6000 165 6050 175
rect 6170 165 6220 175
rect 6340 165 6390 175
rect 6510 165 6560 175
rect 6680 165 6730 175
rect 6850 165 6900 175
rect 7020 165 7070 175
rect 7190 165 7240 175
rect 7360 165 7410 175
rect 7530 165 7580 175
rect 7700 165 7750 175
rect 7850 165 7900 175
rect 8020 165 8070 175
rect 8190 165 8240 175
rect 8360 165 8410 175
rect 8530 165 8580 175
rect 8700 165 8750 175
rect 8870 165 8920 175
rect 9040 165 9090 175
rect 9210 165 9260 175
rect 9380 165 9430 175
rect 9550 165 9600 175
rect 9720 165 9770 175
rect 9890 165 9940 175
rect 10060 165 10110 175
rect 10230 165 10280 175
rect 10400 165 10450 175
rect 10570 165 10620 175
rect 10740 165 10790 175
rect 10910 165 10960 175
rect 11080 165 11130 175
rect 11250 165 11300 175
rect 11420 165 11470 175
rect 11590 165 11640 175
rect 11760 165 11810 175
rect 11930 165 11980 175
rect 12100 165 12150 175
rect 12270 165 12320 175
rect 12440 165 12490 175
rect 12610 165 12660 175
rect 12780 165 12830 175
rect 12950 165 13000 175
rect 13120 165 13170 175
rect 13290 165 13340 175
rect 13460 165 13510 175
rect 13630 165 13680 175
rect 13800 165 13850 175
rect 13970 165 14020 175
rect 14140 165 14190 175
rect 14310 165 14360 175
rect 14480 165 14530 175
rect 14650 165 14700 175
rect 14820 165 14870 175
rect 14990 165 15040 175
rect 15160 165 15210 175
rect 15330 165 15380 175
rect 15500 165 15550 175
rect 15670 165 15720 175
rect 15840 165 15890 175
rect 16010 165 16060 175
rect 16180 165 16230 175
rect 16350 165 16400 175
rect 16520 165 16570 175
rect 16690 165 16740 175
rect 16860 165 16910 175
rect 17030 165 17080 175
rect 17200 165 17250 175
rect 17370 165 17420 175
rect 17540 165 17590 175
rect 17710 165 17760 175
rect 17880 165 17930 175
rect 18050 165 18100 175
rect 18220 165 18270 175
rect 18390 165 18440 175
rect 18560 165 18610 175
rect 18730 165 18780 175
rect 18900 165 18950 175
rect 19070 165 19120 175
rect 19240 165 19290 175
rect 19410 165 19460 175
rect 19580 165 19630 175
rect 19750 165 19800 175
rect 19920 165 19970 175
rect 20090 165 20140 175
rect 20260 165 20310 175
rect 20430 165 20480 175
rect 20600 165 20650 175
rect 20770 165 20820 175
rect 20940 165 20990 175
rect 21110 165 21160 175
rect 21280 165 21330 175
rect 21450 165 21500 175
rect 21620 165 21670 175
rect 21790 165 21840 175
rect 21960 165 22010 175
rect 22130 165 22180 175
rect 22300 165 22350 175
rect 22470 165 22520 175
rect 22640 165 22690 175
rect 22810 165 22860 175
rect 22980 165 23030 175
rect 23150 165 23200 175
rect 23320 165 23370 175
rect 23490 165 23540 175
rect 23660 165 23710 175
rect 23830 165 23880 175
rect 24000 165 24050 175
rect 24170 165 24220 175
rect 24340 165 24390 175
rect 24510 165 24560 175
rect 24680 165 24730 175
rect 24850 165 24900 175
rect 25020 165 25070 175
rect 25190 165 25240 175
rect 25360 165 25410 175
rect 25530 165 25580 175
rect 25700 165 25750 175
rect 25870 165 25920 175
rect 26040 165 26090 175
rect 26210 165 26260 175
rect 26380 165 26430 175
rect 26550 165 26600 175
rect 26720 165 26770 175
rect 26890 165 26940 175
rect 27060 165 27110 175
rect 27230 165 27280 175
rect 27400 165 27450 175
rect 27570 165 27620 175
rect 27740 165 27790 175
rect 27910 165 27960 175
rect 28080 165 28130 175
rect 28250 165 28300 175
rect 28420 165 28470 175
rect 28590 165 28640 175
rect 28760 165 28810 175
rect 28930 165 28980 175
rect 29100 165 29150 175
rect 29270 165 29320 175
rect 29440 165 29490 175
rect 29610 165 29660 175
rect 305 100 345 105
rect 305 65 310 100
rect 340 65 345 100
rect -470 55 75 65
rect 305 60 345 65
rect 475 100 515 105
rect 475 65 480 100
rect 510 65 515 100
rect 475 60 515 65
rect 840 100 880 105
rect 840 65 845 100
rect 875 65 880 100
rect 840 60 880 65
rect 1010 100 1050 105
rect 1010 65 1015 100
rect 1045 65 1050 100
rect 1010 60 1050 65
rect 1180 100 1220 105
rect 1180 65 1185 100
rect 1215 65 1220 100
rect 1180 60 1220 65
rect 1350 100 1390 105
rect 1350 65 1355 100
rect 1385 65 1390 100
rect 1350 60 1390 65
rect 1520 100 1560 105
rect 1520 65 1525 100
rect 1555 65 1560 100
rect 1520 60 1560 65
rect 1690 100 1730 105
rect 1690 65 1695 100
rect 1725 65 1730 100
rect 1690 60 1730 65
rect 1860 100 1900 105
rect 1860 65 1865 100
rect 1895 65 1900 100
rect 1860 60 1900 65
rect 2030 100 2070 105
rect 2030 65 2035 100
rect 2065 65 2070 100
rect 2030 60 2070 65
rect 2350 100 2390 105
rect 2350 65 2355 100
rect 2385 65 2390 100
rect 2350 60 2390 65
rect 2520 100 2560 105
rect 2520 65 2525 100
rect 2555 65 2560 100
rect 2520 60 2560 65
rect 2690 100 2730 105
rect 2690 65 2695 100
rect 2725 65 2730 100
rect 2690 60 2730 65
rect 2860 100 2900 105
rect 2860 65 2865 100
rect 2895 65 2900 100
rect 2860 60 2900 65
rect 3030 100 3070 105
rect 3030 65 3035 100
rect 3065 65 3070 100
rect 3030 60 3070 65
rect 3200 100 3240 105
rect 3200 65 3205 100
rect 3235 65 3240 100
rect 3200 60 3240 65
rect 3370 100 3410 105
rect 3370 65 3375 100
rect 3405 65 3410 100
rect 3370 60 3410 65
rect 3540 100 3580 105
rect 3540 65 3545 100
rect 3575 65 3580 100
rect 3540 60 3580 65
rect 3710 100 3750 105
rect 3710 65 3715 100
rect 3745 65 3750 100
rect 3710 60 3750 65
rect 3880 100 3920 105
rect 3880 65 3885 100
rect 3915 65 3920 100
rect 3880 60 3920 65
rect 4050 100 4090 105
rect 4050 65 4055 100
rect 4085 65 4090 100
rect 4050 60 4090 65
rect 4220 100 4260 105
rect 4220 65 4225 100
rect 4255 65 4260 100
rect 4220 60 4260 65
rect 4390 100 4430 105
rect 4390 65 4395 100
rect 4425 65 4430 100
rect 4390 60 4430 65
rect 4560 100 4600 105
rect 4560 65 4565 100
rect 4595 65 4600 100
rect 4560 60 4600 65
rect 4730 100 4770 105
rect 4730 65 4735 100
rect 4765 65 4770 100
rect 4730 60 4770 65
rect 4900 100 4940 105
rect 4900 65 4905 100
rect 4935 65 4940 100
rect 4900 60 4940 65
rect 5070 100 5110 105
rect 5070 65 5075 100
rect 5105 65 5110 100
rect 5070 60 5110 65
rect 5240 100 5280 105
rect 5240 65 5245 100
rect 5275 65 5280 100
rect 5240 60 5280 65
rect 5410 100 5450 105
rect 5410 65 5415 100
rect 5445 65 5450 100
rect 5410 60 5450 65
rect 5580 100 5620 105
rect 5580 65 5585 100
rect 5615 65 5620 100
rect 5580 60 5620 65
rect 5750 100 5790 105
rect 5750 65 5755 100
rect 5785 65 5790 100
rect 5750 60 5790 65
rect 5920 100 5960 105
rect 5920 65 5925 100
rect 5955 65 5960 100
rect 5920 60 5960 65
rect 6090 100 6130 105
rect 6090 65 6095 100
rect 6125 65 6130 100
rect 6090 60 6130 65
rect 6260 100 6300 105
rect 6260 65 6265 100
rect 6295 65 6300 100
rect 6260 60 6300 65
rect 6430 100 6470 105
rect 6430 65 6435 100
rect 6465 65 6470 100
rect 6430 60 6470 65
rect 6600 100 6640 105
rect 6600 65 6605 100
rect 6635 65 6640 100
rect 6600 60 6640 65
rect 6770 100 6810 105
rect 6770 65 6775 100
rect 6805 65 6810 100
rect 6770 60 6810 65
rect 6940 100 6980 105
rect 6940 65 6945 100
rect 6975 65 6980 100
rect 6940 60 6980 65
rect 7110 100 7150 105
rect 7110 65 7115 100
rect 7145 65 7150 100
rect 7110 60 7150 65
rect 7280 100 7320 105
rect 7280 65 7285 100
rect 7315 65 7320 100
rect 7280 60 7320 65
rect 7450 100 7490 105
rect 7450 65 7455 100
rect 7485 65 7490 100
rect 7450 60 7490 65
rect 7620 100 7660 105
rect 7620 65 7625 100
rect 7655 65 7660 100
rect 7620 60 7660 65
rect 7940 100 7980 105
rect 7940 65 7945 100
rect 7975 65 7980 100
rect 7940 60 7980 65
rect 8110 100 8150 105
rect 8110 65 8115 100
rect 8145 65 8150 100
rect 8110 60 8150 65
rect 8280 100 8320 105
rect 8280 65 8285 100
rect 8315 65 8320 100
rect 8280 60 8320 65
rect 8450 100 8490 105
rect 8450 65 8455 100
rect 8485 65 8490 100
rect 8450 60 8490 65
rect 8620 100 8660 105
rect 8620 65 8625 100
rect 8655 65 8660 100
rect 8620 60 8660 65
rect 8790 100 8830 105
rect 8790 65 8795 100
rect 8825 65 8830 100
rect 8790 60 8830 65
rect 8960 100 9000 105
rect 8960 65 8965 100
rect 8995 65 9000 100
rect 8960 60 9000 65
rect 9130 100 9170 105
rect 9130 65 9135 100
rect 9165 65 9170 100
rect 9130 60 9170 65
rect 9300 100 9340 105
rect 9300 65 9305 100
rect 9335 65 9340 100
rect 9300 60 9340 65
rect 9470 100 9510 105
rect 9470 65 9475 100
rect 9505 65 9510 100
rect 9470 60 9510 65
rect 9640 100 9680 105
rect 9640 65 9645 100
rect 9675 65 9680 100
rect 9640 60 9680 65
rect 9810 100 9850 105
rect 9810 65 9815 100
rect 9845 65 9850 100
rect 9810 60 9850 65
rect 9980 100 10020 105
rect 9980 65 9985 100
rect 10015 65 10020 100
rect 9980 60 10020 65
rect 10150 100 10190 105
rect 10150 65 10155 100
rect 10185 65 10190 100
rect 10150 60 10190 65
rect 10320 100 10360 105
rect 10320 65 10325 100
rect 10355 65 10360 100
rect 10320 60 10360 65
rect 10490 100 10530 105
rect 10490 65 10495 100
rect 10525 65 10530 100
rect 10490 60 10530 65
rect 10660 100 10700 105
rect 10660 65 10665 100
rect 10695 65 10700 100
rect 10660 60 10700 65
rect 10830 100 10870 105
rect 10830 65 10835 100
rect 10865 65 10870 100
rect 10830 60 10870 65
rect 11000 100 11040 105
rect 11000 65 11005 100
rect 11035 65 11040 100
rect 11000 60 11040 65
rect 11170 100 11210 105
rect 11170 65 11175 100
rect 11205 65 11210 100
rect 11170 60 11210 65
rect 11340 100 11380 105
rect 11340 65 11345 100
rect 11375 65 11380 100
rect 11340 60 11380 65
rect 11510 100 11550 105
rect 11510 65 11515 100
rect 11545 65 11550 100
rect 11510 60 11550 65
rect 11680 100 11720 105
rect 11680 65 11685 100
rect 11715 65 11720 100
rect 11680 60 11720 65
rect 11850 100 11890 105
rect 11850 65 11855 100
rect 11885 65 11890 100
rect 11850 60 11890 65
rect 12020 100 12060 105
rect 12020 65 12025 100
rect 12055 65 12060 100
rect 12020 60 12060 65
rect 12190 100 12230 105
rect 12190 65 12195 100
rect 12225 65 12230 100
rect 12190 60 12230 65
rect 12360 100 12400 105
rect 12360 65 12365 100
rect 12395 65 12400 100
rect 12360 60 12400 65
rect 12530 100 12570 105
rect 12530 65 12535 100
rect 12565 65 12570 100
rect 12530 60 12570 65
rect 12700 100 12740 105
rect 12700 65 12705 100
rect 12735 65 12740 100
rect 12700 60 12740 65
rect 12870 100 12910 105
rect 12870 65 12875 100
rect 12905 65 12910 100
rect 12870 60 12910 65
rect 13040 100 13080 105
rect 13040 65 13045 100
rect 13075 65 13080 100
rect 13040 60 13080 65
rect 13210 100 13250 105
rect 13210 65 13215 100
rect 13245 65 13250 100
rect 13210 60 13250 65
rect 13380 100 13420 105
rect 13380 65 13385 100
rect 13415 65 13420 100
rect 13380 60 13420 65
rect 13550 100 13590 105
rect 13550 65 13555 100
rect 13585 65 13590 100
rect 13550 60 13590 65
rect 13720 100 13760 105
rect 13720 65 13725 100
rect 13755 65 13760 100
rect 13720 60 13760 65
rect 13890 100 13930 105
rect 13890 65 13895 100
rect 13925 65 13930 100
rect 13890 60 13930 65
rect 14060 100 14100 105
rect 14060 65 14065 100
rect 14095 65 14100 100
rect 14060 60 14100 65
rect 14230 100 14270 105
rect 14230 65 14235 100
rect 14265 65 14270 100
rect 14230 60 14270 65
rect 14400 100 14440 105
rect 14400 65 14405 100
rect 14435 65 14440 100
rect 14400 60 14440 65
rect 14570 100 14610 105
rect 14570 65 14575 100
rect 14605 65 14610 100
rect 14570 60 14610 65
rect 14740 100 14780 105
rect 14740 65 14745 100
rect 14775 65 14780 100
rect 14740 60 14780 65
rect 14910 100 14950 105
rect 14910 65 14915 100
rect 14945 65 14950 100
rect 14910 60 14950 65
rect 15080 100 15120 105
rect 15080 65 15085 100
rect 15115 65 15120 100
rect 15080 60 15120 65
rect 15250 100 15290 105
rect 15250 65 15255 100
rect 15285 65 15290 100
rect 15250 60 15290 65
rect 15420 100 15460 105
rect 15420 65 15425 100
rect 15455 65 15460 100
rect 15420 60 15460 65
rect 15590 100 15630 105
rect 15590 65 15595 100
rect 15625 65 15630 100
rect 15590 60 15630 65
rect 15760 100 15800 105
rect 15760 65 15765 100
rect 15795 65 15800 100
rect 15760 60 15800 65
rect 15930 100 15970 105
rect 15930 65 15935 100
rect 15965 65 15970 100
rect 15930 60 15970 65
rect 16100 100 16140 105
rect 16100 65 16105 100
rect 16135 65 16140 100
rect 16100 60 16140 65
rect 16270 100 16310 105
rect 16270 65 16275 100
rect 16305 65 16310 100
rect 16270 60 16310 65
rect 16440 100 16480 105
rect 16440 65 16445 100
rect 16475 65 16480 100
rect 16440 60 16480 65
rect 16610 100 16650 105
rect 16610 65 16615 100
rect 16645 65 16650 100
rect 16610 60 16650 65
rect 16780 100 16820 105
rect 16780 65 16785 100
rect 16815 65 16820 100
rect 16780 60 16820 65
rect 16950 100 16990 105
rect 16950 65 16955 100
rect 16985 65 16990 100
rect 16950 60 16990 65
rect 17120 100 17160 105
rect 17120 65 17125 100
rect 17155 65 17160 100
rect 17120 60 17160 65
rect 17290 100 17330 105
rect 17290 65 17295 100
rect 17325 65 17330 100
rect 17290 60 17330 65
rect 17460 100 17500 105
rect 17460 65 17465 100
rect 17495 65 17500 100
rect 17460 60 17500 65
rect 17630 100 17670 105
rect 17630 65 17635 100
rect 17665 65 17670 100
rect 17630 60 17670 65
rect 17800 100 17840 105
rect 17800 65 17805 100
rect 17835 65 17840 100
rect 17800 60 17840 65
rect 17970 100 18010 105
rect 17970 65 17975 100
rect 18005 65 18010 100
rect 17970 60 18010 65
rect 18140 100 18180 105
rect 18140 65 18145 100
rect 18175 65 18180 100
rect 18140 60 18180 65
rect 18310 100 18350 105
rect 18310 65 18315 100
rect 18345 65 18350 100
rect 18310 60 18350 65
rect 18480 100 18520 105
rect 18480 65 18485 100
rect 18515 65 18520 100
rect 18480 60 18520 65
rect 18650 100 18690 105
rect 18650 65 18655 100
rect 18685 65 18690 100
rect 18650 60 18690 65
rect 18820 100 18860 105
rect 18820 65 18825 100
rect 18855 65 18860 100
rect 18820 60 18860 65
rect 18990 100 19030 105
rect 18990 65 18995 100
rect 19025 65 19030 100
rect 18990 60 19030 65
rect 19160 100 19200 105
rect 19160 65 19165 100
rect 19195 65 19200 100
rect 19160 60 19200 65
rect 19330 100 19370 105
rect 19330 65 19335 100
rect 19365 65 19370 100
rect 19330 60 19370 65
rect 19500 100 19540 105
rect 19500 65 19505 100
rect 19535 65 19540 100
rect 19500 60 19540 65
rect 19670 100 19710 105
rect 19670 65 19675 100
rect 19705 65 19710 100
rect 19670 60 19710 65
rect 19840 100 19880 105
rect 19840 65 19845 100
rect 19875 65 19880 100
rect 19840 60 19880 65
rect 20010 100 20050 105
rect 20010 65 20015 100
rect 20045 65 20050 100
rect 20010 60 20050 65
rect 20180 100 20220 105
rect 20180 65 20185 100
rect 20215 65 20220 100
rect 20180 60 20220 65
rect 20350 100 20390 105
rect 20350 65 20355 100
rect 20385 65 20390 100
rect 20350 60 20390 65
rect 20520 100 20560 105
rect 20520 65 20525 100
rect 20555 65 20560 100
rect 20520 60 20560 65
rect 20690 100 20730 105
rect 20690 65 20695 100
rect 20725 65 20730 100
rect 20690 60 20730 65
rect 20860 100 20900 105
rect 20860 65 20865 100
rect 20895 65 20900 100
rect 20860 60 20900 65
rect 21030 100 21070 105
rect 21030 65 21035 100
rect 21065 65 21070 100
rect 21030 60 21070 65
rect 21200 100 21240 105
rect 21200 65 21205 100
rect 21235 65 21240 100
rect 21200 60 21240 65
rect 21370 100 21410 105
rect 21370 65 21375 100
rect 21405 65 21410 100
rect 21370 60 21410 65
rect 21540 100 21580 105
rect 21540 65 21545 100
rect 21575 65 21580 100
rect 21540 60 21580 65
rect 21710 100 21750 105
rect 21710 65 21715 100
rect 21745 65 21750 100
rect 21710 60 21750 65
rect 21880 100 21920 105
rect 21880 65 21885 100
rect 21915 65 21920 100
rect 21880 60 21920 65
rect 22050 100 22090 105
rect 22050 65 22055 100
rect 22085 65 22090 100
rect 22050 60 22090 65
rect 22220 100 22260 105
rect 22220 65 22225 100
rect 22255 65 22260 100
rect 22220 60 22260 65
rect 22390 100 22430 105
rect 22390 65 22395 100
rect 22425 65 22430 100
rect 22390 60 22430 65
rect 22560 100 22600 105
rect 22560 65 22565 100
rect 22595 65 22600 100
rect 22560 60 22600 65
rect 22730 100 22770 105
rect 22730 65 22735 100
rect 22765 65 22770 100
rect 22730 60 22770 65
rect 22900 100 22940 105
rect 22900 65 22905 100
rect 22935 65 22940 100
rect 22900 60 22940 65
rect 23070 100 23110 105
rect 23070 65 23075 100
rect 23105 65 23110 100
rect 23070 60 23110 65
rect 23240 100 23280 105
rect 23240 65 23245 100
rect 23275 65 23280 100
rect 23240 60 23280 65
rect 23410 100 23450 105
rect 23410 65 23415 100
rect 23445 65 23450 100
rect 23410 60 23450 65
rect 23580 100 23620 105
rect 23580 65 23585 100
rect 23615 65 23620 100
rect 23580 60 23620 65
rect 23750 100 23790 105
rect 23750 65 23755 100
rect 23785 65 23790 100
rect 23750 60 23790 65
rect 23920 100 23960 105
rect 23920 65 23925 100
rect 23955 65 23960 100
rect 23920 60 23960 65
rect 24090 100 24130 105
rect 24090 65 24095 100
rect 24125 65 24130 100
rect 24090 60 24130 65
rect 24260 100 24300 105
rect 24260 65 24265 100
rect 24295 65 24300 100
rect 24260 60 24300 65
rect 24430 100 24470 105
rect 24430 65 24435 100
rect 24465 65 24470 100
rect 24430 60 24470 65
rect 24600 100 24640 105
rect 24600 65 24605 100
rect 24635 65 24640 100
rect 24600 60 24640 65
rect 24770 100 24810 105
rect 24770 65 24775 100
rect 24805 65 24810 100
rect 24770 60 24810 65
rect 24940 100 24980 105
rect 24940 65 24945 100
rect 24975 65 24980 100
rect 24940 60 24980 65
rect 25110 100 25150 105
rect 25110 65 25115 100
rect 25145 65 25150 100
rect 25110 60 25150 65
rect 25280 100 25320 105
rect 25280 65 25285 100
rect 25315 65 25320 100
rect 25280 60 25320 65
rect 25450 100 25490 105
rect 25450 65 25455 100
rect 25485 65 25490 100
rect 25450 60 25490 65
rect 25620 100 25660 105
rect 25620 65 25625 100
rect 25655 65 25660 100
rect 25620 60 25660 65
rect 25790 100 25830 105
rect 25790 65 25795 100
rect 25825 65 25830 100
rect 25790 60 25830 65
rect 25960 100 26000 105
rect 25960 65 25965 100
rect 25995 65 26000 100
rect 25960 60 26000 65
rect 26130 100 26170 105
rect 26130 65 26135 100
rect 26165 65 26170 100
rect 26130 60 26170 65
rect 26300 100 26340 105
rect 26300 65 26305 100
rect 26335 65 26340 100
rect 26300 60 26340 65
rect 26470 100 26510 105
rect 26470 65 26475 100
rect 26505 65 26510 100
rect 26470 60 26510 65
rect 26640 100 26680 105
rect 26640 65 26645 100
rect 26675 65 26680 100
rect 26640 60 26680 65
rect 26810 100 26850 105
rect 26810 65 26815 100
rect 26845 65 26850 100
rect 26810 60 26850 65
rect 26980 100 27020 105
rect 26980 65 26985 100
rect 27015 65 27020 100
rect 26980 60 27020 65
rect 27150 100 27190 105
rect 27150 65 27155 100
rect 27185 65 27190 100
rect 27150 60 27190 65
rect 27320 100 27360 105
rect 27320 65 27325 100
rect 27355 65 27360 100
rect 27320 60 27360 65
rect 27490 100 27530 105
rect 27490 65 27495 100
rect 27525 65 27530 100
rect 27490 60 27530 65
rect 27660 100 27700 105
rect 27660 65 27665 100
rect 27695 65 27700 100
rect 27660 60 27700 65
rect 27830 100 27870 105
rect 27830 65 27835 100
rect 27865 65 27870 100
rect 27830 60 27870 65
rect 28000 100 28040 105
rect 28000 65 28005 100
rect 28035 65 28040 100
rect 28000 60 28040 65
rect 28170 100 28210 105
rect 28170 65 28175 100
rect 28205 65 28210 100
rect 28170 60 28210 65
rect 28340 100 28380 105
rect 28340 65 28345 100
rect 28375 65 28380 100
rect 28340 60 28380 65
rect 28510 100 28550 105
rect 28510 65 28515 100
rect 28545 65 28550 100
rect 28510 60 28550 65
rect 28680 100 28720 105
rect 28680 65 28685 100
rect 28715 65 28720 100
rect 28680 60 28720 65
rect 28850 100 28890 105
rect 28850 65 28855 100
rect 28885 65 28890 100
rect 28850 60 28890 65
rect 29020 100 29060 105
rect 29020 65 29025 100
rect 29055 65 29060 100
rect 29020 60 29060 65
rect 29190 100 29230 105
rect 29190 65 29195 100
rect 29225 65 29230 100
rect 29190 60 29230 65
rect 29360 100 29400 105
rect 29360 65 29365 100
rect 29395 65 29400 100
rect 29360 60 29400 65
rect 29530 100 29570 105
rect 29530 65 29535 100
rect 29565 65 29570 100
rect 29530 60 29570 65
rect -470 15 35 55
rect 65 15 75 55
rect -470 5 75 15
rect 215 40 265 50
rect 385 40 435 50
rect 555 40 605 50
rect 215 10 225 40
rect 255 10 395 40
rect 425 10 565 40
rect 595 10 605 40
rect 215 0 265 10
rect 385 0 435 10
rect 555 0 605 10
rect 750 40 800 50
rect 920 40 970 50
rect 1090 40 1140 50
rect 1260 40 1310 50
rect 1430 40 1480 50
rect 1600 40 1650 50
rect 1770 40 1820 50
rect 1940 40 1990 50
rect 2110 40 2160 50
rect 750 10 760 40
rect 790 10 930 40
rect 960 10 1100 40
rect 1130 10 1270 40
rect 1300 10 1440 40
rect 1470 10 1610 40
rect 1640 10 1780 40
rect 1810 10 1950 40
rect 1980 10 2120 40
rect 2150 10 2160 40
rect 750 0 800 10
rect 920 0 970 10
rect 1090 0 1140 10
rect 1260 0 1310 10
rect 1430 0 1480 10
rect 1600 0 1650 10
rect 1770 0 1820 10
rect 1940 0 1990 10
rect 2110 0 2160 10
rect 2260 40 2310 50
rect 2430 40 2480 50
rect 2600 40 2650 50
rect 2770 40 2820 50
rect 2940 40 2990 50
rect 3110 40 3160 50
rect 3280 40 3330 50
rect 3450 40 3500 50
rect 3620 40 3670 50
rect 3790 40 3840 50
rect 3960 40 4010 50
rect 4130 40 4180 50
rect 4300 40 4350 50
rect 4470 40 4520 50
rect 4640 40 4690 50
rect 4810 40 4860 50
rect 4980 40 5030 50
rect 5150 40 5200 50
rect 5320 40 5370 50
rect 5490 40 5540 50
rect 5660 40 5710 50
rect 5830 40 5880 50
rect 6000 40 6050 50
rect 6170 40 6220 50
rect 6340 40 6390 50
rect 6510 40 6560 50
rect 6680 40 6730 50
rect 6850 40 6900 50
rect 7020 40 7070 50
rect 7190 40 7240 50
rect 7360 40 7410 50
rect 7530 40 7580 50
rect 7700 40 7750 50
rect 2260 10 2270 40
rect 2300 10 2440 40
rect 2470 10 2610 40
rect 2640 10 2780 40
rect 2810 10 2950 40
rect 2980 10 3120 40
rect 3150 10 3290 40
rect 3320 10 3460 40
rect 3490 10 3630 40
rect 3660 10 3800 40
rect 3830 10 3970 40
rect 4000 10 4140 40
rect 4170 10 4310 40
rect 4340 10 4480 40
rect 4510 10 4650 40
rect 4680 10 4820 40
rect 4850 10 4990 40
rect 5020 10 5160 40
rect 5190 10 5330 40
rect 5360 10 5500 40
rect 5530 10 5670 40
rect 5700 10 5840 40
rect 5870 10 6010 40
rect 6040 10 6180 40
rect 6210 10 6350 40
rect 6380 10 6520 40
rect 6550 10 6690 40
rect 6720 10 6860 40
rect 6890 10 7030 40
rect 7060 10 7200 40
rect 7230 10 7370 40
rect 7400 10 7540 40
rect 7570 10 7710 40
rect 7740 10 7750 40
rect 2260 0 2310 10
rect 2430 0 2480 10
rect 2600 0 2650 10
rect 2770 0 2820 10
rect 2940 0 2990 10
rect 3110 0 3160 10
rect 3280 0 3330 10
rect 3450 0 3500 10
rect 3620 0 3670 10
rect 3790 0 3840 10
rect 3960 0 4010 10
rect 4130 0 4180 10
rect 4300 0 4350 10
rect 4470 0 4520 10
rect 4640 0 4690 10
rect 4810 0 4860 10
rect 4980 0 5030 10
rect 5150 0 5200 10
rect 5320 0 5370 10
rect 5490 0 5540 10
rect 5660 0 5710 10
rect 5830 0 5880 10
rect 6000 0 6050 10
rect 6170 0 6220 10
rect 6340 0 6390 10
rect 6510 0 6560 10
rect 6680 0 6730 10
rect 6850 0 6900 10
rect 7020 0 7070 10
rect 7190 0 7240 10
rect 7360 0 7410 10
rect 7530 0 7580 10
rect 7700 0 7750 10
rect 7850 40 7900 50
rect 8020 40 8070 50
rect 8190 40 8240 50
rect 8360 40 8410 50
rect 8530 40 8580 50
rect 8700 40 8750 50
rect 8870 40 8920 50
rect 9040 40 9090 50
rect 9210 40 9260 50
rect 9380 40 9430 50
rect 9550 40 9600 50
rect 9720 40 9770 50
rect 9890 40 9940 50
rect 10060 40 10110 50
rect 10230 40 10280 50
rect 10400 40 10450 50
rect 10570 40 10620 50
rect 10740 40 10790 50
rect 10910 40 10960 50
rect 11080 40 11130 50
rect 11250 40 11300 50
rect 11420 40 11470 50
rect 11590 40 11640 50
rect 11760 40 11810 50
rect 11930 40 11980 50
rect 12100 40 12150 50
rect 12270 40 12320 50
rect 12440 40 12490 50
rect 12610 40 12660 50
rect 12780 40 12830 50
rect 12950 40 13000 50
rect 13120 40 13170 50
rect 13290 40 13340 50
rect 13460 40 13510 50
rect 13630 40 13680 50
rect 13800 40 13850 50
rect 13970 40 14020 50
rect 14140 40 14190 50
rect 14310 40 14360 50
rect 14480 40 14530 50
rect 14650 40 14700 50
rect 14820 40 14870 50
rect 14990 40 15040 50
rect 15160 40 15210 50
rect 15330 40 15380 50
rect 15500 40 15550 50
rect 15670 40 15720 50
rect 15840 40 15890 50
rect 16010 40 16060 50
rect 16180 40 16230 50
rect 16350 40 16400 50
rect 16520 40 16570 50
rect 16690 40 16740 50
rect 16860 40 16910 50
rect 17030 40 17080 50
rect 17200 40 17250 50
rect 17370 40 17420 50
rect 17540 40 17590 50
rect 17710 40 17760 50
rect 17880 40 17930 50
rect 18050 40 18100 50
rect 18220 40 18270 50
rect 18390 40 18440 50
rect 18560 40 18610 50
rect 18730 40 18780 50
rect 18900 40 18950 50
rect 19070 40 19120 50
rect 19240 40 19290 50
rect 19410 40 19460 50
rect 19580 40 19630 50
rect 19750 40 19800 50
rect 19920 40 19970 50
rect 20090 40 20140 50
rect 20260 40 20310 50
rect 20430 40 20480 50
rect 20600 40 20650 50
rect 20770 40 20820 50
rect 20940 40 20990 50
rect 21110 40 21160 50
rect 21280 40 21330 50
rect 21450 40 21500 50
rect 21620 40 21670 50
rect 21790 40 21840 50
rect 21960 40 22010 50
rect 22130 40 22180 50
rect 22300 40 22350 50
rect 22470 40 22520 50
rect 22640 40 22690 50
rect 22810 40 22860 50
rect 22980 40 23030 50
rect 23150 40 23200 50
rect 23320 40 23370 50
rect 23490 40 23540 50
rect 23660 40 23710 50
rect 23830 40 23880 50
rect 24000 40 24050 50
rect 24170 40 24220 50
rect 24340 40 24390 50
rect 24510 40 24560 50
rect 24680 40 24730 50
rect 24850 40 24900 50
rect 25020 40 25070 50
rect 25190 40 25240 50
rect 25360 40 25410 50
rect 25530 40 25580 50
rect 25700 40 25750 50
rect 25870 40 25920 50
rect 26040 40 26090 50
rect 26210 40 26260 50
rect 26380 40 26430 50
rect 26550 40 26600 50
rect 26720 40 26770 50
rect 26890 40 26940 50
rect 27060 40 27110 50
rect 27230 40 27280 50
rect 27400 40 27450 50
rect 27570 40 27620 50
rect 27740 40 27790 50
rect 27910 40 27960 50
rect 28080 40 28130 50
rect 28250 40 28300 50
rect 28420 40 28470 50
rect 28590 40 28640 50
rect 28760 40 28810 50
rect 28930 40 28980 50
rect 29100 40 29150 50
rect 29270 40 29320 50
rect 29440 40 29490 50
rect 29610 40 29660 50
rect 7850 10 7860 40
rect 7890 10 8030 40
rect 8060 10 8200 40
rect 8230 10 8370 40
rect 8400 10 8540 40
rect 8570 10 8710 40
rect 8740 10 8880 40
rect 8910 10 9050 40
rect 9080 10 9220 40
rect 9250 10 9390 40
rect 9420 10 9560 40
rect 9590 10 9730 40
rect 9760 10 9900 40
rect 9930 10 10070 40
rect 10100 10 10240 40
rect 10270 10 10410 40
rect 10440 10 10580 40
rect 10610 10 10750 40
rect 10780 10 10920 40
rect 10950 10 11090 40
rect 11120 10 11260 40
rect 11290 10 11430 40
rect 11460 10 11600 40
rect 11630 10 11770 40
rect 11800 10 11940 40
rect 11970 10 12110 40
rect 12140 10 12280 40
rect 12310 10 12450 40
rect 12480 10 12620 40
rect 12650 10 12790 40
rect 12820 10 12960 40
rect 12990 10 13130 40
rect 13160 10 13300 40
rect 13330 10 13470 40
rect 13500 10 13640 40
rect 13670 10 13810 40
rect 13840 10 13980 40
rect 14010 10 14150 40
rect 14180 10 14320 40
rect 14350 10 14490 40
rect 14520 10 14660 40
rect 14690 10 14830 40
rect 14860 10 15000 40
rect 15030 10 15170 40
rect 15200 10 15340 40
rect 15370 10 15510 40
rect 15540 10 15680 40
rect 15710 10 15850 40
rect 15880 10 16020 40
rect 16050 10 16190 40
rect 16220 10 16360 40
rect 16390 10 16530 40
rect 16560 10 16700 40
rect 16730 10 16870 40
rect 16900 10 17040 40
rect 17070 10 17210 40
rect 17240 10 17380 40
rect 17410 10 17550 40
rect 17580 10 17720 40
rect 17750 10 17890 40
rect 17920 10 18060 40
rect 18090 10 18230 40
rect 18260 10 18400 40
rect 18430 10 18570 40
rect 18600 10 18740 40
rect 18770 10 18910 40
rect 18940 10 19080 40
rect 19110 10 19250 40
rect 19280 10 19420 40
rect 19450 10 19590 40
rect 19620 10 19760 40
rect 19790 10 19930 40
rect 19960 10 20100 40
rect 20130 10 20270 40
rect 20300 10 20440 40
rect 20470 10 20610 40
rect 20640 10 20780 40
rect 20810 10 20950 40
rect 20980 10 21120 40
rect 21150 10 21290 40
rect 21320 10 21460 40
rect 21490 10 21630 40
rect 21660 10 21800 40
rect 21830 10 21970 40
rect 22000 10 22140 40
rect 22170 10 22310 40
rect 22340 10 22480 40
rect 22510 10 22650 40
rect 22680 10 22820 40
rect 22850 10 22990 40
rect 23020 10 23160 40
rect 23190 10 23330 40
rect 23360 10 23500 40
rect 23530 10 23670 40
rect 23700 10 23840 40
rect 23870 10 24010 40
rect 24040 10 24180 40
rect 24210 10 24350 40
rect 24380 10 24520 40
rect 24550 10 24690 40
rect 24720 10 24860 40
rect 24890 10 25030 40
rect 25060 10 25200 40
rect 25230 10 25370 40
rect 25400 10 25540 40
rect 25570 10 25710 40
rect 25740 10 25880 40
rect 25910 10 26050 40
rect 26080 10 26220 40
rect 26250 10 26390 40
rect 26420 10 26560 40
rect 26590 10 26730 40
rect 26760 10 26900 40
rect 26930 10 27070 40
rect 27100 10 27240 40
rect 27270 10 27410 40
rect 27440 10 27580 40
rect 27610 10 27750 40
rect 27780 10 27920 40
rect 27950 10 28090 40
rect 28120 10 28260 40
rect 28290 10 28430 40
rect 28460 10 28600 40
rect 28630 10 28770 40
rect 28800 10 28940 40
rect 28970 10 29110 40
rect 29140 10 29280 40
rect 29310 10 29450 40
rect 29480 10 29620 40
rect 29650 10 29660 40
rect 7850 0 7900 10
rect 8020 0 8070 10
rect 8190 0 8240 10
rect 8360 0 8410 10
rect 8530 0 8580 10
rect 8700 0 8750 10
rect 8870 0 8920 10
rect 9040 0 9090 10
rect 9210 0 9260 10
rect 9380 0 9430 10
rect 9550 0 9600 10
rect 9720 0 9770 10
rect 9890 0 9940 10
rect 10060 0 10110 10
rect 10230 0 10280 10
rect 10400 0 10450 10
rect 10570 0 10620 10
rect 10740 0 10790 10
rect 10910 0 10960 10
rect 11080 0 11130 10
rect 11250 0 11300 10
rect 11420 0 11470 10
rect 11590 0 11640 10
rect 11760 0 11810 10
rect 11930 0 11980 10
rect 12100 0 12150 10
rect 12270 0 12320 10
rect 12440 0 12490 10
rect 12610 0 12660 10
rect 12780 0 12830 10
rect 12950 0 13000 10
rect 13120 0 13170 10
rect 13290 0 13340 10
rect 13460 0 13510 10
rect 13630 0 13680 10
rect 13800 0 13850 10
rect 13970 0 14020 10
rect 14140 0 14190 10
rect 14310 0 14360 10
rect 14480 0 14530 10
rect 14650 0 14700 10
rect 14820 0 14870 10
rect 14990 0 15040 10
rect 15160 0 15210 10
rect 15330 0 15380 10
rect 15500 0 15550 10
rect 15670 0 15720 10
rect 15840 0 15890 10
rect 16010 0 16060 10
rect 16180 0 16230 10
rect 16350 0 16400 10
rect 16520 0 16570 10
rect 16690 0 16740 10
rect 16860 0 16910 10
rect 17030 0 17080 10
rect 17200 0 17250 10
rect 17370 0 17420 10
rect 17540 0 17590 10
rect 17710 0 17760 10
rect 17880 0 17930 10
rect 18050 0 18100 10
rect 18220 0 18270 10
rect 18390 0 18440 10
rect 18560 0 18610 10
rect 18730 0 18780 10
rect 18900 0 18950 10
rect 19070 0 19120 10
rect 19240 0 19290 10
rect 19410 0 19460 10
rect 19580 0 19630 10
rect 19750 0 19800 10
rect 19920 0 19970 10
rect 20090 0 20140 10
rect 20260 0 20310 10
rect 20430 0 20480 10
rect 20600 0 20650 10
rect 20770 0 20820 10
rect 20940 0 20990 10
rect 21110 0 21160 10
rect 21280 0 21330 10
rect 21450 0 21500 10
rect 21620 0 21670 10
rect 21790 0 21840 10
rect 21960 0 22010 10
rect 22130 0 22180 10
rect 22300 0 22350 10
rect 22470 0 22520 10
rect 22640 0 22690 10
rect 22810 0 22860 10
rect 22980 0 23030 10
rect 23150 0 23200 10
rect 23320 0 23370 10
rect 23490 0 23540 10
rect 23660 0 23710 10
rect 23830 0 23880 10
rect 24000 0 24050 10
rect 24170 0 24220 10
rect 24340 0 24390 10
rect 24510 0 24560 10
rect 24680 0 24730 10
rect 24850 0 24900 10
rect 25020 0 25070 10
rect 25190 0 25240 10
rect 25360 0 25410 10
rect 25530 0 25580 10
rect 25700 0 25750 10
rect 25870 0 25920 10
rect 26040 0 26090 10
rect 26210 0 26260 10
rect 26380 0 26430 10
rect 26550 0 26600 10
rect 26720 0 26770 10
rect 26890 0 26940 10
rect 27060 0 27110 10
rect 27230 0 27280 10
rect 27400 0 27450 10
rect 27570 0 27620 10
rect 27740 0 27790 10
rect 27910 0 27960 10
rect 28080 0 28130 10
rect 28250 0 28300 10
rect 28420 0 28470 10
rect 28590 0 28640 10
rect 28760 0 28810 10
rect 28930 0 28980 10
rect 29100 0 29150 10
rect 29270 0 29320 10
rect 29440 0 29490 10
rect 29610 0 29660 10
rect 90 -30 565 -20
rect 90 -60 100 -30
rect 130 -60 265 -30
rect 300 -60 350 -30
rect 385 -60 435 -30
rect 470 -60 520 -30
rect 555 -60 565 -30
rect 90 -70 565 -60
rect 645 -25 2120 -20
rect 645 -65 650 -25
rect 700 -30 2120 -25
rect 700 -60 800 -30
rect 835 -60 885 -30
rect 920 -60 970 -30
rect 1005 -60 1055 -30
rect 1090 -60 1140 -30
rect 1175 -60 1225 -30
rect 1260 -60 1310 -30
rect 1345 -60 1395 -30
rect 1430 -60 1480 -30
rect 1515 -60 1565 -30
rect 1600 -60 1650 -30
rect 1685 -60 1735 -30
rect 1770 -60 1820 -30
rect 1855 -60 1905 -30
rect 1940 -60 1990 -30
rect 2025 -60 2075 -30
rect 2110 -60 2120 -30
rect 700 -65 2120 -60
rect 645 -70 2120 -65
rect 2185 -25 7710 -20
rect 2185 -65 2190 -25
rect 2240 -30 7710 -25
rect 2240 -60 2310 -30
rect 2345 -60 2395 -30
rect 2430 -60 2480 -30
rect 2515 -60 2565 -30
rect 2600 -60 2650 -30
rect 2685 -60 2735 -30
rect 2770 -60 2820 -30
rect 2855 -60 2905 -30
rect 2940 -60 2990 -30
rect 3025 -60 3075 -30
rect 3110 -60 3160 -30
rect 3195 -60 3245 -30
rect 3280 -60 3330 -30
rect 3365 -60 3415 -30
rect 3450 -60 3500 -30
rect 3535 -60 3585 -30
rect 3620 -60 3670 -30
rect 3705 -60 3755 -30
rect 3790 -60 3840 -30
rect 3875 -60 3925 -30
rect 3960 -60 4010 -30
rect 4045 -60 4095 -30
rect 4130 -60 4180 -30
rect 4215 -60 4265 -30
rect 4300 -60 4350 -30
rect 4385 -60 4435 -30
rect 4470 -60 4520 -30
rect 4555 -60 4605 -30
rect 4640 -60 4690 -30
rect 4725 -60 4775 -30
rect 4810 -60 4860 -30
rect 4895 -60 4945 -30
rect 4980 -60 5030 -30
rect 5065 -60 5115 -30
rect 5150 -60 5200 -30
rect 5235 -60 5285 -30
rect 5320 -60 5370 -30
rect 5405 -60 5455 -30
rect 5490 -60 5540 -30
rect 5575 -60 5625 -30
rect 5660 -60 5710 -30
rect 5745 -60 5795 -30
rect 5830 -60 5880 -30
rect 5915 -60 5965 -30
rect 6000 -60 6050 -30
rect 6085 -60 6135 -30
rect 6170 -60 6220 -30
rect 6255 -60 6305 -30
rect 6340 -60 6390 -30
rect 6425 -60 6475 -30
rect 6510 -60 6560 -30
rect 6595 -60 6645 -30
rect 6680 -60 6730 -30
rect 6765 -60 6815 -30
rect 6850 -60 6900 -30
rect 6935 -60 6985 -30
rect 7020 -60 7070 -30
rect 7105 -60 7155 -30
rect 7190 -60 7240 -30
rect 7275 -60 7325 -30
rect 7360 -60 7410 -30
rect 7445 -60 7495 -30
rect 7530 -60 7580 -30
rect 7615 -60 7665 -30
rect 7700 -60 7710 -30
rect 2240 -65 7710 -60
rect 2185 -70 7710 -65
rect 7775 -25 29620 -20
rect 7775 -65 7780 -25
rect 7830 -30 29620 -25
rect 7830 -60 7900 -30
rect 7935 -60 7985 -30
rect 8020 -60 8070 -30
rect 8105 -60 8155 -30
rect 8190 -60 8240 -30
rect 8275 -60 8325 -30
rect 8360 -60 8410 -30
rect 8445 -60 8495 -30
rect 8530 -60 8580 -30
rect 8615 -60 8665 -30
rect 8700 -60 8750 -30
rect 8785 -60 8835 -30
rect 8870 -60 8920 -30
rect 8955 -60 9005 -30
rect 9040 -60 9090 -30
rect 9125 -60 9175 -30
rect 9210 -60 9260 -30
rect 9295 -60 9345 -30
rect 9380 -60 9430 -30
rect 9465 -60 9515 -30
rect 9550 -60 9600 -30
rect 9635 -60 9685 -30
rect 9720 -60 9770 -30
rect 9805 -60 9855 -30
rect 9890 -60 9940 -30
rect 9975 -60 10025 -30
rect 10060 -60 10110 -30
rect 10145 -60 10195 -30
rect 10230 -60 10280 -30
rect 10315 -60 10365 -30
rect 10400 -60 10450 -30
rect 10485 -60 10535 -30
rect 10570 -60 10620 -30
rect 10655 -60 10705 -30
rect 10740 -60 10790 -30
rect 10825 -60 10875 -30
rect 10910 -60 10960 -30
rect 10995 -60 11045 -30
rect 11080 -60 11130 -30
rect 11165 -60 11215 -30
rect 11250 -60 11300 -30
rect 11335 -60 11385 -30
rect 11420 -60 11470 -30
rect 11505 -60 11555 -30
rect 11590 -60 11640 -30
rect 11675 -60 11725 -30
rect 11760 -60 11810 -30
rect 11845 -60 11895 -30
rect 11930 -60 11980 -30
rect 12015 -60 12065 -30
rect 12100 -60 12150 -30
rect 12185 -60 12235 -30
rect 12270 -60 12320 -30
rect 12355 -60 12405 -30
rect 12440 -60 12490 -30
rect 12525 -60 12575 -30
rect 12610 -60 12660 -30
rect 12695 -60 12745 -30
rect 12780 -60 12830 -30
rect 12865 -60 12915 -30
rect 12950 -60 13000 -30
rect 13035 -60 13085 -30
rect 13120 -60 13170 -30
rect 13205 -60 13255 -30
rect 13290 -60 13340 -30
rect 13375 -60 13425 -30
rect 13460 -60 13510 -30
rect 13545 -60 13595 -30
rect 13630 -60 13680 -30
rect 13715 -60 13765 -30
rect 13800 -60 13850 -30
rect 13885 -60 13935 -30
rect 13970 -60 14020 -30
rect 14055 -60 14105 -30
rect 14140 -60 14190 -30
rect 14225 -60 14275 -30
rect 14310 -60 14360 -30
rect 14395 -60 14445 -30
rect 14480 -60 14530 -30
rect 14565 -60 14615 -30
rect 14650 -60 14700 -30
rect 14735 -60 14785 -30
rect 14820 -60 14870 -30
rect 14905 -60 14955 -30
rect 14990 -60 15040 -30
rect 15075 -60 15125 -30
rect 15160 -60 15210 -30
rect 15245 -60 15295 -30
rect 15330 -60 15380 -30
rect 15415 -60 15465 -30
rect 15500 -60 15550 -30
rect 15585 -60 15635 -30
rect 15670 -60 15720 -30
rect 15755 -60 15805 -30
rect 15840 -60 15890 -30
rect 15925 -60 15975 -30
rect 16010 -60 16060 -30
rect 16095 -60 16145 -30
rect 16180 -60 16230 -30
rect 16265 -60 16315 -30
rect 16350 -60 16400 -30
rect 16435 -60 16485 -30
rect 16520 -60 16570 -30
rect 16605 -60 16655 -30
rect 16690 -60 16740 -30
rect 16775 -60 16825 -30
rect 16860 -60 16910 -30
rect 16945 -60 16995 -30
rect 17030 -60 17080 -30
rect 17115 -60 17165 -30
rect 17200 -60 17250 -30
rect 17285 -60 17335 -30
rect 17370 -60 17420 -30
rect 17455 -60 17505 -30
rect 17540 -60 17590 -30
rect 17625 -60 17675 -30
rect 17710 -60 17760 -30
rect 17795 -60 17845 -30
rect 17880 -60 17930 -30
rect 17965 -60 18015 -30
rect 18050 -60 18100 -30
rect 18135 -60 18185 -30
rect 18220 -60 18270 -30
rect 18305 -60 18355 -30
rect 18390 -60 18440 -30
rect 18475 -60 18525 -30
rect 18560 -60 18610 -30
rect 18645 -60 18695 -30
rect 18730 -60 18780 -30
rect 18815 -60 18865 -30
rect 18900 -60 18950 -30
rect 18985 -60 19035 -30
rect 19070 -60 19120 -30
rect 19155 -60 19205 -30
rect 19240 -60 19290 -30
rect 19325 -60 19375 -30
rect 19410 -60 19460 -30
rect 19495 -60 19545 -30
rect 19580 -60 19630 -30
rect 19665 -60 19715 -30
rect 19750 -60 19800 -30
rect 19835 -60 19885 -30
rect 19920 -60 19970 -30
rect 20005 -60 20055 -30
rect 20090 -60 20140 -30
rect 20175 -60 20225 -30
rect 20260 -60 20310 -30
rect 20345 -60 20395 -30
rect 20430 -60 20480 -30
rect 20515 -60 20565 -30
rect 20600 -60 20650 -30
rect 20685 -60 20735 -30
rect 20770 -60 20820 -30
rect 20855 -60 20905 -30
rect 20940 -60 20990 -30
rect 21025 -60 21075 -30
rect 21110 -60 21160 -30
rect 21195 -60 21245 -30
rect 21280 -60 21330 -30
rect 21365 -60 21415 -30
rect 21450 -60 21500 -30
rect 21535 -60 21585 -30
rect 21620 -60 21670 -30
rect 21705 -60 21755 -30
rect 21790 -60 21840 -30
rect 21875 -60 21925 -30
rect 21960 -60 22010 -30
rect 22045 -60 22095 -30
rect 22130 -60 22180 -30
rect 22215 -60 22265 -30
rect 22300 -60 22350 -30
rect 22385 -60 22435 -30
rect 22470 -60 22520 -30
rect 22555 -60 22605 -30
rect 22640 -60 22690 -30
rect 22725 -60 22775 -30
rect 22810 -60 22860 -30
rect 22895 -60 22945 -30
rect 22980 -60 23030 -30
rect 23065 -60 23115 -30
rect 23150 -60 23200 -30
rect 23235 -60 23285 -30
rect 23320 -60 23370 -30
rect 23405 -60 23455 -30
rect 23490 -60 23540 -30
rect 23575 -60 23625 -30
rect 23660 -60 23710 -30
rect 23745 -60 23795 -30
rect 23830 -60 23880 -30
rect 23915 -60 23965 -30
rect 24000 -60 24050 -30
rect 24085 -60 24135 -30
rect 24170 -60 24220 -30
rect 24255 -60 24305 -30
rect 24340 -60 24390 -30
rect 24425 -60 24475 -30
rect 24510 -60 24560 -30
rect 24595 -60 24645 -30
rect 24680 -60 24730 -30
rect 24765 -60 24815 -30
rect 24850 -60 24900 -30
rect 24935 -60 24985 -30
rect 25020 -60 25070 -30
rect 25105 -60 25155 -30
rect 25190 -60 25240 -30
rect 25275 -60 25325 -30
rect 25360 -60 25410 -30
rect 25445 -60 25495 -30
rect 25530 -60 25580 -30
rect 25615 -60 25665 -30
rect 25700 -60 25750 -30
rect 25785 -60 25835 -30
rect 25870 -60 25920 -30
rect 25955 -60 26005 -30
rect 26040 -60 26090 -30
rect 26125 -60 26175 -30
rect 26210 -60 26260 -30
rect 26295 -60 26345 -30
rect 26380 -60 26430 -30
rect 26465 -60 26515 -30
rect 26550 -60 26600 -30
rect 26635 -60 26685 -30
rect 26720 -60 26770 -30
rect 26805 -60 26855 -30
rect 26890 -60 26940 -30
rect 26975 -60 27025 -30
rect 27060 -60 27110 -30
rect 27145 -60 27195 -30
rect 27230 -60 27280 -30
rect 27315 -60 27365 -30
rect 27400 -60 27450 -30
rect 27485 -60 27535 -30
rect 27570 -60 27620 -30
rect 27655 -60 27705 -30
rect 27740 -60 27790 -30
rect 27825 -60 27875 -30
rect 27910 -60 27960 -30
rect 27995 -60 28045 -30
rect 28080 -60 28130 -30
rect 28165 -60 28215 -30
rect 28250 -60 28300 -30
rect 28335 -60 28385 -30
rect 28420 -60 28470 -30
rect 28505 -60 28555 -30
rect 28590 -60 28640 -30
rect 28675 -60 28725 -30
rect 28760 -60 28810 -30
rect 28845 -60 28895 -30
rect 28930 -60 28980 -30
rect 29015 -60 29065 -30
rect 29100 -60 29150 -30
rect 29185 -60 29235 -30
rect 29270 -60 29320 -30
rect 29355 -60 29405 -30
rect 29440 -60 29490 -30
rect 29525 -60 29575 -30
rect 29610 -60 29620 -30
rect 7830 -65 29620 -60
rect 7775 -70 29620 -65
rect 7925 -230 8005 -225
rect 7925 -255 7965 -230
rect 105 -260 7965 -255
rect 8000 -255 8005 -230
rect 15575 -230 15655 -225
rect 15575 -255 15615 -230
rect 8000 -260 15615 -255
rect 15650 -255 15655 -230
rect 29515 -230 29595 -225
rect 29515 -255 29555 -230
rect 15650 -260 29555 -255
rect 29590 -255 29595 -230
rect 29590 -260 43625 -255
rect 105 -265 43625 -260
rect 105 -295 115 -265
rect 150 -295 200 -265
rect 235 -295 285 -265
rect 320 -295 370 -265
rect 405 -295 455 -265
rect 490 -295 540 -265
rect 575 -295 625 -265
rect 660 -295 710 -265
rect 745 -295 795 -265
rect 830 -295 880 -265
rect 915 -295 965 -265
rect 1000 -295 1050 -265
rect 1085 -295 1135 -265
rect 1170 -295 1220 -265
rect 1255 -295 1305 -265
rect 1340 -295 1390 -265
rect 1425 -295 1475 -265
rect 1510 -295 1560 -265
rect 1595 -295 1645 -265
rect 1680 -295 1730 -265
rect 1765 -295 1815 -265
rect 1850 -295 1900 -265
rect 1935 -295 1985 -265
rect 2020 -295 2070 -265
rect 2105 -295 2155 -265
rect 2190 -295 2240 -265
rect 2275 -295 2325 -265
rect 2360 -295 2410 -265
rect 2445 -295 2495 -265
rect 2530 -295 2580 -265
rect 2615 -295 2665 -265
rect 2700 -295 2750 -265
rect 2785 -295 2835 -265
rect 2870 -295 2920 -265
rect 2955 -295 3005 -265
rect 3040 -295 3090 -265
rect 3125 -295 3175 -265
rect 3210 -295 3260 -265
rect 3295 -295 3345 -265
rect 3380 -295 3430 -265
rect 3465 -295 3515 -265
rect 3550 -295 3600 -265
rect 3635 -295 3685 -265
rect 3720 -295 3770 -265
rect 3805 -295 3855 -265
rect 3890 -295 3940 -265
rect 3975 -295 4025 -265
rect 4060 -295 4110 -265
rect 4145 -295 4195 -265
rect 4230 -295 4280 -265
rect 4315 -295 4365 -265
rect 4400 -295 4450 -265
rect 4485 -295 4535 -265
rect 4570 -295 4620 -265
rect 4655 -295 4705 -265
rect 4740 -295 4790 -265
rect 4825 -295 4875 -265
rect 4910 -295 4960 -265
rect 4995 -295 5045 -265
rect 5080 -295 5130 -265
rect 5165 -295 5215 -265
rect 5250 -295 5300 -265
rect 5335 -295 5385 -265
rect 5420 -295 5470 -265
rect 5505 -295 5555 -265
rect 5590 -295 5640 -265
rect 5675 -295 5725 -265
rect 5760 -295 5810 -265
rect 5845 -295 5895 -265
rect 5930 -295 5980 -265
rect 6015 -295 6065 -265
rect 6100 -295 6150 -265
rect 6185 -295 6235 -265
rect 6270 -295 6320 -265
rect 6355 -295 6405 -265
rect 6440 -295 6490 -265
rect 6525 -295 6575 -265
rect 6610 -295 6660 -265
rect 6695 -295 6745 -265
rect 6780 -295 6830 -265
rect 6865 -295 6915 -265
rect 6950 -295 7000 -265
rect 7035 -295 7085 -265
rect 7120 -295 7170 -265
rect 7205 -295 7255 -265
rect 7290 -295 7340 -265
rect 7375 -295 7425 -265
rect 7460 -295 7510 -265
rect 7545 -295 7595 -265
rect 7630 -295 7680 -265
rect 7715 -295 7765 -265
rect 7800 -295 7850 -265
rect 7885 -295 7935 -265
rect 7970 -295 8020 -265
rect 8055 -295 8105 -265
rect 8140 -295 8190 -265
rect 8225 -295 8275 -265
rect 8310 -295 8360 -265
rect 8395 -295 8445 -265
rect 8480 -295 8530 -265
rect 8565 -295 8615 -265
rect 8650 -295 8700 -265
rect 8735 -295 8785 -265
rect 8820 -295 8870 -265
rect 8905 -295 8955 -265
rect 8990 -295 9040 -265
rect 9075 -295 9125 -265
rect 9160 -295 9210 -265
rect 9245 -295 9295 -265
rect 9330 -295 9380 -265
rect 9415 -295 9465 -265
rect 9500 -295 9550 -265
rect 9585 -295 9635 -265
rect 9670 -295 9720 -265
rect 9755 -295 9805 -265
rect 9840 -295 9890 -265
rect 9925 -295 9975 -265
rect 10010 -295 10060 -265
rect 10095 -295 10145 -265
rect 10180 -295 10230 -265
rect 10265 -295 10315 -265
rect 10350 -295 10400 -265
rect 10435 -295 10485 -265
rect 10520 -295 10570 -265
rect 10605 -295 10655 -265
rect 10690 -295 10740 -265
rect 10775 -295 10825 -265
rect 10860 -295 10910 -265
rect 10945 -295 10995 -265
rect 11030 -295 11080 -265
rect 11115 -295 11165 -265
rect 11200 -295 11250 -265
rect 11285 -295 11335 -265
rect 11370 -295 11420 -265
rect 11455 -295 11505 -265
rect 11540 -295 11590 -265
rect 11625 -295 11675 -265
rect 11710 -295 11760 -265
rect 11795 -295 11845 -265
rect 11880 -295 11930 -265
rect 11965 -295 12015 -265
rect 12050 -295 12100 -265
rect 12135 -295 12185 -265
rect 12220 -295 12270 -265
rect 12305 -295 12355 -265
rect 12390 -295 12440 -265
rect 12475 -295 12525 -265
rect 12560 -295 12610 -265
rect 12645 -295 12695 -265
rect 12730 -295 12780 -265
rect 12815 -295 12865 -265
rect 12900 -295 12950 -265
rect 12985 -295 13035 -265
rect 13070 -295 13120 -265
rect 13155 -295 13205 -265
rect 13240 -295 13290 -265
rect 13325 -295 13375 -265
rect 13410 -295 13460 -265
rect 13495 -295 13545 -265
rect 13580 -295 13630 -265
rect 13665 -295 13715 -265
rect 13750 -295 13800 -265
rect 13835 -295 13885 -265
rect 13920 -295 13970 -265
rect 14005 -295 14055 -265
rect 14090 -295 14140 -265
rect 14175 -295 14225 -265
rect 14260 -295 14310 -265
rect 14345 -295 14395 -265
rect 14430 -295 14480 -265
rect 14515 -295 14565 -265
rect 14600 -295 14650 -265
rect 14685 -295 14735 -265
rect 14770 -295 14820 -265
rect 14855 -295 14905 -265
rect 14940 -295 14990 -265
rect 15025 -295 15075 -265
rect 15110 -295 15160 -265
rect 15195 -295 15245 -265
rect 15280 -295 15330 -265
rect 15365 -295 15415 -265
rect 15450 -295 15500 -265
rect 15535 -295 15585 -265
rect 15620 -295 15670 -265
rect 15705 -295 15755 -265
rect 15790 -295 15840 -265
rect 15875 -295 15925 -265
rect 15960 -295 16010 -265
rect 16045 -295 16095 -265
rect 16130 -295 16180 -265
rect 16215 -295 16265 -265
rect 16300 -295 16350 -265
rect 16385 -295 16435 -265
rect 16470 -295 16520 -265
rect 16555 -295 16605 -265
rect 16640 -295 16690 -265
rect 16725 -295 16775 -265
rect 16810 -295 16860 -265
rect 16895 -295 16945 -265
rect 16980 -295 17030 -265
rect 17065 -295 17115 -265
rect 17150 -295 17200 -265
rect 17235 -295 17285 -265
rect 17320 -295 17370 -265
rect 17405 -295 17455 -265
rect 17490 -295 17540 -265
rect 17575 -295 17625 -265
rect 17660 -295 17710 -265
rect 17745 -295 17795 -265
rect 17830 -295 17880 -265
rect 17915 -295 17965 -265
rect 18000 -295 18050 -265
rect 18085 -295 18135 -265
rect 18170 -295 18220 -265
rect 18255 -295 18305 -265
rect 18340 -295 18390 -265
rect 18425 -295 18475 -265
rect 18510 -295 18560 -265
rect 18595 -295 18645 -265
rect 18680 -295 18730 -265
rect 18765 -295 18815 -265
rect 18850 -295 18900 -265
rect 18935 -295 18985 -265
rect 19020 -295 19070 -265
rect 19105 -295 19155 -265
rect 19190 -295 19240 -265
rect 19275 -295 19325 -265
rect 19360 -295 19410 -265
rect 19445 -295 19495 -265
rect 19530 -295 19580 -265
rect 19615 -295 19665 -265
rect 19700 -295 19750 -265
rect 19785 -295 19835 -265
rect 19870 -295 19920 -265
rect 19955 -295 20005 -265
rect 20040 -295 20090 -265
rect 20125 -295 20175 -265
rect 20210 -295 20260 -265
rect 20295 -295 20345 -265
rect 20380 -295 20430 -265
rect 20465 -295 20515 -265
rect 20550 -295 20600 -265
rect 20635 -295 20685 -265
rect 20720 -295 20770 -265
rect 20805 -295 20855 -265
rect 20890 -295 20940 -265
rect 20975 -295 21025 -265
rect 21060 -295 21110 -265
rect 21145 -295 21195 -265
rect 21230 -295 21280 -265
rect 21315 -295 21365 -265
rect 21400 -295 21450 -265
rect 21485 -295 21535 -265
rect 21570 -295 21620 -265
rect 21655 -295 21705 -265
rect 21740 -295 21790 -265
rect 21825 -295 21875 -265
rect 21910 -295 21960 -265
rect 21995 -295 22045 -265
rect 22080 -295 22130 -265
rect 22165 -295 22215 -265
rect 22250 -295 22300 -265
rect 22335 -295 22385 -265
rect 22420 -295 22470 -265
rect 22505 -295 22555 -265
rect 22590 -295 22640 -265
rect 22675 -295 22725 -265
rect 22760 -295 22810 -265
rect 22845 -295 22895 -265
rect 22930 -295 22980 -265
rect 23015 -295 23065 -265
rect 23100 -295 23150 -265
rect 23185 -295 23235 -265
rect 23270 -295 23320 -265
rect 23355 -295 23405 -265
rect 23440 -295 23490 -265
rect 23525 -295 23575 -265
rect 23610 -295 23660 -265
rect 23695 -295 23745 -265
rect 23780 -295 23830 -265
rect 23865 -295 23915 -265
rect 23950 -295 24000 -265
rect 24035 -295 24085 -265
rect 24120 -295 24170 -265
rect 24205 -295 24255 -265
rect 24290 -295 24340 -265
rect 24375 -295 24425 -265
rect 24460 -295 24510 -265
rect 24545 -295 24595 -265
rect 24630 -295 24680 -265
rect 24715 -295 24765 -265
rect 24800 -295 24850 -265
rect 24885 -295 24935 -265
rect 24970 -295 25020 -265
rect 25055 -295 25105 -265
rect 25140 -295 25190 -265
rect 25225 -295 25275 -265
rect 25310 -295 25360 -265
rect 25395 -295 25445 -265
rect 25480 -295 25530 -265
rect 25565 -295 25615 -265
rect 25650 -295 25700 -265
rect 25735 -295 25785 -265
rect 25820 -295 25870 -265
rect 25905 -295 25955 -265
rect 25990 -295 26040 -265
rect 26075 -295 26125 -265
rect 26160 -295 26210 -265
rect 26245 -295 26295 -265
rect 26330 -295 26380 -265
rect 26415 -295 26465 -265
rect 26500 -295 26550 -265
rect 26585 -295 26635 -265
rect 26670 -295 26720 -265
rect 26755 -295 26805 -265
rect 26840 -295 26890 -265
rect 26925 -295 26975 -265
rect 27010 -295 27060 -265
rect 27095 -295 27145 -265
rect 27180 -295 27230 -265
rect 27265 -295 27315 -265
rect 27350 -295 27400 -265
rect 27435 -295 27485 -265
rect 27520 -295 27570 -265
rect 27605 -295 27655 -265
rect 27690 -295 27740 -265
rect 27775 -295 27825 -265
rect 27860 -295 27910 -265
rect 27945 -295 27995 -265
rect 28030 -295 28080 -265
rect 28115 -295 28165 -265
rect 28200 -295 28250 -265
rect 28285 -295 28335 -265
rect 28370 -295 28420 -265
rect 28455 -295 28505 -265
rect 28540 -295 28590 -265
rect 28625 -295 28675 -265
rect 28710 -295 28760 -265
rect 28795 -295 28845 -265
rect 28880 -295 28930 -265
rect 28965 -295 29015 -265
rect 29050 -295 29100 -265
rect 29135 -295 29185 -265
rect 29220 -295 29270 -265
rect 29305 -295 29355 -265
rect 29390 -295 29440 -265
rect 29475 -295 29525 -265
rect 29560 -295 29610 -265
rect 29645 -295 29695 -265
rect 29730 -295 29780 -265
rect 29815 -295 29865 -265
rect 29900 -295 29950 -265
rect 29985 -295 30035 -265
rect 30070 -295 30120 -265
rect 30155 -295 30205 -265
rect 30240 -295 30290 -265
rect 30325 -295 30375 -265
rect 30410 -295 30460 -265
rect 30495 -295 30545 -265
rect 30580 -295 30630 -265
rect 30665 -295 30715 -265
rect 30750 -295 30800 -265
rect 30835 -295 30885 -265
rect 30920 -295 30970 -265
rect 31005 -295 31055 -265
rect 31090 -295 31140 -265
rect 31175 -295 31225 -265
rect 31260 -295 31310 -265
rect 31345 -295 31395 -265
rect 31430 -295 31480 -265
rect 31515 -295 31565 -265
rect 31600 -295 31650 -265
rect 31685 -295 31735 -265
rect 31770 -295 31820 -265
rect 31855 -295 31905 -265
rect 31940 -295 31990 -265
rect 32025 -295 32075 -265
rect 32110 -295 32160 -265
rect 32195 -295 32245 -265
rect 32280 -295 32330 -265
rect 32365 -295 32415 -265
rect 32450 -295 32500 -265
rect 32535 -295 32585 -265
rect 32620 -295 32670 -265
rect 32705 -295 32755 -265
rect 32790 -295 32840 -265
rect 32875 -295 32925 -265
rect 32960 -295 33010 -265
rect 33045 -295 33095 -265
rect 33130 -295 33180 -265
rect 33215 -295 33265 -265
rect 33300 -295 33350 -265
rect 33385 -295 33435 -265
rect 33470 -295 33520 -265
rect 33555 -295 33605 -265
rect 33640 -295 33690 -265
rect 33725 -295 33775 -265
rect 33810 -295 33860 -265
rect 33895 -295 33945 -265
rect 33980 -295 34030 -265
rect 34065 -295 34115 -265
rect 34150 -295 34200 -265
rect 34235 -295 34285 -265
rect 34320 -295 34370 -265
rect 34405 -295 34455 -265
rect 34490 -295 34540 -265
rect 34575 -295 34625 -265
rect 34660 -295 34710 -265
rect 34745 -295 34795 -265
rect 34830 -295 34880 -265
rect 34915 -295 34965 -265
rect 35000 -295 35050 -265
rect 35085 -295 35135 -265
rect 35170 -295 35220 -265
rect 35255 -295 35305 -265
rect 35340 -295 35390 -265
rect 35425 -295 35475 -265
rect 35510 -295 35560 -265
rect 35595 -295 35645 -265
rect 35680 -295 35730 -265
rect 35765 -295 35815 -265
rect 35850 -295 35900 -265
rect 35935 -295 35985 -265
rect 36020 -295 36070 -265
rect 36105 -295 36155 -265
rect 36190 -295 36240 -265
rect 36275 -295 36325 -265
rect 36360 -295 36410 -265
rect 36445 -295 36495 -265
rect 36530 -295 36580 -265
rect 36615 -295 36665 -265
rect 36700 -295 36750 -265
rect 36785 -295 36835 -265
rect 36870 -295 36920 -265
rect 36955 -295 37005 -265
rect 37040 -295 37090 -265
rect 37125 -295 37175 -265
rect 37210 -295 37260 -265
rect 37295 -295 37345 -265
rect 37380 -295 37430 -265
rect 37465 -295 37515 -265
rect 37550 -295 37600 -265
rect 37635 -295 37685 -265
rect 37720 -295 37770 -265
rect 37805 -295 37855 -265
rect 37890 -295 37940 -265
rect 37975 -295 38025 -265
rect 38060 -295 38110 -265
rect 38145 -295 38195 -265
rect 38230 -295 38280 -265
rect 38315 -295 38365 -265
rect 38400 -295 38450 -265
rect 38485 -295 38535 -265
rect 38570 -295 38620 -265
rect 38655 -295 38705 -265
rect 38740 -295 38790 -265
rect 38825 -295 38875 -265
rect 38910 -295 38960 -265
rect 38995 -295 39045 -265
rect 39080 -295 39130 -265
rect 39165 -295 39215 -265
rect 39250 -295 39300 -265
rect 39335 -295 39385 -265
rect 39420 -295 39470 -265
rect 39505 -295 39555 -265
rect 39590 -295 39640 -265
rect 39675 -295 39725 -265
rect 39760 -295 39810 -265
rect 39845 -295 39895 -265
rect 39930 -295 39980 -265
rect 40015 -295 40065 -265
rect 40100 -295 40150 -265
rect 40185 -295 40235 -265
rect 40270 -295 40320 -265
rect 40355 -295 40405 -265
rect 40440 -295 40490 -265
rect 40525 -295 40575 -265
rect 40610 -295 40660 -265
rect 40695 -295 40745 -265
rect 40780 -295 40830 -265
rect 40865 -295 40915 -265
rect 40950 -295 41000 -265
rect 41035 -295 41085 -265
rect 41120 -295 41170 -265
rect 41205 -295 41255 -265
rect 41290 -295 41340 -265
rect 41375 -295 41425 -265
rect 41460 -295 41510 -265
rect 41545 -295 41595 -265
rect 41630 -295 41680 -265
rect 41715 -295 41765 -265
rect 41800 -295 41850 -265
rect 41885 -295 41935 -265
rect 41970 -295 42020 -265
rect 42055 -295 42105 -265
rect 42140 -295 42190 -265
rect 42225 -295 42275 -265
rect 42310 -295 42360 -265
rect 42395 -295 42445 -265
rect 42480 -295 42530 -265
rect 42565 -295 42615 -265
rect 42650 -295 42700 -265
rect 42735 -295 42785 -265
rect 42820 -295 42870 -265
rect 42905 -295 42955 -265
rect 42990 -295 43040 -265
rect 43075 -295 43125 -265
rect 43160 -295 43210 -265
rect 43245 -295 43295 -265
rect 43330 -295 43380 -265
rect 43415 -295 43465 -265
rect 43500 -295 43550 -265
rect 43585 -295 43625 -265
rect 105 -305 43625 -295
rect 65 -335 115 -325
rect 235 -335 285 -325
rect 405 -335 455 -325
rect 575 -335 625 -325
rect 745 -335 795 -325
rect 915 -335 965 -325
rect 1085 -335 1135 -325
rect 1255 -335 1305 -325
rect 1425 -335 1475 -325
rect 1595 -335 1645 -325
rect 1765 -335 1815 -325
rect 1935 -335 1985 -325
rect 2105 -335 2155 -325
rect 2275 -335 2325 -325
rect 2445 -335 2495 -325
rect 2615 -335 2665 -325
rect 2785 -335 2835 -325
rect 2955 -335 3005 -325
rect 3125 -335 3175 -325
rect 3295 -335 3345 -325
rect 3465 -335 3515 -325
rect 3635 -335 3685 -325
rect 3805 -335 3855 -325
rect 3975 -335 4025 -325
rect 4145 -335 4195 -325
rect 4315 -335 4365 -325
rect 4485 -335 4535 -325
rect 4655 -335 4705 -325
rect 4825 -335 4875 -325
rect 4995 -335 5045 -325
rect 5165 -335 5215 -325
rect 5335 -335 5385 -325
rect 5505 -335 5555 -325
rect 5675 -335 5725 -325
rect 5845 -335 5895 -325
rect 6015 -335 6065 -325
rect 6185 -335 6235 -325
rect 6355 -335 6405 -325
rect 6525 -335 6575 -325
rect 6695 -335 6745 -325
rect 6865 -335 6915 -325
rect 7035 -335 7085 -325
rect 7205 -335 7255 -325
rect 7375 -335 7425 -325
rect 7545 -335 7595 -325
rect 7715 -335 7765 -325
rect 7885 -335 7935 -325
rect 8055 -335 8105 -325
rect 8225 -335 8275 -325
rect 8395 -335 8445 -325
rect 8565 -335 8615 -325
rect 8735 -335 8785 -325
rect 8905 -335 8955 -325
rect 9075 -335 9125 -325
rect 9245 -335 9295 -325
rect 9415 -335 9465 -325
rect 9585 -335 9635 -325
rect 9755 -335 9805 -325
rect 9925 -335 9975 -325
rect 10095 -335 10145 -325
rect 10265 -335 10315 -325
rect 10435 -335 10485 -325
rect 10605 -335 10655 -325
rect 10775 -335 10825 -325
rect 10945 -335 10995 -325
rect 11115 -335 11165 -325
rect 11285 -335 11335 -325
rect 11455 -335 11505 -325
rect 11625 -335 11675 -325
rect 11795 -335 11845 -325
rect 11965 -335 12015 -325
rect 12135 -335 12185 -325
rect 12305 -335 12355 -325
rect 12475 -335 12525 -325
rect 12645 -335 12695 -325
rect 12815 -335 12865 -325
rect 12985 -335 13035 -325
rect 13155 -335 13205 -325
rect 13325 -335 13375 -325
rect 13495 -335 13545 -325
rect 13665 -335 13715 -325
rect 13835 -335 13885 -325
rect 14005 -335 14055 -325
rect 14175 -335 14225 -325
rect 14345 -335 14395 -325
rect 14515 -335 14565 -325
rect 14685 -335 14735 -325
rect 14855 -335 14905 -325
rect 15025 -335 15075 -325
rect 15195 -335 15245 -325
rect 15365 -335 15415 -325
rect 15535 -335 15585 -325
rect 15705 -335 15755 -325
rect 15875 -335 15925 -325
rect 16045 -335 16095 -325
rect 16215 -335 16265 -325
rect 16385 -335 16435 -325
rect 16555 -335 16605 -325
rect 16725 -335 16775 -325
rect 16895 -335 16945 -325
rect 17065 -335 17115 -325
rect 17235 -335 17285 -325
rect 17405 -335 17455 -325
rect 17575 -335 17625 -325
rect 17745 -335 17795 -325
rect 17915 -335 17965 -325
rect 18085 -335 18135 -325
rect 18255 -335 18305 -325
rect 18425 -335 18475 -325
rect 18595 -335 18645 -325
rect 18765 -335 18815 -325
rect 18935 -335 18985 -325
rect 19105 -335 19155 -325
rect 19275 -335 19325 -325
rect 19445 -335 19495 -325
rect 19615 -335 19665 -325
rect 19785 -335 19835 -325
rect 19955 -335 20005 -325
rect 20125 -335 20175 -325
rect 20295 -335 20345 -325
rect 20465 -335 20515 -325
rect 20635 -335 20685 -325
rect 20805 -335 20855 -325
rect 20975 -335 21025 -325
rect 21145 -335 21195 -325
rect 21315 -335 21365 -325
rect 21485 -335 21535 -325
rect 21655 -335 21705 -325
rect 21825 -335 21875 -325
rect 21995 -335 22045 -325
rect 22165 -335 22215 -325
rect 22335 -335 22385 -325
rect 22505 -335 22555 -325
rect 22675 -335 22725 -325
rect 22845 -335 22895 -325
rect 23015 -335 23065 -325
rect 23185 -335 23235 -325
rect 23355 -335 23405 -325
rect 23525 -335 23575 -325
rect 23695 -335 23745 -325
rect 23865 -335 23915 -325
rect 24035 -335 24085 -325
rect 24205 -335 24255 -325
rect 24375 -335 24425 -325
rect 24545 -335 24595 -325
rect 24715 -335 24765 -325
rect 24885 -335 24935 -325
rect 25055 -335 25105 -325
rect 25225 -335 25275 -325
rect 25395 -335 25445 -325
rect 25565 -335 25615 -325
rect 25735 -335 25785 -325
rect 25905 -335 25955 -325
rect 26075 -335 26125 -325
rect 26245 -335 26295 -325
rect 26415 -335 26465 -325
rect 26585 -335 26635 -325
rect 26755 -335 26805 -325
rect 26925 -335 26975 -325
rect 27095 -335 27145 -325
rect 27265 -335 27315 -325
rect 27435 -335 27485 -325
rect 27605 -335 27655 -325
rect 27775 -335 27825 -325
rect 27945 -335 27995 -325
rect 28115 -335 28165 -325
rect 28285 -335 28335 -325
rect 28455 -335 28505 -325
rect 28625 -335 28675 -325
rect 28795 -335 28845 -325
rect 28965 -335 29015 -325
rect 29135 -335 29185 -325
rect 29305 -335 29355 -325
rect 29475 -335 29525 -325
rect 29645 -335 29695 -325
rect 29815 -335 29865 -325
rect 29985 -335 30035 -325
rect 30155 -335 30205 -325
rect 30325 -335 30375 -325
rect 30495 -335 30545 -325
rect 30665 -335 30715 -325
rect 30835 -335 30885 -325
rect 31005 -335 31055 -325
rect 31175 -335 31225 -325
rect 31345 -335 31395 -325
rect 31515 -335 31565 -325
rect 31685 -335 31735 -325
rect 31855 -335 31905 -325
rect 32025 -335 32075 -325
rect 32195 -335 32245 -325
rect 32365 -335 32415 -325
rect 32535 -335 32585 -325
rect 32705 -335 32755 -325
rect 32875 -335 32925 -325
rect 33045 -335 33095 -325
rect 33215 -335 33265 -325
rect 33385 -335 33435 -325
rect 33555 -335 33605 -325
rect 33725 -335 33775 -325
rect 33895 -335 33945 -325
rect 34065 -335 34115 -325
rect 34235 -335 34285 -325
rect 34405 -335 34455 -325
rect 34575 -335 34625 -325
rect 34745 -335 34795 -325
rect 34915 -335 34965 -325
rect 35085 -335 35135 -325
rect 35255 -335 35305 -325
rect 35425 -335 35475 -325
rect 35595 -335 35645 -325
rect 35765 -335 35815 -325
rect 35935 -335 35985 -325
rect 36105 -335 36155 -325
rect 36275 -335 36325 -325
rect 36445 -335 36495 -325
rect 36615 -335 36665 -325
rect 36785 -335 36835 -325
rect 36955 -335 37005 -325
rect 37125 -335 37175 -325
rect 37295 -335 37345 -325
rect 37465 -335 37515 -325
rect 37635 -335 37685 -325
rect 37805 -335 37855 -325
rect 37975 -335 38025 -325
rect 38145 -335 38195 -325
rect 38315 -335 38365 -325
rect 38485 -335 38535 -325
rect 38655 -335 38705 -325
rect 38825 -335 38875 -325
rect 38995 -335 39045 -325
rect 39165 -335 39215 -325
rect 39335 -335 39385 -325
rect 39505 -335 39555 -325
rect 39675 -335 39725 -325
rect 39845 -335 39895 -325
rect 40015 -335 40065 -325
rect 40185 -335 40235 -325
rect 40355 -335 40405 -325
rect 40525 -335 40575 -325
rect 40695 -335 40745 -325
rect 40865 -335 40915 -325
rect 41035 -335 41085 -325
rect 41205 -335 41255 -325
rect 41375 -335 41425 -325
rect 41545 -335 41595 -325
rect 41715 -335 41765 -325
rect 41885 -335 41935 -325
rect 42055 -335 42105 -325
rect 42225 -335 42275 -325
rect 42395 -335 42445 -325
rect 42565 -335 42615 -325
rect 42735 -335 42785 -325
rect 42905 -335 42955 -325
rect 43075 -335 43125 -325
rect 43245 -335 43295 -325
rect 43415 -335 43465 -325
rect 43585 -335 43635 -325
rect 65 -365 75 -335
rect 105 -365 245 -335
rect 275 -365 415 -335
rect 445 -365 585 -335
rect 615 -365 755 -335
rect 785 -365 925 -335
rect 955 -365 1095 -335
rect 1125 -365 1265 -335
rect 1295 -365 1435 -335
rect 1465 -365 1605 -335
rect 1635 -365 1775 -335
rect 1805 -365 1945 -335
rect 1975 -365 2115 -335
rect 2145 -365 2285 -335
rect 2315 -365 2455 -335
rect 2485 -365 2625 -335
rect 2655 -365 2795 -335
rect 2825 -365 2965 -335
rect 2995 -365 3135 -335
rect 3165 -365 3305 -335
rect 3335 -365 3475 -335
rect 3505 -365 3645 -335
rect 3675 -365 3815 -335
rect 3845 -365 3985 -335
rect 4015 -365 4155 -335
rect 4185 -365 4325 -335
rect 4355 -365 4495 -335
rect 4525 -365 4665 -335
rect 4695 -365 4835 -335
rect 4865 -365 5005 -335
rect 5035 -365 5175 -335
rect 5205 -365 5345 -335
rect 5375 -365 5515 -335
rect 5545 -365 5685 -335
rect 5715 -365 5855 -335
rect 5885 -365 6025 -335
rect 6055 -365 6195 -335
rect 6225 -365 6365 -335
rect 6395 -365 6535 -335
rect 6565 -365 6705 -335
rect 6735 -365 6875 -335
rect 6905 -365 7045 -335
rect 7075 -365 7215 -335
rect 7245 -365 7385 -335
rect 7415 -365 7555 -335
rect 7585 -365 7725 -335
rect 7755 -365 7895 -335
rect 7925 -365 8065 -335
rect 8095 -365 8235 -335
rect 8265 -365 8405 -335
rect 8435 -365 8575 -335
rect 8605 -365 8745 -335
rect 8775 -365 8915 -335
rect 8945 -365 9085 -335
rect 9115 -365 9255 -335
rect 9285 -365 9425 -335
rect 9455 -365 9595 -335
rect 9625 -365 9765 -335
rect 9795 -365 9935 -335
rect 9965 -365 10105 -335
rect 10135 -365 10275 -335
rect 10305 -365 10445 -335
rect 10475 -365 10615 -335
rect 10645 -365 10785 -335
rect 10815 -365 10955 -335
rect 10985 -365 11125 -335
rect 11155 -365 11295 -335
rect 11325 -365 11465 -335
rect 11495 -365 11635 -335
rect 11665 -365 11805 -335
rect 11835 -365 11975 -335
rect 12005 -365 12145 -335
rect 12175 -365 12315 -335
rect 12345 -365 12485 -335
rect 12515 -365 12655 -335
rect 12685 -365 12825 -335
rect 12855 -365 12995 -335
rect 13025 -365 13165 -335
rect 13195 -365 13335 -335
rect 13365 -365 13505 -335
rect 13535 -365 13675 -335
rect 13705 -365 13845 -335
rect 13875 -365 14015 -335
rect 14045 -365 14185 -335
rect 14215 -365 14355 -335
rect 14385 -365 14525 -335
rect 14555 -365 14695 -335
rect 14725 -365 14865 -335
rect 14895 -365 15035 -335
rect 15065 -365 15205 -335
rect 15235 -365 15375 -335
rect 15405 -365 15545 -335
rect 15575 -365 15715 -335
rect 15745 -365 15885 -335
rect 15915 -365 16055 -335
rect 16085 -365 16225 -335
rect 16255 -365 16395 -335
rect 16425 -365 16565 -335
rect 16595 -365 16735 -335
rect 16765 -365 16905 -335
rect 16935 -365 17075 -335
rect 17105 -365 17245 -335
rect 17275 -365 17415 -335
rect 17445 -365 17585 -335
rect 17615 -365 17755 -335
rect 17785 -365 17925 -335
rect 17955 -365 18095 -335
rect 18125 -365 18265 -335
rect 18295 -365 18435 -335
rect 18465 -365 18605 -335
rect 18635 -365 18775 -335
rect 18805 -365 18945 -335
rect 18975 -365 19115 -335
rect 19145 -365 19285 -335
rect 19315 -365 19455 -335
rect 19485 -365 19625 -335
rect 19655 -365 19795 -335
rect 19825 -365 19965 -335
rect 19995 -365 20135 -335
rect 20165 -365 20305 -335
rect 20335 -365 20475 -335
rect 20505 -365 20645 -335
rect 20675 -365 20815 -335
rect 20845 -365 20985 -335
rect 21015 -365 21155 -335
rect 21185 -365 21325 -335
rect 21355 -365 21495 -335
rect 21525 -365 21665 -335
rect 21695 -365 21835 -335
rect 21865 -365 22005 -335
rect 22035 -365 22175 -335
rect 22205 -365 22345 -335
rect 22375 -365 22515 -335
rect 22545 -365 22685 -335
rect 22715 -365 22855 -335
rect 22885 -365 23025 -335
rect 23055 -365 23195 -335
rect 23225 -365 23365 -335
rect 23395 -365 23535 -335
rect 23565 -365 23705 -335
rect 23735 -365 23875 -335
rect 23905 -365 24045 -335
rect 24075 -365 24215 -335
rect 24245 -365 24385 -335
rect 24415 -365 24555 -335
rect 24585 -365 24725 -335
rect 24755 -365 24895 -335
rect 24925 -365 25065 -335
rect 25095 -365 25235 -335
rect 25265 -365 25405 -335
rect 25435 -365 25575 -335
rect 25605 -365 25745 -335
rect 25775 -365 25915 -335
rect 25945 -365 26085 -335
rect 26115 -365 26255 -335
rect 26285 -365 26425 -335
rect 26455 -365 26595 -335
rect 26625 -365 26765 -335
rect 26795 -365 26935 -335
rect 26965 -365 27105 -335
rect 27135 -365 27275 -335
rect 27305 -365 27445 -335
rect 27475 -365 27615 -335
rect 27645 -365 27785 -335
rect 27815 -365 27955 -335
rect 27985 -365 28125 -335
rect 28155 -365 28295 -335
rect 28325 -365 28465 -335
rect 28495 -365 28635 -335
rect 28665 -365 28805 -335
rect 28835 -365 28975 -335
rect 29005 -365 29145 -335
rect 29175 -365 29315 -335
rect 29345 -365 29485 -335
rect 29515 -365 29655 -335
rect 29685 -365 29825 -335
rect 29855 -365 29995 -335
rect 30025 -365 30165 -335
rect 30195 -365 30335 -335
rect 30365 -365 30505 -335
rect 30535 -365 30675 -335
rect 30705 -365 30845 -335
rect 30875 -365 31015 -335
rect 31045 -365 31185 -335
rect 31215 -365 31355 -335
rect 31385 -365 31525 -335
rect 31555 -365 31695 -335
rect 31725 -365 31865 -335
rect 31895 -365 32035 -335
rect 32065 -365 32205 -335
rect 32235 -365 32375 -335
rect 32405 -365 32545 -335
rect 32575 -365 32715 -335
rect 32745 -365 32885 -335
rect 32915 -365 33055 -335
rect 33085 -365 33225 -335
rect 33255 -365 33395 -335
rect 33425 -365 33565 -335
rect 33595 -365 33735 -335
rect 33765 -365 33905 -335
rect 33935 -365 34075 -335
rect 34105 -365 34245 -335
rect 34275 -365 34415 -335
rect 34445 -365 34585 -335
rect 34615 -365 34755 -335
rect 34785 -365 34925 -335
rect 34955 -365 35095 -335
rect 35125 -365 35265 -335
rect 35295 -365 35435 -335
rect 35465 -365 35605 -335
rect 35635 -365 35775 -335
rect 35805 -365 35945 -335
rect 35975 -365 36115 -335
rect 36145 -365 36285 -335
rect 36315 -365 36455 -335
rect 36485 -365 36625 -335
rect 36655 -365 36795 -335
rect 36825 -365 36965 -335
rect 36995 -365 37135 -335
rect 37165 -365 37305 -335
rect 37335 -365 37475 -335
rect 37505 -365 37645 -335
rect 37675 -365 37815 -335
rect 37845 -365 37985 -335
rect 38015 -365 38155 -335
rect 38185 -365 38325 -335
rect 38355 -365 38495 -335
rect 38525 -365 38665 -335
rect 38695 -365 38835 -335
rect 38865 -365 39005 -335
rect 39035 -365 39175 -335
rect 39205 -365 39345 -335
rect 39375 -365 39515 -335
rect 39545 -365 39685 -335
rect 39715 -365 39855 -335
rect 39885 -365 40025 -335
rect 40055 -365 40195 -335
rect 40225 -365 40365 -335
rect 40395 -365 40535 -335
rect 40565 -365 40705 -335
rect 40735 -365 40875 -335
rect 40905 -365 41045 -335
rect 41075 -365 41215 -335
rect 41245 -365 41385 -335
rect 41415 -365 41555 -335
rect 41585 -365 41725 -335
rect 41755 -365 41895 -335
rect 41925 -365 42065 -335
rect 42095 -365 42235 -335
rect 42265 -365 42405 -335
rect 42435 -365 42575 -335
rect 42605 -365 42745 -335
rect 42775 -365 42915 -335
rect 42945 -365 43085 -335
rect 43115 -365 43255 -335
rect 43285 -365 43425 -335
rect 43455 -365 43595 -335
rect 43625 -365 43645 -335
rect 65 -375 115 -365
rect 235 -375 285 -365
rect 405 -375 455 -365
rect 575 -375 625 -365
rect 745 -375 795 -365
rect 915 -375 965 -365
rect 1085 -375 1135 -365
rect 1255 -375 1305 -365
rect 1425 -375 1475 -365
rect 1595 -375 1645 -365
rect 1765 -375 1815 -365
rect 1935 -375 1985 -365
rect 2105 -375 2155 -365
rect 2275 -375 2325 -365
rect 2445 -375 2495 -365
rect 2615 -375 2665 -365
rect 2785 -375 2835 -365
rect 2955 -375 3005 -365
rect 3125 -375 3175 -365
rect 3295 -375 3345 -365
rect 3465 -375 3515 -365
rect 3635 -375 3685 -365
rect 3805 -375 3855 -365
rect 3975 -375 4025 -365
rect 4145 -375 4195 -365
rect 4315 -375 4365 -365
rect 4485 -375 4535 -365
rect 4655 -375 4705 -365
rect 4825 -375 4875 -365
rect 4995 -375 5045 -365
rect 5165 -375 5215 -365
rect 5335 -375 5385 -365
rect 5505 -375 5555 -365
rect 5675 -375 5725 -365
rect 5845 -375 5895 -365
rect 6015 -375 6065 -365
rect 6185 -375 6235 -365
rect 6355 -375 6405 -365
rect 6525 -375 6575 -365
rect 6695 -375 6745 -365
rect 6865 -375 6915 -365
rect 7035 -375 7085 -365
rect 7205 -375 7255 -365
rect 7375 -375 7425 -365
rect 7545 -375 7595 -365
rect 7715 -375 7765 -365
rect 7885 -375 7935 -365
rect 8055 -375 8105 -365
rect 8225 -375 8275 -365
rect 8395 -375 8445 -365
rect 8565 -375 8615 -365
rect 8735 -375 8785 -365
rect 8905 -375 8955 -365
rect 9075 -375 9125 -365
rect 9245 -375 9295 -365
rect 9415 -375 9465 -365
rect 9585 -375 9635 -365
rect 9755 -375 9805 -365
rect 9925 -375 9975 -365
rect 10095 -375 10145 -365
rect 10265 -375 10315 -365
rect 10435 -375 10485 -365
rect 10605 -375 10655 -365
rect 10775 -375 10825 -365
rect 10945 -375 10995 -365
rect 11115 -375 11165 -365
rect 11285 -375 11335 -365
rect 11455 -375 11505 -365
rect 11625 -375 11675 -365
rect 11795 -375 11845 -365
rect 11965 -375 12015 -365
rect 12135 -375 12185 -365
rect 12305 -375 12355 -365
rect 12475 -375 12525 -365
rect 12645 -375 12695 -365
rect 12815 -375 12865 -365
rect 12985 -375 13035 -365
rect 13155 -375 13205 -365
rect 13325 -375 13375 -365
rect 13495 -375 13545 -365
rect 13665 -375 13715 -365
rect 13835 -375 13885 -365
rect 14005 -375 14055 -365
rect 14175 -375 14225 -365
rect 14345 -375 14395 -365
rect 14515 -375 14565 -365
rect 14685 -375 14735 -365
rect 14855 -375 14905 -365
rect 15025 -375 15075 -365
rect 15195 -375 15245 -365
rect 15365 -375 15415 -365
rect 15535 -375 15585 -365
rect 15705 -375 15755 -365
rect 15875 -375 15925 -365
rect 16045 -375 16095 -365
rect 16215 -375 16265 -365
rect 16385 -375 16435 -365
rect 16555 -375 16605 -365
rect 16725 -375 16775 -365
rect 16895 -375 16945 -365
rect 17065 -375 17115 -365
rect 17235 -375 17285 -365
rect 17405 -375 17455 -365
rect 17575 -375 17625 -365
rect 17745 -375 17795 -365
rect 17915 -375 17965 -365
rect 18085 -375 18135 -365
rect 18255 -375 18305 -365
rect 18425 -375 18475 -365
rect 18595 -375 18645 -365
rect 18765 -375 18815 -365
rect 18935 -375 18985 -365
rect 19105 -375 19155 -365
rect 19275 -375 19325 -365
rect 19445 -375 19495 -365
rect 19615 -375 19665 -365
rect 19785 -375 19835 -365
rect 19955 -375 20005 -365
rect 20125 -375 20175 -365
rect 20295 -375 20345 -365
rect 20465 -375 20515 -365
rect 20635 -375 20685 -365
rect 20805 -375 20855 -365
rect 20975 -375 21025 -365
rect 21145 -375 21195 -365
rect 21315 -375 21365 -365
rect 21485 -375 21535 -365
rect 21655 -375 21705 -365
rect 21825 -375 21875 -365
rect 21995 -375 22045 -365
rect 22165 -375 22215 -365
rect 22335 -375 22385 -365
rect 22505 -375 22555 -365
rect 22675 -375 22725 -365
rect 22845 -375 22895 -365
rect 23015 -375 23065 -365
rect 23185 -375 23235 -365
rect 23355 -375 23405 -365
rect 23525 -375 23575 -365
rect 23695 -375 23745 -365
rect 23865 -375 23915 -365
rect 24035 -375 24085 -365
rect 24205 -375 24255 -365
rect 24375 -375 24425 -365
rect 24545 -375 24595 -365
rect 24715 -375 24765 -365
rect 24885 -375 24935 -365
rect 25055 -375 25105 -365
rect 25225 -375 25275 -365
rect 25395 -375 25445 -365
rect 25565 -375 25615 -365
rect 25735 -375 25785 -365
rect 25905 -375 25955 -365
rect 26075 -375 26125 -365
rect 26245 -375 26295 -365
rect 26415 -375 26465 -365
rect 26585 -375 26635 -365
rect 26755 -375 26805 -365
rect 26925 -375 26975 -365
rect 27095 -375 27145 -365
rect 27265 -375 27315 -365
rect 27435 -375 27485 -365
rect 27605 -375 27655 -365
rect 27775 -375 27825 -365
rect 27945 -375 27995 -365
rect 28115 -375 28165 -365
rect 28285 -375 28335 -365
rect 28455 -375 28505 -365
rect 28625 -375 28675 -365
rect 28795 -375 28845 -365
rect 28965 -375 29015 -365
rect 29135 -375 29185 -365
rect 29305 -375 29355 -365
rect 29475 -375 29525 -365
rect 29645 -375 29695 -365
rect 29815 -375 29865 -365
rect 29985 -375 30035 -365
rect 30155 -375 30205 -365
rect 30325 -375 30375 -365
rect 30495 -375 30545 -365
rect 30665 -375 30715 -365
rect 30835 -375 30885 -365
rect 31005 -375 31055 -365
rect 31175 -375 31225 -365
rect 31345 -375 31395 -365
rect 31515 -375 31565 -365
rect 31685 -375 31735 -365
rect 31855 -375 31905 -365
rect 32025 -375 32075 -365
rect 32195 -375 32245 -365
rect 32365 -375 32415 -365
rect 32535 -375 32585 -365
rect 32705 -375 32755 -365
rect 32875 -375 32925 -365
rect 33045 -375 33095 -365
rect 33215 -375 33265 -365
rect 33385 -375 33435 -365
rect 33555 -375 33605 -365
rect 33725 -375 33775 -365
rect 33895 -375 33945 -365
rect 34065 -375 34115 -365
rect 34235 -375 34285 -365
rect 34405 -375 34455 -365
rect 34575 -375 34625 -365
rect 34745 -375 34795 -365
rect 34915 -375 34965 -365
rect 35085 -375 35135 -365
rect 35255 -375 35305 -365
rect 35425 -375 35475 -365
rect 35595 -375 35645 -365
rect 35765 -375 35815 -365
rect 35935 -375 35985 -365
rect 36105 -375 36155 -365
rect 36275 -375 36325 -365
rect 36445 -375 36495 -365
rect 36615 -375 36665 -365
rect 36785 -375 36835 -365
rect 36955 -375 37005 -365
rect 37125 -375 37175 -365
rect 37295 -375 37345 -365
rect 37465 -375 37515 -365
rect 37635 -375 37685 -365
rect 37805 -375 37855 -365
rect 37975 -375 38025 -365
rect 38145 -375 38195 -365
rect 38315 -375 38365 -365
rect 38485 -375 38535 -365
rect 38655 -375 38705 -365
rect 38825 -375 38875 -365
rect 38995 -375 39045 -365
rect 39165 -375 39215 -365
rect 39335 -375 39385 -365
rect 39505 -375 39555 -365
rect 39675 -375 39725 -365
rect 39845 -375 39895 -365
rect 40015 -375 40065 -365
rect 40185 -375 40235 -365
rect 40355 -375 40405 -365
rect 40525 -375 40575 -365
rect 40695 -375 40745 -365
rect 40865 -375 40915 -365
rect 41035 -375 41085 -365
rect 41205 -375 41255 -365
rect 41375 -375 41425 -365
rect 41545 -375 41595 -365
rect 41715 -375 41765 -365
rect 41885 -375 41935 -365
rect 42055 -375 42105 -365
rect 42225 -375 42275 -365
rect 42395 -375 42445 -365
rect 42565 -375 42615 -365
rect 42735 -375 42785 -365
rect 42905 -375 42955 -365
rect 43075 -375 43125 -365
rect 43245 -375 43295 -365
rect 43415 -375 43465 -365
rect 43585 -375 43635 -365
rect 155 -440 195 -435
rect 155 -475 160 -440
rect 190 -475 195 -440
rect 155 -480 195 -475
rect 325 -440 365 -435
rect 325 -475 330 -440
rect 360 -475 365 -440
rect 325 -480 365 -475
rect 495 -440 535 -435
rect 495 -475 500 -440
rect 530 -475 535 -440
rect 495 -480 535 -475
rect 665 -440 705 -435
rect 665 -475 670 -440
rect 700 -475 705 -440
rect 665 -480 705 -475
rect 835 -440 875 -435
rect 835 -475 840 -440
rect 870 -475 875 -440
rect 835 -480 875 -475
rect 1005 -440 1045 -435
rect 1005 -475 1010 -440
rect 1040 -475 1045 -440
rect 1005 -480 1045 -475
rect 1175 -440 1215 -435
rect 1175 -475 1180 -440
rect 1210 -475 1215 -440
rect 1175 -480 1215 -475
rect 1345 -440 1385 -435
rect 1345 -475 1350 -440
rect 1380 -475 1385 -440
rect 1345 -480 1385 -475
rect 1515 -440 1555 -435
rect 1515 -475 1520 -440
rect 1550 -475 1555 -440
rect 1515 -480 1555 -475
rect 1685 -440 1725 -435
rect 1685 -475 1690 -440
rect 1720 -475 1725 -440
rect 1685 -480 1725 -475
rect 1855 -440 1895 -435
rect 1855 -475 1860 -440
rect 1890 -475 1895 -440
rect 1855 -480 1895 -475
rect 2025 -440 2065 -435
rect 2025 -475 2030 -440
rect 2060 -475 2065 -440
rect 2025 -480 2065 -475
rect 2195 -440 2235 -435
rect 2195 -475 2200 -440
rect 2230 -475 2235 -440
rect 2195 -480 2235 -475
rect 2365 -440 2405 -435
rect 2365 -475 2370 -440
rect 2400 -475 2405 -440
rect 2365 -480 2405 -475
rect 2535 -440 2575 -435
rect 2535 -475 2540 -440
rect 2570 -475 2575 -440
rect 2535 -480 2575 -475
rect 2705 -440 2745 -435
rect 2705 -475 2710 -440
rect 2740 -475 2745 -440
rect 2705 -480 2745 -475
rect 2875 -440 2915 -435
rect 2875 -475 2880 -440
rect 2910 -475 2915 -440
rect 2875 -480 2915 -475
rect 3045 -440 3085 -435
rect 3045 -475 3050 -440
rect 3080 -475 3085 -440
rect 3045 -480 3085 -475
rect 3215 -440 3255 -435
rect 3215 -475 3220 -440
rect 3250 -475 3255 -440
rect 3215 -480 3255 -475
rect 3385 -440 3425 -435
rect 3385 -475 3390 -440
rect 3420 -475 3425 -440
rect 3385 -480 3425 -475
rect 3555 -440 3595 -435
rect 3555 -475 3560 -440
rect 3590 -475 3595 -440
rect 3555 -480 3595 -475
rect 3725 -440 3765 -435
rect 3725 -475 3730 -440
rect 3760 -475 3765 -440
rect 3725 -480 3765 -475
rect 3895 -440 3935 -435
rect 3895 -475 3900 -440
rect 3930 -475 3935 -440
rect 3895 -480 3935 -475
rect 4065 -440 4105 -435
rect 4065 -475 4070 -440
rect 4100 -475 4105 -440
rect 4065 -480 4105 -475
rect 4235 -440 4275 -435
rect 4235 -475 4240 -440
rect 4270 -475 4275 -440
rect 4235 -480 4275 -475
rect 4405 -440 4445 -435
rect 4405 -475 4410 -440
rect 4440 -475 4445 -440
rect 4405 -480 4445 -475
rect 4575 -440 4615 -435
rect 4575 -475 4580 -440
rect 4610 -475 4615 -440
rect 4575 -480 4615 -475
rect 4745 -440 4785 -435
rect 4745 -475 4750 -440
rect 4780 -475 4785 -440
rect 4745 -480 4785 -475
rect 4915 -440 4955 -435
rect 4915 -475 4920 -440
rect 4950 -475 4955 -440
rect 4915 -480 4955 -475
rect 5085 -440 5125 -435
rect 5085 -475 5090 -440
rect 5120 -475 5125 -440
rect 5085 -480 5125 -475
rect 5255 -440 5295 -435
rect 5255 -475 5260 -440
rect 5290 -475 5295 -440
rect 5255 -480 5295 -475
rect 5425 -440 5465 -435
rect 5425 -475 5430 -440
rect 5460 -475 5465 -440
rect 5425 -480 5465 -475
rect 5595 -440 5635 -435
rect 5595 -475 5600 -440
rect 5630 -475 5635 -440
rect 5595 -480 5635 -475
rect 5765 -440 5805 -435
rect 5765 -475 5770 -440
rect 5800 -475 5805 -440
rect 5765 -480 5805 -475
rect 5935 -440 5975 -435
rect 5935 -475 5940 -440
rect 5970 -475 5975 -440
rect 5935 -480 5975 -475
rect 6105 -440 6145 -435
rect 6105 -475 6110 -440
rect 6140 -475 6145 -440
rect 6105 -480 6145 -475
rect 6275 -440 6315 -435
rect 6275 -475 6280 -440
rect 6310 -475 6315 -440
rect 6275 -480 6315 -475
rect 6445 -440 6485 -435
rect 6445 -475 6450 -440
rect 6480 -475 6485 -440
rect 6445 -480 6485 -475
rect 6615 -440 6655 -435
rect 6615 -475 6620 -440
rect 6650 -475 6655 -440
rect 6615 -480 6655 -475
rect 6785 -440 6825 -435
rect 6785 -475 6790 -440
rect 6820 -475 6825 -440
rect 6785 -480 6825 -475
rect 6955 -440 6995 -435
rect 6955 -475 6960 -440
rect 6990 -475 6995 -440
rect 6955 -480 6995 -475
rect 7125 -440 7165 -435
rect 7125 -475 7130 -440
rect 7160 -475 7165 -440
rect 7125 -480 7165 -475
rect 7295 -440 7335 -435
rect 7295 -475 7300 -440
rect 7330 -475 7335 -440
rect 7295 -480 7335 -475
rect 7465 -440 7505 -435
rect 7465 -475 7470 -440
rect 7500 -475 7505 -440
rect 7465 -480 7505 -475
rect 7635 -440 7675 -435
rect 7635 -475 7640 -440
rect 7670 -475 7675 -440
rect 7635 -480 7675 -475
rect 7805 -440 7845 -435
rect 7805 -475 7810 -440
rect 7840 -475 7845 -440
rect 7805 -480 7845 -475
rect 7975 -440 8015 -435
rect 7975 -475 7980 -440
rect 8010 -475 8015 -440
rect 7975 -480 8015 -475
rect 8145 -440 8185 -435
rect 8145 -475 8150 -440
rect 8180 -475 8185 -440
rect 8145 -480 8185 -475
rect 8315 -440 8355 -435
rect 8315 -475 8320 -440
rect 8350 -475 8355 -440
rect 8315 -480 8355 -475
rect 8485 -440 8525 -435
rect 8485 -475 8490 -440
rect 8520 -475 8525 -440
rect 8485 -480 8525 -475
rect 8655 -440 8695 -435
rect 8655 -475 8660 -440
rect 8690 -475 8695 -440
rect 8655 -480 8695 -475
rect 8825 -440 8865 -435
rect 8825 -475 8830 -440
rect 8860 -475 8865 -440
rect 8825 -480 8865 -475
rect 8995 -440 9035 -435
rect 8995 -475 9000 -440
rect 9030 -475 9035 -440
rect 8995 -480 9035 -475
rect 9165 -440 9205 -435
rect 9165 -475 9170 -440
rect 9200 -475 9205 -440
rect 9165 -480 9205 -475
rect 9335 -440 9375 -435
rect 9335 -475 9340 -440
rect 9370 -475 9375 -440
rect 9335 -480 9375 -475
rect 9505 -440 9545 -435
rect 9505 -475 9510 -440
rect 9540 -475 9545 -440
rect 9505 -480 9545 -475
rect 9675 -440 9715 -435
rect 9675 -475 9680 -440
rect 9710 -475 9715 -440
rect 9675 -480 9715 -475
rect 9845 -440 9885 -435
rect 9845 -475 9850 -440
rect 9880 -475 9885 -440
rect 9845 -480 9885 -475
rect 10015 -440 10055 -435
rect 10015 -475 10020 -440
rect 10050 -475 10055 -440
rect 10015 -480 10055 -475
rect 10185 -440 10225 -435
rect 10185 -475 10190 -440
rect 10220 -475 10225 -440
rect 10185 -480 10225 -475
rect 10355 -440 10395 -435
rect 10355 -475 10360 -440
rect 10390 -475 10395 -440
rect 10355 -480 10395 -475
rect 10525 -440 10565 -435
rect 10525 -475 10530 -440
rect 10560 -475 10565 -440
rect 10525 -480 10565 -475
rect 10695 -440 10735 -435
rect 10695 -475 10700 -440
rect 10730 -475 10735 -440
rect 10695 -480 10735 -475
rect 10865 -440 10905 -435
rect 10865 -475 10870 -440
rect 10900 -475 10905 -440
rect 10865 -480 10905 -475
rect 11035 -440 11075 -435
rect 11035 -475 11040 -440
rect 11070 -475 11075 -440
rect 11035 -480 11075 -475
rect 11205 -440 11245 -435
rect 11205 -475 11210 -440
rect 11240 -475 11245 -440
rect 11205 -480 11245 -475
rect 11375 -440 11415 -435
rect 11375 -475 11380 -440
rect 11410 -475 11415 -440
rect 11375 -480 11415 -475
rect 11545 -440 11585 -435
rect 11545 -475 11550 -440
rect 11580 -475 11585 -440
rect 11545 -480 11585 -475
rect 11715 -440 11755 -435
rect 11715 -475 11720 -440
rect 11750 -475 11755 -440
rect 11715 -480 11755 -475
rect 11885 -440 11925 -435
rect 11885 -475 11890 -440
rect 11920 -475 11925 -440
rect 11885 -480 11925 -475
rect 12055 -440 12095 -435
rect 12055 -475 12060 -440
rect 12090 -475 12095 -440
rect 12055 -480 12095 -475
rect 12225 -440 12265 -435
rect 12225 -475 12230 -440
rect 12260 -475 12265 -440
rect 12225 -480 12265 -475
rect 12395 -440 12435 -435
rect 12395 -475 12400 -440
rect 12430 -475 12435 -440
rect 12395 -480 12435 -475
rect 12565 -440 12605 -435
rect 12565 -475 12570 -440
rect 12600 -475 12605 -440
rect 12565 -480 12605 -475
rect 12735 -440 12775 -435
rect 12735 -475 12740 -440
rect 12770 -475 12775 -440
rect 12735 -480 12775 -475
rect 12905 -440 12945 -435
rect 12905 -475 12910 -440
rect 12940 -475 12945 -440
rect 12905 -480 12945 -475
rect 13075 -440 13115 -435
rect 13075 -475 13080 -440
rect 13110 -475 13115 -440
rect 13075 -480 13115 -475
rect 13245 -440 13285 -435
rect 13245 -475 13250 -440
rect 13280 -475 13285 -440
rect 13245 -480 13285 -475
rect 13415 -440 13455 -435
rect 13415 -475 13420 -440
rect 13450 -475 13455 -440
rect 13415 -480 13455 -475
rect 13585 -440 13625 -435
rect 13585 -475 13590 -440
rect 13620 -475 13625 -440
rect 13585 -480 13625 -475
rect 13755 -440 13795 -435
rect 13755 -475 13760 -440
rect 13790 -475 13795 -440
rect 13755 -480 13795 -475
rect 13925 -440 13965 -435
rect 13925 -475 13930 -440
rect 13960 -475 13965 -440
rect 13925 -480 13965 -475
rect 14095 -440 14135 -435
rect 14095 -475 14100 -440
rect 14130 -475 14135 -440
rect 14095 -480 14135 -475
rect 14265 -440 14305 -435
rect 14265 -475 14270 -440
rect 14300 -475 14305 -440
rect 14265 -480 14305 -475
rect 14435 -440 14475 -435
rect 14435 -475 14440 -440
rect 14470 -475 14475 -440
rect 14435 -480 14475 -475
rect 14605 -440 14645 -435
rect 14605 -475 14610 -440
rect 14640 -475 14645 -440
rect 14605 -480 14645 -475
rect 14775 -440 14815 -435
rect 14775 -475 14780 -440
rect 14810 -475 14815 -440
rect 14775 -480 14815 -475
rect 14945 -440 14985 -435
rect 14945 -475 14950 -440
rect 14980 -475 14985 -440
rect 14945 -480 14985 -475
rect 15115 -440 15155 -435
rect 15115 -475 15120 -440
rect 15150 -475 15155 -440
rect 15115 -480 15155 -475
rect 15285 -440 15325 -435
rect 15285 -475 15290 -440
rect 15320 -475 15325 -440
rect 15285 -480 15325 -475
rect 15455 -440 15495 -435
rect 15455 -475 15460 -440
rect 15490 -475 15495 -440
rect 15455 -480 15495 -475
rect 15625 -440 15665 -435
rect 15625 -475 15630 -440
rect 15660 -475 15665 -440
rect 15625 -480 15665 -475
rect 15795 -440 15835 -435
rect 15795 -475 15800 -440
rect 15830 -475 15835 -440
rect 15795 -480 15835 -475
rect 15965 -440 16005 -435
rect 15965 -475 15970 -440
rect 16000 -475 16005 -440
rect 15965 -480 16005 -475
rect 16135 -440 16175 -435
rect 16135 -475 16140 -440
rect 16170 -475 16175 -440
rect 16135 -480 16175 -475
rect 16305 -440 16345 -435
rect 16305 -475 16310 -440
rect 16340 -475 16345 -440
rect 16305 -480 16345 -475
rect 16475 -440 16515 -435
rect 16475 -475 16480 -440
rect 16510 -475 16515 -440
rect 16475 -480 16515 -475
rect 16645 -440 16685 -435
rect 16645 -475 16650 -440
rect 16680 -475 16685 -440
rect 16645 -480 16685 -475
rect 16815 -440 16855 -435
rect 16815 -475 16820 -440
rect 16850 -475 16855 -440
rect 16815 -480 16855 -475
rect 16985 -440 17025 -435
rect 16985 -475 16990 -440
rect 17020 -475 17025 -440
rect 16985 -480 17025 -475
rect 17155 -440 17195 -435
rect 17155 -475 17160 -440
rect 17190 -475 17195 -440
rect 17155 -480 17195 -475
rect 17325 -440 17365 -435
rect 17325 -475 17330 -440
rect 17360 -475 17365 -440
rect 17325 -480 17365 -475
rect 17495 -440 17535 -435
rect 17495 -475 17500 -440
rect 17530 -475 17535 -440
rect 17495 -480 17535 -475
rect 17665 -440 17705 -435
rect 17665 -475 17670 -440
rect 17700 -475 17705 -440
rect 17665 -480 17705 -475
rect 17835 -440 17875 -435
rect 17835 -475 17840 -440
rect 17870 -475 17875 -440
rect 17835 -480 17875 -475
rect 18005 -440 18045 -435
rect 18005 -475 18010 -440
rect 18040 -475 18045 -440
rect 18005 -480 18045 -475
rect 18175 -440 18215 -435
rect 18175 -475 18180 -440
rect 18210 -475 18215 -440
rect 18175 -480 18215 -475
rect 18345 -440 18385 -435
rect 18345 -475 18350 -440
rect 18380 -475 18385 -440
rect 18345 -480 18385 -475
rect 18515 -440 18555 -435
rect 18515 -475 18520 -440
rect 18550 -475 18555 -440
rect 18515 -480 18555 -475
rect 18685 -440 18725 -435
rect 18685 -475 18690 -440
rect 18720 -475 18725 -440
rect 18685 -480 18725 -475
rect 18855 -440 18895 -435
rect 18855 -475 18860 -440
rect 18890 -475 18895 -440
rect 18855 -480 18895 -475
rect 19025 -440 19065 -435
rect 19025 -475 19030 -440
rect 19060 -475 19065 -440
rect 19025 -480 19065 -475
rect 19195 -440 19235 -435
rect 19195 -475 19200 -440
rect 19230 -475 19235 -440
rect 19195 -480 19235 -475
rect 19365 -440 19405 -435
rect 19365 -475 19370 -440
rect 19400 -475 19405 -440
rect 19365 -480 19405 -475
rect 19535 -440 19575 -435
rect 19535 -475 19540 -440
rect 19570 -475 19575 -440
rect 19535 -480 19575 -475
rect 19705 -440 19745 -435
rect 19705 -475 19710 -440
rect 19740 -475 19745 -440
rect 19705 -480 19745 -475
rect 19875 -440 19915 -435
rect 19875 -475 19880 -440
rect 19910 -475 19915 -440
rect 19875 -480 19915 -475
rect 20045 -440 20085 -435
rect 20045 -475 20050 -440
rect 20080 -475 20085 -440
rect 20045 -480 20085 -475
rect 20215 -440 20255 -435
rect 20215 -475 20220 -440
rect 20250 -475 20255 -440
rect 20215 -480 20255 -475
rect 20385 -440 20425 -435
rect 20385 -475 20390 -440
rect 20420 -475 20425 -440
rect 20385 -480 20425 -475
rect 20555 -440 20595 -435
rect 20555 -475 20560 -440
rect 20590 -475 20595 -440
rect 20555 -480 20595 -475
rect 20725 -440 20765 -435
rect 20725 -475 20730 -440
rect 20760 -475 20765 -440
rect 20725 -480 20765 -475
rect 20895 -440 20935 -435
rect 20895 -475 20900 -440
rect 20930 -475 20935 -440
rect 20895 -480 20935 -475
rect 21065 -440 21105 -435
rect 21065 -475 21070 -440
rect 21100 -475 21105 -440
rect 21065 -480 21105 -475
rect 21235 -440 21275 -435
rect 21235 -475 21240 -440
rect 21270 -475 21275 -440
rect 21235 -480 21275 -475
rect 21405 -440 21445 -435
rect 21405 -475 21410 -440
rect 21440 -475 21445 -440
rect 21405 -480 21445 -475
rect 21575 -440 21615 -435
rect 21575 -475 21580 -440
rect 21610 -475 21615 -440
rect 21575 -480 21615 -475
rect 21745 -440 21785 -435
rect 21745 -475 21750 -440
rect 21780 -475 21785 -440
rect 21745 -480 21785 -475
rect 21915 -440 21955 -435
rect 21915 -475 21920 -440
rect 21950 -475 21955 -440
rect 21915 -480 21955 -475
rect 22085 -440 22125 -435
rect 22085 -475 22090 -440
rect 22120 -475 22125 -440
rect 22085 -480 22125 -475
rect 22255 -440 22295 -435
rect 22255 -475 22260 -440
rect 22290 -475 22295 -440
rect 22255 -480 22295 -475
rect 22425 -440 22465 -435
rect 22425 -475 22430 -440
rect 22460 -475 22465 -440
rect 22425 -480 22465 -475
rect 22595 -440 22635 -435
rect 22595 -475 22600 -440
rect 22630 -475 22635 -440
rect 22595 -480 22635 -475
rect 22765 -440 22805 -435
rect 22765 -475 22770 -440
rect 22800 -475 22805 -440
rect 22765 -480 22805 -475
rect 22935 -440 22975 -435
rect 22935 -475 22940 -440
rect 22970 -475 22975 -440
rect 22935 -480 22975 -475
rect 23105 -440 23145 -435
rect 23105 -475 23110 -440
rect 23140 -475 23145 -440
rect 23105 -480 23145 -475
rect 23275 -440 23315 -435
rect 23275 -475 23280 -440
rect 23310 -475 23315 -440
rect 23275 -480 23315 -475
rect 23445 -440 23485 -435
rect 23445 -475 23450 -440
rect 23480 -475 23485 -440
rect 23445 -480 23485 -475
rect 23615 -440 23655 -435
rect 23615 -475 23620 -440
rect 23650 -475 23655 -440
rect 23615 -480 23655 -475
rect 23785 -440 23825 -435
rect 23785 -475 23790 -440
rect 23820 -475 23825 -440
rect 23785 -480 23825 -475
rect 23955 -440 23995 -435
rect 23955 -475 23960 -440
rect 23990 -475 23995 -440
rect 23955 -480 23995 -475
rect 24125 -440 24165 -435
rect 24125 -475 24130 -440
rect 24160 -475 24165 -440
rect 24125 -480 24165 -475
rect 24295 -440 24335 -435
rect 24295 -475 24300 -440
rect 24330 -475 24335 -440
rect 24295 -480 24335 -475
rect 24465 -440 24505 -435
rect 24465 -475 24470 -440
rect 24500 -475 24505 -440
rect 24465 -480 24505 -475
rect 24635 -440 24675 -435
rect 24635 -475 24640 -440
rect 24670 -475 24675 -440
rect 24635 -480 24675 -475
rect 24805 -440 24845 -435
rect 24805 -475 24810 -440
rect 24840 -475 24845 -440
rect 24805 -480 24845 -475
rect 24975 -440 25015 -435
rect 24975 -475 24980 -440
rect 25010 -475 25015 -440
rect 24975 -480 25015 -475
rect 25145 -440 25185 -435
rect 25145 -475 25150 -440
rect 25180 -475 25185 -440
rect 25145 -480 25185 -475
rect 25315 -440 25355 -435
rect 25315 -475 25320 -440
rect 25350 -475 25355 -440
rect 25315 -480 25355 -475
rect 25485 -440 25525 -435
rect 25485 -475 25490 -440
rect 25520 -475 25525 -440
rect 25485 -480 25525 -475
rect 25655 -440 25695 -435
rect 25655 -475 25660 -440
rect 25690 -475 25695 -440
rect 25655 -480 25695 -475
rect 25825 -440 25865 -435
rect 25825 -475 25830 -440
rect 25860 -475 25865 -440
rect 25825 -480 25865 -475
rect 25995 -440 26035 -435
rect 25995 -475 26000 -440
rect 26030 -475 26035 -440
rect 25995 -480 26035 -475
rect 26165 -440 26205 -435
rect 26165 -475 26170 -440
rect 26200 -475 26205 -440
rect 26165 -480 26205 -475
rect 26335 -440 26375 -435
rect 26335 -475 26340 -440
rect 26370 -475 26375 -440
rect 26335 -480 26375 -475
rect 26505 -440 26545 -435
rect 26505 -475 26510 -440
rect 26540 -475 26545 -440
rect 26505 -480 26545 -475
rect 26675 -440 26715 -435
rect 26675 -475 26680 -440
rect 26710 -475 26715 -440
rect 26675 -480 26715 -475
rect 26845 -440 26885 -435
rect 26845 -475 26850 -440
rect 26880 -475 26885 -440
rect 26845 -480 26885 -475
rect 27015 -440 27055 -435
rect 27015 -475 27020 -440
rect 27050 -475 27055 -440
rect 27015 -480 27055 -475
rect 27185 -440 27225 -435
rect 27185 -475 27190 -440
rect 27220 -475 27225 -440
rect 27185 -480 27225 -475
rect 27355 -440 27395 -435
rect 27355 -475 27360 -440
rect 27390 -475 27395 -440
rect 27355 -480 27395 -475
rect 27525 -440 27565 -435
rect 27525 -475 27530 -440
rect 27560 -475 27565 -440
rect 27525 -480 27565 -475
rect 27695 -440 27735 -435
rect 27695 -475 27700 -440
rect 27730 -475 27735 -440
rect 27695 -480 27735 -475
rect 27865 -440 27905 -435
rect 27865 -475 27870 -440
rect 27900 -475 27905 -440
rect 27865 -480 27905 -475
rect 28035 -440 28075 -435
rect 28035 -475 28040 -440
rect 28070 -475 28075 -440
rect 28035 -480 28075 -475
rect 28205 -440 28245 -435
rect 28205 -475 28210 -440
rect 28240 -475 28245 -440
rect 28205 -480 28245 -475
rect 28375 -440 28415 -435
rect 28375 -475 28380 -440
rect 28410 -475 28415 -440
rect 28375 -480 28415 -475
rect 28545 -440 28585 -435
rect 28545 -475 28550 -440
rect 28580 -475 28585 -440
rect 28545 -480 28585 -475
rect 28715 -440 28755 -435
rect 28715 -475 28720 -440
rect 28750 -475 28755 -440
rect 28715 -480 28755 -475
rect 28885 -440 28925 -435
rect 28885 -475 28890 -440
rect 28920 -475 28925 -440
rect 28885 -480 28925 -475
rect 29055 -440 29095 -435
rect 29055 -475 29060 -440
rect 29090 -475 29095 -440
rect 29055 -480 29095 -475
rect 29225 -440 29265 -435
rect 29225 -475 29230 -440
rect 29260 -475 29265 -440
rect 29225 -480 29265 -475
rect 29395 -440 29435 -435
rect 29395 -475 29400 -440
rect 29430 -475 29435 -440
rect 29395 -480 29435 -475
rect 29565 -440 29605 -435
rect 29565 -475 29570 -440
rect 29600 -475 29605 -440
rect 29565 -480 29605 -475
rect 29735 -440 29775 -435
rect 29735 -475 29740 -440
rect 29770 -475 29775 -440
rect 29735 -480 29775 -475
rect 29905 -440 29945 -435
rect 29905 -475 29910 -440
rect 29940 -475 29945 -440
rect 29905 -480 29945 -475
rect 30075 -440 30115 -435
rect 30075 -475 30080 -440
rect 30110 -475 30115 -440
rect 30075 -480 30115 -475
rect 30245 -440 30285 -435
rect 30245 -475 30250 -440
rect 30280 -475 30285 -440
rect 30245 -480 30285 -475
rect 30415 -440 30455 -435
rect 30415 -475 30420 -440
rect 30450 -475 30455 -440
rect 30415 -480 30455 -475
rect 30585 -440 30625 -435
rect 30585 -475 30590 -440
rect 30620 -475 30625 -440
rect 30585 -480 30625 -475
rect 30755 -440 30795 -435
rect 30755 -475 30760 -440
rect 30790 -475 30795 -440
rect 30755 -480 30795 -475
rect 30925 -440 30965 -435
rect 30925 -475 30930 -440
rect 30960 -475 30965 -440
rect 30925 -480 30965 -475
rect 31095 -440 31135 -435
rect 31095 -475 31100 -440
rect 31130 -475 31135 -440
rect 31095 -480 31135 -475
rect 31265 -440 31305 -435
rect 31265 -475 31270 -440
rect 31300 -475 31305 -440
rect 31265 -480 31305 -475
rect 31435 -440 31475 -435
rect 31435 -475 31440 -440
rect 31470 -475 31475 -440
rect 31435 -480 31475 -475
rect 31605 -440 31645 -435
rect 31605 -475 31610 -440
rect 31640 -475 31645 -440
rect 31605 -480 31645 -475
rect 31775 -440 31815 -435
rect 31775 -475 31780 -440
rect 31810 -475 31815 -440
rect 31775 -480 31815 -475
rect 31945 -440 31985 -435
rect 31945 -475 31950 -440
rect 31980 -475 31985 -440
rect 31945 -480 31985 -475
rect 32115 -440 32155 -435
rect 32115 -475 32120 -440
rect 32150 -475 32155 -440
rect 32115 -480 32155 -475
rect 32285 -440 32325 -435
rect 32285 -475 32290 -440
rect 32320 -475 32325 -440
rect 32285 -480 32325 -475
rect 32455 -440 32495 -435
rect 32455 -475 32460 -440
rect 32490 -475 32495 -440
rect 32455 -480 32495 -475
rect 32625 -440 32665 -435
rect 32625 -475 32630 -440
rect 32660 -475 32665 -440
rect 32625 -480 32665 -475
rect 32795 -440 32835 -435
rect 32795 -475 32800 -440
rect 32830 -475 32835 -440
rect 32795 -480 32835 -475
rect 32965 -440 33005 -435
rect 32965 -475 32970 -440
rect 33000 -475 33005 -440
rect 32965 -480 33005 -475
rect 33135 -440 33175 -435
rect 33135 -475 33140 -440
rect 33170 -475 33175 -440
rect 33135 -480 33175 -475
rect 33305 -440 33345 -435
rect 33305 -475 33310 -440
rect 33340 -475 33345 -440
rect 33305 -480 33345 -475
rect 33475 -440 33515 -435
rect 33475 -475 33480 -440
rect 33510 -475 33515 -440
rect 33475 -480 33515 -475
rect 33645 -440 33685 -435
rect 33645 -475 33650 -440
rect 33680 -475 33685 -440
rect 33645 -480 33685 -475
rect 33815 -440 33855 -435
rect 33815 -475 33820 -440
rect 33850 -475 33855 -440
rect 33815 -480 33855 -475
rect 33985 -440 34025 -435
rect 33985 -475 33990 -440
rect 34020 -475 34025 -440
rect 33985 -480 34025 -475
rect 34155 -440 34195 -435
rect 34155 -475 34160 -440
rect 34190 -475 34195 -440
rect 34155 -480 34195 -475
rect 34325 -440 34365 -435
rect 34325 -475 34330 -440
rect 34360 -475 34365 -440
rect 34325 -480 34365 -475
rect 34495 -440 34535 -435
rect 34495 -475 34500 -440
rect 34530 -475 34535 -440
rect 34495 -480 34535 -475
rect 34665 -440 34705 -435
rect 34665 -475 34670 -440
rect 34700 -475 34705 -440
rect 34665 -480 34705 -475
rect 34835 -440 34875 -435
rect 34835 -475 34840 -440
rect 34870 -475 34875 -440
rect 34835 -480 34875 -475
rect 35005 -440 35045 -435
rect 35005 -475 35010 -440
rect 35040 -475 35045 -440
rect 35005 -480 35045 -475
rect 35175 -440 35215 -435
rect 35175 -475 35180 -440
rect 35210 -475 35215 -440
rect 35175 -480 35215 -475
rect 35345 -440 35385 -435
rect 35345 -475 35350 -440
rect 35380 -475 35385 -440
rect 35345 -480 35385 -475
rect 35515 -440 35555 -435
rect 35515 -475 35520 -440
rect 35550 -475 35555 -440
rect 35515 -480 35555 -475
rect 35685 -440 35725 -435
rect 35685 -475 35690 -440
rect 35720 -475 35725 -440
rect 35685 -480 35725 -475
rect 35855 -440 35895 -435
rect 35855 -475 35860 -440
rect 35890 -475 35895 -440
rect 35855 -480 35895 -475
rect 36025 -440 36065 -435
rect 36025 -475 36030 -440
rect 36060 -475 36065 -440
rect 36025 -480 36065 -475
rect 36195 -440 36235 -435
rect 36195 -475 36200 -440
rect 36230 -475 36235 -440
rect 36195 -480 36235 -475
rect 36365 -440 36405 -435
rect 36365 -475 36370 -440
rect 36400 -475 36405 -440
rect 36365 -480 36405 -475
rect 36535 -440 36575 -435
rect 36535 -475 36540 -440
rect 36570 -475 36575 -440
rect 36535 -480 36575 -475
rect 36705 -440 36745 -435
rect 36705 -475 36710 -440
rect 36740 -475 36745 -440
rect 36705 -480 36745 -475
rect 36875 -440 36915 -435
rect 36875 -475 36880 -440
rect 36910 -475 36915 -440
rect 36875 -480 36915 -475
rect 37045 -440 37085 -435
rect 37045 -475 37050 -440
rect 37080 -475 37085 -440
rect 37045 -480 37085 -475
rect 37215 -440 37255 -435
rect 37215 -475 37220 -440
rect 37250 -475 37255 -440
rect 37215 -480 37255 -475
rect 37385 -440 37425 -435
rect 37385 -475 37390 -440
rect 37420 -475 37425 -440
rect 37385 -480 37425 -475
rect 37555 -440 37595 -435
rect 37555 -475 37560 -440
rect 37590 -475 37595 -440
rect 37555 -480 37595 -475
rect 37725 -440 37765 -435
rect 37725 -475 37730 -440
rect 37760 -475 37765 -440
rect 37725 -480 37765 -475
rect 37895 -440 37935 -435
rect 37895 -475 37900 -440
rect 37930 -475 37935 -440
rect 37895 -480 37935 -475
rect 38065 -440 38105 -435
rect 38065 -475 38070 -440
rect 38100 -475 38105 -440
rect 38065 -480 38105 -475
rect 38235 -440 38275 -435
rect 38235 -475 38240 -440
rect 38270 -475 38275 -440
rect 38235 -480 38275 -475
rect 38405 -440 38445 -435
rect 38405 -475 38410 -440
rect 38440 -475 38445 -440
rect 38405 -480 38445 -475
rect 38575 -440 38615 -435
rect 38575 -475 38580 -440
rect 38610 -475 38615 -440
rect 38575 -480 38615 -475
rect 38745 -440 38785 -435
rect 38745 -475 38750 -440
rect 38780 -475 38785 -440
rect 38745 -480 38785 -475
rect 38915 -440 38955 -435
rect 38915 -475 38920 -440
rect 38950 -475 38955 -440
rect 38915 -480 38955 -475
rect 39085 -440 39125 -435
rect 39085 -475 39090 -440
rect 39120 -475 39125 -440
rect 39085 -480 39125 -475
rect 39255 -440 39295 -435
rect 39255 -475 39260 -440
rect 39290 -475 39295 -440
rect 39255 -480 39295 -475
rect 39425 -440 39465 -435
rect 39425 -475 39430 -440
rect 39460 -475 39465 -440
rect 39425 -480 39465 -475
rect 39595 -440 39635 -435
rect 39595 -475 39600 -440
rect 39630 -475 39635 -440
rect 39595 -480 39635 -475
rect 39765 -440 39805 -435
rect 39765 -475 39770 -440
rect 39800 -475 39805 -440
rect 39765 -480 39805 -475
rect 39935 -440 39975 -435
rect 39935 -475 39940 -440
rect 39970 -475 39975 -440
rect 39935 -480 39975 -475
rect 40105 -440 40145 -435
rect 40105 -475 40110 -440
rect 40140 -475 40145 -440
rect 40105 -480 40145 -475
rect 40275 -440 40315 -435
rect 40275 -475 40280 -440
rect 40310 -475 40315 -440
rect 40275 -480 40315 -475
rect 40445 -440 40485 -435
rect 40445 -475 40450 -440
rect 40480 -475 40485 -440
rect 40445 -480 40485 -475
rect 40615 -440 40655 -435
rect 40615 -475 40620 -440
rect 40650 -475 40655 -440
rect 40615 -480 40655 -475
rect 40785 -440 40825 -435
rect 40785 -475 40790 -440
rect 40820 -475 40825 -440
rect 40785 -480 40825 -475
rect 40955 -440 40995 -435
rect 40955 -475 40960 -440
rect 40990 -475 40995 -440
rect 40955 -480 40995 -475
rect 41125 -440 41165 -435
rect 41125 -475 41130 -440
rect 41160 -475 41165 -440
rect 41125 -480 41165 -475
rect 41295 -440 41335 -435
rect 41295 -475 41300 -440
rect 41330 -475 41335 -440
rect 41295 -480 41335 -475
rect 41465 -440 41505 -435
rect 41465 -475 41470 -440
rect 41500 -475 41505 -440
rect 41465 -480 41505 -475
rect 41635 -440 41675 -435
rect 41635 -475 41640 -440
rect 41670 -475 41675 -440
rect 41635 -480 41675 -475
rect 41805 -440 41845 -435
rect 41805 -475 41810 -440
rect 41840 -475 41845 -440
rect 41805 -480 41845 -475
rect 41975 -440 42015 -435
rect 41975 -475 41980 -440
rect 42010 -475 42015 -440
rect 41975 -480 42015 -475
rect 42145 -440 42185 -435
rect 42145 -475 42150 -440
rect 42180 -475 42185 -440
rect 42145 -480 42185 -475
rect 42315 -440 42355 -435
rect 42315 -475 42320 -440
rect 42350 -475 42355 -440
rect 42315 -480 42355 -475
rect 42485 -440 42525 -435
rect 42485 -475 42490 -440
rect 42520 -475 42525 -440
rect 42485 -480 42525 -475
rect 42655 -440 42695 -435
rect 42655 -475 42660 -440
rect 42690 -475 42695 -440
rect 42655 -480 42695 -475
rect 42825 -440 42865 -435
rect 42825 -475 42830 -440
rect 42860 -475 42865 -440
rect 42825 -480 42865 -475
rect 42995 -440 43035 -435
rect 42995 -475 43000 -440
rect 43030 -475 43035 -440
rect 42995 -480 43035 -475
rect 43165 -440 43205 -435
rect 43165 -475 43170 -440
rect 43200 -475 43205 -440
rect 43165 -480 43205 -475
rect 43335 -440 43375 -435
rect 43335 -475 43340 -440
rect 43370 -475 43375 -440
rect 43335 -480 43375 -475
rect 43505 -440 43545 -435
rect 43505 -475 43510 -440
rect 43540 -475 43545 -440
rect 43505 -480 43545 -475
rect 65 -550 115 -540
rect 235 -550 285 -540
rect 405 -550 455 -540
rect 575 -550 625 -540
rect 745 -550 795 -540
rect 915 -550 965 -540
rect 1085 -550 1135 -540
rect 1255 -550 1305 -540
rect 1425 -550 1475 -540
rect 1595 -550 1645 -540
rect 1765 -550 1815 -540
rect 1935 -550 1985 -540
rect 2105 -550 2155 -540
rect 2275 -550 2325 -540
rect 2445 -550 2495 -540
rect 2615 -550 2665 -540
rect 2785 -550 2835 -540
rect 2955 -550 3005 -540
rect 3125 -550 3175 -540
rect 3295 -550 3345 -540
rect 3465 -550 3515 -540
rect 3635 -550 3685 -540
rect 3805 -550 3855 -540
rect 3975 -550 4025 -540
rect 4145 -550 4195 -540
rect 4315 -550 4365 -540
rect 4485 -550 4535 -540
rect 4655 -550 4705 -540
rect 4825 -550 4875 -540
rect 4995 -550 5045 -540
rect 5165 -550 5215 -540
rect 5335 -550 5385 -540
rect 5505 -550 5555 -540
rect 5675 -550 5725 -540
rect 5845 -550 5895 -540
rect 6015 -550 6065 -540
rect 6185 -550 6235 -540
rect 6355 -550 6405 -540
rect 6525 -550 6575 -540
rect 6695 -550 6745 -540
rect 6865 -550 6915 -540
rect 7035 -550 7085 -540
rect 7205 -550 7255 -540
rect 7375 -550 7425 -540
rect 7545 -550 7595 -540
rect 7715 -550 7765 -540
rect 7885 -550 7935 -540
rect 8055 -550 8105 -540
rect 8225 -550 8275 -540
rect 8395 -550 8445 -540
rect 8565 -550 8615 -540
rect 8735 -550 8785 -540
rect 8905 -550 8955 -540
rect 9075 -550 9125 -540
rect 9245 -550 9295 -540
rect 9415 -550 9465 -540
rect 9585 -550 9635 -540
rect 9755 -550 9805 -540
rect 9925 -550 9975 -540
rect 10095 -550 10145 -540
rect 10265 -550 10315 -540
rect 10435 -550 10485 -540
rect 10605 -550 10655 -540
rect 10775 -550 10825 -540
rect 10945 -550 10995 -540
rect 11115 -550 11165 -540
rect 11285 -550 11335 -540
rect 11455 -550 11505 -540
rect 11625 -550 11675 -540
rect 11795 -550 11845 -540
rect 11965 -550 12015 -540
rect 12135 -550 12185 -540
rect 12305 -550 12355 -540
rect 12475 -550 12525 -540
rect 12645 -550 12695 -540
rect 12815 -550 12865 -540
rect 12985 -550 13035 -540
rect 13155 -550 13205 -540
rect 13325 -550 13375 -540
rect 13495 -550 13545 -540
rect 13665 -550 13715 -540
rect 13835 -550 13885 -540
rect 14005 -550 14055 -540
rect 14175 -550 14225 -540
rect 14345 -550 14395 -540
rect 14515 -550 14565 -540
rect 14685 -550 14735 -540
rect 14855 -550 14905 -540
rect 15025 -550 15075 -540
rect 15195 -550 15245 -540
rect 15365 -550 15415 -540
rect 15535 -550 15585 -540
rect 15705 -550 15755 -540
rect 15875 -550 15925 -540
rect 16045 -550 16095 -540
rect 16215 -550 16265 -540
rect 16385 -550 16435 -540
rect 16555 -550 16605 -540
rect 16725 -550 16775 -540
rect 16895 -550 16945 -540
rect 17065 -550 17115 -540
rect 17235 -550 17285 -540
rect 17405 -550 17455 -540
rect 17575 -550 17625 -540
rect 17745 -550 17795 -540
rect 17915 -550 17965 -540
rect 18085 -550 18135 -540
rect 18255 -550 18305 -540
rect 18425 -550 18475 -540
rect 18595 -550 18645 -540
rect 18765 -550 18815 -540
rect 18935 -550 18985 -540
rect 19105 -550 19155 -540
rect 19275 -550 19325 -540
rect 19445 -550 19495 -540
rect 19615 -550 19665 -540
rect 19785 -550 19835 -540
rect 19955 -550 20005 -540
rect 20125 -550 20175 -540
rect 20295 -550 20345 -540
rect 20465 -550 20515 -540
rect 20635 -550 20685 -540
rect 20805 -550 20855 -540
rect 20975 -550 21025 -540
rect 21145 -550 21195 -540
rect 21315 -550 21365 -540
rect 21485 -550 21535 -540
rect 21655 -550 21705 -540
rect 21825 -550 21875 -540
rect 21995 -550 22045 -540
rect 22165 -550 22215 -540
rect 22335 -550 22385 -540
rect 22505 -550 22555 -540
rect 22675 -550 22725 -540
rect 22845 -550 22895 -540
rect 23015 -550 23065 -540
rect 23185 -550 23235 -540
rect 23355 -550 23405 -540
rect 23525 -550 23575 -540
rect 23695 -550 23745 -540
rect 23865 -550 23915 -540
rect 24035 -550 24085 -540
rect 24205 -550 24255 -540
rect 24375 -550 24425 -540
rect 24545 -550 24595 -540
rect 24715 -550 24765 -540
rect 24885 -550 24935 -540
rect 25055 -550 25105 -540
rect 25225 -550 25275 -540
rect 25395 -550 25445 -540
rect 25565 -550 25615 -540
rect 25735 -550 25785 -540
rect 25905 -550 25955 -540
rect 26075 -550 26125 -540
rect 26245 -550 26295 -540
rect 26415 -550 26465 -540
rect 26585 -550 26635 -540
rect 26755 -550 26805 -540
rect 26925 -550 26975 -540
rect 27095 -550 27145 -540
rect 27265 -550 27315 -540
rect 27435 -550 27485 -540
rect 27605 -550 27655 -540
rect 27775 -550 27825 -540
rect 27945 -550 27995 -540
rect 28115 -550 28165 -540
rect 28285 -550 28335 -540
rect 28455 -550 28505 -540
rect 28625 -550 28675 -540
rect 28795 -550 28845 -540
rect 28965 -550 29015 -540
rect 29135 -550 29185 -540
rect 29305 -550 29355 -540
rect 29475 -550 29525 -540
rect 29645 -550 29695 -540
rect 29815 -550 29865 -540
rect 29985 -550 30035 -540
rect 30155 -550 30205 -540
rect 30325 -550 30375 -540
rect 30495 -550 30545 -540
rect 30665 -550 30715 -540
rect 30835 -550 30885 -540
rect 31005 -550 31055 -540
rect 31175 -550 31225 -540
rect 31345 -550 31395 -540
rect 31515 -550 31565 -540
rect 31685 -550 31735 -540
rect 31855 -550 31905 -540
rect 32025 -550 32075 -540
rect 32195 -550 32245 -540
rect 32365 -550 32415 -540
rect 32535 -550 32585 -540
rect 32705 -550 32755 -540
rect 32875 -550 32925 -540
rect 33045 -550 33095 -540
rect 33215 -550 33265 -540
rect 33385 -550 33435 -540
rect 33555 -550 33605 -540
rect 33725 -550 33775 -540
rect 33895 -550 33945 -540
rect 34065 -550 34115 -540
rect 34235 -550 34285 -540
rect 34405 -550 34455 -540
rect 34575 -550 34625 -540
rect 34745 -550 34795 -540
rect 34915 -550 34965 -540
rect 35085 -550 35135 -540
rect 35255 -550 35305 -540
rect 35425 -550 35475 -540
rect 35595 -550 35645 -540
rect 35765 -550 35815 -540
rect 35935 -550 35985 -540
rect 36105 -550 36155 -540
rect 36275 -550 36325 -540
rect 36445 -550 36495 -540
rect 36615 -550 36665 -540
rect 36785 -550 36835 -540
rect 36955 -550 37005 -540
rect 37125 -550 37175 -540
rect 37295 -550 37345 -540
rect 37465 -550 37515 -540
rect 37635 -550 37685 -540
rect 37805 -550 37855 -540
rect 37975 -550 38025 -540
rect 38145 -550 38195 -540
rect 38315 -550 38365 -540
rect 38485 -550 38535 -540
rect 38655 -550 38705 -540
rect 38825 -550 38875 -540
rect 38995 -550 39045 -540
rect 39165 -550 39215 -540
rect 39335 -550 39385 -540
rect 39505 -550 39555 -540
rect 39675 -550 39725 -540
rect 39845 -550 39895 -540
rect 40015 -550 40065 -540
rect 40185 -550 40235 -540
rect 40355 -550 40405 -540
rect 40525 -550 40575 -540
rect 40695 -550 40745 -540
rect 40865 -550 40915 -540
rect 41035 -550 41085 -540
rect 41205 -550 41255 -540
rect 41375 -550 41425 -540
rect 41545 -550 41595 -540
rect 41715 -550 41765 -540
rect 41885 -550 41935 -540
rect 42055 -550 42105 -540
rect 42225 -550 42275 -540
rect 42395 -550 42445 -540
rect 42565 -550 42615 -540
rect 42735 -550 42785 -540
rect 42905 -550 42955 -540
rect 43075 -550 43125 -540
rect 43245 -550 43295 -540
rect 43415 -550 43465 -540
rect 43585 -550 43635 -540
rect 55 -580 75 -550
rect 105 -580 245 -550
rect 275 -580 415 -550
rect 445 -580 585 -550
rect 615 -580 755 -550
rect 785 -580 925 -550
rect 955 -580 1095 -550
rect 1125 -580 1265 -550
rect 1295 -580 1435 -550
rect 1465 -580 1605 -550
rect 1635 -580 1775 -550
rect 1805 -580 1945 -550
rect 1975 -580 2115 -550
rect 2145 -580 2285 -550
rect 2315 -580 2455 -550
rect 2485 -580 2625 -550
rect 2655 -580 2795 -550
rect 2825 -580 2965 -550
rect 2995 -580 3135 -550
rect 3165 -580 3305 -550
rect 3335 -580 3475 -550
rect 3505 -580 3645 -550
rect 3675 -580 3815 -550
rect 3845 -580 3985 -550
rect 4015 -580 4155 -550
rect 4185 -580 4325 -550
rect 4355 -580 4495 -550
rect 4525 -580 4665 -550
rect 4695 -580 4835 -550
rect 4865 -580 5005 -550
rect 5035 -580 5175 -550
rect 5205 -580 5345 -550
rect 5375 -580 5515 -550
rect 5545 -580 5685 -550
rect 5715 -580 5855 -550
rect 5885 -580 6025 -550
rect 6055 -580 6195 -550
rect 6225 -580 6365 -550
rect 6395 -580 6535 -550
rect 6565 -580 6705 -550
rect 6735 -580 6875 -550
rect 6905 -580 7045 -550
rect 7075 -580 7215 -550
rect 7245 -580 7385 -550
rect 7415 -580 7555 -550
rect 7585 -580 7725 -550
rect 7755 -580 7895 -550
rect 7925 -580 8065 -550
rect 8095 -580 8235 -550
rect 8265 -580 8405 -550
rect 8435 -580 8575 -550
rect 8605 -580 8745 -550
rect 8775 -580 8915 -550
rect 8945 -580 9085 -550
rect 9115 -580 9255 -550
rect 9285 -580 9425 -550
rect 9455 -580 9595 -550
rect 9625 -580 9765 -550
rect 9795 -580 9935 -550
rect 9965 -580 10105 -550
rect 10135 -580 10275 -550
rect 10305 -580 10445 -550
rect 10475 -580 10615 -550
rect 10645 -580 10785 -550
rect 10815 -580 10955 -550
rect 10985 -580 11125 -550
rect 11155 -580 11295 -550
rect 11325 -580 11465 -550
rect 11495 -580 11635 -550
rect 11665 -580 11805 -550
rect 11835 -580 11975 -550
rect 12005 -580 12145 -550
rect 12175 -580 12315 -550
rect 12345 -580 12485 -550
rect 12515 -580 12655 -550
rect 12685 -580 12825 -550
rect 12855 -580 12995 -550
rect 13025 -580 13165 -550
rect 13195 -580 13335 -550
rect 13365 -580 13505 -550
rect 13535 -580 13675 -550
rect 13705 -580 13845 -550
rect 13875 -580 14015 -550
rect 14045 -580 14185 -550
rect 14215 -580 14355 -550
rect 14385 -580 14525 -550
rect 14555 -580 14695 -550
rect 14725 -580 14865 -550
rect 14895 -580 15035 -550
rect 15065 -580 15205 -550
rect 15235 -580 15375 -550
rect 15405 -580 15545 -550
rect 15575 -580 15715 -550
rect 15745 -580 15885 -550
rect 15915 -580 16055 -550
rect 16085 -580 16225 -550
rect 16255 -580 16395 -550
rect 16425 -580 16565 -550
rect 16595 -580 16735 -550
rect 16765 -580 16905 -550
rect 16935 -580 17075 -550
rect 17105 -580 17245 -550
rect 17275 -580 17415 -550
rect 17445 -580 17585 -550
rect 17615 -580 17755 -550
rect 17785 -580 17925 -550
rect 17955 -580 18095 -550
rect 18125 -580 18265 -550
rect 18295 -580 18435 -550
rect 18465 -580 18605 -550
rect 18635 -580 18775 -550
rect 18805 -580 18945 -550
rect 18975 -580 19115 -550
rect 19145 -580 19285 -550
rect 19315 -580 19455 -550
rect 19485 -580 19625 -550
rect 19655 -580 19795 -550
rect 19825 -580 19965 -550
rect 19995 -580 20135 -550
rect 20165 -580 20305 -550
rect 20335 -580 20475 -550
rect 20505 -580 20645 -550
rect 20675 -580 20815 -550
rect 20845 -580 20985 -550
rect 21015 -580 21155 -550
rect 21185 -580 21325 -550
rect 21355 -580 21495 -550
rect 21525 -580 21665 -550
rect 21695 -580 21835 -550
rect 21865 -580 22005 -550
rect 22035 -580 22175 -550
rect 22205 -580 22345 -550
rect 22375 -580 22515 -550
rect 22545 -580 22685 -550
rect 22715 -580 22855 -550
rect 22885 -580 23025 -550
rect 23055 -580 23195 -550
rect 23225 -580 23365 -550
rect 23395 -580 23535 -550
rect 23565 -580 23705 -550
rect 23735 -580 23875 -550
rect 23905 -580 24045 -550
rect 24075 -580 24215 -550
rect 24245 -580 24385 -550
rect 24415 -580 24555 -550
rect 24585 -580 24725 -550
rect 24755 -580 24895 -550
rect 24925 -580 25065 -550
rect 25095 -580 25235 -550
rect 25265 -580 25405 -550
rect 25435 -580 25575 -550
rect 25605 -580 25745 -550
rect 25775 -580 25915 -550
rect 25945 -580 26085 -550
rect 26115 -580 26255 -550
rect 26285 -580 26425 -550
rect 26455 -580 26595 -550
rect 26625 -580 26765 -550
rect 26795 -580 26935 -550
rect 26965 -580 27105 -550
rect 27135 -580 27275 -550
rect 27305 -580 27445 -550
rect 27475 -580 27615 -550
rect 27645 -580 27785 -550
rect 27815 -580 27955 -550
rect 27985 -580 28125 -550
rect 28155 -580 28295 -550
rect 28325 -580 28465 -550
rect 28495 -580 28635 -550
rect 28665 -580 28805 -550
rect 28835 -580 28975 -550
rect 29005 -580 29145 -550
rect 29175 -580 29315 -550
rect 29345 -580 29485 -550
rect 29515 -580 29655 -550
rect 29685 -580 29825 -550
rect 29855 -580 29995 -550
rect 30025 -580 30165 -550
rect 30195 -580 30335 -550
rect 30365 -580 30505 -550
rect 30535 -580 30675 -550
rect 30705 -580 30845 -550
rect 30875 -580 31015 -550
rect 31045 -580 31185 -550
rect 31215 -580 31355 -550
rect 31385 -580 31525 -550
rect 31555 -580 31695 -550
rect 31725 -580 31865 -550
rect 31895 -580 32035 -550
rect 32065 -580 32205 -550
rect 32235 -580 32375 -550
rect 32405 -580 32545 -550
rect 32575 -580 32715 -550
rect 32745 -580 32885 -550
rect 32915 -580 33055 -550
rect 33085 -580 33225 -550
rect 33255 -580 33395 -550
rect 33425 -580 33565 -550
rect 33595 -580 33735 -550
rect 33765 -580 33905 -550
rect 33935 -580 34075 -550
rect 34105 -580 34245 -550
rect 34275 -580 34415 -550
rect 34445 -580 34585 -550
rect 34615 -580 34755 -550
rect 34785 -580 34925 -550
rect 34955 -580 35095 -550
rect 35125 -580 35265 -550
rect 35295 -580 35435 -550
rect 35465 -580 35605 -550
rect 35635 -580 35775 -550
rect 35805 -580 35945 -550
rect 35975 -580 36115 -550
rect 36145 -580 36285 -550
rect 36315 -580 36455 -550
rect 36485 -580 36625 -550
rect 36655 -580 36795 -550
rect 36825 -580 36965 -550
rect 36995 -580 37135 -550
rect 37165 -580 37305 -550
rect 37335 -580 37475 -550
rect 37505 -580 37645 -550
rect 37675 -580 37815 -550
rect 37845 -580 37985 -550
rect 38015 -580 38155 -550
rect 38185 -580 38325 -550
rect 38355 -580 38495 -550
rect 38525 -580 38665 -550
rect 38695 -580 38835 -550
rect 38865 -580 39005 -550
rect 39035 -580 39175 -550
rect 39205 -580 39345 -550
rect 39375 -580 39515 -550
rect 39545 -580 39685 -550
rect 39715 -580 39855 -550
rect 39885 -580 40025 -550
rect 40055 -580 40195 -550
rect 40225 -580 40365 -550
rect 40395 -580 40535 -550
rect 40565 -580 40705 -550
rect 40735 -580 40875 -550
rect 40905 -580 41045 -550
rect 41075 -580 41215 -550
rect 41245 -580 41385 -550
rect 41415 -580 41555 -550
rect 41585 -580 41725 -550
rect 41755 -580 41895 -550
rect 41925 -580 42065 -550
rect 42095 -580 42235 -550
rect 42265 -580 42405 -550
rect 42435 -580 42575 -550
rect 42605 -580 42745 -550
rect 42775 -580 42915 -550
rect 42945 -580 43085 -550
rect 43115 -580 43255 -550
rect 43285 -580 43425 -550
rect 43455 -580 43595 -550
rect 43625 -580 43635 -550
rect 65 -590 115 -580
rect 235 -590 285 -580
rect 405 -590 455 -580
rect 575 -590 625 -580
rect 745 -590 795 -580
rect 915 -590 965 -580
rect 1085 -590 1135 -580
rect 1255 -590 1305 -580
rect 1425 -590 1475 -580
rect 1595 -590 1645 -580
rect 1765 -590 1815 -580
rect 1935 -590 1985 -580
rect 2105 -590 2155 -580
rect 2275 -590 2325 -580
rect 2445 -590 2495 -580
rect 2615 -590 2665 -580
rect 2785 -590 2835 -580
rect 2955 -590 3005 -580
rect 3125 -590 3175 -580
rect 3295 -590 3345 -580
rect 3465 -590 3515 -580
rect 3635 -590 3685 -580
rect 3805 -590 3855 -580
rect 3975 -590 4025 -580
rect 4145 -590 4195 -580
rect 4315 -590 4365 -580
rect 4485 -590 4535 -580
rect 4655 -590 4705 -580
rect 4825 -590 4875 -580
rect 4995 -590 5045 -580
rect 5165 -590 5215 -580
rect 5335 -590 5385 -580
rect 5505 -590 5555 -580
rect 5675 -590 5725 -580
rect 5845 -590 5895 -580
rect 6015 -590 6065 -580
rect 6185 -590 6235 -580
rect 6355 -590 6405 -580
rect 6525 -590 6575 -580
rect 6695 -590 6745 -580
rect 6865 -590 6915 -580
rect 7035 -590 7085 -580
rect 7205 -590 7255 -580
rect 7375 -590 7425 -580
rect 7545 -590 7595 -580
rect 7715 -590 7765 -580
rect 7885 -590 7935 -580
rect 8055 -590 8105 -580
rect 8225 -590 8275 -580
rect 8395 -590 8445 -580
rect 8565 -590 8615 -580
rect 8735 -590 8785 -580
rect 8905 -590 8955 -580
rect 9075 -590 9125 -580
rect 9245 -590 9295 -580
rect 9415 -590 9465 -580
rect 9585 -590 9635 -580
rect 9755 -590 9805 -580
rect 9925 -590 9975 -580
rect 10095 -590 10145 -580
rect 10265 -590 10315 -580
rect 10435 -590 10485 -580
rect 10605 -590 10655 -580
rect 10775 -590 10825 -580
rect 10945 -590 10995 -580
rect 11115 -590 11165 -580
rect 11285 -590 11335 -580
rect 11455 -590 11505 -580
rect 11625 -590 11675 -580
rect 11795 -590 11845 -580
rect 11965 -590 12015 -580
rect 12135 -590 12185 -580
rect 12305 -590 12355 -580
rect 12475 -590 12525 -580
rect 12645 -590 12695 -580
rect 12815 -590 12865 -580
rect 12985 -590 13035 -580
rect 13155 -590 13205 -580
rect 13325 -590 13375 -580
rect 13495 -590 13545 -580
rect 13665 -590 13715 -580
rect 13835 -590 13885 -580
rect 14005 -590 14055 -580
rect 14175 -590 14225 -580
rect 14345 -590 14395 -580
rect 14515 -590 14565 -580
rect 14685 -590 14735 -580
rect 14855 -590 14905 -580
rect 15025 -590 15075 -580
rect 15195 -590 15245 -580
rect 15365 -590 15415 -580
rect 15535 -590 15585 -580
rect 15705 -590 15755 -580
rect 15875 -590 15925 -580
rect 16045 -590 16095 -580
rect 16215 -590 16265 -580
rect 16385 -590 16435 -580
rect 16555 -590 16605 -580
rect 16725 -590 16775 -580
rect 16895 -590 16945 -580
rect 17065 -590 17115 -580
rect 17235 -590 17285 -580
rect 17405 -590 17455 -580
rect 17575 -590 17625 -580
rect 17745 -590 17795 -580
rect 17915 -590 17965 -580
rect 18085 -590 18135 -580
rect 18255 -590 18305 -580
rect 18425 -590 18475 -580
rect 18595 -590 18645 -580
rect 18765 -590 18815 -580
rect 18935 -590 18985 -580
rect 19105 -590 19155 -580
rect 19275 -590 19325 -580
rect 19445 -590 19495 -580
rect 19615 -590 19665 -580
rect 19785 -590 19835 -580
rect 19955 -590 20005 -580
rect 20125 -590 20175 -580
rect 20295 -590 20345 -580
rect 20465 -590 20515 -580
rect 20635 -590 20685 -580
rect 20805 -590 20855 -580
rect 20975 -590 21025 -580
rect 21145 -590 21195 -580
rect 21315 -590 21365 -580
rect 21485 -590 21535 -580
rect 21655 -590 21705 -580
rect 21825 -590 21875 -580
rect 21995 -590 22045 -580
rect 22165 -590 22215 -580
rect 22335 -590 22385 -580
rect 22505 -590 22555 -580
rect 22675 -590 22725 -580
rect 22845 -590 22895 -580
rect 23015 -590 23065 -580
rect 23185 -590 23235 -580
rect 23355 -590 23405 -580
rect 23525 -590 23575 -580
rect 23695 -590 23745 -580
rect 23865 -590 23915 -580
rect 24035 -590 24085 -580
rect 24205 -590 24255 -580
rect 24375 -590 24425 -580
rect 24545 -590 24595 -580
rect 24715 -590 24765 -580
rect 24885 -590 24935 -580
rect 25055 -590 25105 -580
rect 25225 -590 25275 -580
rect 25395 -590 25445 -580
rect 25565 -590 25615 -580
rect 25735 -590 25785 -580
rect 25905 -590 25955 -580
rect 26075 -590 26125 -580
rect 26245 -590 26295 -580
rect 26415 -590 26465 -580
rect 26585 -590 26635 -580
rect 26755 -590 26805 -580
rect 26925 -590 26975 -580
rect 27095 -590 27145 -580
rect 27265 -590 27315 -580
rect 27435 -590 27485 -580
rect 27605 -590 27655 -580
rect 27775 -590 27825 -580
rect 27945 -590 27995 -580
rect 28115 -590 28165 -580
rect 28285 -590 28335 -580
rect 28455 -590 28505 -580
rect 28625 -590 28675 -580
rect 28795 -590 28845 -580
rect 28965 -590 29015 -580
rect 29135 -590 29185 -580
rect 29305 -590 29355 -580
rect 29475 -590 29525 -580
rect 29645 -590 29695 -580
rect 29815 -590 29865 -580
rect 29985 -590 30035 -580
rect 30155 -590 30205 -580
rect 30325 -590 30375 -580
rect 30495 -590 30545 -580
rect 30665 -590 30715 -580
rect 30835 -590 30885 -580
rect 31005 -590 31055 -580
rect 31175 -590 31225 -580
rect 31345 -590 31395 -580
rect 31515 -590 31565 -580
rect 31685 -590 31735 -580
rect 31855 -590 31905 -580
rect 32025 -590 32075 -580
rect 32195 -590 32245 -580
rect 32365 -590 32415 -580
rect 32535 -590 32585 -580
rect 32705 -590 32755 -580
rect 32875 -590 32925 -580
rect 33045 -590 33095 -580
rect 33215 -590 33265 -580
rect 33385 -590 33435 -580
rect 33555 -590 33605 -580
rect 33725 -590 33775 -580
rect 33895 -590 33945 -580
rect 34065 -590 34115 -580
rect 34235 -590 34285 -580
rect 34405 -590 34455 -580
rect 34575 -590 34625 -580
rect 34745 -590 34795 -580
rect 34915 -590 34965 -580
rect 35085 -590 35135 -580
rect 35255 -590 35305 -580
rect 35425 -590 35475 -580
rect 35595 -590 35645 -580
rect 35765 -590 35815 -580
rect 35935 -590 35985 -580
rect 36105 -590 36155 -580
rect 36275 -590 36325 -580
rect 36445 -590 36495 -580
rect 36615 -590 36665 -580
rect 36785 -590 36835 -580
rect 36955 -590 37005 -580
rect 37125 -590 37175 -580
rect 37295 -590 37345 -580
rect 37465 -590 37515 -580
rect 37635 -590 37685 -580
rect 37805 -590 37855 -580
rect 37975 -590 38025 -580
rect 38145 -590 38195 -580
rect 38315 -590 38365 -580
rect 38485 -590 38535 -580
rect 38655 -590 38705 -580
rect 38825 -590 38875 -580
rect 38995 -590 39045 -580
rect 39165 -590 39215 -580
rect 39335 -590 39385 -580
rect 39505 -590 39555 -580
rect 39675 -590 39725 -580
rect 39845 -590 39895 -580
rect 40015 -590 40065 -580
rect 40185 -590 40235 -580
rect 40355 -590 40405 -580
rect 40525 -590 40575 -580
rect 40695 -590 40745 -580
rect 40865 -590 40915 -580
rect 41035 -590 41085 -580
rect 41205 -590 41255 -580
rect 41375 -590 41425 -580
rect 41545 -590 41595 -580
rect 41715 -590 41765 -580
rect 41885 -590 41935 -580
rect 42055 -590 42105 -580
rect 42225 -590 42275 -580
rect 42395 -590 42445 -580
rect 42565 -590 42615 -580
rect 42735 -590 42785 -580
rect 42905 -590 42955 -580
rect 43075 -590 43125 -580
rect 43245 -590 43295 -580
rect 43415 -590 43465 -580
rect 43585 -590 43635 -580
rect 65 -650 115 -640
rect 235 -650 285 -640
rect 405 -650 455 -640
rect 575 -650 625 -640
rect 745 -650 795 -640
rect 915 -650 965 -640
rect 1085 -650 1135 -640
rect 1255 -650 1305 -640
rect 1425 -650 1475 -640
rect 1595 -650 1645 -640
rect 1765 -650 1815 -640
rect 1935 -650 1985 -640
rect 2105 -650 2155 -640
rect 2275 -650 2325 -640
rect 2445 -650 2495 -640
rect 2615 -650 2665 -640
rect 2785 -650 2835 -640
rect 2955 -650 3005 -640
rect 3125 -650 3175 -640
rect 3295 -650 3345 -640
rect 3465 -650 3515 -640
rect 3635 -650 3685 -640
rect 3805 -650 3855 -640
rect 3975 -650 4025 -640
rect 4145 -650 4195 -640
rect 4315 -650 4365 -640
rect 4485 -650 4535 -640
rect 4655 -650 4705 -640
rect 4825 -650 4875 -640
rect 4995 -650 5045 -640
rect 5165 -650 5215 -640
rect 5335 -650 5385 -640
rect 5505 -650 5555 -640
rect 5675 -650 5725 -640
rect 5845 -650 5895 -640
rect 6015 -650 6065 -640
rect 6185 -650 6235 -640
rect 6355 -650 6405 -640
rect 6525 -650 6575 -640
rect 6695 -650 6745 -640
rect 6865 -650 6915 -640
rect 7035 -650 7085 -640
rect 7205 -650 7255 -640
rect 7375 -650 7425 -640
rect 7545 -650 7595 -640
rect 7715 -650 7765 -640
rect 7885 -650 7935 -640
rect 8055 -650 8105 -640
rect 8225 -650 8275 -640
rect 8395 -650 8445 -640
rect 8565 -650 8615 -640
rect 8735 -650 8785 -640
rect 8905 -650 8955 -640
rect 9075 -650 9125 -640
rect 9245 -650 9295 -640
rect 9415 -650 9465 -640
rect 9585 -650 9635 -640
rect 9755 -650 9805 -640
rect 9925 -650 9975 -640
rect 10095 -650 10145 -640
rect 10265 -650 10315 -640
rect 10435 -650 10485 -640
rect 10605 -650 10655 -640
rect 10775 -650 10825 -640
rect 10945 -650 10995 -640
rect 11115 -650 11165 -640
rect 11285 -650 11335 -640
rect 11455 -650 11505 -640
rect 11625 -650 11675 -640
rect 11795 -650 11845 -640
rect 11965 -650 12015 -640
rect 12135 -650 12185 -640
rect 12305 -650 12355 -640
rect 12475 -650 12525 -640
rect 12645 -650 12695 -640
rect 12815 -650 12865 -640
rect 12985 -650 13035 -640
rect 13155 -650 13205 -640
rect 13325 -650 13375 -640
rect 13495 -650 13545 -640
rect 13665 -650 13715 -640
rect 13835 -650 13885 -640
rect 14005 -650 14055 -640
rect 14175 -650 14225 -640
rect 14345 -650 14395 -640
rect 14515 -650 14565 -640
rect 14685 -650 14735 -640
rect 14855 -650 14905 -640
rect 15025 -650 15075 -640
rect 15195 -650 15245 -640
rect 15365 -650 15415 -640
rect 15535 -650 15585 -640
rect 15705 -650 15755 -640
rect 15875 -650 15925 -640
rect 16045 -650 16095 -640
rect 16215 -650 16265 -640
rect 16385 -650 16435 -640
rect 16555 -650 16605 -640
rect 16725 -650 16775 -640
rect 16895 -650 16945 -640
rect 17065 -650 17115 -640
rect 17235 -650 17285 -640
rect 17405 -650 17455 -640
rect 17575 -650 17625 -640
rect 17745 -650 17795 -640
rect 17915 -650 17965 -640
rect 18085 -650 18135 -640
rect 18255 -650 18305 -640
rect 18425 -650 18475 -640
rect 18595 -650 18645 -640
rect 18765 -650 18815 -640
rect 18935 -650 18985 -640
rect 19105 -650 19155 -640
rect 19275 -650 19325 -640
rect 19445 -650 19495 -640
rect 19615 -650 19665 -640
rect 19785 -650 19835 -640
rect 19955 -650 20005 -640
rect 20125 -650 20175 -640
rect 20295 -650 20345 -640
rect 20465 -650 20515 -640
rect 20635 -650 20685 -640
rect 20805 -650 20855 -640
rect 20975 -650 21025 -640
rect 21145 -650 21195 -640
rect 21315 -650 21365 -640
rect 21485 -650 21535 -640
rect 21655 -650 21705 -640
rect 21825 -650 21875 -640
rect 21995 -650 22045 -640
rect 22165 -650 22215 -640
rect 22335 -650 22385 -640
rect 22505 -650 22555 -640
rect 22675 -650 22725 -640
rect 22845 -650 22895 -640
rect 23015 -650 23065 -640
rect 23185 -650 23235 -640
rect 23355 -650 23405 -640
rect 23525 -650 23575 -640
rect 23695 -650 23745 -640
rect 23865 -650 23915 -640
rect 24035 -650 24085 -640
rect 24205 -650 24255 -640
rect 24375 -650 24425 -640
rect 24545 -650 24595 -640
rect 24715 -650 24765 -640
rect 24885 -650 24935 -640
rect 25055 -650 25105 -640
rect 25225 -650 25275 -640
rect 25395 -650 25445 -640
rect 25565 -650 25615 -640
rect 25735 -650 25785 -640
rect 25905 -650 25955 -640
rect 26075 -650 26125 -640
rect 26245 -650 26295 -640
rect 26415 -650 26465 -640
rect 26585 -650 26635 -640
rect 26755 -650 26805 -640
rect 26925 -650 26975 -640
rect 27095 -650 27145 -640
rect 27265 -650 27315 -640
rect 27435 -650 27485 -640
rect 27605 -650 27655 -640
rect 27775 -650 27825 -640
rect 27945 -650 27995 -640
rect 28115 -650 28165 -640
rect 28285 -650 28335 -640
rect 28455 -650 28505 -640
rect 28625 -650 28675 -640
rect 28795 -650 28845 -640
rect 28965 -650 29015 -640
rect 29135 -650 29185 -640
rect 29305 -650 29355 -640
rect 29475 -650 29525 -640
rect 29645 -650 29695 -640
rect 29815 -650 29865 -640
rect 29985 -650 30035 -640
rect 30155 -650 30205 -640
rect 30325 -650 30375 -640
rect 30495 -650 30545 -640
rect 30665 -650 30715 -640
rect 30835 -650 30885 -640
rect 31005 -650 31055 -640
rect 31175 -650 31225 -640
rect 31345 -650 31395 -640
rect 31515 -650 31565 -640
rect 31685 -650 31735 -640
rect 31855 -650 31905 -640
rect 32025 -650 32075 -640
rect 32195 -650 32245 -640
rect 32365 -650 32415 -640
rect 32535 -650 32585 -640
rect 32705 -650 32755 -640
rect 32875 -650 32925 -640
rect 33045 -650 33095 -640
rect 33215 -650 33265 -640
rect 33385 -650 33435 -640
rect 33555 -650 33605 -640
rect 33725 -650 33775 -640
rect 33895 -650 33945 -640
rect 34065 -650 34115 -640
rect 34235 -650 34285 -640
rect 34405 -650 34455 -640
rect 34575 -650 34625 -640
rect 34745 -650 34795 -640
rect 34915 -650 34965 -640
rect 35085 -650 35135 -640
rect 35255 -650 35305 -640
rect 35425 -650 35475 -640
rect 35595 -650 35645 -640
rect 35765 -650 35815 -640
rect 35935 -650 35985 -640
rect 36105 -650 36155 -640
rect 36275 -650 36325 -640
rect 36445 -650 36495 -640
rect 36615 -650 36665 -640
rect 36785 -650 36835 -640
rect 36955 -650 37005 -640
rect 37125 -650 37175 -640
rect 37295 -650 37345 -640
rect 37465 -650 37515 -640
rect 37635 -650 37685 -640
rect 37805 -650 37855 -640
rect 37975 -650 38025 -640
rect 38145 -650 38195 -640
rect 38315 -650 38365 -640
rect 38485 -650 38535 -640
rect 38655 -650 38705 -640
rect 38825 -650 38875 -640
rect 38995 -650 39045 -640
rect 39165 -650 39215 -640
rect 39335 -650 39385 -640
rect 39505 -650 39555 -640
rect 39675 -650 39725 -640
rect 39845 -650 39895 -640
rect 40015 -650 40065 -640
rect 40185 -650 40235 -640
rect 40355 -650 40405 -640
rect 40525 -650 40575 -640
rect 40695 -650 40745 -640
rect 40865 -650 40915 -640
rect 41035 -650 41085 -640
rect 41205 -650 41255 -640
rect 41375 -650 41425 -640
rect 41545 -650 41595 -640
rect 41715 -650 41765 -640
rect 41885 -650 41935 -640
rect 42055 -650 42105 -640
rect 42225 -650 42275 -640
rect 42395 -650 42445 -640
rect 42565 -650 42615 -640
rect 42735 -650 42785 -640
rect 42905 -650 42955 -640
rect 43075 -650 43125 -640
rect 43245 -650 43295 -640
rect 43415 -650 43465 -640
rect 43585 -650 43635 -640
rect 55 -680 75 -650
rect 105 -680 245 -650
rect 275 -680 415 -650
rect 445 -680 585 -650
rect 615 -680 755 -650
rect 785 -680 925 -650
rect 955 -680 1095 -650
rect 1125 -680 1265 -650
rect 1295 -680 1435 -650
rect 1465 -680 1605 -650
rect 1635 -680 1775 -650
rect 1805 -680 1945 -650
rect 1975 -680 2115 -650
rect 2145 -680 2285 -650
rect 2315 -680 2455 -650
rect 2485 -680 2625 -650
rect 2655 -680 2795 -650
rect 2825 -680 2965 -650
rect 2995 -680 3135 -650
rect 3165 -680 3305 -650
rect 3335 -680 3475 -650
rect 3505 -680 3645 -650
rect 3675 -680 3815 -650
rect 3845 -680 3985 -650
rect 4015 -680 4155 -650
rect 4185 -680 4325 -650
rect 4355 -680 4495 -650
rect 4525 -680 4665 -650
rect 4695 -680 4835 -650
rect 4865 -680 5005 -650
rect 5035 -680 5175 -650
rect 5205 -680 5345 -650
rect 5375 -680 5515 -650
rect 5545 -680 5685 -650
rect 5715 -680 5855 -650
rect 5885 -680 6025 -650
rect 6055 -680 6195 -650
rect 6225 -680 6365 -650
rect 6395 -680 6535 -650
rect 6565 -680 6705 -650
rect 6735 -680 6875 -650
rect 6905 -680 7045 -650
rect 7075 -680 7215 -650
rect 7245 -680 7385 -650
rect 7415 -680 7555 -650
rect 7585 -680 7725 -650
rect 7755 -680 7895 -650
rect 7925 -680 8065 -650
rect 8095 -680 8235 -650
rect 8265 -680 8405 -650
rect 8435 -680 8575 -650
rect 8605 -680 8745 -650
rect 8775 -680 8915 -650
rect 8945 -680 9085 -650
rect 9115 -680 9255 -650
rect 9285 -680 9425 -650
rect 9455 -680 9595 -650
rect 9625 -680 9765 -650
rect 9795 -680 9935 -650
rect 9965 -680 10105 -650
rect 10135 -680 10275 -650
rect 10305 -680 10445 -650
rect 10475 -680 10615 -650
rect 10645 -680 10785 -650
rect 10815 -680 10955 -650
rect 10985 -680 11125 -650
rect 11155 -680 11295 -650
rect 11325 -680 11465 -650
rect 11495 -680 11635 -650
rect 11665 -680 11805 -650
rect 11835 -680 11975 -650
rect 12005 -680 12145 -650
rect 12175 -680 12315 -650
rect 12345 -680 12485 -650
rect 12515 -680 12655 -650
rect 12685 -680 12825 -650
rect 12855 -680 12995 -650
rect 13025 -680 13165 -650
rect 13195 -680 13335 -650
rect 13365 -680 13505 -650
rect 13535 -680 13675 -650
rect 13705 -680 13845 -650
rect 13875 -680 14015 -650
rect 14045 -680 14185 -650
rect 14215 -680 14355 -650
rect 14385 -680 14525 -650
rect 14555 -680 14695 -650
rect 14725 -680 14865 -650
rect 14895 -680 15035 -650
rect 15065 -680 15205 -650
rect 15235 -680 15375 -650
rect 15405 -680 15545 -650
rect 15575 -680 15715 -650
rect 15745 -680 15885 -650
rect 15915 -680 16055 -650
rect 16085 -680 16225 -650
rect 16255 -680 16395 -650
rect 16425 -680 16565 -650
rect 16595 -680 16735 -650
rect 16765 -680 16905 -650
rect 16935 -680 17075 -650
rect 17105 -680 17245 -650
rect 17275 -680 17415 -650
rect 17445 -680 17585 -650
rect 17615 -680 17755 -650
rect 17785 -680 17925 -650
rect 17955 -680 18095 -650
rect 18125 -680 18265 -650
rect 18295 -680 18435 -650
rect 18465 -680 18605 -650
rect 18635 -680 18775 -650
rect 18805 -680 18945 -650
rect 18975 -680 19115 -650
rect 19145 -680 19285 -650
rect 19315 -680 19455 -650
rect 19485 -680 19625 -650
rect 19655 -680 19795 -650
rect 19825 -680 19965 -650
rect 19995 -680 20135 -650
rect 20165 -680 20305 -650
rect 20335 -680 20475 -650
rect 20505 -680 20645 -650
rect 20675 -680 20815 -650
rect 20845 -680 20985 -650
rect 21015 -680 21155 -650
rect 21185 -680 21325 -650
rect 21355 -680 21495 -650
rect 21525 -680 21665 -650
rect 21695 -680 21835 -650
rect 21865 -680 22005 -650
rect 22035 -680 22175 -650
rect 22205 -680 22345 -650
rect 22375 -680 22515 -650
rect 22545 -680 22685 -650
rect 22715 -680 22855 -650
rect 22885 -680 23025 -650
rect 23055 -680 23195 -650
rect 23225 -680 23365 -650
rect 23395 -680 23535 -650
rect 23565 -680 23705 -650
rect 23735 -680 23875 -650
rect 23905 -680 24045 -650
rect 24075 -680 24215 -650
rect 24245 -680 24385 -650
rect 24415 -680 24555 -650
rect 24585 -680 24725 -650
rect 24755 -680 24895 -650
rect 24925 -680 25065 -650
rect 25095 -680 25235 -650
rect 25265 -680 25405 -650
rect 25435 -680 25575 -650
rect 25605 -680 25745 -650
rect 25775 -680 25915 -650
rect 25945 -680 26085 -650
rect 26115 -680 26255 -650
rect 26285 -680 26425 -650
rect 26455 -680 26595 -650
rect 26625 -680 26765 -650
rect 26795 -680 26935 -650
rect 26965 -680 27105 -650
rect 27135 -680 27275 -650
rect 27305 -680 27445 -650
rect 27475 -680 27615 -650
rect 27645 -680 27785 -650
rect 27815 -680 27955 -650
rect 27985 -680 28125 -650
rect 28155 -680 28295 -650
rect 28325 -680 28465 -650
rect 28495 -680 28635 -650
rect 28665 -680 28805 -650
rect 28835 -680 28975 -650
rect 29005 -680 29145 -650
rect 29175 -680 29315 -650
rect 29345 -680 29485 -650
rect 29515 -680 29655 -650
rect 29685 -680 29825 -650
rect 29855 -680 29995 -650
rect 30025 -680 30165 -650
rect 30195 -680 30335 -650
rect 30365 -680 30505 -650
rect 30535 -680 30675 -650
rect 30705 -680 30845 -650
rect 30875 -680 31015 -650
rect 31045 -680 31185 -650
rect 31215 -680 31355 -650
rect 31385 -680 31525 -650
rect 31555 -680 31695 -650
rect 31725 -680 31865 -650
rect 31895 -680 32035 -650
rect 32065 -680 32205 -650
rect 32235 -680 32375 -650
rect 32405 -680 32545 -650
rect 32575 -680 32715 -650
rect 32745 -680 32885 -650
rect 32915 -680 33055 -650
rect 33085 -680 33225 -650
rect 33255 -680 33395 -650
rect 33425 -680 33565 -650
rect 33595 -680 33735 -650
rect 33765 -680 33905 -650
rect 33935 -680 34075 -650
rect 34105 -680 34245 -650
rect 34275 -680 34415 -650
rect 34445 -680 34585 -650
rect 34615 -680 34755 -650
rect 34785 -680 34925 -650
rect 34955 -680 35095 -650
rect 35125 -680 35265 -650
rect 35295 -680 35435 -650
rect 35465 -680 35605 -650
rect 35635 -680 35775 -650
rect 35805 -680 35945 -650
rect 35975 -680 36115 -650
rect 36145 -680 36285 -650
rect 36315 -680 36455 -650
rect 36485 -680 36625 -650
rect 36655 -680 36795 -650
rect 36825 -680 36965 -650
rect 36995 -680 37135 -650
rect 37165 -680 37305 -650
rect 37335 -680 37475 -650
rect 37505 -680 37645 -650
rect 37675 -680 37815 -650
rect 37845 -680 37985 -650
rect 38015 -680 38155 -650
rect 38185 -680 38325 -650
rect 38355 -680 38495 -650
rect 38525 -680 38665 -650
rect 38695 -680 38835 -650
rect 38865 -680 39005 -650
rect 39035 -680 39175 -650
rect 39205 -680 39345 -650
rect 39375 -680 39515 -650
rect 39545 -680 39685 -650
rect 39715 -680 39855 -650
rect 39885 -680 40025 -650
rect 40055 -680 40195 -650
rect 40225 -680 40365 -650
rect 40395 -680 40535 -650
rect 40565 -680 40705 -650
rect 40735 -680 40875 -650
rect 40905 -680 41045 -650
rect 41075 -680 41215 -650
rect 41245 -680 41385 -650
rect 41415 -680 41555 -650
rect 41585 -680 41725 -650
rect 41755 -680 41895 -650
rect 41925 -680 42065 -650
rect 42095 -680 42235 -650
rect 42265 -680 42405 -650
rect 42435 -680 42575 -650
rect 42605 -680 42745 -650
rect 42775 -680 42915 -650
rect 42945 -680 43085 -650
rect 43115 -680 43255 -650
rect 43285 -680 43425 -650
rect 43455 -680 43595 -650
rect 43625 -680 43635 -650
rect 65 -690 115 -680
rect 235 -690 285 -680
rect 405 -690 455 -680
rect 575 -690 625 -680
rect 745 -690 795 -680
rect 915 -690 965 -680
rect 1085 -690 1135 -680
rect 1255 -690 1305 -680
rect 1425 -690 1475 -680
rect 1595 -690 1645 -680
rect 1765 -690 1815 -680
rect 1935 -690 1985 -680
rect 2105 -690 2155 -680
rect 2275 -690 2325 -680
rect 2445 -690 2495 -680
rect 2615 -690 2665 -680
rect 2785 -690 2835 -680
rect 2955 -690 3005 -680
rect 3125 -690 3175 -680
rect 3295 -690 3345 -680
rect 3465 -690 3515 -680
rect 3635 -690 3685 -680
rect 3805 -690 3855 -680
rect 3975 -690 4025 -680
rect 4145 -690 4195 -680
rect 4315 -690 4365 -680
rect 4485 -690 4535 -680
rect 4655 -690 4705 -680
rect 4825 -690 4875 -680
rect 4995 -690 5045 -680
rect 5165 -690 5215 -680
rect 5335 -690 5385 -680
rect 5505 -690 5555 -680
rect 5675 -690 5725 -680
rect 5845 -690 5895 -680
rect 6015 -690 6065 -680
rect 6185 -690 6235 -680
rect 6355 -690 6405 -680
rect 6525 -690 6575 -680
rect 6695 -690 6745 -680
rect 6865 -690 6915 -680
rect 7035 -690 7085 -680
rect 7205 -690 7255 -680
rect 7375 -690 7425 -680
rect 7545 -690 7595 -680
rect 7715 -690 7765 -680
rect 7885 -690 7935 -680
rect 8055 -690 8105 -680
rect 8225 -690 8275 -680
rect 8395 -690 8445 -680
rect 8565 -690 8615 -680
rect 8735 -690 8785 -680
rect 8905 -690 8955 -680
rect 9075 -690 9125 -680
rect 9245 -690 9295 -680
rect 9415 -690 9465 -680
rect 9585 -690 9635 -680
rect 9755 -690 9805 -680
rect 9925 -690 9975 -680
rect 10095 -690 10145 -680
rect 10265 -690 10315 -680
rect 10435 -690 10485 -680
rect 10605 -690 10655 -680
rect 10775 -690 10825 -680
rect 10945 -690 10995 -680
rect 11115 -690 11165 -680
rect 11285 -690 11335 -680
rect 11455 -690 11505 -680
rect 11625 -690 11675 -680
rect 11795 -690 11845 -680
rect 11965 -690 12015 -680
rect 12135 -690 12185 -680
rect 12305 -690 12355 -680
rect 12475 -690 12525 -680
rect 12645 -690 12695 -680
rect 12815 -690 12865 -680
rect 12985 -690 13035 -680
rect 13155 -690 13205 -680
rect 13325 -690 13375 -680
rect 13495 -690 13545 -680
rect 13665 -690 13715 -680
rect 13835 -690 13885 -680
rect 14005 -690 14055 -680
rect 14175 -690 14225 -680
rect 14345 -690 14395 -680
rect 14515 -690 14565 -680
rect 14685 -690 14735 -680
rect 14855 -690 14905 -680
rect 15025 -690 15075 -680
rect 15195 -690 15245 -680
rect 15365 -690 15415 -680
rect 15535 -690 15585 -680
rect 15705 -690 15755 -680
rect 15875 -690 15925 -680
rect 16045 -690 16095 -680
rect 16215 -690 16265 -680
rect 16385 -690 16435 -680
rect 16555 -690 16605 -680
rect 16725 -690 16775 -680
rect 16895 -690 16945 -680
rect 17065 -690 17115 -680
rect 17235 -690 17285 -680
rect 17405 -690 17455 -680
rect 17575 -690 17625 -680
rect 17745 -690 17795 -680
rect 17915 -690 17965 -680
rect 18085 -690 18135 -680
rect 18255 -690 18305 -680
rect 18425 -690 18475 -680
rect 18595 -690 18645 -680
rect 18765 -690 18815 -680
rect 18935 -690 18985 -680
rect 19105 -690 19155 -680
rect 19275 -690 19325 -680
rect 19445 -690 19495 -680
rect 19615 -690 19665 -680
rect 19785 -690 19835 -680
rect 19955 -690 20005 -680
rect 20125 -690 20175 -680
rect 20295 -690 20345 -680
rect 20465 -690 20515 -680
rect 20635 -690 20685 -680
rect 20805 -690 20855 -680
rect 20975 -690 21025 -680
rect 21145 -690 21195 -680
rect 21315 -690 21365 -680
rect 21485 -690 21535 -680
rect 21655 -690 21705 -680
rect 21825 -690 21875 -680
rect 21995 -690 22045 -680
rect 22165 -690 22215 -680
rect 22335 -690 22385 -680
rect 22505 -690 22555 -680
rect 22675 -690 22725 -680
rect 22845 -690 22895 -680
rect 23015 -690 23065 -680
rect 23185 -690 23235 -680
rect 23355 -690 23405 -680
rect 23525 -690 23575 -680
rect 23695 -690 23745 -680
rect 23865 -690 23915 -680
rect 24035 -690 24085 -680
rect 24205 -690 24255 -680
rect 24375 -690 24425 -680
rect 24545 -690 24595 -680
rect 24715 -690 24765 -680
rect 24885 -690 24935 -680
rect 25055 -690 25105 -680
rect 25225 -690 25275 -680
rect 25395 -690 25445 -680
rect 25565 -690 25615 -680
rect 25735 -690 25785 -680
rect 25905 -690 25955 -680
rect 26075 -690 26125 -680
rect 26245 -690 26295 -680
rect 26415 -690 26465 -680
rect 26585 -690 26635 -680
rect 26755 -690 26805 -680
rect 26925 -690 26975 -680
rect 27095 -690 27145 -680
rect 27265 -690 27315 -680
rect 27435 -690 27485 -680
rect 27605 -690 27655 -680
rect 27775 -690 27825 -680
rect 27945 -690 27995 -680
rect 28115 -690 28165 -680
rect 28285 -690 28335 -680
rect 28455 -690 28505 -680
rect 28625 -690 28675 -680
rect 28795 -690 28845 -680
rect 28965 -690 29015 -680
rect 29135 -690 29185 -680
rect 29305 -690 29355 -680
rect 29475 -690 29525 -680
rect 29645 -690 29695 -680
rect 29815 -690 29865 -680
rect 29985 -690 30035 -680
rect 30155 -690 30205 -680
rect 30325 -690 30375 -680
rect 30495 -690 30545 -680
rect 30665 -690 30715 -680
rect 30835 -690 30885 -680
rect 31005 -690 31055 -680
rect 31175 -690 31225 -680
rect 31345 -690 31395 -680
rect 31515 -690 31565 -680
rect 31685 -690 31735 -680
rect 31855 -690 31905 -680
rect 32025 -690 32075 -680
rect 32195 -690 32245 -680
rect 32365 -690 32415 -680
rect 32535 -690 32585 -680
rect 32705 -690 32755 -680
rect 32875 -690 32925 -680
rect 33045 -690 33095 -680
rect 33215 -690 33265 -680
rect 33385 -690 33435 -680
rect 33555 -690 33605 -680
rect 33725 -690 33775 -680
rect 33895 -690 33945 -680
rect 34065 -690 34115 -680
rect 34235 -690 34285 -680
rect 34405 -690 34455 -680
rect 34575 -690 34625 -680
rect 34745 -690 34795 -680
rect 34915 -690 34965 -680
rect 35085 -690 35135 -680
rect 35255 -690 35305 -680
rect 35425 -690 35475 -680
rect 35595 -690 35645 -680
rect 35765 -690 35815 -680
rect 35935 -690 35985 -680
rect 36105 -690 36155 -680
rect 36275 -690 36325 -680
rect 36445 -690 36495 -680
rect 36615 -690 36665 -680
rect 36785 -690 36835 -680
rect 36955 -690 37005 -680
rect 37125 -690 37175 -680
rect 37295 -690 37345 -680
rect 37465 -690 37515 -680
rect 37635 -690 37685 -680
rect 37805 -690 37855 -680
rect 37975 -690 38025 -680
rect 38145 -690 38195 -680
rect 38315 -690 38365 -680
rect 38485 -690 38535 -680
rect 38655 -690 38705 -680
rect 38825 -690 38875 -680
rect 38995 -690 39045 -680
rect 39165 -690 39215 -680
rect 39335 -690 39385 -680
rect 39505 -690 39555 -680
rect 39675 -690 39725 -680
rect 39845 -690 39895 -680
rect 40015 -690 40065 -680
rect 40185 -690 40235 -680
rect 40355 -690 40405 -680
rect 40525 -690 40575 -680
rect 40695 -690 40745 -680
rect 40865 -690 40915 -680
rect 41035 -690 41085 -680
rect 41205 -690 41255 -680
rect 41375 -690 41425 -680
rect 41545 -690 41595 -680
rect 41715 -690 41765 -680
rect 41885 -690 41935 -680
rect 42055 -690 42105 -680
rect 42225 -690 42275 -680
rect 42395 -690 42445 -680
rect 42565 -690 42615 -680
rect 42735 -690 42785 -680
rect 42905 -690 42955 -680
rect 43075 -690 43125 -680
rect 43245 -690 43295 -680
rect 43415 -690 43465 -680
rect 43585 -690 43635 -680
<< via2 >>
rect 225 175 255 205
rect 565 175 595 205
rect 760 175 790 205
rect 1440 175 1470 205
rect 2120 175 2150 205
rect 2270 175 2300 205
rect 2950 175 2980 205
rect 3630 175 3660 205
rect 4310 175 4340 205
rect 4990 175 5020 205
rect 5670 175 5700 205
rect 6350 175 6380 205
rect 7030 175 7060 205
rect 7710 175 7740 205
rect 7860 175 7890 205
rect 8540 175 8570 205
rect 9220 175 9250 205
rect 9900 175 9930 205
rect 10580 175 10610 205
rect 11260 175 11290 205
rect 11940 175 11970 205
rect 12620 175 12650 205
rect 13300 175 13330 205
rect 13980 175 14010 205
rect 14660 175 14690 205
rect 15340 175 15370 205
rect 16020 175 16050 205
rect 16700 175 16730 205
rect 17380 175 17410 205
rect 18060 175 18090 205
rect 18740 175 18770 205
rect 19420 175 19450 205
rect 20100 175 20130 205
rect 20780 175 20810 205
rect 21460 175 21490 205
rect 22140 175 22170 205
rect 22820 175 22850 205
rect 23500 175 23530 205
rect 24180 175 24210 205
rect 24860 175 24890 205
rect 25540 175 25570 205
rect 26220 175 26250 205
rect 26900 175 26930 205
rect 27580 175 27610 205
rect 28260 175 28290 205
rect 28940 175 28970 205
rect 29620 175 29650 205
rect 310 65 340 100
rect 480 65 510 100
rect 845 65 875 100
rect 1015 65 1045 100
rect 1185 65 1215 100
rect 1355 65 1385 100
rect 1525 65 1555 100
rect 1695 65 1725 100
rect 1865 65 1895 100
rect 2035 65 2065 100
rect 2355 65 2385 100
rect 2525 65 2555 100
rect 2695 65 2725 100
rect 2865 65 2895 100
rect 3035 65 3065 100
rect 3205 65 3235 100
rect 3375 65 3405 100
rect 3545 65 3575 100
rect 3715 65 3745 100
rect 3885 65 3915 100
rect 4055 65 4085 100
rect 4225 65 4255 100
rect 4395 65 4425 100
rect 4565 65 4595 100
rect 4735 65 4765 100
rect 4905 65 4935 100
rect 5075 65 5105 100
rect 5245 65 5275 100
rect 5415 65 5445 100
rect 5585 65 5615 100
rect 5755 65 5785 100
rect 5925 65 5955 100
rect 6095 65 6125 100
rect 6265 65 6295 100
rect 6435 65 6465 100
rect 6605 65 6635 100
rect 6775 65 6805 100
rect 6945 65 6975 100
rect 7115 65 7145 100
rect 7285 65 7315 100
rect 7455 65 7485 100
rect 7625 65 7655 100
rect 7945 65 7975 100
rect 8115 65 8145 100
rect 8285 65 8315 100
rect 8455 65 8485 100
rect 8625 65 8655 100
rect 8795 65 8825 100
rect 8965 65 8995 100
rect 9135 65 9165 100
rect 9305 65 9335 100
rect 9475 65 9505 100
rect 9645 65 9675 100
rect 9815 65 9845 100
rect 9985 65 10015 100
rect 10155 65 10185 100
rect 10325 65 10355 100
rect 10495 65 10525 100
rect 10665 65 10695 100
rect 10835 65 10865 100
rect 11005 65 11035 100
rect 11175 65 11205 100
rect 11345 65 11375 100
rect 11515 65 11545 100
rect 11685 65 11715 100
rect 11855 65 11885 100
rect 12025 65 12055 100
rect 12195 65 12225 100
rect 12365 65 12395 100
rect 12535 65 12565 100
rect 12705 65 12735 100
rect 12875 65 12905 100
rect 13045 65 13075 100
rect 13215 65 13245 100
rect 13385 65 13415 100
rect 13555 65 13585 100
rect 13725 65 13755 100
rect 13895 65 13925 100
rect 14065 65 14095 100
rect 14235 65 14265 100
rect 14405 65 14435 100
rect 14575 65 14605 100
rect 14745 65 14775 100
rect 14915 65 14945 100
rect 15085 65 15115 100
rect 15255 65 15285 100
rect 15425 65 15455 100
rect 15595 65 15625 100
rect 15765 65 15795 100
rect 15935 65 15965 100
rect 16105 65 16135 100
rect 16275 65 16305 100
rect 16445 65 16475 100
rect 16615 65 16645 100
rect 16785 65 16815 100
rect 16955 65 16985 100
rect 17125 65 17155 100
rect 17295 65 17325 100
rect 17465 65 17495 100
rect 17635 65 17665 100
rect 17805 65 17835 100
rect 17975 65 18005 100
rect 18145 65 18175 100
rect 18315 65 18345 100
rect 18485 65 18515 100
rect 18655 65 18685 100
rect 18825 65 18855 100
rect 18995 65 19025 100
rect 19165 65 19195 100
rect 19335 65 19365 100
rect 19505 65 19535 100
rect 19675 65 19705 100
rect 19845 65 19875 100
rect 20015 65 20045 100
rect 20185 65 20215 100
rect 20355 65 20385 100
rect 20525 65 20555 100
rect 20695 65 20725 100
rect 20865 65 20895 100
rect 21035 65 21065 100
rect 21205 65 21235 100
rect 21375 65 21405 100
rect 21545 65 21575 100
rect 21715 65 21745 100
rect 21885 65 21915 100
rect 22055 65 22085 100
rect 22225 65 22255 100
rect 22395 65 22425 100
rect 22565 65 22595 100
rect 22735 65 22765 100
rect 22905 65 22935 100
rect 23075 65 23105 100
rect 23245 65 23275 100
rect 23415 65 23445 100
rect 23585 65 23615 100
rect 23755 65 23785 100
rect 23925 65 23955 100
rect 24095 65 24125 100
rect 24265 65 24295 100
rect 24435 65 24465 100
rect 24605 65 24635 100
rect 24775 65 24805 100
rect 24945 65 24975 100
rect 25115 65 25145 100
rect 25285 65 25315 100
rect 25455 65 25485 100
rect 25625 65 25655 100
rect 25795 65 25825 100
rect 25965 65 25995 100
rect 26135 65 26165 100
rect 26305 65 26335 100
rect 26475 65 26505 100
rect 26645 65 26675 100
rect 26815 65 26845 100
rect 26985 65 27015 100
rect 27155 65 27185 100
rect 27325 65 27355 100
rect 27495 65 27525 100
rect 27665 65 27695 100
rect 27835 65 27865 100
rect 28005 65 28035 100
rect 28175 65 28205 100
rect 28345 65 28375 100
rect 28515 65 28545 100
rect 28685 65 28715 100
rect 28855 65 28885 100
rect 29025 65 29055 100
rect 29195 65 29225 100
rect 29365 65 29395 100
rect 29535 65 29565 100
rect 225 10 255 40
rect 565 10 595 40
rect 760 10 790 40
rect 1440 10 1470 40
rect 2440 10 2470 40
rect 3120 10 3150 40
rect 3630 10 3660 40
rect 4310 10 4340 40
rect 4990 10 5020 40
rect 5500 10 5530 40
rect 8200 10 8230 40
rect 8880 10 8910 40
rect 9390 10 9420 40
rect 10070 10 10100 40
rect 10750 10 10780 40
rect 11260 10 11290 40
rect 11940 10 11970 40
rect 12280 10 12310 40
rect 14150 10 14180 40
rect 14830 10 14860 40
rect 15340 10 15370 40
rect 16020 10 16050 40
rect 16700 10 16730 40
rect 17210 10 17240 40
rect 17890 10 17920 40
rect 18230 10 18260 40
rect 21290 10 21320 40
rect 22310 10 22340 40
rect 24180 10 24210 40
rect 24860 10 24890 40
rect 25370 10 25400 40
rect 26050 10 26080 40
rect 26730 10 26760 40
rect 27750 10 27780 40
rect 650 -65 700 -25
rect 2190 -65 2240 -25
rect 7780 -65 7830 -25
rect 7965 -260 8000 -230
rect 15615 -260 15650 -230
rect 29555 -260 29590 -230
rect 75 -365 105 -335
rect 755 -365 785 -335
rect 1435 -365 1465 -335
rect 2285 -365 2315 -335
rect 2965 -365 2995 -335
rect 3475 -365 3505 -335
rect 4155 -365 4185 -335
rect 4835 -365 4865 -335
rect 5345 -365 5375 -335
rect 5855 -365 5885 -335
rect 6535 -365 6565 -335
rect 7215 -365 7245 -335
rect 8065 -365 8095 -335
rect 8745 -365 8775 -335
rect 9255 -365 9285 -335
rect 9935 -365 9965 -335
rect 10615 -365 10645 -335
rect 11125 -365 11155 -335
rect 11805 -365 11835 -335
rect 12485 -365 12515 -335
rect 13165 -365 13195 -335
rect 14015 -365 14045 -335
rect 14695 -365 14725 -335
rect 15205 -365 15235 -335
rect 15885 -365 15915 -335
rect 16565 -365 16595 -335
rect 17075 -365 17105 -335
rect 17755 -365 17785 -335
rect 18435 -365 18465 -335
rect 19115 -365 19145 -335
rect 19965 -365 19995 -335
rect 20645 -365 20675 -335
rect 21155 -365 21185 -335
rect 21835 -365 21865 -335
rect 22515 -365 22545 -335
rect 23195 -365 23225 -335
rect 24045 -365 24075 -335
rect 24725 -365 24755 -335
rect 25235 -365 25265 -335
rect 25915 -365 25945 -335
rect 26595 -365 26625 -335
rect 27105 -365 27135 -335
rect 27615 -365 27645 -335
rect 28295 -365 28325 -335
rect 28975 -365 29005 -335
rect 29825 -365 29855 -335
rect 30505 -365 30535 -335
rect 31015 -365 31045 -335
rect 31695 -365 31725 -335
rect 32375 -365 32405 -335
rect 32885 -365 32915 -335
rect 33565 -365 33595 -335
rect 34245 -365 34275 -335
rect 34925 -365 34955 -335
rect 35775 -365 35805 -335
rect 36455 -365 36485 -335
rect 36965 -365 36995 -335
rect 37645 -365 37675 -335
rect 38325 -365 38355 -335
rect 38835 -365 38865 -335
rect 39515 -365 39545 -335
rect 40195 -365 40225 -335
rect 40875 -365 40905 -335
rect 41725 -365 41755 -335
rect 42405 -365 42435 -335
rect 42915 -365 42945 -335
rect 43595 -365 43625 -335
rect 160 -475 190 -440
rect 330 -475 360 -440
rect 500 -475 530 -440
rect 670 -475 700 -440
rect 840 -475 870 -440
rect 1010 -475 1040 -440
rect 1180 -475 1210 -440
rect 1350 -475 1380 -440
rect 1520 -475 1550 -440
rect 1690 -475 1720 -440
rect 1860 -475 1890 -440
rect 2030 -475 2060 -440
rect 2200 -475 2230 -440
rect 2370 -475 2400 -440
rect 2540 -475 2570 -440
rect 2710 -475 2740 -440
rect 2880 -475 2910 -440
rect 3050 -475 3080 -440
rect 3220 -475 3250 -440
rect 3390 -475 3420 -440
rect 3560 -475 3590 -440
rect 3730 -475 3760 -440
rect 3900 -475 3930 -440
rect 4070 -475 4100 -440
rect 4240 -475 4270 -440
rect 4410 -475 4440 -440
rect 4580 -475 4610 -440
rect 4750 -475 4780 -440
rect 4920 -475 4950 -440
rect 5090 -475 5120 -440
rect 5260 -475 5290 -440
rect 5430 -475 5460 -440
rect 5600 -475 5630 -440
rect 5770 -475 5800 -440
rect 5940 -475 5970 -440
rect 6110 -475 6140 -440
rect 6280 -475 6310 -440
rect 6450 -475 6480 -440
rect 6620 -475 6650 -440
rect 6790 -475 6820 -440
rect 6960 -475 6990 -440
rect 7130 -475 7160 -440
rect 7300 -475 7330 -440
rect 7470 -475 7500 -440
rect 7640 -475 7670 -440
rect 7810 -475 7840 -440
rect 7980 -475 8010 -440
rect 8150 -475 8180 -440
rect 8320 -475 8350 -440
rect 8490 -475 8520 -440
rect 8660 -475 8690 -440
rect 8830 -475 8860 -440
rect 9000 -475 9030 -440
rect 9170 -475 9200 -440
rect 9340 -475 9370 -440
rect 9510 -475 9540 -440
rect 9680 -475 9710 -440
rect 9850 -475 9880 -440
rect 10020 -475 10050 -440
rect 10190 -475 10220 -440
rect 10360 -475 10390 -440
rect 10530 -475 10560 -440
rect 10700 -475 10730 -440
rect 10870 -475 10900 -440
rect 11040 -475 11070 -440
rect 11210 -475 11240 -440
rect 11380 -475 11410 -440
rect 11550 -475 11580 -440
rect 11720 -475 11750 -440
rect 11890 -475 11920 -440
rect 12060 -475 12090 -440
rect 12230 -475 12260 -440
rect 12400 -475 12430 -440
rect 12570 -475 12600 -440
rect 12740 -475 12770 -440
rect 12910 -475 12940 -440
rect 13080 -475 13110 -440
rect 13250 -475 13280 -440
rect 13420 -475 13450 -440
rect 13590 -475 13620 -440
rect 13760 -475 13790 -440
rect 13930 -475 13960 -440
rect 14100 -475 14130 -440
rect 14270 -475 14300 -440
rect 14440 -475 14470 -440
rect 14610 -475 14640 -440
rect 14780 -475 14810 -440
rect 14950 -475 14980 -440
rect 15120 -475 15150 -440
rect 15290 -475 15320 -440
rect 15460 -475 15490 -440
rect 15630 -475 15660 -440
rect 15800 -475 15830 -440
rect 15970 -475 16000 -440
rect 16140 -475 16170 -440
rect 16310 -475 16340 -440
rect 16480 -475 16510 -440
rect 16650 -475 16680 -440
rect 16820 -475 16850 -440
rect 16990 -475 17020 -440
rect 17160 -475 17190 -440
rect 17330 -475 17360 -440
rect 17500 -475 17530 -440
rect 17670 -475 17700 -440
rect 17840 -475 17870 -440
rect 18010 -475 18040 -440
rect 18180 -475 18210 -440
rect 18350 -475 18380 -440
rect 18520 -475 18550 -440
rect 18690 -475 18720 -440
rect 18860 -475 18890 -440
rect 19030 -475 19060 -440
rect 19200 -475 19230 -440
rect 19370 -475 19400 -440
rect 19540 -475 19570 -440
rect 19710 -475 19740 -440
rect 19880 -475 19910 -440
rect 20050 -475 20080 -440
rect 20220 -475 20250 -440
rect 20390 -475 20420 -440
rect 20560 -475 20590 -440
rect 20730 -475 20760 -440
rect 20900 -475 20930 -440
rect 21070 -475 21100 -440
rect 21240 -475 21270 -440
rect 21410 -475 21440 -440
rect 21580 -475 21610 -440
rect 21750 -475 21780 -440
rect 21920 -475 21950 -440
rect 22090 -475 22120 -440
rect 22260 -475 22290 -440
rect 22430 -475 22460 -440
rect 22600 -475 22630 -440
rect 22770 -475 22800 -440
rect 22940 -475 22970 -440
rect 23110 -475 23140 -440
rect 23280 -475 23310 -440
rect 23450 -475 23480 -440
rect 23620 -475 23650 -440
rect 23790 -475 23820 -440
rect 23960 -475 23990 -440
rect 24130 -475 24160 -440
rect 24300 -475 24330 -440
rect 24470 -475 24500 -440
rect 24640 -475 24670 -440
rect 24810 -475 24840 -440
rect 24980 -475 25010 -440
rect 25150 -475 25180 -440
rect 25320 -475 25350 -440
rect 25490 -475 25520 -440
rect 25660 -475 25690 -440
rect 25830 -475 25860 -440
rect 26000 -475 26030 -440
rect 26170 -475 26200 -440
rect 26340 -475 26370 -440
rect 26510 -475 26540 -440
rect 26680 -475 26710 -440
rect 26850 -475 26880 -440
rect 27020 -475 27050 -440
rect 27190 -475 27220 -440
rect 27360 -475 27390 -440
rect 27530 -475 27560 -440
rect 27700 -475 27730 -440
rect 27870 -475 27900 -440
rect 28040 -475 28070 -440
rect 28210 -475 28240 -440
rect 28380 -475 28410 -440
rect 28550 -475 28580 -440
rect 28720 -475 28750 -440
rect 28890 -475 28920 -440
rect 29060 -475 29090 -440
rect 29230 -475 29260 -440
rect 29400 -475 29430 -440
rect 29570 -475 29600 -440
rect 29740 -475 29770 -440
rect 29910 -475 29940 -440
rect 30080 -475 30110 -440
rect 30250 -475 30280 -440
rect 30420 -475 30450 -440
rect 30590 -475 30620 -440
rect 30760 -475 30790 -440
rect 30930 -475 30960 -440
rect 31100 -475 31130 -440
rect 31270 -475 31300 -440
rect 31440 -475 31470 -440
rect 31610 -475 31640 -440
rect 31780 -475 31810 -440
rect 31950 -475 31980 -440
rect 32120 -475 32150 -440
rect 32290 -475 32320 -440
rect 32460 -475 32490 -440
rect 32630 -475 32660 -440
rect 32800 -475 32830 -440
rect 32970 -475 33000 -440
rect 33140 -475 33170 -440
rect 33310 -475 33340 -440
rect 33480 -475 33510 -440
rect 33650 -475 33680 -440
rect 33820 -475 33850 -440
rect 33990 -475 34020 -440
rect 34160 -475 34190 -440
rect 34330 -475 34360 -440
rect 34500 -475 34530 -440
rect 34670 -475 34700 -440
rect 34840 -475 34870 -440
rect 35010 -475 35040 -440
rect 35180 -475 35210 -440
rect 35350 -475 35380 -440
rect 35520 -475 35550 -440
rect 35690 -475 35720 -440
rect 35860 -475 35890 -440
rect 36030 -475 36060 -440
rect 36200 -475 36230 -440
rect 36370 -475 36400 -440
rect 36540 -475 36570 -440
rect 36710 -475 36740 -440
rect 36880 -475 36910 -440
rect 37050 -475 37080 -440
rect 37220 -475 37250 -440
rect 37390 -475 37420 -440
rect 37560 -475 37590 -440
rect 37730 -475 37760 -440
rect 37900 -475 37930 -440
rect 38070 -475 38100 -440
rect 38240 -475 38270 -440
rect 38410 -475 38440 -440
rect 38580 -475 38610 -440
rect 38750 -475 38780 -440
rect 38920 -475 38950 -440
rect 39090 -475 39120 -440
rect 39260 -475 39290 -440
rect 39430 -475 39460 -440
rect 39600 -475 39630 -440
rect 39770 -475 39800 -440
rect 39940 -475 39970 -440
rect 40110 -475 40140 -440
rect 40280 -475 40310 -440
rect 40450 -475 40480 -440
rect 40620 -475 40650 -440
rect 40790 -475 40820 -440
rect 40960 -475 40990 -440
rect 41130 -475 41160 -440
rect 41300 -475 41330 -440
rect 41470 -475 41500 -440
rect 41640 -475 41670 -440
rect 41810 -475 41840 -440
rect 41980 -475 42010 -440
rect 42150 -475 42180 -440
rect 42320 -475 42350 -440
rect 42490 -475 42520 -440
rect 42660 -475 42690 -440
rect 42830 -475 42860 -440
rect 43000 -475 43030 -440
rect 43170 -475 43200 -440
rect 43340 -475 43370 -440
rect 43510 -475 43540 -440
rect 75 -580 105 -550
rect 755 -580 785 -550
rect 1435 -580 1465 -550
rect 2115 -580 2145 -550
rect 2795 -580 2825 -550
rect 3475 -580 3505 -550
rect 4155 -580 4185 -550
rect 4835 -580 4865 -550
rect 5515 -580 5545 -550
rect 6195 -580 6225 -550
rect 6875 -580 6905 -550
rect 7555 -580 7585 -550
rect 8235 -580 8265 -550
rect 8915 -580 8945 -550
rect 9595 -580 9625 -550
rect 10275 -580 10305 -550
rect 10955 -580 10985 -550
rect 11635 -580 11665 -550
rect 12315 -580 12345 -550
rect 12995 -580 13025 -550
rect 13675 -580 13705 -550
rect 14355 -580 14385 -550
rect 15035 -580 15065 -550
rect 15715 -580 15745 -550
rect 16395 -580 16425 -550
rect 17075 -580 17105 -550
rect 17755 -580 17785 -550
rect 18435 -580 18465 -550
rect 19115 -580 19145 -550
rect 19795 -580 19825 -550
rect 20475 -580 20505 -550
rect 21155 -580 21185 -550
rect 21835 -580 21865 -550
rect 22515 -580 22545 -550
rect 23195 -580 23225 -550
rect 23875 -580 23905 -550
rect 24555 -580 24585 -550
rect 25235 -580 25265 -550
rect 25915 -580 25945 -550
rect 26595 -580 26625 -550
rect 27275 -580 27305 -550
rect 27955 -580 27985 -550
rect 28635 -580 28665 -550
rect 29315 -580 29345 -550
rect 29995 -580 30025 -550
rect 30675 -580 30705 -550
rect 31355 -580 31385 -550
rect 32035 -580 32065 -550
rect 32715 -580 32745 -550
rect 33395 -580 33425 -550
rect 34075 -580 34105 -550
rect 34755 -580 34785 -550
rect 35435 -580 35465 -550
rect 36115 -580 36145 -550
rect 36795 -580 36825 -550
rect 37475 -580 37505 -550
rect 38155 -580 38185 -550
rect 38835 -580 38865 -550
rect 39515 -580 39545 -550
rect 40195 -580 40225 -550
rect 40875 -580 40905 -550
rect 41555 -580 41585 -550
rect 42235 -580 42265 -550
rect 42915 -580 42945 -550
rect 75 -680 105 -650
rect 755 -680 785 -650
rect 1435 -680 1465 -650
rect 2115 -680 2145 -650
rect 2795 -680 2825 -650
rect 3475 -680 3505 -650
rect 4155 -680 4185 -650
rect 4835 -680 4865 -650
rect 5515 -680 5545 -650
rect 6195 -680 6225 -650
rect 6875 -680 6905 -650
rect 7555 -680 7585 -650
rect 8235 -680 8265 -650
rect 8915 -680 8945 -650
rect 9595 -680 9625 -650
rect 10275 -680 10305 -650
rect 10955 -680 10985 -650
rect 11635 -680 11665 -650
rect 12315 -680 12345 -650
rect 12995 -680 13025 -650
rect 13675 -680 13705 -650
rect 14355 -680 14385 -650
rect 15035 -680 15065 -650
rect 15715 -680 15745 -650
rect 16395 -680 16425 -650
rect 17075 -680 17105 -650
rect 17755 -680 17785 -650
rect 18435 -680 18465 -650
rect 19115 -680 19145 -650
rect 19795 -680 19825 -650
rect 20475 -680 20505 -650
rect 21155 -680 21185 -650
rect 21835 -680 21865 -650
rect 22515 -680 22545 -650
rect 23195 -680 23225 -650
rect 23875 -680 23905 -650
rect 24555 -680 24585 -650
rect 25235 -680 25265 -650
rect 25915 -680 25945 -650
rect 26595 -680 26625 -650
rect 27275 -680 27305 -650
rect 27955 -680 27985 -650
rect 28635 -680 28665 -650
rect 29315 -680 29345 -650
rect 29995 -680 30025 -650
rect 30675 -680 30705 -650
rect 31355 -680 31385 -650
rect 32035 -680 32065 -650
rect 32715 -680 32745 -650
rect 33395 -680 33425 -650
rect 34075 -680 34105 -650
rect 34755 -680 34785 -650
rect 35435 -680 35465 -650
rect 36115 -680 36145 -650
rect 36795 -680 36825 -650
rect 37475 -680 37505 -650
rect 38155 -680 38185 -650
rect 38835 -680 38865 -650
rect 39515 -680 39545 -650
rect 40195 -680 40225 -650
rect 40875 -680 40905 -650
rect 41555 -680 41585 -650
rect 42235 -680 42265 -650
rect 42915 -680 42945 -650
<< metal3 >>
rect 200 285 280 290
rect 200 240 210 285
rect 270 240 280 285
rect 200 235 280 240
rect 540 285 620 290
rect 540 240 550 285
rect 610 240 620 285
rect 540 235 620 240
rect 735 285 815 290
rect 735 240 745 285
rect 805 240 815 285
rect 735 235 815 240
rect 1415 285 1495 290
rect 1415 240 1425 285
rect 1485 240 1495 285
rect 1415 235 1495 240
rect 2095 285 2175 290
rect 2095 240 2105 285
rect 2165 240 2175 285
rect 2095 235 2175 240
rect 2245 285 2325 290
rect 2245 240 2255 285
rect 2315 240 2325 285
rect 2245 235 2325 240
rect 2925 285 3005 290
rect 2925 240 2935 285
rect 2995 240 3005 285
rect 2925 235 3005 240
rect 3605 285 3685 290
rect 3605 240 3615 285
rect 3675 240 3685 285
rect 3605 235 3685 240
rect 4285 285 4365 290
rect 4285 240 4295 285
rect 4355 240 4365 285
rect 4285 235 4365 240
rect 4965 285 5045 290
rect 4965 240 4975 285
rect 5035 240 5045 285
rect 4965 235 5045 240
rect 5645 285 5725 290
rect 5645 240 5655 285
rect 5715 240 5725 285
rect 5645 235 5725 240
rect 6325 285 6405 290
rect 6325 240 6335 285
rect 6395 240 6405 285
rect 6325 235 6405 240
rect 7005 285 7085 290
rect 7005 240 7015 285
rect 7075 240 7085 285
rect 7005 235 7085 240
rect 7685 285 7765 290
rect 7685 240 7695 285
rect 7755 240 7765 285
rect 7685 235 7765 240
rect 7835 285 7915 290
rect 7835 240 7845 285
rect 7905 240 7915 285
rect 7835 235 7915 240
rect 8515 285 8595 290
rect 8515 240 8525 285
rect 8585 240 8595 285
rect 8515 235 8595 240
rect 9195 285 9275 290
rect 9195 240 9205 285
rect 9265 240 9275 285
rect 9195 235 9275 240
rect 9875 285 9955 290
rect 9875 240 9885 285
rect 9945 240 9955 285
rect 9875 235 9955 240
rect 10555 285 10635 290
rect 10555 240 10565 285
rect 10625 240 10635 285
rect 10555 235 10635 240
rect 11235 285 11315 290
rect 11235 240 11245 285
rect 11305 240 11315 285
rect 11235 235 11315 240
rect 11915 285 11995 290
rect 11915 240 11925 285
rect 11985 240 11995 285
rect 11915 235 11995 240
rect 12595 285 12675 290
rect 12595 240 12605 285
rect 12665 240 12675 285
rect 12595 235 12675 240
rect 13275 285 13355 290
rect 13275 240 13285 285
rect 13345 240 13355 285
rect 13275 235 13355 240
rect 13955 285 14035 290
rect 13955 240 13965 285
rect 14025 240 14035 285
rect 13955 235 14035 240
rect 14635 285 14715 290
rect 14635 240 14645 285
rect 14705 240 14715 285
rect 14635 235 14715 240
rect 15315 285 15395 290
rect 15315 240 15325 285
rect 15385 240 15395 285
rect 15315 235 15395 240
rect 15995 285 16075 290
rect 15995 240 16005 285
rect 16065 240 16075 285
rect 15995 235 16075 240
rect 16675 285 16755 290
rect 16675 240 16685 285
rect 16745 240 16755 285
rect 16675 235 16755 240
rect 17355 285 17435 290
rect 17355 240 17365 285
rect 17425 240 17435 285
rect 17355 235 17435 240
rect 18035 285 18115 290
rect 18035 240 18045 285
rect 18105 240 18115 285
rect 18035 235 18115 240
rect 18715 285 18795 290
rect 18715 240 18725 285
rect 18785 240 18795 285
rect 18715 235 18795 240
rect 19395 285 19475 290
rect 19395 240 19405 285
rect 19465 240 19475 285
rect 19395 235 19475 240
rect 20075 285 20155 290
rect 20075 240 20085 285
rect 20145 240 20155 285
rect 20075 235 20155 240
rect 20755 285 20835 290
rect 20755 240 20765 285
rect 20825 240 20835 285
rect 20755 235 20835 240
rect 21435 285 21515 290
rect 21435 240 21445 285
rect 21505 240 21515 285
rect 21435 235 21515 240
rect 22115 285 22195 290
rect 22115 240 22125 285
rect 22185 240 22195 285
rect 22115 235 22195 240
rect 22795 285 22875 290
rect 22795 240 22805 285
rect 22865 240 22875 285
rect 22795 235 22875 240
rect 23475 285 23555 290
rect 23475 240 23485 285
rect 23545 240 23555 285
rect 23475 235 23555 240
rect 24155 285 24235 290
rect 24155 240 24165 285
rect 24225 240 24235 285
rect 24155 235 24235 240
rect 24835 285 24915 290
rect 24835 240 24845 285
rect 24905 240 24915 285
rect 24835 235 24915 240
rect 25515 285 25595 290
rect 25515 240 25525 285
rect 25585 240 25595 285
rect 25515 235 25595 240
rect 26195 285 26275 290
rect 26195 240 26205 285
rect 26265 240 26275 285
rect 26195 235 26275 240
rect 26875 285 26955 290
rect 26875 240 26885 285
rect 26945 240 26955 285
rect 26875 235 26955 240
rect 27555 285 27635 290
rect 27555 240 27565 285
rect 27625 240 27635 285
rect 27555 235 27635 240
rect 28235 285 28315 290
rect 28235 240 28245 285
rect 28305 240 28315 285
rect 28235 235 28315 240
rect 28915 285 28995 290
rect 28915 240 28925 285
rect 28985 240 28995 285
rect 28915 235 28995 240
rect 29595 285 29670 290
rect 29595 240 29605 285
rect 29665 240 29670 285
rect 29595 235 29670 240
rect 215 205 265 235
rect 215 175 225 205
rect 255 175 265 205
rect 215 165 265 175
rect 555 205 605 235
rect 555 175 565 205
rect 595 175 605 205
rect 555 165 605 175
rect 750 205 800 235
rect 750 175 760 205
rect 790 175 800 205
rect 750 165 800 175
rect 1430 205 1480 235
rect 1430 175 1440 205
rect 1470 175 1480 205
rect 1430 165 1480 175
rect 2110 205 2160 235
rect 2110 175 2120 205
rect 2150 175 2160 205
rect 2110 165 2160 175
rect 2260 205 2310 235
rect 2260 175 2270 205
rect 2300 175 2310 205
rect 2260 165 2310 175
rect 2940 205 2990 235
rect 2940 175 2950 205
rect 2980 175 2990 205
rect 2940 165 2990 175
rect 3620 205 3670 235
rect 3620 175 3630 205
rect 3660 175 3670 205
rect 3620 165 3670 175
rect 4300 205 4350 235
rect 4300 175 4310 205
rect 4340 175 4350 205
rect 4300 165 4350 175
rect 4980 205 5030 235
rect 4980 175 4990 205
rect 5020 175 5030 205
rect 4980 165 5030 175
rect 5660 205 5710 235
rect 5660 175 5670 205
rect 5700 175 5710 205
rect 5660 165 5710 175
rect 6340 205 6390 235
rect 6340 175 6350 205
rect 6380 175 6390 205
rect 6340 165 6390 175
rect 7020 205 7070 235
rect 7020 175 7030 205
rect 7060 175 7070 205
rect 7020 165 7070 175
rect 7700 205 7750 235
rect 7700 175 7710 205
rect 7740 175 7750 205
rect 7700 165 7750 175
rect 7850 205 7900 235
rect 7850 175 7860 205
rect 7890 175 7900 205
rect 7850 165 7900 175
rect 8530 205 8580 235
rect 8530 175 8540 205
rect 8570 175 8580 205
rect 8530 165 8580 175
rect 9210 205 9260 235
rect 9210 175 9220 205
rect 9250 175 9260 205
rect 9210 165 9260 175
rect 9890 205 9940 235
rect 9890 175 9900 205
rect 9930 175 9940 205
rect 9890 165 9940 175
rect 10570 205 10620 235
rect 10570 175 10580 205
rect 10610 175 10620 205
rect 10570 165 10620 175
rect 11250 205 11300 235
rect 11250 175 11260 205
rect 11290 175 11300 205
rect 11250 165 11300 175
rect 11930 205 11980 235
rect 11930 175 11940 205
rect 11970 175 11980 205
rect 11930 165 11980 175
rect 12610 205 12660 235
rect 12610 175 12620 205
rect 12650 175 12660 205
rect 12610 165 12660 175
rect 13290 205 13340 235
rect 13290 175 13300 205
rect 13330 175 13340 205
rect 13290 165 13340 175
rect 13970 205 14020 235
rect 13970 175 13980 205
rect 14010 175 14020 205
rect 13970 165 14020 175
rect 14650 205 14700 235
rect 14650 175 14660 205
rect 14690 175 14700 205
rect 14650 165 14700 175
rect 15330 205 15380 235
rect 15330 175 15340 205
rect 15370 175 15380 205
rect 15330 165 15380 175
rect 16010 205 16060 235
rect 16010 175 16020 205
rect 16050 175 16060 205
rect 16010 165 16060 175
rect 16690 205 16740 235
rect 16690 175 16700 205
rect 16730 175 16740 205
rect 16690 165 16740 175
rect 17370 205 17420 235
rect 17370 175 17380 205
rect 17410 175 17420 205
rect 17370 165 17420 175
rect 18050 205 18100 235
rect 18050 175 18060 205
rect 18090 175 18100 205
rect 18050 165 18100 175
rect 18730 205 18780 235
rect 18730 175 18740 205
rect 18770 175 18780 205
rect 18730 165 18780 175
rect 19410 205 19460 235
rect 19410 175 19420 205
rect 19450 175 19460 205
rect 19410 165 19460 175
rect 20090 205 20140 235
rect 20090 175 20100 205
rect 20130 175 20140 205
rect 20090 165 20140 175
rect 20770 205 20820 235
rect 20770 175 20780 205
rect 20810 175 20820 205
rect 20770 165 20820 175
rect 21450 205 21500 235
rect 21450 175 21460 205
rect 21490 175 21500 205
rect 21450 165 21500 175
rect 22130 205 22180 235
rect 22130 175 22140 205
rect 22170 175 22180 205
rect 22130 165 22180 175
rect 22810 205 22860 235
rect 22810 175 22820 205
rect 22850 175 22860 205
rect 22810 165 22860 175
rect 23490 205 23540 235
rect 23490 175 23500 205
rect 23530 175 23540 205
rect 23490 165 23540 175
rect 24170 205 24220 235
rect 24170 175 24180 205
rect 24210 175 24220 205
rect 24170 165 24220 175
rect 24850 205 24900 235
rect 24850 175 24860 205
rect 24890 175 24900 205
rect 24850 165 24900 175
rect 25530 205 25580 235
rect 25530 175 25540 205
rect 25570 175 25580 205
rect 25530 165 25580 175
rect 26210 205 26260 235
rect 26210 175 26220 205
rect 26250 175 26260 205
rect 26210 165 26260 175
rect 26890 205 26940 235
rect 26890 175 26900 205
rect 26930 175 26940 205
rect 26890 165 26940 175
rect 27570 205 27620 235
rect 27570 175 27580 205
rect 27610 175 27620 205
rect 27570 165 27620 175
rect 28250 205 28300 235
rect 28250 175 28260 205
rect 28290 175 28300 205
rect 28250 165 28300 175
rect 28930 205 28980 235
rect 28930 175 28940 205
rect 28970 175 28980 205
rect 28930 165 28980 175
rect 29610 205 29660 235
rect 29610 175 29620 205
rect 29650 175 29660 205
rect 29610 165 29660 175
rect 295 105 355 110
rect 295 60 305 105
rect 345 60 355 105
rect 295 55 355 60
rect 465 105 525 110
rect 465 60 475 105
rect 515 60 525 105
rect 465 55 525 60
rect 640 105 705 115
rect 640 60 645 105
rect 700 60 705 105
rect 215 40 265 50
rect 215 10 225 40
rect 255 10 265 40
rect 45 -135 135 -125
rect 215 -130 265 10
rect 555 40 605 50
rect 555 10 565 40
rect 595 10 605 40
rect 555 -130 605 10
rect 640 -25 705 60
rect 830 105 890 110
rect 830 60 840 105
rect 880 60 890 105
rect 830 55 890 60
rect 1000 105 1060 110
rect 1000 60 1010 105
rect 1050 60 1060 105
rect 1000 55 1060 60
rect 1170 105 1230 110
rect 1170 60 1180 105
rect 1220 60 1230 105
rect 1170 55 1230 60
rect 1340 105 1400 110
rect 1340 60 1350 105
rect 1390 60 1400 105
rect 1340 55 1400 60
rect 1510 105 1570 110
rect 1510 60 1520 105
rect 1560 60 1570 105
rect 1510 55 1570 60
rect 1680 105 1740 110
rect 1680 60 1690 105
rect 1730 60 1740 105
rect 1680 55 1740 60
rect 1850 105 1910 110
rect 1850 60 1860 105
rect 1900 60 1910 105
rect 1850 55 1910 60
rect 2020 105 2080 110
rect 2020 60 2030 105
rect 2070 60 2080 105
rect 2020 55 2080 60
rect 2180 105 2245 115
rect 2180 60 2185 105
rect 2240 60 2245 105
rect 640 -65 650 -25
rect 700 -65 705 -25
rect 640 -80 705 -65
rect 750 40 800 50
rect 750 10 760 40
rect 790 10 800 40
rect 750 -130 800 10
rect 1430 40 1480 50
rect 1430 10 1440 40
rect 1470 10 1480 40
rect 1430 0 1480 10
rect 1440 -130 1470 0
rect 2180 -25 2245 60
rect 2340 105 2400 110
rect 2340 60 2350 105
rect 2390 60 2400 105
rect 2340 55 2400 60
rect 2510 105 2570 110
rect 2510 60 2520 105
rect 2560 60 2570 105
rect 2510 55 2570 60
rect 2680 105 2740 110
rect 2680 60 2690 105
rect 2730 60 2740 105
rect 2680 55 2740 60
rect 2850 105 2910 110
rect 2850 60 2860 105
rect 2900 60 2910 105
rect 2850 55 2910 60
rect 3020 105 3080 110
rect 3020 60 3030 105
rect 3070 60 3080 105
rect 3020 55 3080 60
rect 3190 105 3250 110
rect 3190 60 3200 105
rect 3240 60 3250 105
rect 3190 55 3250 60
rect 3360 105 3420 110
rect 3360 60 3370 105
rect 3410 60 3420 105
rect 3360 55 3420 60
rect 3530 105 3590 110
rect 3530 60 3540 105
rect 3580 60 3590 105
rect 3530 55 3590 60
rect 3700 105 3760 110
rect 3700 60 3710 105
rect 3750 60 3760 105
rect 3700 55 3760 60
rect 3870 105 3930 110
rect 3870 60 3880 105
rect 3920 60 3930 105
rect 3870 55 3930 60
rect 4040 105 4100 110
rect 4040 60 4050 105
rect 4090 60 4100 105
rect 4040 55 4100 60
rect 4210 105 4270 110
rect 4210 60 4220 105
rect 4260 60 4270 105
rect 4210 55 4270 60
rect 4380 105 4440 110
rect 4380 60 4390 105
rect 4430 60 4440 105
rect 4380 55 4440 60
rect 4550 105 4610 110
rect 4550 60 4560 105
rect 4600 60 4610 105
rect 4550 55 4610 60
rect 4720 105 4780 110
rect 4720 60 4730 105
rect 4770 60 4780 105
rect 4720 55 4780 60
rect 4890 105 4950 110
rect 4890 60 4900 105
rect 4940 60 4950 105
rect 4890 55 4950 60
rect 5060 105 5120 110
rect 5060 60 5070 105
rect 5110 60 5120 105
rect 5060 55 5120 60
rect 5230 105 5290 110
rect 5230 60 5240 105
rect 5280 60 5290 105
rect 5230 55 5290 60
rect 5400 105 5460 110
rect 5400 60 5410 105
rect 5450 60 5460 105
rect 5400 55 5460 60
rect 5570 105 5630 110
rect 5570 60 5580 105
rect 5620 60 5630 105
rect 5570 55 5630 60
rect 5740 105 5800 110
rect 5740 60 5750 105
rect 5790 60 5800 105
rect 5740 55 5800 60
rect 5910 105 5970 110
rect 5910 60 5920 105
rect 5960 60 5970 105
rect 5910 55 5970 60
rect 6080 105 6140 110
rect 6080 60 6090 105
rect 6130 60 6140 105
rect 6080 55 6140 60
rect 6250 105 6310 110
rect 6250 60 6260 105
rect 6300 60 6310 105
rect 6250 55 6310 60
rect 6420 105 6480 110
rect 6420 60 6430 105
rect 6470 60 6480 105
rect 6420 55 6480 60
rect 6590 105 6650 110
rect 6590 60 6600 105
rect 6640 60 6650 105
rect 6590 55 6650 60
rect 6760 105 6820 110
rect 6760 60 6770 105
rect 6810 60 6820 105
rect 6760 55 6820 60
rect 6930 105 6990 110
rect 6930 60 6940 105
rect 6980 60 6990 105
rect 6930 55 6990 60
rect 7100 105 7160 110
rect 7100 60 7110 105
rect 7150 60 7160 105
rect 7100 55 7160 60
rect 7270 105 7330 110
rect 7270 60 7280 105
rect 7320 60 7330 105
rect 7270 55 7330 60
rect 7440 105 7500 110
rect 7440 60 7450 105
rect 7490 60 7500 105
rect 7440 55 7500 60
rect 7610 105 7670 110
rect 7610 60 7620 105
rect 7660 60 7670 105
rect 7610 55 7670 60
rect 7770 105 7835 115
rect 7770 60 7775 105
rect 7830 60 7835 105
rect 2430 40 2480 50
rect 2430 10 2440 40
rect 2470 10 2480 40
rect 2430 0 2480 10
rect 3110 40 3160 50
rect 3110 10 3120 40
rect 3150 10 3160 40
rect 3110 0 3160 10
rect 3620 40 3670 50
rect 3620 10 3630 40
rect 3660 10 3670 40
rect 3620 0 3670 10
rect 4300 40 4350 50
rect 4300 10 4310 40
rect 4340 10 4350 40
rect 4300 0 4350 10
rect 4980 40 5030 50
rect 4980 10 4990 40
rect 5020 10 5030 40
rect 4980 0 5030 10
rect 5490 40 5540 50
rect 5490 10 5500 40
rect 5530 10 5540 40
rect 5490 0 5540 10
rect 2180 -65 2190 -25
rect 2240 -65 2245 -25
rect 2180 -70 2245 -65
rect 2440 -125 2470 0
rect 3120 -125 3150 0
rect 2285 -130 2315 -125
rect 45 -185 65 -135
rect 115 -185 135 -135
rect 45 -195 135 -185
rect 195 -140 285 -130
rect 195 -190 215 -140
rect 265 -190 285 -140
rect 65 -335 115 -195
rect 195 -200 285 -190
rect 535 -140 625 -130
rect 535 -190 555 -140
rect 605 -190 625 -140
rect 535 -200 625 -190
rect 725 -135 815 -130
rect 725 -185 745 -135
rect 795 -185 815 -135
rect 725 -195 815 -185
rect 1410 -140 1500 -130
rect 1410 -190 1430 -140
rect 1480 -190 1500 -140
rect 65 -365 75 -335
rect 105 -365 115 -335
rect 65 -375 115 -365
rect 745 -335 795 -195
rect 1410 -200 1500 -190
rect 2255 -140 2345 -130
rect 2255 -190 2275 -140
rect 2325 -190 2345 -140
rect 2255 -200 2345 -190
rect 2410 -135 2500 -125
rect 2410 -185 2430 -135
rect 2480 -185 2500 -135
rect 2410 -195 2500 -185
rect 2935 -135 3025 -125
rect 2935 -185 2955 -135
rect 3005 -185 3025 -135
rect 2935 -195 3025 -185
rect 3090 -135 3180 -125
rect 3090 -185 3110 -135
rect 3160 -185 3180 -135
rect 3090 -195 3180 -185
rect 3445 -135 3535 -125
rect 3630 -130 3660 0
rect 4310 -125 4340 0
rect 4990 -125 5020 0
rect 4155 -130 4185 -125
rect 3445 -185 3465 -135
rect 3515 -185 3535 -135
rect 3445 -195 3535 -185
rect 3600 -140 3690 -130
rect 3600 -190 3620 -140
rect 3670 -190 3690 -140
rect 2435 -200 2465 -195
rect 1435 -325 1465 -200
rect 2280 -205 2320 -200
rect 2285 -325 2315 -205
rect 2965 -325 2995 -195
rect 3475 -325 3505 -195
rect 3600 -200 3690 -190
rect 4125 -140 4215 -130
rect 4125 -190 4145 -140
rect 4195 -190 4215 -140
rect 4125 -200 4215 -190
rect 4280 -135 4370 -125
rect 4280 -185 4300 -135
rect 4350 -185 4370 -135
rect 4280 -195 4370 -185
rect 4805 -135 4895 -125
rect 4805 -185 4825 -135
rect 4875 -185 4895 -135
rect 4805 -195 4895 -185
rect 4960 -135 5050 -125
rect 4960 -185 4980 -135
rect 5030 -185 5050 -135
rect 4960 -195 5050 -185
rect 5315 -135 5405 -125
rect 5500 -130 5530 0
rect 7770 -25 7835 60
rect 7930 105 7990 110
rect 7930 60 7940 105
rect 7980 60 7990 105
rect 7930 55 7990 60
rect 8100 105 8160 110
rect 8100 60 8110 105
rect 8150 60 8160 105
rect 8100 55 8160 60
rect 8270 105 8330 110
rect 8270 60 8280 105
rect 8320 60 8330 105
rect 8270 55 8330 60
rect 8440 105 8500 110
rect 8440 60 8450 105
rect 8490 60 8500 105
rect 8440 55 8500 60
rect 8610 105 8670 110
rect 8610 60 8620 105
rect 8660 60 8670 105
rect 8610 55 8670 60
rect 8780 105 8840 110
rect 8780 60 8790 105
rect 8830 60 8840 105
rect 8780 55 8840 60
rect 8950 105 9010 110
rect 8950 60 8960 105
rect 9000 60 9010 105
rect 8950 55 9010 60
rect 9120 105 9180 110
rect 9120 60 9130 105
rect 9170 60 9180 105
rect 9120 55 9180 60
rect 9290 105 9350 110
rect 9290 60 9300 105
rect 9340 60 9350 105
rect 9290 55 9350 60
rect 9460 105 9520 110
rect 9460 60 9470 105
rect 9510 60 9520 105
rect 9460 55 9520 60
rect 9630 105 9690 110
rect 9630 60 9640 105
rect 9680 60 9690 105
rect 9630 55 9690 60
rect 9800 105 9860 110
rect 9800 60 9810 105
rect 9850 60 9860 105
rect 9800 55 9860 60
rect 9970 105 10030 110
rect 9970 60 9980 105
rect 10020 60 10030 105
rect 9970 55 10030 60
rect 10140 105 10200 110
rect 10140 60 10150 105
rect 10190 60 10200 105
rect 10140 55 10200 60
rect 10310 105 10370 110
rect 10310 60 10320 105
rect 10360 60 10370 105
rect 10310 55 10370 60
rect 10480 105 10540 110
rect 10480 60 10490 105
rect 10530 60 10540 105
rect 10480 55 10540 60
rect 10650 105 10710 110
rect 10650 60 10660 105
rect 10700 60 10710 105
rect 10650 55 10710 60
rect 10820 105 10880 110
rect 10820 60 10830 105
rect 10870 60 10880 105
rect 10820 55 10880 60
rect 10990 105 11050 110
rect 10990 60 11000 105
rect 11040 60 11050 105
rect 10990 55 11050 60
rect 11160 105 11220 110
rect 11160 60 11170 105
rect 11210 60 11220 105
rect 11160 55 11220 60
rect 11330 105 11390 110
rect 11330 60 11340 105
rect 11380 60 11390 105
rect 11330 55 11390 60
rect 11500 105 11560 110
rect 11500 60 11510 105
rect 11550 60 11560 105
rect 11500 55 11560 60
rect 11670 105 11730 110
rect 11670 60 11680 105
rect 11720 60 11730 105
rect 11670 55 11730 60
rect 11840 105 11900 110
rect 11840 60 11850 105
rect 11890 60 11900 105
rect 11840 55 11900 60
rect 12010 105 12070 110
rect 12010 60 12020 105
rect 12060 60 12070 105
rect 12010 55 12070 60
rect 12180 105 12240 110
rect 12180 60 12190 105
rect 12230 60 12240 105
rect 12180 55 12240 60
rect 12350 105 12410 110
rect 12350 60 12360 105
rect 12400 60 12410 105
rect 12350 55 12410 60
rect 12520 105 12580 110
rect 12520 60 12530 105
rect 12570 60 12580 105
rect 12520 55 12580 60
rect 12690 105 12750 110
rect 12690 60 12700 105
rect 12740 60 12750 105
rect 12690 55 12750 60
rect 12860 105 12920 110
rect 12860 60 12870 105
rect 12910 60 12920 105
rect 12860 55 12920 60
rect 13030 105 13090 110
rect 13030 60 13040 105
rect 13080 60 13090 105
rect 13030 55 13090 60
rect 13200 105 13260 110
rect 13200 60 13210 105
rect 13250 60 13260 105
rect 13200 55 13260 60
rect 13370 105 13430 110
rect 13370 60 13380 105
rect 13420 60 13430 105
rect 13370 55 13430 60
rect 13540 105 13600 110
rect 13540 60 13550 105
rect 13590 60 13600 105
rect 13540 55 13600 60
rect 13710 105 13770 110
rect 13710 60 13720 105
rect 13760 60 13770 105
rect 13710 55 13770 60
rect 13880 105 13940 110
rect 13880 60 13890 105
rect 13930 60 13940 105
rect 13880 55 13940 60
rect 14050 105 14110 110
rect 14050 60 14060 105
rect 14100 60 14110 105
rect 14050 55 14110 60
rect 14220 105 14280 110
rect 14220 60 14230 105
rect 14270 60 14280 105
rect 14220 55 14280 60
rect 14390 105 14450 110
rect 14390 60 14400 105
rect 14440 60 14450 105
rect 14390 55 14450 60
rect 14560 105 14620 110
rect 14560 60 14570 105
rect 14610 60 14620 105
rect 14560 55 14620 60
rect 14730 105 14790 110
rect 14730 60 14740 105
rect 14780 60 14790 105
rect 14730 55 14790 60
rect 14900 105 14960 110
rect 14900 60 14910 105
rect 14950 60 14960 105
rect 14900 55 14960 60
rect 15070 105 15130 110
rect 15070 60 15080 105
rect 15120 60 15130 105
rect 15070 55 15130 60
rect 15240 105 15300 110
rect 15240 60 15250 105
rect 15290 60 15300 105
rect 15240 55 15300 60
rect 15410 105 15470 110
rect 15410 60 15420 105
rect 15460 60 15470 105
rect 15410 55 15470 60
rect 15580 105 15640 110
rect 15580 60 15590 105
rect 15630 60 15640 105
rect 15580 55 15640 60
rect 15750 105 15810 110
rect 15750 60 15760 105
rect 15800 60 15810 105
rect 15750 55 15810 60
rect 15920 105 15980 110
rect 15920 60 15930 105
rect 15970 60 15980 105
rect 15920 55 15980 60
rect 16090 105 16150 110
rect 16090 60 16100 105
rect 16140 60 16150 105
rect 16090 55 16150 60
rect 16260 105 16320 110
rect 16260 60 16270 105
rect 16310 60 16320 105
rect 16260 55 16320 60
rect 16430 105 16490 110
rect 16430 60 16440 105
rect 16480 60 16490 105
rect 16430 55 16490 60
rect 16600 105 16660 110
rect 16600 60 16610 105
rect 16650 60 16660 105
rect 16600 55 16660 60
rect 16770 105 16830 110
rect 16770 60 16780 105
rect 16820 60 16830 105
rect 16770 55 16830 60
rect 16940 105 17000 110
rect 16940 60 16950 105
rect 16990 60 17000 105
rect 16940 55 17000 60
rect 17110 105 17170 110
rect 17110 60 17120 105
rect 17160 60 17170 105
rect 17110 55 17170 60
rect 17280 105 17340 110
rect 17280 60 17290 105
rect 17330 60 17340 105
rect 17280 55 17340 60
rect 17450 105 17510 110
rect 17450 60 17460 105
rect 17500 60 17510 105
rect 17450 55 17510 60
rect 17620 105 17680 110
rect 17620 60 17630 105
rect 17670 60 17680 105
rect 17620 55 17680 60
rect 17790 105 17850 110
rect 17790 60 17800 105
rect 17840 60 17850 105
rect 17790 55 17850 60
rect 17960 105 18020 110
rect 17960 60 17970 105
rect 18010 60 18020 105
rect 17960 55 18020 60
rect 18130 105 18190 110
rect 18130 60 18140 105
rect 18180 60 18190 105
rect 18130 55 18190 60
rect 18300 105 18360 110
rect 18300 60 18310 105
rect 18350 60 18360 105
rect 18300 55 18360 60
rect 18470 105 18530 110
rect 18470 60 18480 105
rect 18520 60 18530 105
rect 18470 55 18530 60
rect 18640 105 18700 110
rect 18640 60 18650 105
rect 18690 60 18700 105
rect 18640 55 18700 60
rect 18810 105 18870 110
rect 18810 60 18820 105
rect 18860 60 18870 105
rect 18810 55 18870 60
rect 18980 105 19040 110
rect 18980 60 18990 105
rect 19030 60 19040 105
rect 18980 55 19040 60
rect 19150 105 19210 110
rect 19150 60 19160 105
rect 19200 60 19210 105
rect 19150 55 19210 60
rect 19320 105 19380 110
rect 19320 60 19330 105
rect 19370 60 19380 105
rect 19320 55 19380 60
rect 19490 105 19550 110
rect 19490 60 19500 105
rect 19540 60 19550 105
rect 19490 55 19550 60
rect 19660 105 19720 110
rect 19660 60 19670 105
rect 19710 60 19720 105
rect 19660 55 19720 60
rect 19830 105 19890 110
rect 19830 60 19840 105
rect 19880 60 19890 105
rect 19830 55 19890 60
rect 20000 105 20060 110
rect 20000 60 20010 105
rect 20050 60 20060 105
rect 20000 55 20060 60
rect 20170 105 20230 110
rect 20170 60 20180 105
rect 20220 60 20230 105
rect 20170 55 20230 60
rect 20340 105 20400 110
rect 20340 60 20350 105
rect 20390 60 20400 105
rect 20340 55 20400 60
rect 20510 105 20570 110
rect 20510 60 20520 105
rect 20560 60 20570 105
rect 20510 55 20570 60
rect 20680 105 20740 110
rect 20680 60 20690 105
rect 20730 60 20740 105
rect 20680 55 20740 60
rect 20850 105 20910 110
rect 20850 60 20860 105
rect 20900 60 20910 105
rect 20850 55 20910 60
rect 21020 105 21080 110
rect 21020 60 21030 105
rect 21070 60 21080 105
rect 21020 55 21080 60
rect 21190 105 21250 110
rect 21190 60 21200 105
rect 21240 60 21250 105
rect 21190 55 21250 60
rect 21360 105 21420 110
rect 21360 60 21370 105
rect 21410 60 21420 105
rect 21360 55 21420 60
rect 21530 105 21590 110
rect 21530 60 21540 105
rect 21580 60 21590 105
rect 21530 55 21590 60
rect 21700 105 21760 110
rect 21700 60 21710 105
rect 21750 60 21760 105
rect 21700 55 21760 60
rect 21870 105 21930 110
rect 21870 60 21880 105
rect 21920 60 21930 105
rect 21870 55 21930 60
rect 22040 105 22100 110
rect 22040 60 22050 105
rect 22090 60 22100 105
rect 22040 55 22100 60
rect 22210 105 22270 110
rect 22210 60 22220 105
rect 22260 60 22270 105
rect 22210 55 22270 60
rect 22380 105 22440 110
rect 22380 60 22390 105
rect 22430 60 22440 105
rect 22380 55 22440 60
rect 22550 105 22610 110
rect 22550 60 22560 105
rect 22600 60 22610 105
rect 22550 55 22610 60
rect 22720 105 22780 110
rect 22720 60 22730 105
rect 22770 60 22780 105
rect 22720 55 22780 60
rect 22890 105 22950 110
rect 22890 60 22900 105
rect 22940 60 22950 105
rect 22890 55 22950 60
rect 23060 105 23120 110
rect 23060 60 23070 105
rect 23110 60 23120 105
rect 23060 55 23120 60
rect 23230 105 23290 110
rect 23230 60 23240 105
rect 23280 60 23290 105
rect 23230 55 23290 60
rect 23400 105 23460 110
rect 23400 60 23410 105
rect 23450 60 23460 105
rect 23400 55 23460 60
rect 23570 105 23630 110
rect 23570 60 23580 105
rect 23620 60 23630 105
rect 23570 55 23630 60
rect 23740 105 23800 110
rect 23740 60 23750 105
rect 23790 60 23800 105
rect 23740 55 23800 60
rect 23910 105 23970 110
rect 23910 60 23920 105
rect 23960 60 23970 105
rect 23910 55 23970 60
rect 24080 105 24140 110
rect 24080 60 24090 105
rect 24130 60 24140 105
rect 24080 55 24140 60
rect 24250 105 24310 110
rect 24250 60 24260 105
rect 24300 60 24310 105
rect 24250 55 24310 60
rect 24420 105 24480 110
rect 24420 60 24430 105
rect 24470 60 24480 105
rect 24420 55 24480 60
rect 24590 105 24650 110
rect 24590 60 24600 105
rect 24640 60 24650 105
rect 24590 55 24650 60
rect 24760 105 24820 110
rect 24760 60 24770 105
rect 24810 60 24820 105
rect 24760 55 24820 60
rect 24930 105 24990 110
rect 24930 60 24940 105
rect 24980 60 24990 105
rect 24930 55 24990 60
rect 25100 105 25160 110
rect 25100 60 25110 105
rect 25150 60 25160 105
rect 25100 55 25160 60
rect 25270 105 25330 110
rect 25270 60 25280 105
rect 25320 60 25330 105
rect 25270 55 25330 60
rect 25440 105 25500 110
rect 25440 60 25450 105
rect 25490 60 25500 105
rect 25440 55 25500 60
rect 25610 105 25670 110
rect 25610 60 25620 105
rect 25660 60 25670 105
rect 25610 55 25670 60
rect 25780 105 25840 110
rect 25780 60 25790 105
rect 25830 60 25840 105
rect 25780 55 25840 60
rect 25950 105 26010 110
rect 25950 60 25960 105
rect 26000 60 26010 105
rect 25950 55 26010 60
rect 26120 105 26180 110
rect 26120 60 26130 105
rect 26170 60 26180 105
rect 26120 55 26180 60
rect 26290 105 26350 110
rect 26290 60 26300 105
rect 26340 60 26350 105
rect 26290 55 26350 60
rect 26460 105 26520 110
rect 26460 60 26470 105
rect 26510 60 26520 105
rect 26460 55 26520 60
rect 26630 105 26690 110
rect 26630 60 26640 105
rect 26680 60 26690 105
rect 26630 55 26690 60
rect 26800 105 26860 110
rect 26800 60 26810 105
rect 26850 60 26860 105
rect 26800 55 26860 60
rect 26970 105 27030 110
rect 26970 60 26980 105
rect 27020 60 27030 105
rect 26970 55 27030 60
rect 27140 105 27200 110
rect 27140 60 27150 105
rect 27190 60 27200 105
rect 27140 55 27200 60
rect 27310 105 27370 110
rect 27310 60 27320 105
rect 27360 60 27370 105
rect 27310 55 27370 60
rect 27480 105 27540 110
rect 27480 60 27490 105
rect 27530 60 27540 105
rect 27480 55 27540 60
rect 27650 105 27710 110
rect 27650 60 27660 105
rect 27700 60 27710 105
rect 27650 55 27710 60
rect 27820 105 27880 110
rect 27820 60 27830 105
rect 27870 60 27880 105
rect 27820 55 27880 60
rect 27990 105 28050 110
rect 27990 60 28000 105
rect 28040 60 28050 105
rect 27990 55 28050 60
rect 28160 105 28220 110
rect 28160 60 28170 105
rect 28210 60 28220 105
rect 28160 55 28220 60
rect 28330 105 28390 110
rect 28330 60 28340 105
rect 28380 60 28390 105
rect 28330 55 28390 60
rect 28500 105 28560 110
rect 28500 60 28510 105
rect 28550 60 28560 105
rect 28500 55 28560 60
rect 28670 105 28730 110
rect 28670 60 28680 105
rect 28720 60 28730 105
rect 28670 55 28730 60
rect 28840 105 28900 110
rect 28840 60 28850 105
rect 28890 60 28900 105
rect 28840 55 28900 60
rect 29010 105 29070 110
rect 29010 60 29020 105
rect 29060 60 29070 105
rect 29010 55 29070 60
rect 29180 105 29240 110
rect 29180 60 29190 105
rect 29230 60 29240 105
rect 29180 55 29240 60
rect 29350 105 29410 110
rect 29350 60 29360 105
rect 29400 60 29410 105
rect 29350 55 29410 60
rect 29520 105 29580 110
rect 29520 60 29530 105
rect 29570 60 29580 105
rect 29520 55 29580 60
rect 7770 -65 7780 -25
rect 7830 -65 7835 -25
rect 7770 -70 7835 -65
rect 5315 -185 5335 -135
rect 5385 -185 5405 -135
rect 5315 -195 5405 -185
rect 5470 -140 5560 -130
rect 5470 -190 5490 -140
rect 5540 -190 5560 -140
rect 4305 -200 4335 -195
rect 4150 -205 4190 -200
rect 4155 -325 4185 -205
rect 4835 -325 4865 -195
rect 5345 -325 5375 -195
rect 5470 -200 5560 -190
rect 5845 -135 5915 -125
rect 5995 -130 6045 -110
rect 6335 -130 6385 -110
rect 6530 -130 6580 -110
rect 7220 -130 7250 -110
rect 5895 -185 5915 -135
rect 5845 -195 5915 -185
rect 5975 -140 6065 -130
rect 5975 -190 5995 -140
rect 6045 -190 6065 -140
rect 745 -365 755 -335
rect 785 -365 795 -335
rect 745 -375 795 -365
rect 1425 -335 1475 -325
rect 1425 -365 1435 -335
rect 1465 -365 1475 -335
rect 1425 -375 1475 -365
rect 2275 -335 2325 -325
rect 2275 -365 2285 -335
rect 2315 -365 2325 -335
rect 2275 -375 2325 -365
rect 2955 -335 3005 -325
rect 2955 -365 2965 -335
rect 2995 -365 3005 -335
rect 2955 -375 3005 -365
rect 3465 -335 3515 -325
rect 3465 -365 3475 -335
rect 3505 -365 3515 -335
rect 3465 -375 3515 -365
rect 4145 -335 4195 -325
rect 4145 -365 4155 -335
rect 4185 -365 4195 -335
rect 4145 -375 4195 -365
rect 4825 -335 4875 -325
rect 4825 -365 4835 -335
rect 4865 -365 4875 -335
rect 4825 -375 4875 -365
rect 5335 -335 5385 -325
rect 5335 -365 5345 -335
rect 5375 -365 5385 -335
rect 5335 -375 5385 -365
rect 5845 -335 5895 -195
rect 5975 -200 6065 -190
rect 6315 -140 6405 -130
rect 6315 -190 6335 -140
rect 6385 -190 6405 -140
rect 6315 -200 6405 -190
rect 6505 -135 6595 -130
rect 6505 -185 6525 -135
rect 6575 -185 6595 -135
rect 6505 -195 6595 -185
rect 7190 -140 7280 -130
rect 7190 -190 7210 -140
rect 7260 -190 7280 -140
rect 5845 -365 5855 -335
rect 5885 -365 5895 -335
rect 5845 -375 5895 -365
rect 6525 -335 6575 -195
rect 7190 -200 7280 -190
rect 7215 -325 7245 -200
rect 7935 -225 7985 55
rect 8190 40 8240 50
rect 8190 10 8200 40
rect 8230 10 8240 40
rect 8190 0 8240 10
rect 8870 40 8920 50
rect 8870 10 8880 40
rect 8910 10 8920 40
rect 8870 0 8920 10
rect 9380 40 9430 50
rect 9380 10 9390 40
rect 9420 10 9430 40
rect 9380 0 9430 10
rect 10060 40 10110 50
rect 10060 10 10070 40
rect 10100 10 10110 40
rect 10060 0 10110 10
rect 10740 40 10790 50
rect 10740 10 10750 40
rect 10780 10 10790 40
rect 10740 0 10790 10
rect 11250 40 11300 50
rect 11250 10 11260 40
rect 11290 10 11300 40
rect 11250 0 11300 10
rect 11930 40 11980 50
rect 11930 10 11940 40
rect 11970 10 11980 40
rect 11930 0 11980 10
rect 12270 40 12320 50
rect 12270 10 12280 40
rect 12310 10 12320 40
rect 12270 0 12320 10
rect 14140 40 14190 50
rect 14140 10 14150 40
rect 14180 10 14190 40
rect 14140 0 14190 10
rect 14820 40 14870 50
rect 14820 10 14830 40
rect 14860 10 14870 40
rect 14820 0 14870 10
rect 15330 40 15380 50
rect 15330 10 15340 40
rect 15370 10 15380 40
rect 15330 0 15380 10
rect 8200 -125 8230 0
rect 8880 -125 8910 0
rect 8065 -130 8095 -125
rect 8035 -140 8125 -130
rect 8035 -190 8055 -140
rect 8105 -190 8125 -140
rect 8035 -200 8125 -190
rect 8170 -135 8260 -125
rect 8170 -185 8190 -135
rect 8240 -185 8260 -135
rect 8170 -195 8260 -185
rect 8715 -135 8805 -125
rect 8715 -185 8735 -135
rect 8785 -185 8805 -135
rect 8715 -195 8805 -185
rect 8850 -135 8940 -125
rect 8850 -185 8870 -135
rect 8920 -185 8940 -135
rect 8850 -195 8940 -185
rect 9225 -135 9315 -125
rect 9390 -130 9420 0
rect 10070 -125 10100 0
rect 10750 -125 10780 0
rect 9935 -130 9965 -125
rect 9225 -185 9245 -135
rect 9295 -185 9315 -135
rect 9225 -195 9315 -185
rect 9360 -140 9450 -130
rect 9360 -190 9380 -140
rect 9430 -190 9450 -140
rect 8195 -200 8225 -195
rect 8060 -205 8100 -200
rect 7925 -230 8005 -225
rect 7925 -260 7965 -230
rect 8000 -260 8005 -230
rect 7925 -305 8005 -260
rect 8065 -325 8095 -205
rect 8745 -325 8775 -195
rect 9255 -325 9285 -195
rect 9360 -200 9450 -190
rect 9905 -140 9995 -130
rect 9905 -190 9925 -140
rect 9975 -190 9995 -140
rect 9905 -200 9995 -190
rect 10040 -135 10130 -125
rect 10040 -185 10060 -135
rect 10110 -185 10130 -135
rect 10040 -195 10130 -185
rect 10585 -135 10675 -125
rect 10585 -185 10605 -135
rect 10655 -185 10675 -135
rect 10585 -195 10675 -185
rect 10720 -135 10810 -125
rect 10720 -185 10740 -135
rect 10790 -185 10810 -135
rect 10720 -195 10810 -185
rect 11095 -135 11185 -125
rect 11260 -130 11290 0
rect 11940 -110 11970 0
rect 12280 -110 12310 0
rect 11095 -185 11115 -135
rect 11165 -185 11185 -135
rect 11095 -195 11185 -185
rect 11230 -140 11320 -130
rect 11230 -190 11250 -140
rect 11300 -190 11320 -140
rect 10065 -200 10095 -195
rect 9930 -205 9970 -200
rect 9935 -325 9965 -205
rect 10615 -325 10645 -195
rect 11125 -325 11155 -195
rect 11230 -200 11320 -190
rect 11795 -135 11865 -125
rect 11930 -130 11980 -110
rect 12265 -130 12315 -110
rect 12480 -130 12530 -110
rect 13170 -130 13200 -110
rect 14150 -125 14180 0
rect 14830 -125 14860 0
rect 14015 -130 14045 -125
rect 11845 -185 11865 -135
rect 11795 -195 11865 -185
rect 11910 -140 12000 -130
rect 11910 -190 11930 -140
rect 11980 -190 12000 -140
rect 6525 -365 6535 -335
rect 6565 -365 6575 -335
rect 6525 -375 6575 -365
rect 7205 -335 7255 -325
rect 7205 -365 7215 -335
rect 7245 -365 7255 -335
rect 7205 -375 7255 -365
rect 8055 -335 8105 -325
rect 8055 -365 8065 -335
rect 8095 -365 8105 -335
rect 8055 -375 8105 -365
rect 8735 -335 8785 -325
rect 8735 -365 8745 -335
rect 8775 -365 8785 -335
rect 8735 -375 8785 -365
rect 9245 -335 9295 -325
rect 9245 -365 9255 -335
rect 9285 -365 9295 -335
rect 9245 -375 9295 -365
rect 9925 -335 9975 -325
rect 9925 -365 9935 -335
rect 9965 -365 9975 -335
rect 9925 -375 9975 -365
rect 10605 -335 10655 -325
rect 10605 -365 10615 -335
rect 10645 -365 10655 -335
rect 10605 -375 10655 -365
rect 11115 -335 11165 -325
rect 11115 -365 11125 -335
rect 11155 -365 11165 -335
rect 11115 -375 11165 -365
rect 11795 -335 11845 -195
rect 11910 -200 12000 -190
rect 12245 -140 12335 -130
rect 12245 -190 12265 -140
rect 12315 -190 12335 -140
rect 12245 -200 12335 -190
rect 12455 -135 12545 -130
rect 12455 -185 12475 -135
rect 12525 -185 12545 -135
rect 12455 -195 12545 -185
rect 13140 -140 13230 -130
rect 13140 -190 13160 -140
rect 13210 -190 13230 -140
rect 11795 -365 11805 -335
rect 11835 -365 11845 -335
rect 11795 -375 11845 -365
rect 12475 -335 12525 -195
rect 13140 -200 13230 -190
rect 13985 -140 14075 -130
rect 13985 -190 14005 -140
rect 14055 -190 14075 -140
rect 13985 -200 14075 -190
rect 14120 -135 14210 -125
rect 14120 -185 14140 -135
rect 14190 -185 14210 -135
rect 14120 -195 14210 -185
rect 14665 -135 14755 -125
rect 14665 -185 14685 -135
rect 14735 -185 14755 -135
rect 14665 -195 14755 -185
rect 14800 -135 14890 -125
rect 14800 -185 14820 -135
rect 14870 -185 14890 -135
rect 14800 -195 14890 -185
rect 15175 -135 15265 -125
rect 15340 -130 15370 0
rect 15175 -185 15195 -135
rect 15245 -185 15265 -135
rect 15175 -195 15265 -185
rect 15310 -140 15400 -130
rect 15310 -190 15330 -140
rect 15380 -190 15400 -140
rect 14145 -200 14175 -195
rect 13165 -325 13195 -200
rect 14010 -205 14050 -200
rect 14015 -325 14045 -205
rect 14695 -325 14725 -195
rect 15205 -325 15235 -195
rect 15310 -200 15400 -190
rect 15585 -225 15635 55
rect 16010 40 16060 50
rect 16010 10 16020 40
rect 16050 10 16060 40
rect 16010 0 16060 10
rect 16690 40 16740 50
rect 16690 10 16700 40
rect 16730 10 16740 40
rect 16690 0 16740 10
rect 17200 40 17250 50
rect 17200 10 17210 40
rect 17240 10 17250 40
rect 17200 0 17250 10
rect 17880 40 17930 50
rect 17880 10 17890 40
rect 17920 10 17930 40
rect 17880 0 17930 10
rect 18220 40 18270 50
rect 18220 10 18230 40
rect 18260 10 18270 40
rect 18220 0 18270 10
rect 21280 40 21330 50
rect 21280 10 21290 40
rect 21320 10 21330 40
rect 21280 0 21330 10
rect 22300 40 22350 50
rect 22300 10 22310 40
rect 22340 10 22350 40
rect 22300 0 22350 10
rect 24170 40 24220 50
rect 24170 10 24180 40
rect 24210 10 24220 40
rect 24170 0 24220 10
rect 24850 40 24900 50
rect 24850 10 24860 40
rect 24890 10 24900 40
rect 24850 0 24900 10
rect 25360 40 25410 50
rect 25360 10 25370 40
rect 25400 10 25410 40
rect 25360 0 25410 10
rect 26040 40 26090 50
rect 26040 10 26050 40
rect 26080 10 26090 40
rect 26040 0 26090 10
rect 26720 40 26770 50
rect 26720 10 26730 40
rect 26760 10 26770 40
rect 26720 0 26770 10
rect 27740 40 27790 50
rect 27740 10 27750 40
rect 27780 10 27790 40
rect 27740 0 27790 10
rect 16020 -125 16050 0
rect 16700 -125 16730 0
rect 15885 -130 15915 -125
rect 15855 -140 15945 -130
rect 15855 -190 15875 -140
rect 15925 -190 15945 -140
rect 15855 -200 15945 -190
rect 15990 -135 16080 -125
rect 15990 -185 16010 -135
rect 16060 -185 16080 -135
rect 15990 -195 16080 -185
rect 16535 -135 16625 -125
rect 16535 -185 16555 -135
rect 16605 -185 16625 -135
rect 16535 -195 16625 -185
rect 16670 -135 16760 -125
rect 16670 -185 16690 -135
rect 16740 -185 16760 -135
rect 16670 -195 16760 -185
rect 17045 -135 17135 -125
rect 17210 -130 17240 0
rect 17890 -110 17920 0
rect 18230 -110 18260 0
rect 17045 -185 17065 -135
rect 17115 -185 17135 -135
rect 17045 -195 17135 -185
rect 17180 -140 17270 -130
rect 17180 -190 17200 -140
rect 17250 -190 17270 -140
rect 16015 -200 16045 -195
rect 15880 -205 15920 -200
rect 15575 -230 15655 -225
rect 15575 -260 15615 -230
rect 15650 -260 15655 -230
rect 15575 -305 15655 -260
rect 15885 -325 15915 -205
rect 16565 -325 16595 -195
rect 17075 -325 17105 -195
rect 17180 -200 17270 -190
rect 17745 -135 17815 -125
rect 17880 -130 17930 -110
rect 18215 -130 18265 -110
rect 18430 -130 18480 -110
rect 19120 -130 19150 -110
rect 19965 -130 19995 -125
rect 17795 -185 17815 -135
rect 17745 -195 17815 -185
rect 17860 -140 17950 -130
rect 17860 -190 17880 -140
rect 17930 -190 17950 -140
rect 12475 -365 12485 -335
rect 12515 -365 12525 -335
rect 12475 -375 12525 -365
rect 13155 -335 13205 -325
rect 13155 -365 13165 -335
rect 13195 -365 13205 -335
rect 13155 -375 13205 -365
rect 14005 -335 14055 -325
rect 14005 -365 14015 -335
rect 14045 -365 14055 -335
rect 14005 -375 14055 -365
rect 14685 -335 14735 -325
rect 14685 -365 14695 -335
rect 14725 -365 14735 -335
rect 14685 -375 14735 -365
rect 15195 -335 15245 -325
rect 15195 -365 15205 -335
rect 15235 -365 15245 -335
rect 15195 -375 15245 -365
rect 15875 -335 15925 -325
rect 15875 -365 15885 -335
rect 15915 -365 15925 -335
rect 15875 -375 15925 -365
rect 16555 -335 16605 -325
rect 16555 -365 16565 -335
rect 16595 -365 16605 -335
rect 16555 -375 16605 -365
rect 17065 -335 17115 -325
rect 17065 -365 17075 -335
rect 17105 -365 17115 -335
rect 17065 -375 17115 -365
rect 17745 -335 17795 -195
rect 17860 -200 17950 -190
rect 18195 -140 18285 -130
rect 18195 -190 18215 -140
rect 18265 -190 18285 -140
rect 18195 -200 18285 -190
rect 18405 -135 18495 -130
rect 18405 -185 18425 -135
rect 18475 -185 18495 -135
rect 18405 -195 18495 -185
rect 19090 -140 19180 -130
rect 19090 -190 19110 -140
rect 19160 -190 19180 -140
rect 17745 -365 17755 -335
rect 17785 -365 17795 -335
rect 17745 -375 17795 -365
rect 18425 -335 18475 -195
rect 19090 -200 19180 -190
rect 19935 -140 20025 -130
rect 19935 -190 19955 -140
rect 20005 -190 20025 -140
rect 19935 -200 20025 -190
rect 20615 -135 20705 -125
rect 20615 -185 20635 -135
rect 20685 -185 20705 -135
rect 20615 -195 20705 -185
rect 21125 -135 21215 -125
rect 21290 -130 21320 0
rect 22310 -110 22340 0
rect 21815 -130 21895 -125
rect 22300 -130 22350 -110
rect 24180 -125 24210 0
rect 24860 -125 24890 0
rect 24045 -130 24075 -125
rect 21125 -185 21145 -135
rect 21195 -185 21215 -135
rect 21125 -195 21215 -185
rect 21260 -140 21350 -130
rect 21260 -190 21280 -140
rect 21330 -190 21350 -140
rect 19115 -325 19145 -200
rect 19960 -205 20000 -200
rect 19965 -325 19995 -205
rect 20645 -325 20675 -195
rect 21155 -325 21185 -195
rect 21260 -200 21350 -190
rect 21805 -135 21895 -130
rect 21805 -190 21825 -135
rect 21875 -190 21895 -135
rect 21805 -200 21895 -190
rect 22280 -140 22370 -130
rect 22280 -190 22300 -140
rect 22350 -190 22370 -140
rect 22280 -200 22370 -190
rect 22485 -135 22575 -130
rect 22485 -185 22505 -135
rect 22555 -185 22575 -135
rect 22485 -195 22575 -185
rect 23170 -140 23260 -130
rect 23170 -190 23190 -140
rect 23240 -190 23260 -140
rect 18425 -365 18435 -335
rect 18465 -365 18475 -335
rect 18425 -375 18475 -365
rect 19105 -335 19155 -325
rect 19105 -365 19115 -335
rect 19145 -365 19155 -335
rect 19105 -375 19155 -365
rect 19955 -335 20005 -325
rect 19955 -365 19965 -335
rect 19995 -365 20005 -335
rect 19955 -375 20005 -365
rect 20635 -335 20685 -325
rect 20635 -365 20645 -335
rect 20675 -365 20685 -335
rect 20635 -375 20685 -365
rect 21145 -335 21195 -325
rect 21145 -365 21155 -335
rect 21185 -365 21195 -335
rect 21145 -375 21195 -365
rect 21825 -335 21875 -200
rect 21825 -365 21835 -335
rect 21865 -365 21875 -335
rect 21825 -375 21875 -365
rect 22505 -335 22555 -195
rect 23170 -200 23260 -190
rect 24015 -140 24105 -130
rect 24015 -190 24035 -140
rect 24085 -190 24105 -140
rect 24015 -200 24105 -190
rect 24150 -135 24240 -125
rect 24150 -185 24170 -135
rect 24220 -185 24240 -135
rect 24150 -195 24240 -185
rect 24695 -135 24785 -125
rect 24695 -185 24715 -135
rect 24765 -185 24785 -135
rect 24695 -195 24785 -185
rect 24830 -135 24920 -125
rect 24830 -185 24850 -135
rect 24900 -185 24920 -135
rect 24830 -195 24920 -185
rect 25205 -135 25295 -125
rect 25370 -130 25400 0
rect 26050 -125 26080 0
rect 26730 -125 26760 0
rect 27750 -110 27780 0
rect 25915 -130 25945 -125
rect 25205 -185 25225 -135
rect 25275 -185 25295 -135
rect 25205 -195 25295 -185
rect 25340 -140 25430 -130
rect 25340 -190 25360 -140
rect 25410 -190 25430 -140
rect 24175 -200 24205 -195
rect 23195 -325 23225 -200
rect 24040 -205 24080 -200
rect 24045 -325 24075 -205
rect 24725 -325 24755 -195
rect 25235 -325 25265 -195
rect 25340 -200 25430 -190
rect 25885 -140 25975 -130
rect 25885 -190 25905 -140
rect 25955 -190 25975 -140
rect 25885 -200 25975 -190
rect 26020 -135 26110 -125
rect 26020 -185 26040 -135
rect 26090 -185 26110 -135
rect 26020 -195 26110 -185
rect 26565 -135 26655 -125
rect 26565 -185 26585 -135
rect 26635 -185 26655 -135
rect 26565 -195 26655 -185
rect 26700 -135 26790 -125
rect 26700 -185 26720 -135
rect 26770 -185 26790 -135
rect 26700 -195 26790 -185
rect 27075 -135 27165 -125
rect 27075 -185 27095 -135
rect 27145 -185 27165 -135
rect 27075 -195 27165 -185
rect 27605 -135 27675 -125
rect 27740 -130 27790 -110
rect 28290 -130 28340 -110
rect 28980 -130 29010 -110
rect 27655 -185 27675 -135
rect 27605 -195 27675 -185
rect 27720 -140 27810 -130
rect 27720 -190 27740 -140
rect 27790 -190 27810 -140
rect 26045 -200 26075 -195
rect 25910 -205 25950 -200
rect 25915 -325 25945 -205
rect 26595 -325 26625 -195
rect 27105 -325 27135 -195
rect 22505 -365 22515 -335
rect 22545 -365 22555 -335
rect 22505 -375 22555 -365
rect 23185 -335 23235 -325
rect 23185 -365 23195 -335
rect 23225 -365 23235 -335
rect 23185 -375 23235 -365
rect 24035 -335 24085 -325
rect 24035 -365 24045 -335
rect 24075 -365 24085 -335
rect 24035 -375 24085 -365
rect 24715 -335 24765 -325
rect 24715 -365 24725 -335
rect 24755 -365 24765 -335
rect 24715 -375 24765 -365
rect 25225 -335 25275 -325
rect 25225 -365 25235 -335
rect 25265 -365 25275 -335
rect 25225 -375 25275 -365
rect 25905 -335 25955 -325
rect 25905 -365 25915 -335
rect 25945 -365 25955 -335
rect 25905 -375 25955 -365
rect 26585 -335 26635 -325
rect 26585 -365 26595 -335
rect 26625 -365 26635 -335
rect 26585 -375 26635 -365
rect 27095 -335 27145 -325
rect 27095 -365 27105 -335
rect 27135 -365 27145 -335
rect 27095 -375 27145 -365
rect 27605 -335 27655 -195
rect 27720 -200 27810 -190
rect 28265 -135 28355 -130
rect 28265 -185 28285 -135
rect 28335 -185 28355 -135
rect 28265 -195 28355 -185
rect 28950 -140 29040 -130
rect 28950 -190 28970 -140
rect 29020 -190 29040 -140
rect 27605 -365 27615 -335
rect 27645 -365 27655 -335
rect 27605 -375 27655 -365
rect 28285 -335 28335 -195
rect 28950 -200 29040 -190
rect 28975 -325 29005 -200
rect 29530 -225 29570 55
rect 29825 -130 29855 -125
rect 29795 -140 29885 -130
rect 29795 -190 29815 -140
rect 29865 -190 29885 -140
rect 29795 -200 29885 -190
rect 30475 -135 30565 -125
rect 30475 -185 30495 -135
rect 30545 -185 30565 -135
rect 30475 -195 30565 -185
rect 30985 -135 31075 -125
rect 31695 -130 31725 -125
rect 30985 -185 31005 -135
rect 31055 -185 31075 -135
rect 30985 -195 31075 -185
rect 31665 -140 31755 -130
rect 31665 -190 31685 -140
rect 31735 -190 31755 -140
rect 29820 -205 29860 -200
rect 29515 -230 29595 -225
rect 29515 -260 29555 -230
rect 29590 -260 29595 -230
rect 29515 -305 29595 -260
rect 29825 -325 29855 -205
rect 30505 -325 30535 -195
rect 31015 -325 31045 -195
rect 31665 -200 31755 -190
rect 32345 -135 32435 -125
rect 32345 -185 32365 -135
rect 32415 -185 32435 -135
rect 32345 -195 32435 -185
rect 32855 -135 32945 -125
rect 32855 -185 32875 -135
rect 32925 -185 32945 -135
rect 32855 -195 32945 -185
rect 33555 -135 33625 -125
rect 34240 -130 34290 -110
rect 34930 -130 34960 -110
rect 35775 -130 35805 -125
rect 33605 -185 33625 -135
rect 33555 -195 33625 -185
rect 34215 -135 34305 -130
rect 34215 -185 34235 -135
rect 34285 -185 34305 -135
rect 34215 -195 34305 -185
rect 34900 -140 34990 -130
rect 34900 -190 34920 -140
rect 34970 -190 34990 -140
rect 31690 -205 31730 -200
rect 31695 -325 31725 -205
rect 32375 -325 32405 -195
rect 32885 -325 32915 -195
rect 28285 -365 28295 -335
rect 28325 -365 28335 -335
rect 28285 -375 28335 -365
rect 28965 -335 29015 -325
rect 28965 -365 28975 -335
rect 29005 -365 29015 -335
rect 28965 -375 29015 -365
rect 29815 -335 29865 -325
rect 29815 -365 29825 -335
rect 29855 -365 29865 -335
rect 29815 -375 29865 -365
rect 30495 -335 30545 -325
rect 30495 -365 30505 -335
rect 30535 -365 30545 -335
rect 30495 -375 30545 -365
rect 31005 -335 31055 -325
rect 31005 -365 31015 -335
rect 31045 -365 31055 -335
rect 31005 -375 31055 -365
rect 31685 -335 31735 -325
rect 31685 -365 31695 -335
rect 31725 -365 31735 -335
rect 31685 -375 31735 -365
rect 32365 -335 32415 -325
rect 32365 -365 32375 -335
rect 32405 -365 32415 -335
rect 32365 -375 32415 -365
rect 32875 -335 32925 -325
rect 32875 -365 32885 -335
rect 32915 -365 32925 -335
rect 32875 -375 32925 -365
rect 33555 -335 33605 -195
rect 33555 -365 33565 -335
rect 33595 -365 33605 -335
rect 33555 -375 33605 -365
rect 34235 -335 34285 -195
rect 34900 -200 34990 -190
rect 35745 -140 35835 -130
rect 35745 -190 35765 -140
rect 35815 -190 35835 -140
rect 35745 -200 35835 -190
rect 36425 -135 36515 -125
rect 36425 -185 36445 -135
rect 36495 -185 36515 -135
rect 36425 -195 36515 -185
rect 36935 -135 37025 -125
rect 37645 -130 37675 -125
rect 36935 -185 36955 -135
rect 37005 -185 37025 -135
rect 36935 -195 37025 -185
rect 37615 -140 37705 -130
rect 37615 -190 37635 -140
rect 37685 -190 37705 -140
rect 34925 -325 34955 -200
rect 35770 -205 35810 -200
rect 35775 -325 35805 -205
rect 36455 -325 36485 -195
rect 36965 -325 36995 -195
rect 37615 -200 37705 -190
rect 38295 -135 38385 -125
rect 38295 -185 38315 -135
rect 38365 -185 38385 -135
rect 38295 -195 38385 -185
rect 38805 -135 38895 -125
rect 38805 -185 38825 -135
rect 38875 -185 38895 -135
rect 38805 -195 38895 -185
rect 39505 -135 39575 -125
rect 40190 -130 40240 -110
rect 40880 -130 40910 -110
rect 41725 -130 41755 -125
rect 39555 -185 39575 -135
rect 39505 -195 39575 -185
rect 40165 -135 40255 -130
rect 40165 -185 40185 -135
rect 40235 -185 40255 -135
rect 40165 -195 40255 -185
rect 40850 -140 40940 -130
rect 40850 -190 40870 -140
rect 40920 -190 40940 -140
rect 37640 -205 37680 -200
rect 37645 -325 37675 -205
rect 38325 -325 38355 -195
rect 38835 -325 38865 -195
rect 34235 -365 34245 -335
rect 34275 -365 34285 -335
rect 34235 -375 34285 -365
rect 34915 -335 34965 -325
rect 34915 -365 34925 -335
rect 34955 -365 34965 -335
rect 34915 -375 34965 -365
rect 35765 -335 35815 -325
rect 35765 -365 35775 -335
rect 35805 -365 35815 -335
rect 35765 -375 35815 -365
rect 36445 -335 36495 -325
rect 36445 -365 36455 -335
rect 36485 -365 36495 -335
rect 36445 -375 36495 -365
rect 36955 -335 37005 -325
rect 36955 -365 36965 -335
rect 36995 -365 37005 -335
rect 36955 -375 37005 -365
rect 37635 -335 37685 -325
rect 37635 -365 37645 -335
rect 37675 -365 37685 -335
rect 37635 -375 37685 -365
rect 38315 -335 38365 -325
rect 38315 -365 38325 -335
rect 38355 -365 38365 -335
rect 38315 -375 38365 -365
rect 38825 -335 38875 -325
rect 38825 -365 38835 -335
rect 38865 -365 38875 -335
rect 38825 -375 38875 -365
rect 39505 -335 39555 -195
rect 39505 -365 39515 -335
rect 39545 -365 39555 -335
rect 39505 -375 39555 -365
rect 40185 -335 40235 -195
rect 40850 -200 40940 -190
rect 41695 -140 41785 -130
rect 41695 -190 41715 -140
rect 41765 -190 41785 -140
rect 41695 -200 41785 -190
rect 42375 -135 42465 -125
rect 42375 -185 42395 -135
rect 42445 -185 42465 -135
rect 42375 -195 42465 -185
rect 42885 -135 42975 -125
rect 43595 -130 43625 -125
rect 42885 -185 42905 -135
rect 42955 -185 42975 -135
rect 42885 -195 42975 -185
rect 43565 -140 43655 -130
rect 43565 -190 43585 -140
rect 43635 -190 43655 -140
rect 40875 -325 40905 -200
rect 41720 -205 41760 -200
rect 41725 -325 41755 -205
rect 42405 -325 42435 -195
rect 42915 -325 42945 -195
rect 43565 -200 43655 -190
rect 43590 -205 43630 -200
rect 43595 -325 43625 -205
rect 40185 -365 40195 -335
rect 40225 -365 40235 -335
rect 40185 -375 40235 -365
rect 40865 -335 40915 -325
rect 40865 -365 40875 -335
rect 40905 -365 40915 -335
rect 40865 -375 40915 -365
rect 41715 -335 41765 -325
rect 41715 -365 41725 -335
rect 41755 -365 41765 -335
rect 41715 -375 41765 -365
rect 42395 -335 42445 -325
rect 42395 -365 42405 -335
rect 42435 -365 42445 -335
rect 42395 -375 42445 -365
rect 42905 -335 42955 -325
rect 42905 -365 42915 -335
rect 42945 -365 42955 -335
rect 42905 -375 42955 -365
rect 43585 -335 43635 -325
rect 43585 -365 43595 -335
rect 43625 -365 43635 -335
rect 43585 -375 43635 -365
rect 145 -435 205 -430
rect 145 -480 155 -435
rect 195 -480 205 -435
rect 145 -485 205 -480
rect 315 -435 375 -430
rect 315 -480 325 -435
rect 365 -480 375 -435
rect 315 -485 375 -480
rect 485 -435 545 -430
rect 485 -480 495 -435
rect 535 -480 545 -435
rect 485 -485 545 -480
rect 655 -435 715 -430
rect 655 -480 665 -435
rect 705 -480 715 -435
rect 655 -485 715 -480
rect 825 -435 885 -430
rect 825 -480 835 -435
rect 875 -480 885 -435
rect 825 -485 885 -480
rect 995 -435 1055 -430
rect 995 -480 1005 -435
rect 1045 -480 1055 -435
rect 995 -485 1055 -480
rect 1165 -435 1225 -430
rect 1165 -480 1175 -435
rect 1215 -480 1225 -435
rect 1165 -485 1225 -480
rect 1335 -435 1395 -430
rect 1335 -480 1345 -435
rect 1385 -480 1395 -435
rect 1335 -485 1395 -480
rect 1505 -435 1565 -430
rect 1505 -480 1515 -435
rect 1555 -480 1565 -435
rect 1505 -485 1565 -480
rect 1675 -435 1735 -430
rect 1675 -480 1685 -435
rect 1725 -480 1735 -435
rect 1675 -485 1735 -480
rect 1845 -435 1905 -430
rect 1845 -480 1855 -435
rect 1895 -480 1905 -435
rect 1845 -485 1905 -480
rect 2015 -435 2075 -430
rect 2015 -480 2025 -435
rect 2065 -480 2075 -435
rect 2015 -485 2075 -480
rect 2185 -435 2245 -430
rect 2185 -480 2195 -435
rect 2235 -480 2245 -435
rect 2185 -485 2245 -480
rect 2355 -435 2415 -430
rect 2355 -480 2365 -435
rect 2405 -480 2415 -435
rect 2355 -485 2415 -480
rect 2525 -435 2585 -430
rect 2525 -480 2535 -435
rect 2575 -480 2585 -435
rect 2525 -485 2585 -480
rect 2695 -435 2755 -430
rect 2695 -480 2705 -435
rect 2745 -480 2755 -435
rect 2695 -485 2755 -480
rect 2865 -435 2925 -430
rect 2865 -480 2875 -435
rect 2915 -480 2925 -435
rect 2865 -485 2925 -480
rect 3035 -435 3095 -430
rect 3035 -480 3045 -435
rect 3085 -480 3095 -435
rect 3035 -485 3095 -480
rect 3205 -435 3265 -430
rect 3205 -480 3215 -435
rect 3255 -480 3265 -435
rect 3205 -485 3265 -480
rect 3375 -435 3435 -430
rect 3375 -480 3385 -435
rect 3425 -480 3435 -435
rect 3375 -485 3435 -480
rect 3545 -435 3605 -430
rect 3545 -480 3555 -435
rect 3595 -480 3605 -435
rect 3545 -485 3605 -480
rect 3715 -435 3775 -430
rect 3715 -480 3725 -435
rect 3765 -480 3775 -435
rect 3715 -485 3775 -480
rect 3885 -435 3945 -430
rect 3885 -480 3895 -435
rect 3935 -480 3945 -435
rect 3885 -485 3945 -480
rect 4055 -435 4115 -430
rect 4055 -480 4065 -435
rect 4105 -480 4115 -435
rect 4055 -485 4115 -480
rect 4225 -435 4285 -430
rect 4225 -480 4235 -435
rect 4275 -480 4285 -435
rect 4225 -485 4285 -480
rect 4395 -435 4455 -430
rect 4395 -480 4405 -435
rect 4445 -480 4455 -435
rect 4395 -485 4455 -480
rect 4565 -435 4625 -430
rect 4565 -480 4575 -435
rect 4615 -480 4625 -435
rect 4565 -485 4625 -480
rect 4735 -435 4795 -430
rect 4735 -480 4745 -435
rect 4785 -480 4795 -435
rect 4735 -485 4795 -480
rect 4905 -435 4965 -430
rect 4905 -480 4915 -435
rect 4955 -480 4965 -435
rect 4905 -485 4965 -480
rect 5075 -435 5135 -430
rect 5075 -480 5085 -435
rect 5125 -480 5135 -435
rect 5075 -485 5135 -480
rect 5245 -435 5305 -430
rect 5245 -480 5255 -435
rect 5295 -480 5305 -435
rect 5245 -485 5305 -480
rect 5415 -435 5475 -430
rect 5415 -480 5425 -435
rect 5465 -480 5475 -435
rect 5415 -485 5475 -480
rect 5585 -435 5645 -430
rect 5585 -480 5595 -435
rect 5635 -480 5645 -435
rect 5585 -485 5645 -480
rect 5755 -435 5815 -430
rect 5755 -480 5765 -435
rect 5805 -480 5815 -435
rect 5755 -485 5815 -480
rect 5925 -435 5985 -430
rect 5925 -480 5935 -435
rect 5975 -480 5985 -435
rect 5925 -485 5985 -480
rect 6095 -435 6155 -430
rect 6095 -480 6105 -435
rect 6145 -480 6155 -435
rect 6095 -485 6155 -480
rect 6265 -435 6325 -430
rect 6265 -480 6275 -435
rect 6315 -480 6325 -435
rect 6265 -485 6325 -480
rect 6435 -435 6495 -430
rect 6435 -480 6445 -435
rect 6485 -480 6495 -435
rect 6435 -485 6495 -480
rect 6605 -435 6665 -430
rect 6605 -480 6615 -435
rect 6655 -480 6665 -435
rect 6605 -485 6665 -480
rect 6775 -435 6835 -430
rect 6775 -480 6785 -435
rect 6825 -480 6835 -435
rect 6775 -485 6835 -480
rect 6945 -435 7005 -430
rect 6945 -480 6955 -435
rect 6995 -480 7005 -435
rect 6945 -485 7005 -480
rect 7115 -435 7175 -430
rect 7115 -480 7125 -435
rect 7165 -480 7175 -435
rect 7115 -485 7175 -480
rect 7285 -435 7345 -430
rect 7285 -480 7295 -435
rect 7335 -480 7345 -435
rect 7285 -485 7345 -480
rect 7455 -435 7515 -430
rect 7455 -480 7465 -435
rect 7505 -480 7515 -435
rect 7455 -485 7515 -480
rect 7625 -435 7685 -430
rect 7625 -480 7635 -435
rect 7675 -480 7685 -435
rect 7625 -485 7685 -480
rect 7795 -435 7855 -430
rect 7795 -480 7805 -435
rect 7845 -480 7855 -435
rect 7795 -485 7855 -480
rect 7965 -435 8025 -430
rect 7965 -480 7975 -435
rect 8015 -480 8025 -435
rect 7965 -485 8025 -480
rect 8135 -435 8195 -430
rect 8135 -480 8145 -435
rect 8185 -480 8195 -435
rect 8135 -485 8195 -480
rect 8305 -435 8365 -430
rect 8305 -480 8315 -435
rect 8355 -480 8365 -435
rect 8305 -485 8365 -480
rect 8475 -435 8535 -430
rect 8475 -480 8485 -435
rect 8525 -480 8535 -435
rect 8475 -485 8535 -480
rect 8645 -435 8705 -430
rect 8645 -480 8655 -435
rect 8695 -480 8705 -435
rect 8645 -485 8705 -480
rect 8815 -435 8875 -430
rect 8815 -480 8825 -435
rect 8865 -480 8875 -435
rect 8815 -485 8875 -480
rect 8985 -435 9045 -430
rect 8985 -480 8995 -435
rect 9035 -480 9045 -435
rect 8985 -485 9045 -480
rect 9155 -435 9215 -430
rect 9155 -480 9165 -435
rect 9205 -480 9215 -435
rect 9155 -485 9215 -480
rect 9325 -435 9385 -430
rect 9325 -480 9335 -435
rect 9375 -480 9385 -435
rect 9325 -485 9385 -480
rect 9495 -435 9555 -430
rect 9495 -480 9505 -435
rect 9545 -480 9555 -435
rect 9495 -485 9555 -480
rect 9665 -435 9725 -430
rect 9665 -480 9675 -435
rect 9715 -480 9725 -435
rect 9665 -485 9725 -480
rect 9835 -435 9895 -430
rect 9835 -480 9845 -435
rect 9885 -480 9895 -435
rect 9835 -485 9895 -480
rect 10005 -435 10065 -430
rect 10005 -480 10015 -435
rect 10055 -480 10065 -435
rect 10005 -485 10065 -480
rect 10175 -435 10235 -430
rect 10175 -480 10185 -435
rect 10225 -480 10235 -435
rect 10175 -485 10235 -480
rect 10345 -435 10405 -430
rect 10345 -480 10355 -435
rect 10395 -480 10405 -435
rect 10345 -485 10405 -480
rect 10515 -435 10575 -430
rect 10515 -480 10525 -435
rect 10565 -480 10575 -435
rect 10515 -485 10575 -480
rect 10685 -435 10745 -430
rect 10685 -480 10695 -435
rect 10735 -480 10745 -435
rect 10685 -485 10745 -480
rect 10855 -435 10915 -430
rect 10855 -480 10865 -435
rect 10905 -480 10915 -435
rect 10855 -485 10915 -480
rect 11025 -435 11085 -430
rect 11025 -480 11035 -435
rect 11075 -480 11085 -435
rect 11025 -485 11085 -480
rect 11195 -435 11255 -430
rect 11195 -480 11205 -435
rect 11245 -480 11255 -435
rect 11195 -485 11255 -480
rect 11365 -435 11425 -430
rect 11365 -480 11375 -435
rect 11415 -480 11425 -435
rect 11365 -485 11425 -480
rect 11535 -435 11595 -430
rect 11535 -480 11545 -435
rect 11585 -480 11595 -435
rect 11535 -485 11595 -480
rect 11705 -435 11765 -430
rect 11705 -480 11715 -435
rect 11755 -480 11765 -435
rect 11705 -485 11765 -480
rect 11875 -435 11935 -430
rect 11875 -480 11885 -435
rect 11925 -480 11935 -435
rect 11875 -485 11935 -480
rect 12045 -435 12105 -430
rect 12045 -480 12055 -435
rect 12095 -480 12105 -435
rect 12045 -485 12105 -480
rect 12215 -435 12275 -430
rect 12215 -480 12225 -435
rect 12265 -480 12275 -435
rect 12215 -485 12275 -480
rect 12385 -435 12445 -430
rect 12385 -480 12395 -435
rect 12435 -480 12445 -435
rect 12385 -485 12445 -480
rect 12555 -435 12615 -430
rect 12555 -480 12565 -435
rect 12605 -480 12615 -435
rect 12555 -485 12615 -480
rect 12725 -435 12785 -430
rect 12725 -480 12735 -435
rect 12775 -480 12785 -435
rect 12725 -485 12785 -480
rect 12895 -435 12955 -430
rect 12895 -480 12905 -435
rect 12945 -480 12955 -435
rect 12895 -485 12955 -480
rect 13065 -435 13125 -430
rect 13065 -480 13075 -435
rect 13115 -480 13125 -435
rect 13065 -485 13125 -480
rect 13235 -435 13295 -430
rect 13235 -480 13245 -435
rect 13285 -480 13295 -435
rect 13235 -485 13295 -480
rect 13405 -435 13465 -430
rect 13405 -480 13415 -435
rect 13455 -480 13465 -435
rect 13405 -485 13465 -480
rect 13575 -435 13635 -430
rect 13575 -480 13585 -435
rect 13625 -480 13635 -435
rect 13575 -485 13635 -480
rect 13745 -435 13805 -430
rect 13745 -480 13755 -435
rect 13795 -480 13805 -435
rect 13745 -485 13805 -480
rect 13915 -435 13975 -430
rect 13915 -480 13925 -435
rect 13965 -480 13975 -435
rect 13915 -485 13975 -480
rect 14085 -435 14145 -430
rect 14085 -480 14095 -435
rect 14135 -480 14145 -435
rect 14085 -485 14145 -480
rect 14255 -435 14315 -430
rect 14255 -480 14265 -435
rect 14305 -480 14315 -435
rect 14255 -485 14315 -480
rect 14425 -435 14485 -430
rect 14425 -480 14435 -435
rect 14475 -480 14485 -435
rect 14425 -485 14485 -480
rect 14595 -435 14655 -430
rect 14595 -480 14605 -435
rect 14645 -480 14655 -435
rect 14595 -485 14655 -480
rect 14765 -435 14825 -430
rect 14765 -480 14775 -435
rect 14815 -480 14825 -435
rect 14765 -485 14825 -480
rect 14935 -435 14995 -430
rect 14935 -480 14945 -435
rect 14985 -480 14995 -435
rect 14935 -485 14995 -480
rect 15105 -435 15165 -430
rect 15105 -480 15115 -435
rect 15155 -480 15165 -435
rect 15105 -485 15165 -480
rect 15275 -435 15335 -430
rect 15275 -480 15285 -435
rect 15325 -480 15335 -435
rect 15275 -485 15335 -480
rect 15445 -435 15505 -430
rect 15445 -480 15455 -435
rect 15495 -480 15505 -435
rect 15445 -485 15505 -480
rect 15615 -435 15675 -430
rect 15615 -480 15625 -435
rect 15665 -480 15675 -435
rect 15615 -485 15675 -480
rect 15785 -435 15845 -430
rect 15785 -480 15795 -435
rect 15835 -480 15845 -435
rect 15785 -485 15845 -480
rect 15955 -435 16015 -430
rect 15955 -480 15965 -435
rect 16005 -480 16015 -435
rect 15955 -485 16015 -480
rect 16125 -435 16185 -430
rect 16125 -480 16135 -435
rect 16175 -480 16185 -435
rect 16125 -485 16185 -480
rect 16295 -435 16355 -430
rect 16295 -480 16305 -435
rect 16345 -480 16355 -435
rect 16295 -485 16355 -480
rect 16465 -435 16525 -430
rect 16465 -480 16475 -435
rect 16515 -480 16525 -435
rect 16465 -485 16525 -480
rect 16635 -435 16695 -430
rect 16635 -480 16645 -435
rect 16685 -480 16695 -435
rect 16635 -485 16695 -480
rect 16805 -435 16865 -430
rect 16805 -480 16815 -435
rect 16855 -480 16865 -435
rect 16805 -485 16865 -480
rect 16975 -435 17035 -430
rect 16975 -480 16985 -435
rect 17025 -480 17035 -435
rect 16975 -485 17035 -480
rect 17145 -435 17205 -430
rect 17145 -480 17155 -435
rect 17195 -480 17205 -435
rect 17145 -485 17205 -480
rect 17315 -435 17375 -430
rect 17315 -480 17325 -435
rect 17365 -480 17375 -435
rect 17315 -485 17375 -480
rect 17485 -435 17545 -430
rect 17485 -480 17495 -435
rect 17535 -480 17545 -435
rect 17485 -485 17545 -480
rect 17655 -435 17715 -430
rect 17655 -480 17665 -435
rect 17705 -480 17715 -435
rect 17655 -485 17715 -480
rect 17825 -435 17885 -430
rect 17825 -480 17835 -435
rect 17875 -480 17885 -435
rect 17825 -485 17885 -480
rect 17995 -435 18055 -430
rect 17995 -480 18005 -435
rect 18045 -480 18055 -435
rect 17995 -485 18055 -480
rect 18165 -435 18225 -430
rect 18165 -480 18175 -435
rect 18215 -480 18225 -435
rect 18165 -485 18225 -480
rect 18335 -435 18395 -430
rect 18335 -480 18345 -435
rect 18385 -480 18395 -435
rect 18335 -485 18395 -480
rect 18505 -435 18565 -430
rect 18505 -480 18515 -435
rect 18555 -480 18565 -435
rect 18505 -485 18565 -480
rect 18675 -435 18735 -430
rect 18675 -480 18685 -435
rect 18725 -480 18735 -435
rect 18675 -485 18735 -480
rect 18845 -435 18905 -430
rect 18845 -480 18855 -435
rect 18895 -480 18905 -435
rect 18845 -485 18905 -480
rect 19015 -435 19075 -430
rect 19015 -480 19025 -435
rect 19065 -480 19075 -435
rect 19015 -485 19075 -480
rect 19185 -435 19245 -430
rect 19185 -480 19195 -435
rect 19235 -480 19245 -435
rect 19185 -485 19245 -480
rect 19355 -435 19415 -430
rect 19355 -480 19365 -435
rect 19405 -480 19415 -435
rect 19355 -485 19415 -480
rect 19525 -435 19585 -430
rect 19525 -480 19535 -435
rect 19575 -480 19585 -435
rect 19525 -485 19585 -480
rect 19695 -435 19755 -430
rect 19695 -480 19705 -435
rect 19745 -480 19755 -435
rect 19695 -485 19755 -480
rect 19865 -435 19925 -430
rect 19865 -480 19875 -435
rect 19915 -480 19925 -435
rect 19865 -485 19925 -480
rect 20035 -435 20095 -430
rect 20035 -480 20045 -435
rect 20085 -480 20095 -435
rect 20035 -485 20095 -480
rect 20205 -435 20265 -430
rect 20205 -480 20215 -435
rect 20255 -480 20265 -435
rect 20205 -485 20265 -480
rect 20375 -435 20435 -430
rect 20375 -480 20385 -435
rect 20425 -480 20435 -435
rect 20375 -485 20435 -480
rect 20545 -435 20605 -430
rect 20545 -480 20555 -435
rect 20595 -480 20605 -435
rect 20545 -485 20605 -480
rect 20715 -435 20775 -430
rect 20715 -480 20725 -435
rect 20765 -480 20775 -435
rect 20715 -485 20775 -480
rect 20885 -435 20945 -430
rect 20885 -480 20895 -435
rect 20935 -480 20945 -435
rect 20885 -485 20945 -480
rect 21055 -435 21115 -430
rect 21055 -480 21065 -435
rect 21105 -480 21115 -435
rect 21055 -485 21115 -480
rect 21225 -435 21285 -430
rect 21225 -480 21235 -435
rect 21275 -480 21285 -435
rect 21225 -485 21285 -480
rect 21395 -435 21455 -430
rect 21395 -480 21405 -435
rect 21445 -480 21455 -435
rect 21395 -485 21455 -480
rect 21565 -435 21625 -430
rect 21565 -480 21575 -435
rect 21615 -480 21625 -435
rect 21565 -485 21625 -480
rect 21735 -435 21795 -430
rect 21735 -480 21745 -435
rect 21785 -480 21795 -435
rect 21735 -485 21795 -480
rect 21905 -435 21965 -430
rect 21905 -480 21915 -435
rect 21955 -480 21965 -435
rect 21905 -485 21965 -480
rect 22075 -435 22135 -430
rect 22075 -480 22085 -435
rect 22125 -480 22135 -435
rect 22075 -485 22135 -480
rect 22245 -435 22305 -430
rect 22245 -480 22255 -435
rect 22295 -480 22305 -435
rect 22245 -485 22305 -480
rect 22415 -435 22475 -430
rect 22415 -480 22425 -435
rect 22465 -480 22475 -435
rect 22415 -485 22475 -480
rect 22585 -435 22645 -430
rect 22585 -480 22595 -435
rect 22635 -480 22645 -435
rect 22585 -485 22645 -480
rect 22755 -435 22815 -430
rect 22755 -480 22765 -435
rect 22805 -480 22815 -435
rect 22755 -485 22815 -480
rect 22925 -435 22985 -430
rect 22925 -480 22935 -435
rect 22975 -480 22985 -435
rect 22925 -485 22985 -480
rect 23095 -435 23155 -430
rect 23095 -480 23105 -435
rect 23145 -480 23155 -435
rect 23095 -485 23155 -480
rect 23265 -435 23325 -430
rect 23265 -480 23275 -435
rect 23315 -480 23325 -435
rect 23265 -485 23325 -480
rect 23435 -435 23495 -430
rect 23435 -480 23445 -435
rect 23485 -480 23495 -435
rect 23435 -485 23495 -480
rect 23605 -435 23665 -430
rect 23605 -480 23615 -435
rect 23655 -480 23665 -435
rect 23605 -485 23665 -480
rect 23775 -435 23835 -430
rect 23775 -480 23785 -435
rect 23825 -480 23835 -435
rect 23775 -485 23835 -480
rect 23945 -435 24005 -430
rect 23945 -480 23955 -435
rect 23995 -480 24005 -435
rect 23945 -485 24005 -480
rect 24115 -435 24175 -430
rect 24115 -480 24125 -435
rect 24165 -480 24175 -435
rect 24115 -485 24175 -480
rect 24285 -435 24345 -430
rect 24285 -480 24295 -435
rect 24335 -480 24345 -435
rect 24285 -485 24345 -480
rect 24455 -435 24515 -430
rect 24455 -480 24465 -435
rect 24505 -480 24515 -435
rect 24455 -485 24515 -480
rect 24625 -435 24685 -430
rect 24625 -480 24635 -435
rect 24675 -480 24685 -435
rect 24625 -485 24685 -480
rect 24795 -435 24855 -430
rect 24795 -480 24805 -435
rect 24845 -480 24855 -435
rect 24795 -485 24855 -480
rect 24965 -435 25025 -430
rect 24965 -480 24975 -435
rect 25015 -480 25025 -435
rect 24965 -485 25025 -480
rect 25135 -435 25195 -430
rect 25135 -480 25145 -435
rect 25185 -480 25195 -435
rect 25135 -485 25195 -480
rect 25305 -435 25365 -430
rect 25305 -480 25315 -435
rect 25355 -480 25365 -435
rect 25305 -485 25365 -480
rect 25475 -435 25535 -430
rect 25475 -480 25485 -435
rect 25525 -480 25535 -435
rect 25475 -485 25535 -480
rect 25645 -435 25705 -430
rect 25645 -480 25655 -435
rect 25695 -480 25705 -435
rect 25645 -485 25705 -480
rect 25815 -435 25875 -430
rect 25815 -480 25825 -435
rect 25865 -480 25875 -435
rect 25815 -485 25875 -480
rect 25985 -435 26045 -430
rect 25985 -480 25995 -435
rect 26035 -480 26045 -435
rect 25985 -485 26045 -480
rect 26155 -435 26215 -430
rect 26155 -480 26165 -435
rect 26205 -480 26215 -435
rect 26155 -485 26215 -480
rect 26325 -435 26385 -430
rect 26325 -480 26335 -435
rect 26375 -480 26385 -435
rect 26325 -485 26385 -480
rect 26495 -435 26555 -430
rect 26495 -480 26505 -435
rect 26545 -480 26555 -435
rect 26495 -485 26555 -480
rect 26665 -435 26725 -430
rect 26665 -480 26675 -435
rect 26715 -480 26725 -435
rect 26665 -485 26725 -480
rect 26835 -435 26895 -430
rect 26835 -480 26845 -435
rect 26885 -480 26895 -435
rect 26835 -485 26895 -480
rect 27005 -435 27065 -430
rect 27005 -480 27015 -435
rect 27055 -480 27065 -435
rect 27005 -485 27065 -480
rect 27175 -435 27235 -430
rect 27175 -480 27185 -435
rect 27225 -480 27235 -435
rect 27175 -485 27235 -480
rect 27345 -435 27405 -430
rect 27345 -480 27355 -435
rect 27395 -480 27405 -435
rect 27345 -485 27405 -480
rect 27515 -435 27575 -430
rect 27515 -480 27525 -435
rect 27565 -480 27575 -435
rect 27515 -485 27575 -480
rect 27685 -435 27745 -430
rect 27685 -480 27695 -435
rect 27735 -480 27745 -435
rect 27685 -485 27745 -480
rect 27855 -435 27915 -430
rect 27855 -480 27865 -435
rect 27905 -480 27915 -435
rect 27855 -485 27915 -480
rect 28025 -435 28085 -430
rect 28025 -480 28035 -435
rect 28075 -480 28085 -435
rect 28025 -485 28085 -480
rect 28195 -435 28255 -430
rect 28195 -480 28205 -435
rect 28245 -480 28255 -435
rect 28195 -485 28255 -480
rect 28365 -435 28425 -430
rect 28365 -480 28375 -435
rect 28415 -480 28425 -435
rect 28365 -485 28425 -480
rect 28535 -435 28595 -430
rect 28535 -480 28545 -435
rect 28585 -480 28595 -435
rect 28535 -485 28595 -480
rect 28705 -435 28765 -430
rect 28705 -480 28715 -435
rect 28755 -480 28765 -435
rect 28705 -485 28765 -480
rect 28875 -435 28935 -430
rect 28875 -480 28885 -435
rect 28925 -480 28935 -435
rect 28875 -485 28935 -480
rect 29045 -435 29105 -430
rect 29045 -480 29055 -435
rect 29095 -480 29105 -435
rect 29045 -485 29105 -480
rect 29215 -435 29275 -430
rect 29215 -480 29225 -435
rect 29265 -480 29275 -435
rect 29215 -485 29275 -480
rect 29385 -435 29445 -430
rect 29385 -480 29395 -435
rect 29435 -480 29445 -435
rect 29385 -485 29445 -480
rect 29555 -435 29615 -430
rect 29555 -480 29565 -435
rect 29605 -480 29615 -435
rect 29555 -485 29615 -480
rect 29725 -435 29785 -430
rect 29725 -480 29735 -435
rect 29775 -480 29785 -435
rect 29725 -485 29785 -480
rect 29895 -435 29955 -430
rect 29895 -480 29905 -435
rect 29945 -480 29955 -435
rect 29895 -485 29955 -480
rect 30065 -435 30125 -430
rect 30065 -480 30075 -435
rect 30115 -480 30125 -435
rect 30065 -485 30125 -480
rect 30235 -435 30295 -430
rect 30235 -480 30245 -435
rect 30285 -480 30295 -435
rect 30235 -485 30295 -480
rect 30405 -435 30465 -430
rect 30405 -480 30415 -435
rect 30455 -480 30465 -435
rect 30405 -485 30465 -480
rect 30575 -435 30635 -430
rect 30575 -480 30585 -435
rect 30625 -480 30635 -435
rect 30575 -485 30635 -480
rect 30745 -435 30805 -430
rect 30745 -480 30755 -435
rect 30795 -480 30805 -435
rect 30745 -485 30805 -480
rect 30915 -435 30975 -430
rect 30915 -480 30925 -435
rect 30965 -480 30975 -435
rect 30915 -485 30975 -480
rect 31085 -435 31145 -430
rect 31085 -480 31095 -435
rect 31135 -480 31145 -435
rect 31085 -485 31145 -480
rect 31255 -435 31315 -430
rect 31255 -480 31265 -435
rect 31305 -480 31315 -435
rect 31255 -485 31315 -480
rect 31425 -435 31485 -430
rect 31425 -480 31435 -435
rect 31475 -480 31485 -435
rect 31425 -485 31485 -480
rect 31595 -435 31655 -430
rect 31595 -480 31605 -435
rect 31645 -480 31655 -435
rect 31595 -485 31655 -480
rect 31765 -435 31825 -430
rect 31765 -480 31775 -435
rect 31815 -480 31825 -435
rect 31765 -485 31825 -480
rect 31935 -435 31995 -430
rect 31935 -480 31945 -435
rect 31985 -480 31995 -435
rect 31935 -485 31995 -480
rect 32105 -435 32165 -430
rect 32105 -480 32115 -435
rect 32155 -480 32165 -435
rect 32105 -485 32165 -480
rect 32275 -435 32335 -430
rect 32275 -480 32285 -435
rect 32325 -480 32335 -435
rect 32275 -485 32335 -480
rect 32445 -435 32505 -430
rect 32445 -480 32455 -435
rect 32495 -480 32505 -435
rect 32445 -485 32505 -480
rect 32615 -435 32675 -430
rect 32615 -480 32625 -435
rect 32665 -480 32675 -435
rect 32615 -485 32675 -480
rect 32785 -435 32845 -430
rect 32785 -480 32795 -435
rect 32835 -480 32845 -435
rect 32785 -485 32845 -480
rect 32955 -435 33015 -430
rect 32955 -480 32965 -435
rect 33005 -480 33015 -435
rect 32955 -485 33015 -480
rect 33125 -435 33185 -430
rect 33125 -480 33135 -435
rect 33175 -480 33185 -435
rect 33125 -485 33185 -480
rect 33295 -435 33355 -430
rect 33295 -480 33305 -435
rect 33345 -480 33355 -435
rect 33295 -485 33355 -480
rect 33465 -435 33525 -430
rect 33465 -480 33475 -435
rect 33515 -480 33525 -435
rect 33465 -485 33525 -480
rect 33635 -435 33695 -430
rect 33635 -480 33645 -435
rect 33685 -480 33695 -435
rect 33635 -485 33695 -480
rect 33805 -435 33865 -430
rect 33805 -480 33815 -435
rect 33855 -480 33865 -435
rect 33805 -485 33865 -480
rect 33975 -435 34035 -430
rect 33975 -480 33985 -435
rect 34025 -480 34035 -435
rect 33975 -485 34035 -480
rect 34145 -435 34205 -430
rect 34145 -480 34155 -435
rect 34195 -480 34205 -435
rect 34145 -485 34205 -480
rect 34315 -435 34375 -430
rect 34315 -480 34325 -435
rect 34365 -480 34375 -435
rect 34315 -485 34375 -480
rect 34485 -435 34545 -430
rect 34485 -480 34495 -435
rect 34535 -480 34545 -435
rect 34485 -485 34545 -480
rect 34655 -435 34715 -430
rect 34655 -480 34665 -435
rect 34705 -480 34715 -435
rect 34655 -485 34715 -480
rect 34825 -435 34885 -430
rect 34825 -480 34835 -435
rect 34875 -480 34885 -435
rect 34825 -485 34885 -480
rect 34995 -435 35055 -430
rect 34995 -480 35005 -435
rect 35045 -480 35055 -435
rect 34995 -485 35055 -480
rect 35165 -435 35225 -430
rect 35165 -480 35175 -435
rect 35215 -480 35225 -435
rect 35165 -485 35225 -480
rect 35335 -435 35395 -430
rect 35335 -480 35345 -435
rect 35385 -480 35395 -435
rect 35335 -485 35395 -480
rect 35505 -435 35565 -430
rect 35505 -480 35515 -435
rect 35555 -480 35565 -435
rect 35505 -485 35565 -480
rect 35675 -435 35735 -430
rect 35675 -480 35685 -435
rect 35725 -480 35735 -435
rect 35675 -485 35735 -480
rect 35845 -435 35905 -430
rect 35845 -480 35855 -435
rect 35895 -480 35905 -435
rect 35845 -485 35905 -480
rect 36015 -435 36075 -430
rect 36015 -480 36025 -435
rect 36065 -480 36075 -435
rect 36015 -485 36075 -480
rect 36185 -435 36245 -430
rect 36185 -480 36195 -435
rect 36235 -480 36245 -435
rect 36185 -485 36245 -480
rect 36355 -435 36415 -430
rect 36355 -480 36365 -435
rect 36405 -480 36415 -435
rect 36355 -485 36415 -480
rect 36525 -435 36585 -430
rect 36525 -480 36535 -435
rect 36575 -480 36585 -435
rect 36525 -485 36585 -480
rect 36695 -435 36755 -430
rect 36695 -480 36705 -435
rect 36745 -480 36755 -435
rect 36695 -485 36755 -480
rect 36865 -435 36925 -430
rect 36865 -480 36875 -435
rect 36915 -480 36925 -435
rect 36865 -485 36925 -480
rect 37035 -435 37095 -430
rect 37035 -480 37045 -435
rect 37085 -480 37095 -435
rect 37035 -485 37095 -480
rect 37205 -435 37265 -430
rect 37205 -480 37215 -435
rect 37255 -480 37265 -435
rect 37205 -485 37265 -480
rect 37375 -435 37435 -430
rect 37375 -480 37385 -435
rect 37425 -480 37435 -435
rect 37375 -485 37435 -480
rect 37545 -435 37605 -430
rect 37545 -480 37555 -435
rect 37595 -480 37605 -435
rect 37545 -485 37605 -480
rect 37715 -435 37775 -430
rect 37715 -480 37725 -435
rect 37765 -480 37775 -435
rect 37715 -485 37775 -480
rect 37885 -435 37945 -430
rect 37885 -480 37895 -435
rect 37935 -480 37945 -435
rect 37885 -485 37945 -480
rect 38055 -435 38115 -430
rect 38055 -480 38065 -435
rect 38105 -480 38115 -435
rect 38055 -485 38115 -480
rect 38225 -435 38285 -430
rect 38225 -480 38235 -435
rect 38275 -480 38285 -435
rect 38225 -485 38285 -480
rect 38395 -435 38455 -430
rect 38395 -480 38405 -435
rect 38445 -480 38455 -435
rect 38395 -485 38455 -480
rect 38565 -435 38625 -430
rect 38565 -480 38575 -435
rect 38615 -480 38625 -435
rect 38565 -485 38625 -480
rect 38735 -435 38795 -430
rect 38735 -480 38745 -435
rect 38785 -480 38795 -435
rect 38735 -485 38795 -480
rect 38905 -435 38965 -430
rect 38905 -480 38915 -435
rect 38955 -480 38965 -435
rect 38905 -485 38965 -480
rect 39075 -435 39135 -430
rect 39075 -480 39085 -435
rect 39125 -480 39135 -435
rect 39075 -485 39135 -480
rect 39245 -435 39305 -430
rect 39245 -480 39255 -435
rect 39295 -480 39305 -435
rect 39245 -485 39305 -480
rect 39415 -435 39475 -430
rect 39415 -480 39425 -435
rect 39465 -480 39475 -435
rect 39415 -485 39475 -480
rect 39585 -435 39645 -430
rect 39585 -480 39595 -435
rect 39635 -480 39645 -435
rect 39585 -485 39645 -480
rect 39755 -435 39815 -430
rect 39755 -480 39765 -435
rect 39805 -480 39815 -435
rect 39755 -485 39815 -480
rect 39925 -435 39985 -430
rect 39925 -480 39935 -435
rect 39975 -480 39985 -435
rect 39925 -485 39985 -480
rect 40095 -435 40155 -430
rect 40095 -480 40105 -435
rect 40145 -480 40155 -435
rect 40095 -485 40155 -480
rect 40265 -435 40325 -430
rect 40265 -480 40275 -435
rect 40315 -480 40325 -435
rect 40265 -485 40325 -480
rect 40435 -435 40495 -430
rect 40435 -480 40445 -435
rect 40485 -480 40495 -435
rect 40435 -485 40495 -480
rect 40605 -435 40665 -430
rect 40605 -480 40615 -435
rect 40655 -480 40665 -435
rect 40605 -485 40665 -480
rect 40775 -435 40835 -430
rect 40775 -480 40785 -435
rect 40825 -480 40835 -435
rect 40775 -485 40835 -480
rect 40945 -435 41005 -430
rect 40945 -480 40955 -435
rect 40995 -480 41005 -435
rect 40945 -485 41005 -480
rect 41115 -435 41175 -430
rect 41115 -480 41125 -435
rect 41165 -480 41175 -435
rect 41115 -485 41175 -480
rect 41285 -435 41345 -430
rect 41285 -480 41295 -435
rect 41335 -480 41345 -435
rect 41285 -485 41345 -480
rect 41455 -435 41515 -430
rect 41455 -480 41465 -435
rect 41505 -480 41515 -435
rect 41455 -485 41515 -480
rect 41625 -435 41685 -430
rect 41625 -480 41635 -435
rect 41675 -480 41685 -435
rect 41625 -485 41685 -480
rect 41795 -435 41855 -430
rect 41795 -480 41805 -435
rect 41845 -480 41855 -435
rect 41795 -485 41855 -480
rect 41965 -435 42025 -430
rect 41965 -480 41975 -435
rect 42015 -480 42025 -435
rect 41965 -485 42025 -480
rect 42135 -435 42195 -430
rect 42135 -480 42145 -435
rect 42185 -480 42195 -435
rect 42135 -485 42195 -480
rect 42305 -435 42365 -430
rect 42305 -480 42315 -435
rect 42355 -480 42365 -435
rect 42305 -485 42365 -480
rect 42475 -435 42535 -430
rect 42475 -480 42485 -435
rect 42525 -480 42535 -435
rect 42475 -485 42535 -480
rect 42645 -435 42705 -430
rect 42645 -480 42655 -435
rect 42695 -480 42705 -435
rect 42645 -485 42705 -480
rect 42815 -435 42875 -430
rect 42815 -480 42825 -435
rect 42865 -480 42875 -435
rect 42815 -485 42875 -480
rect 42985 -435 43045 -430
rect 42985 -480 42995 -435
rect 43035 -480 43045 -435
rect 42985 -485 43045 -480
rect 43155 -435 43215 -430
rect 43155 -480 43165 -435
rect 43205 -480 43215 -435
rect 43155 -485 43215 -480
rect 43325 -435 43385 -430
rect 43325 -480 43335 -435
rect 43375 -480 43385 -435
rect 43325 -485 43385 -480
rect 43495 -435 43555 -430
rect 43495 -480 43505 -435
rect 43545 -480 43555 -435
rect 43495 -485 43555 -480
rect 65 -550 115 -540
rect 65 -580 75 -550
rect 105 -580 115 -550
rect 65 -650 115 -580
rect 65 -680 75 -650
rect 105 -680 115 -650
rect 65 -710 115 -680
rect 745 -550 795 -540
rect 745 -580 755 -550
rect 785 -580 795 -550
rect 745 -650 795 -580
rect 745 -680 755 -650
rect 785 -680 795 -650
rect 745 -710 795 -680
rect 1425 -550 1475 -540
rect 1425 -580 1435 -550
rect 1465 -580 1475 -550
rect 1425 -650 1475 -580
rect 1425 -680 1435 -650
rect 1465 -680 1475 -650
rect 1425 -710 1475 -680
rect 2105 -550 2155 -540
rect 2105 -580 2115 -550
rect 2145 -580 2155 -550
rect 2105 -650 2155 -580
rect 2105 -680 2115 -650
rect 2145 -680 2155 -650
rect 2105 -710 2155 -680
rect 2785 -550 2835 -540
rect 2785 -580 2795 -550
rect 2825 -580 2835 -550
rect 2785 -650 2835 -580
rect 2785 -680 2795 -650
rect 2825 -680 2835 -650
rect 2785 -710 2835 -680
rect 3465 -550 3515 -540
rect 3465 -580 3475 -550
rect 3505 -580 3515 -550
rect 3465 -650 3515 -580
rect 3465 -680 3475 -650
rect 3505 -680 3515 -650
rect 3465 -710 3515 -680
rect 4145 -550 4195 -540
rect 4145 -580 4155 -550
rect 4185 -580 4195 -550
rect 4145 -650 4195 -580
rect 4145 -680 4155 -650
rect 4185 -680 4195 -650
rect 4145 -710 4195 -680
rect 4825 -550 4875 -540
rect 4825 -580 4835 -550
rect 4865 -580 4875 -550
rect 4825 -650 4875 -580
rect 4825 -680 4835 -650
rect 4865 -680 4875 -650
rect 4825 -710 4875 -680
rect 5505 -550 5555 -540
rect 5505 -580 5515 -550
rect 5545 -580 5555 -550
rect 5505 -650 5555 -580
rect 5505 -680 5515 -650
rect 5545 -680 5555 -650
rect 5505 -710 5555 -680
rect 6185 -550 6235 -540
rect 6185 -580 6195 -550
rect 6225 -580 6235 -550
rect 6185 -650 6235 -580
rect 6185 -680 6195 -650
rect 6225 -680 6235 -650
rect 6185 -710 6235 -680
rect 6865 -550 6915 -540
rect 6865 -580 6875 -550
rect 6905 -580 6915 -550
rect 6865 -650 6915 -580
rect 6865 -680 6875 -650
rect 6905 -680 6915 -650
rect 6865 -710 6915 -680
rect 7545 -550 7595 -540
rect 7545 -580 7555 -550
rect 7585 -580 7595 -550
rect 7545 -650 7595 -580
rect 7545 -680 7555 -650
rect 7585 -680 7595 -650
rect 7545 -710 7595 -680
rect 8225 -550 8275 -540
rect 8225 -580 8235 -550
rect 8265 -580 8275 -550
rect 8225 -650 8275 -580
rect 8225 -680 8235 -650
rect 8265 -680 8275 -650
rect 8225 -710 8275 -680
rect 8905 -550 8955 -540
rect 8905 -580 8915 -550
rect 8945 -580 8955 -550
rect 8905 -650 8955 -580
rect 8905 -680 8915 -650
rect 8945 -680 8955 -650
rect 8905 -710 8955 -680
rect 9585 -550 9635 -540
rect 9585 -580 9595 -550
rect 9625 -580 9635 -550
rect 9585 -650 9635 -580
rect 9585 -680 9595 -650
rect 9625 -680 9635 -650
rect 9585 -710 9635 -680
rect 10265 -550 10315 -540
rect 10265 -580 10275 -550
rect 10305 -580 10315 -550
rect 10265 -650 10315 -580
rect 10265 -680 10275 -650
rect 10305 -680 10315 -650
rect 10265 -710 10315 -680
rect 10945 -550 10995 -540
rect 10945 -580 10955 -550
rect 10985 -580 10995 -550
rect 10945 -650 10995 -580
rect 10945 -680 10955 -650
rect 10985 -680 10995 -650
rect 10945 -710 10995 -680
rect 11625 -550 11675 -540
rect 11625 -580 11635 -550
rect 11665 -580 11675 -550
rect 11625 -650 11675 -580
rect 11625 -680 11635 -650
rect 11665 -680 11675 -650
rect 11625 -710 11675 -680
rect 12305 -550 12355 -540
rect 12305 -580 12315 -550
rect 12345 -580 12355 -550
rect 12305 -650 12355 -580
rect 12305 -680 12315 -650
rect 12345 -680 12355 -650
rect 12305 -710 12355 -680
rect 12985 -550 13035 -540
rect 12985 -580 12995 -550
rect 13025 -580 13035 -550
rect 12985 -650 13035 -580
rect 12985 -680 12995 -650
rect 13025 -680 13035 -650
rect 12985 -710 13035 -680
rect 13665 -550 13715 -540
rect 13665 -580 13675 -550
rect 13705 -580 13715 -550
rect 13665 -650 13715 -580
rect 13665 -680 13675 -650
rect 13705 -680 13715 -650
rect 13665 -710 13715 -680
rect 14345 -550 14395 -540
rect 14345 -580 14355 -550
rect 14385 -580 14395 -550
rect 14345 -650 14395 -580
rect 14345 -680 14355 -650
rect 14385 -680 14395 -650
rect 14345 -710 14395 -680
rect 15025 -550 15075 -540
rect 15025 -580 15035 -550
rect 15065 -580 15075 -550
rect 15025 -650 15075 -580
rect 15025 -680 15035 -650
rect 15065 -680 15075 -650
rect 15025 -710 15075 -680
rect 15705 -550 15755 -540
rect 15705 -580 15715 -550
rect 15745 -580 15755 -550
rect 15705 -650 15755 -580
rect 15705 -680 15715 -650
rect 15745 -680 15755 -650
rect 15705 -710 15755 -680
rect 16385 -550 16435 -540
rect 16385 -580 16395 -550
rect 16425 -580 16435 -550
rect 16385 -650 16435 -580
rect 16385 -680 16395 -650
rect 16425 -680 16435 -650
rect 16385 -710 16435 -680
rect 17065 -550 17115 -540
rect 17065 -580 17075 -550
rect 17105 -580 17115 -550
rect 17065 -650 17115 -580
rect 17065 -680 17075 -650
rect 17105 -680 17115 -650
rect 17065 -710 17115 -680
rect 17745 -550 17795 -540
rect 17745 -580 17755 -550
rect 17785 -580 17795 -550
rect 17745 -650 17795 -580
rect 17745 -680 17755 -650
rect 17785 -680 17795 -650
rect 17745 -710 17795 -680
rect 18425 -550 18475 -540
rect 18425 -580 18435 -550
rect 18465 -580 18475 -550
rect 18425 -650 18475 -580
rect 18425 -680 18435 -650
rect 18465 -680 18475 -650
rect 18425 -710 18475 -680
rect 19105 -550 19155 -540
rect 19105 -580 19115 -550
rect 19145 -580 19155 -550
rect 19105 -650 19155 -580
rect 19105 -680 19115 -650
rect 19145 -680 19155 -650
rect 19105 -710 19155 -680
rect 19785 -550 19835 -540
rect 19785 -580 19795 -550
rect 19825 -580 19835 -550
rect 19785 -650 19835 -580
rect 19785 -680 19795 -650
rect 19825 -680 19835 -650
rect 19785 -710 19835 -680
rect 20465 -550 20515 -540
rect 20465 -580 20475 -550
rect 20505 -580 20515 -550
rect 20465 -650 20515 -580
rect 20465 -680 20475 -650
rect 20505 -680 20515 -650
rect 20465 -710 20515 -680
rect 21145 -550 21195 -540
rect 21145 -580 21155 -550
rect 21185 -580 21195 -550
rect 21145 -650 21195 -580
rect 21145 -680 21155 -650
rect 21185 -680 21195 -650
rect 21145 -710 21195 -680
rect 21825 -550 21875 -540
rect 21825 -580 21835 -550
rect 21865 -580 21875 -550
rect 21825 -650 21875 -580
rect 21825 -680 21835 -650
rect 21865 -680 21875 -650
rect 21825 -710 21875 -680
rect 22505 -550 22555 -540
rect 22505 -580 22515 -550
rect 22545 -580 22555 -550
rect 22505 -650 22555 -580
rect 22505 -680 22515 -650
rect 22545 -680 22555 -650
rect 22505 -710 22555 -680
rect 23185 -550 23235 -540
rect 23185 -580 23195 -550
rect 23225 -580 23235 -550
rect 23185 -650 23235 -580
rect 23185 -680 23195 -650
rect 23225 -680 23235 -650
rect 23185 -710 23235 -680
rect 23865 -550 23915 -540
rect 23865 -580 23875 -550
rect 23905 -580 23915 -550
rect 23865 -650 23915 -580
rect 23865 -680 23875 -650
rect 23905 -680 23915 -650
rect 23865 -710 23915 -680
rect 24545 -550 24595 -540
rect 24545 -580 24555 -550
rect 24585 -580 24595 -550
rect 24545 -650 24595 -580
rect 24545 -680 24555 -650
rect 24585 -680 24595 -650
rect 24545 -710 24595 -680
rect 25225 -550 25275 -540
rect 25225 -580 25235 -550
rect 25265 -580 25275 -550
rect 25225 -650 25275 -580
rect 25225 -680 25235 -650
rect 25265 -680 25275 -650
rect 25225 -710 25275 -680
rect 25905 -550 25955 -540
rect 25905 -580 25915 -550
rect 25945 -580 25955 -550
rect 25905 -650 25955 -580
rect 25905 -680 25915 -650
rect 25945 -680 25955 -650
rect 25905 -710 25955 -680
rect 26585 -550 26635 -540
rect 26585 -580 26595 -550
rect 26625 -580 26635 -550
rect 26585 -650 26635 -580
rect 26585 -680 26595 -650
rect 26625 -680 26635 -650
rect 26585 -710 26635 -680
rect 27265 -550 27315 -540
rect 27265 -580 27275 -550
rect 27305 -580 27315 -550
rect 27265 -650 27315 -580
rect 27265 -680 27275 -650
rect 27305 -680 27315 -650
rect 27265 -710 27315 -680
rect 27945 -550 27995 -540
rect 27945 -580 27955 -550
rect 27985 -580 27995 -550
rect 27945 -650 27995 -580
rect 27945 -680 27955 -650
rect 27985 -680 27995 -650
rect 27945 -710 27995 -680
rect 28625 -550 28675 -540
rect 28625 -580 28635 -550
rect 28665 -580 28675 -550
rect 28625 -650 28675 -580
rect 28625 -680 28635 -650
rect 28665 -680 28675 -650
rect 28625 -710 28675 -680
rect 29305 -550 29355 -540
rect 29305 -580 29315 -550
rect 29345 -580 29355 -550
rect 29305 -650 29355 -580
rect 29305 -680 29315 -650
rect 29345 -680 29355 -650
rect 29305 -710 29355 -680
rect 29985 -550 30035 -540
rect 29985 -580 29995 -550
rect 30025 -580 30035 -550
rect 29985 -650 30035 -580
rect 29985 -680 29995 -650
rect 30025 -680 30035 -650
rect 29985 -710 30035 -680
rect 30665 -550 30715 -540
rect 30665 -580 30675 -550
rect 30705 -580 30715 -550
rect 30665 -650 30715 -580
rect 30665 -680 30675 -650
rect 30705 -680 30715 -650
rect 30665 -710 30715 -680
rect 31345 -550 31395 -540
rect 31345 -580 31355 -550
rect 31385 -580 31395 -550
rect 31345 -650 31395 -580
rect 31345 -680 31355 -650
rect 31385 -680 31395 -650
rect 31345 -710 31395 -680
rect 32025 -550 32075 -540
rect 32025 -580 32035 -550
rect 32065 -580 32075 -550
rect 32025 -650 32075 -580
rect 32025 -680 32035 -650
rect 32065 -680 32075 -650
rect 32025 -710 32075 -680
rect 32705 -550 32755 -540
rect 32705 -580 32715 -550
rect 32745 -580 32755 -550
rect 32705 -650 32755 -580
rect 32705 -680 32715 -650
rect 32745 -680 32755 -650
rect 32705 -710 32755 -680
rect 33385 -550 33435 -540
rect 33385 -580 33395 -550
rect 33425 -580 33435 -550
rect 33385 -650 33435 -580
rect 33385 -680 33395 -650
rect 33425 -680 33435 -650
rect 33385 -710 33435 -680
rect 34065 -550 34115 -540
rect 34065 -580 34075 -550
rect 34105 -580 34115 -550
rect 34065 -650 34115 -580
rect 34065 -680 34075 -650
rect 34105 -680 34115 -650
rect 34065 -710 34115 -680
rect 34745 -550 34795 -540
rect 34745 -580 34755 -550
rect 34785 -580 34795 -550
rect 34745 -650 34795 -580
rect 34745 -680 34755 -650
rect 34785 -680 34795 -650
rect 34745 -710 34795 -680
rect 35425 -550 35475 -540
rect 35425 -580 35435 -550
rect 35465 -580 35475 -550
rect 35425 -650 35475 -580
rect 35425 -680 35435 -650
rect 35465 -680 35475 -650
rect 35425 -710 35475 -680
rect 36105 -550 36155 -540
rect 36105 -580 36115 -550
rect 36145 -580 36155 -550
rect 36105 -650 36155 -580
rect 36105 -680 36115 -650
rect 36145 -680 36155 -650
rect 36105 -710 36155 -680
rect 36785 -550 36835 -540
rect 36785 -580 36795 -550
rect 36825 -580 36835 -550
rect 36785 -650 36835 -580
rect 36785 -680 36795 -650
rect 36825 -680 36835 -650
rect 36785 -710 36835 -680
rect 37465 -550 37515 -540
rect 37465 -580 37475 -550
rect 37505 -580 37515 -550
rect 37465 -650 37515 -580
rect 37465 -680 37475 -650
rect 37505 -680 37515 -650
rect 37465 -710 37515 -680
rect 38145 -550 38195 -540
rect 38145 -580 38155 -550
rect 38185 -580 38195 -550
rect 38145 -650 38195 -580
rect 38145 -680 38155 -650
rect 38185 -680 38195 -650
rect 38145 -710 38195 -680
rect 38825 -550 38875 -540
rect 38825 -580 38835 -550
rect 38865 -580 38875 -550
rect 38825 -650 38875 -580
rect 38825 -680 38835 -650
rect 38865 -680 38875 -650
rect 38825 -710 38875 -680
rect 39505 -550 39555 -540
rect 39505 -580 39515 -550
rect 39545 -580 39555 -550
rect 39505 -650 39555 -580
rect 39505 -680 39515 -650
rect 39545 -680 39555 -650
rect 39505 -710 39555 -680
rect 40185 -550 40235 -540
rect 40185 -580 40195 -550
rect 40225 -580 40235 -550
rect 40185 -650 40235 -580
rect 40185 -680 40195 -650
rect 40225 -680 40235 -650
rect 40185 -710 40235 -680
rect 40865 -550 40915 -540
rect 40865 -580 40875 -550
rect 40905 -580 40915 -550
rect 40865 -650 40915 -580
rect 40865 -680 40875 -650
rect 40905 -680 40915 -650
rect 40865 -710 40915 -680
rect 41545 -550 41595 -540
rect 41545 -580 41555 -550
rect 41585 -580 41595 -550
rect 41545 -650 41595 -580
rect 41545 -680 41555 -650
rect 41585 -680 41595 -650
rect 41545 -710 41595 -680
rect 42225 -550 42275 -540
rect 42225 -580 42235 -550
rect 42265 -580 42275 -550
rect 42225 -650 42275 -580
rect 42225 -680 42235 -650
rect 42265 -680 42275 -650
rect 42225 -710 42275 -680
rect 42905 -550 42955 -540
rect 42905 -580 42915 -550
rect 42945 -580 42955 -550
rect 42905 -650 42955 -580
rect 42905 -680 42915 -650
rect 42945 -680 42955 -650
rect 42905 -710 42955 -680
rect 50 -715 130 -710
rect 50 -760 60 -715
rect 120 -760 130 -715
rect 50 -765 130 -760
rect 730 -715 810 -710
rect 730 -760 740 -715
rect 800 -760 810 -715
rect 730 -765 810 -760
rect 1410 -715 1490 -710
rect 1410 -760 1420 -715
rect 1480 -760 1490 -715
rect 1410 -765 1490 -760
rect 2090 -715 2170 -710
rect 2090 -760 2100 -715
rect 2160 -760 2170 -715
rect 2090 -765 2170 -760
rect 2770 -715 2850 -710
rect 2770 -760 2780 -715
rect 2840 -760 2850 -715
rect 2770 -765 2850 -760
rect 3450 -715 3530 -710
rect 3450 -760 3460 -715
rect 3520 -760 3530 -715
rect 3450 -765 3530 -760
rect 4130 -715 4210 -710
rect 4130 -760 4140 -715
rect 4200 -760 4210 -715
rect 4130 -765 4210 -760
rect 4810 -715 4890 -710
rect 4810 -760 4820 -715
rect 4880 -760 4890 -715
rect 4810 -765 4890 -760
rect 5490 -715 5570 -710
rect 5490 -760 5500 -715
rect 5560 -760 5570 -715
rect 5490 -765 5570 -760
rect 6170 -715 6250 -710
rect 6170 -760 6180 -715
rect 6240 -760 6250 -715
rect 6170 -765 6250 -760
rect 6850 -715 6930 -710
rect 6850 -760 6860 -715
rect 6920 -760 6930 -715
rect 6850 -765 6930 -760
rect 7530 -715 7610 -710
rect 7530 -760 7540 -715
rect 7600 -760 7610 -715
rect 7530 -765 7610 -760
rect 8210 -715 8290 -710
rect 8210 -760 8220 -715
rect 8280 -760 8290 -715
rect 8210 -765 8290 -760
rect 8890 -715 8970 -710
rect 8890 -760 8900 -715
rect 8960 -760 8970 -715
rect 8890 -765 8970 -760
rect 9570 -715 9650 -710
rect 9570 -760 9580 -715
rect 9640 -760 9650 -715
rect 9570 -765 9650 -760
rect 10250 -715 10330 -710
rect 10250 -760 10260 -715
rect 10320 -760 10330 -715
rect 10250 -765 10330 -760
rect 10930 -715 11010 -710
rect 10930 -760 10940 -715
rect 11000 -760 11010 -715
rect 10930 -765 11010 -760
rect 11610 -715 11690 -710
rect 11610 -760 11620 -715
rect 11680 -760 11690 -715
rect 11610 -765 11690 -760
rect 12290 -715 12370 -710
rect 12290 -760 12300 -715
rect 12360 -760 12370 -715
rect 12290 -765 12370 -760
rect 12970 -715 13050 -710
rect 12970 -760 12980 -715
rect 13040 -760 13050 -715
rect 12970 -765 13050 -760
rect 13650 -715 13730 -710
rect 13650 -760 13660 -715
rect 13720 -760 13730 -715
rect 13650 -765 13730 -760
rect 14330 -715 14410 -710
rect 14330 -760 14340 -715
rect 14400 -760 14410 -715
rect 14330 -765 14410 -760
rect 15010 -715 15090 -710
rect 15010 -760 15020 -715
rect 15080 -760 15090 -715
rect 15010 -765 15090 -760
rect 15690 -715 15770 -710
rect 15690 -760 15700 -715
rect 15760 -760 15770 -715
rect 15690 -765 15770 -760
rect 16370 -715 16450 -710
rect 16370 -760 16380 -715
rect 16440 -760 16450 -715
rect 16370 -765 16450 -760
rect 17050 -715 17130 -710
rect 17050 -760 17060 -715
rect 17120 -760 17130 -715
rect 17050 -765 17130 -760
rect 17730 -715 17810 -710
rect 17730 -760 17740 -715
rect 17800 -760 17810 -715
rect 17730 -765 17810 -760
rect 18410 -715 18490 -710
rect 18410 -760 18420 -715
rect 18480 -760 18490 -715
rect 18410 -765 18490 -760
rect 19090 -715 19170 -710
rect 19090 -760 19100 -715
rect 19160 -760 19170 -715
rect 19090 -765 19170 -760
rect 19770 -715 19850 -710
rect 19770 -760 19780 -715
rect 19840 -760 19850 -715
rect 19770 -765 19850 -760
rect 20450 -715 20530 -710
rect 20450 -760 20460 -715
rect 20520 -760 20530 -715
rect 20450 -765 20530 -760
rect 21130 -715 21210 -710
rect 21130 -760 21140 -715
rect 21200 -760 21210 -715
rect 21130 -765 21210 -760
rect 21815 -715 21890 -710
rect 21815 -760 21820 -715
rect 21880 -760 21890 -715
rect 21815 -765 21890 -760
rect 22490 -715 22570 -710
rect 22490 -760 22500 -715
rect 22560 -760 22570 -715
rect 22490 -765 22570 -760
rect 23170 -715 23250 -710
rect 23170 -760 23180 -715
rect 23240 -760 23250 -715
rect 23170 -765 23250 -760
rect 23850 -715 23930 -710
rect 23850 -760 23860 -715
rect 23920 -760 23930 -715
rect 23850 -765 23930 -760
rect 24530 -715 24610 -710
rect 24530 -760 24540 -715
rect 24600 -760 24610 -715
rect 24530 -765 24610 -760
rect 25210 -715 25290 -710
rect 25210 -760 25220 -715
rect 25280 -760 25290 -715
rect 25210 -765 25290 -760
rect 25890 -715 25970 -710
rect 25890 -760 25900 -715
rect 25960 -760 25970 -715
rect 25890 -765 25970 -760
rect 26570 -715 26650 -710
rect 26570 -760 26580 -715
rect 26640 -760 26650 -715
rect 26570 -765 26650 -760
rect 27250 -715 27330 -710
rect 27250 -760 27260 -715
rect 27320 -760 27330 -715
rect 27250 -765 27330 -760
rect 27930 -715 28010 -710
rect 27930 -760 27940 -715
rect 28000 -760 28010 -715
rect 27930 -765 28010 -760
rect 28610 -715 28690 -710
rect 28610 -760 28620 -715
rect 28680 -760 28690 -715
rect 28610 -765 28690 -760
rect 29290 -715 29370 -710
rect 29290 -760 29300 -715
rect 29360 -760 29370 -715
rect 29290 -765 29370 -760
rect 29970 -715 30050 -710
rect 29970 -760 29980 -715
rect 30040 -760 30050 -715
rect 29970 -765 30050 -760
rect 30650 -715 30730 -710
rect 30650 -760 30660 -715
rect 30720 -760 30730 -715
rect 30650 -765 30730 -760
rect 31330 -715 31410 -710
rect 31330 -760 31340 -715
rect 31400 -760 31410 -715
rect 31330 -765 31410 -760
rect 32010 -715 32090 -710
rect 32010 -760 32020 -715
rect 32080 -760 32090 -715
rect 32010 -765 32090 -760
rect 32690 -715 32770 -710
rect 32690 -760 32700 -715
rect 32760 -760 32770 -715
rect 32690 -765 32770 -760
rect 33370 -715 33450 -710
rect 33370 -760 33380 -715
rect 33440 -760 33450 -715
rect 33370 -765 33450 -760
rect 34050 -715 34130 -710
rect 34050 -760 34060 -715
rect 34120 -760 34130 -715
rect 34050 -765 34130 -760
rect 34730 -715 34810 -710
rect 34730 -760 34740 -715
rect 34800 -760 34810 -715
rect 34730 -765 34810 -760
rect 35410 -715 35490 -710
rect 35410 -760 35420 -715
rect 35480 -760 35490 -715
rect 35410 -765 35490 -760
rect 36090 -715 36170 -710
rect 36090 -760 36100 -715
rect 36160 -760 36170 -715
rect 36090 -765 36170 -760
rect 36770 -715 36850 -710
rect 36770 -760 36780 -715
rect 36840 -760 36850 -715
rect 36770 -765 36850 -760
rect 37450 -715 37530 -710
rect 37450 -760 37460 -715
rect 37520 -760 37530 -715
rect 37450 -765 37530 -760
rect 38130 -715 38210 -710
rect 38130 -760 38140 -715
rect 38200 -760 38210 -715
rect 38130 -765 38210 -760
rect 38810 -715 38890 -710
rect 38810 -760 38820 -715
rect 38880 -760 38890 -715
rect 38810 -765 38890 -760
rect 39490 -715 39570 -710
rect 39490 -760 39500 -715
rect 39560 -760 39570 -715
rect 39490 -765 39570 -760
rect 40170 -715 40250 -710
rect 40170 -760 40180 -715
rect 40240 -760 40250 -715
rect 40170 -765 40250 -760
rect 40850 -715 40930 -710
rect 40850 -760 40860 -715
rect 40920 -760 40930 -715
rect 40850 -765 40930 -760
rect 41530 -715 41610 -710
rect 41530 -760 41540 -715
rect 41600 -760 41610 -715
rect 41530 -765 41610 -760
rect 42210 -715 42290 -710
rect 42210 -760 42220 -715
rect 42280 -760 42290 -715
rect 42210 -765 42290 -760
rect 42890 -715 42970 -710
rect 42890 -760 42900 -715
rect 42960 -760 42970 -715
rect 42890 -765 42970 -760
<< via3 >>
rect 210 240 270 285
rect 550 240 610 285
rect 745 240 805 285
rect 1425 240 1485 285
rect 2105 240 2165 285
rect 2255 240 2315 285
rect 2935 240 2995 285
rect 3615 240 3675 285
rect 4295 240 4355 285
rect 4975 240 5035 285
rect 5655 240 5715 285
rect 6335 240 6395 285
rect 7015 240 7075 285
rect 7695 240 7755 285
rect 7845 240 7905 285
rect 8525 240 8585 285
rect 9205 240 9265 285
rect 9885 240 9945 285
rect 10565 240 10625 285
rect 11245 240 11305 285
rect 11925 240 11985 285
rect 12605 240 12665 285
rect 13285 240 13345 285
rect 13965 240 14025 285
rect 14645 240 14705 285
rect 15325 240 15385 285
rect 16005 240 16065 285
rect 16685 240 16745 285
rect 17365 240 17425 285
rect 18045 240 18105 285
rect 18725 240 18785 285
rect 19405 240 19465 285
rect 20085 240 20145 285
rect 20765 240 20825 285
rect 21445 240 21505 285
rect 22125 240 22185 285
rect 22805 240 22865 285
rect 23485 240 23545 285
rect 24165 240 24225 285
rect 24845 240 24905 285
rect 25525 240 25585 285
rect 26205 240 26265 285
rect 26885 240 26945 285
rect 27565 240 27625 285
rect 28245 240 28305 285
rect 28925 240 28985 285
rect 29605 240 29665 285
rect 305 100 345 105
rect 305 65 310 100
rect 310 65 340 100
rect 340 65 345 100
rect 305 60 345 65
rect 475 100 515 105
rect 475 65 480 100
rect 480 65 510 100
rect 510 65 515 100
rect 475 60 515 65
rect 645 60 700 105
rect 840 100 880 105
rect 840 65 845 100
rect 845 65 875 100
rect 875 65 880 100
rect 840 60 880 65
rect 1010 100 1050 105
rect 1010 65 1015 100
rect 1015 65 1045 100
rect 1045 65 1050 100
rect 1010 60 1050 65
rect 1180 100 1220 105
rect 1180 65 1185 100
rect 1185 65 1215 100
rect 1215 65 1220 100
rect 1180 60 1220 65
rect 1350 100 1390 105
rect 1350 65 1355 100
rect 1355 65 1385 100
rect 1385 65 1390 100
rect 1350 60 1390 65
rect 1520 100 1560 105
rect 1520 65 1525 100
rect 1525 65 1555 100
rect 1555 65 1560 100
rect 1520 60 1560 65
rect 1690 100 1730 105
rect 1690 65 1695 100
rect 1695 65 1725 100
rect 1725 65 1730 100
rect 1690 60 1730 65
rect 1860 100 1900 105
rect 1860 65 1865 100
rect 1865 65 1895 100
rect 1895 65 1900 100
rect 1860 60 1900 65
rect 2030 100 2070 105
rect 2030 65 2035 100
rect 2035 65 2065 100
rect 2065 65 2070 100
rect 2030 60 2070 65
rect 2185 60 2240 105
rect 2350 100 2390 105
rect 2350 65 2355 100
rect 2355 65 2385 100
rect 2385 65 2390 100
rect 2350 60 2390 65
rect 2520 100 2560 105
rect 2520 65 2525 100
rect 2525 65 2555 100
rect 2555 65 2560 100
rect 2520 60 2560 65
rect 2690 100 2730 105
rect 2690 65 2695 100
rect 2695 65 2725 100
rect 2725 65 2730 100
rect 2690 60 2730 65
rect 2860 100 2900 105
rect 2860 65 2865 100
rect 2865 65 2895 100
rect 2895 65 2900 100
rect 2860 60 2900 65
rect 3030 100 3070 105
rect 3030 65 3035 100
rect 3035 65 3065 100
rect 3065 65 3070 100
rect 3030 60 3070 65
rect 3200 100 3240 105
rect 3200 65 3205 100
rect 3205 65 3235 100
rect 3235 65 3240 100
rect 3200 60 3240 65
rect 3370 100 3410 105
rect 3370 65 3375 100
rect 3375 65 3405 100
rect 3405 65 3410 100
rect 3370 60 3410 65
rect 3540 100 3580 105
rect 3540 65 3545 100
rect 3545 65 3575 100
rect 3575 65 3580 100
rect 3540 60 3580 65
rect 3710 100 3750 105
rect 3710 65 3715 100
rect 3715 65 3745 100
rect 3745 65 3750 100
rect 3710 60 3750 65
rect 3880 100 3920 105
rect 3880 65 3885 100
rect 3885 65 3915 100
rect 3915 65 3920 100
rect 3880 60 3920 65
rect 4050 100 4090 105
rect 4050 65 4055 100
rect 4055 65 4085 100
rect 4085 65 4090 100
rect 4050 60 4090 65
rect 4220 100 4260 105
rect 4220 65 4225 100
rect 4225 65 4255 100
rect 4255 65 4260 100
rect 4220 60 4260 65
rect 4390 100 4430 105
rect 4390 65 4395 100
rect 4395 65 4425 100
rect 4425 65 4430 100
rect 4390 60 4430 65
rect 4560 100 4600 105
rect 4560 65 4565 100
rect 4565 65 4595 100
rect 4595 65 4600 100
rect 4560 60 4600 65
rect 4730 100 4770 105
rect 4730 65 4735 100
rect 4735 65 4765 100
rect 4765 65 4770 100
rect 4730 60 4770 65
rect 4900 100 4940 105
rect 4900 65 4905 100
rect 4905 65 4935 100
rect 4935 65 4940 100
rect 4900 60 4940 65
rect 5070 100 5110 105
rect 5070 65 5075 100
rect 5075 65 5105 100
rect 5105 65 5110 100
rect 5070 60 5110 65
rect 5240 100 5280 105
rect 5240 65 5245 100
rect 5245 65 5275 100
rect 5275 65 5280 100
rect 5240 60 5280 65
rect 5410 100 5450 105
rect 5410 65 5415 100
rect 5415 65 5445 100
rect 5445 65 5450 100
rect 5410 60 5450 65
rect 5580 100 5620 105
rect 5580 65 5585 100
rect 5585 65 5615 100
rect 5615 65 5620 100
rect 5580 60 5620 65
rect 5750 100 5790 105
rect 5750 65 5755 100
rect 5755 65 5785 100
rect 5785 65 5790 100
rect 5750 60 5790 65
rect 5920 100 5960 105
rect 5920 65 5925 100
rect 5925 65 5955 100
rect 5955 65 5960 100
rect 5920 60 5960 65
rect 6090 100 6130 105
rect 6090 65 6095 100
rect 6095 65 6125 100
rect 6125 65 6130 100
rect 6090 60 6130 65
rect 6260 100 6300 105
rect 6260 65 6265 100
rect 6265 65 6295 100
rect 6295 65 6300 100
rect 6260 60 6300 65
rect 6430 100 6470 105
rect 6430 65 6435 100
rect 6435 65 6465 100
rect 6465 65 6470 100
rect 6430 60 6470 65
rect 6600 100 6640 105
rect 6600 65 6605 100
rect 6605 65 6635 100
rect 6635 65 6640 100
rect 6600 60 6640 65
rect 6770 100 6810 105
rect 6770 65 6775 100
rect 6775 65 6805 100
rect 6805 65 6810 100
rect 6770 60 6810 65
rect 6940 100 6980 105
rect 6940 65 6945 100
rect 6945 65 6975 100
rect 6975 65 6980 100
rect 6940 60 6980 65
rect 7110 100 7150 105
rect 7110 65 7115 100
rect 7115 65 7145 100
rect 7145 65 7150 100
rect 7110 60 7150 65
rect 7280 100 7320 105
rect 7280 65 7285 100
rect 7285 65 7315 100
rect 7315 65 7320 100
rect 7280 60 7320 65
rect 7450 100 7490 105
rect 7450 65 7455 100
rect 7455 65 7485 100
rect 7485 65 7490 100
rect 7450 60 7490 65
rect 7620 100 7660 105
rect 7620 65 7625 100
rect 7625 65 7655 100
rect 7655 65 7660 100
rect 7620 60 7660 65
rect 7775 60 7830 105
rect 65 -185 115 -135
rect 215 -190 265 -140
rect 555 -190 605 -140
rect 745 -185 795 -135
rect 1430 -190 1480 -140
rect 2275 -190 2325 -140
rect 2430 -185 2480 -135
rect 2955 -185 3005 -135
rect 3110 -185 3160 -135
rect 3465 -185 3515 -135
rect 3620 -190 3670 -140
rect 4145 -190 4195 -140
rect 4300 -185 4350 -135
rect 4825 -185 4875 -135
rect 4980 -185 5030 -135
rect 7940 100 7980 105
rect 7940 65 7945 100
rect 7945 65 7975 100
rect 7975 65 7980 100
rect 7940 60 7980 65
rect 8110 100 8150 105
rect 8110 65 8115 100
rect 8115 65 8145 100
rect 8145 65 8150 100
rect 8110 60 8150 65
rect 8280 100 8320 105
rect 8280 65 8285 100
rect 8285 65 8315 100
rect 8315 65 8320 100
rect 8280 60 8320 65
rect 8450 100 8490 105
rect 8450 65 8455 100
rect 8455 65 8485 100
rect 8485 65 8490 100
rect 8450 60 8490 65
rect 8620 100 8660 105
rect 8620 65 8625 100
rect 8625 65 8655 100
rect 8655 65 8660 100
rect 8620 60 8660 65
rect 8790 100 8830 105
rect 8790 65 8795 100
rect 8795 65 8825 100
rect 8825 65 8830 100
rect 8790 60 8830 65
rect 8960 100 9000 105
rect 8960 65 8965 100
rect 8965 65 8995 100
rect 8995 65 9000 100
rect 8960 60 9000 65
rect 9130 100 9170 105
rect 9130 65 9135 100
rect 9135 65 9165 100
rect 9165 65 9170 100
rect 9130 60 9170 65
rect 9300 100 9340 105
rect 9300 65 9305 100
rect 9305 65 9335 100
rect 9335 65 9340 100
rect 9300 60 9340 65
rect 9470 100 9510 105
rect 9470 65 9475 100
rect 9475 65 9505 100
rect 9505 65 9510 100
rect 9470 60 9510 65
rect 9640 100 9680 105
rect 9640 65 9645 100
rect 9645 65 9675 100
rect 9675 65 9680 100
rect 9640 60 9680 65
rect 9810 100 9850 105
rect 9810 65 9815 100
rect 9815 65 9845 100
rect 9845 65 9850 100
rect 9810 60 9850 65
rect 9980 100 10020 105
rect 9980 65 9985 100
rect 9985 65 10015 100
rect 10015 65 10020 100
rect 9980 60 10020 65
rect 10150 100 10190 105
rect 10150 65 10155 100
rect 10155 65 10185 100
rect 10185 65 10190 100
rect 10150 60 10190 65
rect 10320 100 10360 105
rect 10320 65 10325 100
rect 10325 65 10355 100
rect 10355 65 10360 100
rect 10320 60 10360 65
rect 10490 100 10530 105
rect 10490 65 10495 100
rect 10495 65 10525 100
rect 10525 65 10530 100
rect 10490 60 10530 65
rect 10660 100 10700 105
rect 10660 65 10665 100
rect 10665 65 10695 100
rect 10695 65 10700 100
rect 10660 60 10700 65
rect 10830 100 10870 105
rect 10830 65 10835 100
rect 10835 65 10865 100
rect 10865 65 10870 100
rect 10830 60 10870 65
rect 11000 100 11040 105
rect 11000 65 11005 100
rect 11005 65 11035 100
rect 11035 65 11040 100
rect 11000 60 11040 65
rect 11170 100 11210 105
rect 11170 65 11175 100
rect 11175 65 11205 100
rect 11205 65 11210 100
rect 11170 60 11210 65
rect 11340 100 11380 105
rect 11340 65 11345 100
rect 11345 65 11375 100
rect 11375 65 11380 100
rect 11340 60 11380 65
rect 11510 100 11550 105
rect 11510 65 11515 100
rect 11515 65 11545 100
rect 11545 65 11550 100
rect 11510 60 11550 65
rect 11680 100 11720 105
rect 11680 65 11685 100
rect 11685 65 11715 100
rect 11715 65 11720 100
rect 11680 60 11720 65
rect 11850 100 11890 105
rect 11850 65 11855 100
rect 11855 65 11885 100
rect 11885 65 11890 100
rect 11850 60 11890 65
rect 12020 100 12060 105
rect 12020 65 12025 100
rect 12025 65 12055 100
rect 12055 65 12060 100
rect 12020 60 12060 65
rect 12190 100 12230 105
rect 12190 65 12195 100
rect 12195 65 12225 100
rect 12225 65 12230 100
rect 12190 60 12230 65
rect 12360 100 12400 105
rect 12360 65 12365 100
rect 12365 65 12395 100
rect 12395 65 12400 100
rect 12360 60 12400 65
rect 12530 100 12570 105
rect 12530 65 12535 100
rect 12535 65 12565 100
rect 12565 65 12570 100
rect 12530 60 12570 65
rect 12700 100 12740 105
rect 12700 65 12705 100
rect 12705 65 12735 100
rect 12735 65 12740 100
rect 12700 60 12740 65
rect 12870 100 12910 105
rect 12870 65 12875 100
rect 12875 65 12905 100
rect 12905 65 12910 100
rect 12870 60 12910 65
rect 13040 100 13080 105
rect 13040 65 13045 100
rect 13045 65 13075 100
rect 13075 65 13080 100
rect 13040 60 13080 65
rect 13210 100 13250 105
rect 13210 65 13215 100
rect 13215 65 13245 100
rect 13245 65 13250 100
rect 13210 60 13250 65
rect 13380 100 13420 105
rect 13380 65 13385 100
rect 13385 65 13415 100
rect 13415 65 13420 100
rect 13380 60 13420 65
rect 13550 100 13590 105
rect 13550 65 13555 100
rect 13555 65 13585 100
rect 13585 65 13590 100
rect 13550 60 13590 65
rect 13720 100 13760 105
rect 13720 65 13725 100
rect 13725 65 13755 100
rect 13755 65 13760 100
rect 13720 60 13760 65
rect 13890 100 13930 105
rect 13890 65 13895 100
rect 13895 65 13925 100
rect 13925 65 13930 100
rect 13890 60 13930 65
rect 14060 100 14100 105
rect 14060 65 14065 100
rect 14065 65 14095 100
rect 14095 65 14100 100
rect 14060 60 14100 65
rect 14230 100 14270 105
rect 14230 65 14235 100
rect 14235 65 14265 100
rect 14265 65 14270 100
rect 14230 60 14270 65
rect 14400 100 14440 105
rect 14400 65 14405 100
rect 14405 65 14435 100
rect 14435 65 14440 100
rect 14400 60 14440 65
rect 14570 100 14610 105
rect 14570 65 14575 100
rect 14575 65 14605 100
rect 14605 65 14610 100
rect 14570 60 14610 65
rect 14740 100 14780 105
rect 14740 65 14745 100
rect 14745 65 14775 100
rect 14775 65 14780 100
rect 14740 60 14780 65
rect 14910 100 14950 105
rect 14910 65 14915 100
rect 14915 65 14945 100
rect 14945 65 14950 100
rect 14910 60 14950 65
rect 15080 100 15120 105
rect 15080 65 15085 100
rect 15085 65 15115 100
rect 15115 65 15120 100
rect 15080 60 15120 65
rect 15250 100 15290 105
rect 15250 65 15255 100
rect 15255 65 15285 100
rect 15285 65 15290 100
rect 15250 60 15290 65
rect 15420 100 15460 105
rect 15420 65 15425 100
rect 15425 65 15455 100
rect 15455 65 15460 100
rect 15420 60 15460 65
rect 15590 100 15630 105
rect 15590 65 15595 100
rect 15595 65 15625 100
rect 15625 65 15630 100
rect 15590 60 15630 65
rect 15760 100 15800 105
rect 15760 65 15765 100
rect 15765 65 15795 100
rect 15795 65 15800 100
rect 15760 60 15800 65
rect 15930 100 15970 105
rect 15930 65 15935 100
rect 15935 65 15965 100
rect 15965 65 15970 100
rect 15930 60 15970 65
rect 16100 100 16140 105
rect 16100 65 16105 100
rect 16105 65 16135 100
rect 16135 65 16140 100
rect 16100 60 16140 65
rect 16270 100 16310 105
rect 16270 65 16275 100
rect 16275 65 16305 100
rect 16305 65 16310 100
rect 16270 60 16310 65
rect 16440 100 16480 105
rect 16440 65 16445 100
rect 16445 65 16475 100
rect 16475 65 16480 100
rect 16440 60 16480 65
rect 16610 100 16650 105
rect 16610 65 16615 100
rect 16615 65 16645 100
rect 16645 65 16650 100
rect 16610 60 16650 65
rect 16780 100 16820 105
rect 16780 65 16785 100
rect 16785 65 16815 100
rect 16815 65 16820 100
rect 16780 60 16820 65
rect 16950 100 16990 105
rect 16950 65 16955 100
rect 16955 65 16985 100
rect 16985 65 16990 100
rect 16950 60 16990 65
rect 17120 100 17160 105
rect 17120 65 17125 100
rect 17125 65 17155 100
rect 17155 65 17160 100
rect 17120 60 17160 65
rect 17290 100 17330 105
rect 17290 65 17295 100
rect 17295 65 17325 100
rect 17325 65 17330 100
rect 17290 60 17330 65
rect 17460 100 17500 105
rect 17460 65 17465 100
rect 17465 65 17495 100
rect 17495 65 17500 100
rect 17460 60 17500 65
rect 17630 100 17670 105
rect 17630 65 17635 100
rect 17635 65 17665 100
rect 17665 65 17670 100
rect 17630 60 17670 65
rect 17800 100 17840 105
rect 17800 65 17805 100
rect 17805 65 17835 100
rect 17835 65 17840 100
rect 17800 60 17840 65
rect 17970 100 18010 105
rect 17970 65 17975 100
rect 17975 65 18005 100
rect 18005 65 18010 100
rect 17970 60 18010 65
rect 18140 100 18180 105
rect 18140 65 18145 100
rect 18145 65 18175 100
rect 18175 65 18180 100
rect 18140 60 18180 65
rect 18310 100 18350 105
rect 18310 65 18315 100
rect 18315 65 18345 100
rect 18345 65 18350 100
rect 18310 60 18350 65
rect 18480 100 18520 105
rect 18480 65 18485 100
rect 18485 65 18515 100
rect 18515 65 18520 100
rect 18480 60 18520 65
rect 18650 100 18690 105
rect 18650 65 18655 100
rect 18655 65 18685 100
rect 18685 65 18690 100
rect 18650 60 18690 65
rect 18820 100 18860 105
rect 18820 65 18825 100
rect 18825 65 18855 100
rect 18855 65 18860 100
rect 18820 60 18860 65
rect 18990 100 19030 105
rect 18990 65 18995 100
rect 18995 65 19025 100
rect 19025 65 19030 100
rect 18990 60 19030 65
rect 19160 100 19200 105
rect 19160 65 19165 100
rect 19165 65 19195 100
rect 19195 65 19200 100
rect 19160 60 19200 65
rect 19330 100 19370 105
rect 19330 65 19335 100
rect 19335 65 19365 100
rect 19365 65 19370 100
rect 19330 60 19370 65
rect 19500 100 19540 105
rect 19500 65 19505 100
rect 19505 65 19535 100
rect 19535 65 19540 100
rect 19500 60 19540 65
rect 19670 100 19710 105
rect 19670 65 19675 100
rect 19675 65 19705 100
rect 19705 65 19710 100
rect 19670 60 19710 65
rect 19840 100 19880 105
rect 19840 65 19845 100
rect 19845 65 19875 100
rect 19875 65 19880 100
rect 19840 60 19880 65
rect 20010 100 20050 105
rect 20010 65 20015 100
rect 20015 65 20045 100
rect 20045 65 20050 100
rect 20010 60 20050 65
rect 20180 100 20220 105
rect 20180 65 20185 100
rect 20185 65 20215 100
rect 20215 65 20220 100
rect 20180 60 20220 65
rect 20350 100 20390 105
rect 20350 65 20355 100
rect 20355 65 20385 100
rect 20385 65 20390 100
rect 20350 60 20390 65
rect 20520 100 20560 105
rect 20520 65 20525 100
rect 20525 65 20555 100
rect 20555 65 20560 100
rect 20520 60 20560 65
rect 20690 100 20730 105
rect 20690 65 20695 100
rect 20695 65 20725 100
rect 20725 65 20730 100
rect 20690 60 20730 65
rect 20860 100 20900 105
rect 20860 65 20865 100
rect 20865 65 20895 100
rect 20895 65 20900 100
rect 20860 60 20900 65
rect 21030 100 21070 105
rect 21030 65 21035 100
rect 21035 65 21065 100
rect 21065 65 21070 100
rect 21030 60 21070 65
rect 21200 100 21240 105
rect 21200 65 21205 100
rect 21205 65 21235 100
rect 21235 65 21240 100
rect 21200 60 21240 65
rect 21370 100 21410 105
rect 21370 65 21375 100
rect 21375 65 21405 100
rect 21405 65 21410 100
rect 21370 60 21410 65
rect 21540 100 21580 105
rect 21540 65 21545 100
rect 21545 65 21575 100
rect 21575 65 21580 100
rect 21540 60 21580 65
rect 21710 100 21750 105
rect 21710 65 21715 100
rect 21715 65 21745 100
rect 21745 65 21750 100
rect 21710 60 21750 65
rect 21880 100 21920 105
rect 21880 65 21885 100
rect 21885 65 21915 100
rect 21915 65 21920 100
rect 21880 60 21920 65
rect 22050 100 22090 105
rect 22050 65 22055 100
rect 22055 65 22085 100
rect 22085 65 22090 100
rect 22050 60 22090 65
rect 22220 100 22260 105
rect 22220 65 22225 100
rect 22225 65 22255 100
rect 22255 65 22260 100
rect 22220 60 22260 65
rect 22390 100 22430 105
rect 22390 65 22395 100
rect 22395 65 22425 100
rect 22425 65 22430 100
rect 22390 60 22430 65
rect 22560 100 22600 105
rect 22560 65 22565 100
rect 22565 65 22595 100
rect 22595 65 22600 100
rect 22560 60 22600 65
rect 22730 100 22770 105
rect 22730 65 22735 100
rect 22735 65 22765 100
rect 22765 65 22770 100
rect 22730 60 22770 65
rect 22900 100 22940 105
rect 22900 65 22905 100
rect 22905 65 22935 100
rect 22935 65 22940 100
rect 22900 60 22940 65
rect 23070 100 23110 105
rect 23070 65 23075 100
rect 23075 65 23105 100
rect 23105 65 23110 100
rect 23070 60 23110 65
rect 23240 100 23280 105
rect 23240 65 23245 100
rect 23245 65 23275 100
rect 23275 65 23280 100
rect 23240 60 23280 65
rect 23410 100 23450 105
rect 23410 65 23415 100
rect 23415 65 23445 100
rect 23445 65 23450 100
rect 23410 60 23450 65
rect 23580 100 23620 105
rect 23580 65 23585 100
rect 23585 65 23615 100
rect 23615 65 23620 100
rect 23580 60 23620 65
rect 23750 100 23790 105
rect 23750 65 23755 100
rect 23755 65 23785 100
rect 23785 65 23790 100
rect 23750 60 23790 65
rect 23920 100 23960 105
rect 23920 65 23925 100
rect 23925 65 23955 100
rect 23955 65 23960 100
rect 23920 60 23960 65
rect 24090 100 24130 105
rect 24090 65 24095 100
rect 24095 65 24125 100
rect 24125 65 24130 100
rect 24090 60 24130 65
rect 24260 100 24300 105
rect 24260 65 24265 100
rect 24265 65 24295 100
rect 24295 65 24300 100
rect 24260 60 24300 65
rect 24430 100 24470 105
rect 24430 65 24435 100
rect 24435 65 24465 100
rect 24465 65 24470 100
rect 24430 60 24470 65
rect 24600 100 24640 105
rect 24600 65 24605 100
rect 24605 65 24635 100
rect 24635 65 24640 100
rect 24600 60 24640 65
rect 24770 100 24810 105
rect 24770 65 24775 100
rect 24775 65 24805 100
rect 24805 65 24810 100
rect 24770 60 24810 65
rect 24940 100 24980 105
rect 24940 65 24945 100
rect 24945 65 24975 100
rect 24975 65 24980 100
rect 24940 60 24980 65
rect 25110 100 25150 105
rect 25110 65 25115 100
rect 25115 65 25145 100
rect 25145 65 25150 100
rect 25110 60 25150 65
rect 25280 100 25320 105
rect 25280 65 25285 100
rect 25285 65 25315 100
rect 25315 65 25320 100
rect 25280 60 25320 65
rect 25450 100 25490 105
rect 25450 65 25455 100
rect 25455 65 25485 100
rect 25485 65 25490 100
rect 25450 60 25490 65
rect 25620 100 25660 105
rect 25620 65 25625 100
rect 25625 65 25655 100
rect 25655 65 25660 100
rect 25620 60 25660 65
rect 25790 100 25830 105
rect 25790 65 25795 100
rect 25795 65 25825 100
rect 25825 65 25830 100
rect 25790 60 25830 65
rect 25960 100 26000 105
rect 25960 65 25965 100
rect 25965 65 25995 100
rect 25995 65 26000 100
rect 25960 60 26000 65
rect 26130 100 26170 105
rect 26130 65 26135 100
rect 26135 65 26165 100
rect 26165 65 26170 100
rect 26130 60 26170 65
rect 26300 100 26340 105
rect 26300 65 26305 100
rect 26305 65 26335 100
rect 26335 65 26340 100
rect 26300 60 26340 65
rect 26470 100 26510 105
rect 26470 65 26475 100
rect 26475 65 26505 100
rect 26505 65 26510 100
rect 26470 60 26510 65
rect 26640 100 26680 105
rect 26640 65 26645 100
rect 26645 65 26675 100
rect 26675 65 26680 100
rect 26640 60 26680 65
rect 26810 100 26850 105
rect 26810 65 26815 100
rect 26815 65 26845 100
rect 26845 65 26850 100
rect 26810 60 26850 65
rect 26980 100 27020 105
rect 26980 65 26985 100
rect 26985 65 27015 100
rect 27015 65 27020 100
rect 26980 60 27020 65
rect 27150 100 27190 105
rect 27150 65 27155 100
rect 27155 65 27185 100
rect 27185 65 27190 100
rect 27150 60 27190 65
rect 27320 100 27360 105
rect 27320 65 27325 100
rect 27325 65 27355 100
rect 27355 65 27360 100
rect 27320 60 27360 65
rect 27490 100 27530 105
rect 27490 65 27495 100
rect 27495 65 27525 100
rect 27525 65 27530 100
rect 27490 60 27530 65
rect 27660 100 27700 105
rect 27660 65 27665 100
rect 27665 65 27695 100
rect 27695 65 27700 100
rect 27660 60 27700 65
rect 27830 100 27870 105
rect 27830 65 27835 100
rect 27835 65 27865 100
rect 27865 65 27870 100
rect 27830 60 27870 65
rect 28000 100 28040 105
rect 28000 65 28005 100
rect 28005 65 28035 100
rect 28035 65 28040 100
rect 28000 60 28040 65
rect 28170 100 28210 105
rect 28170 65 28175 100
rect 28175 65 28205 100
rect 28205 65 28210 100
rect 28170 60 28210 65
rect 28340 100 28380 105
rect 28340 65 28345 100
rect 28345 65 28375 100
rect 28375 65 28380 100
rect 28340 60 28380 65
rect 28510 100 28550 105
rect 28510 65 28515 100
rect 28515 65 28545 100
rect 28545 65 28550 100
rect 28510 60 28550 65
rect 28680 100 28720 105
rect 28680 65 28685 100
rect 28685 65 28715 100
rect 28715 65 28720 100
rect 28680 60 28720 65
rect 28850 100 28890 105
rect 28850 65 28855 100
rect 28855 65 28885 100
rect 28885 65 28890 100
rect 28850 60 28890 65
rect 29020 100 29060 105
rect 29020 65 29025 100
rect 29025 65 29055 100
rect 29055 65 29060 100
rect 29020 60 29060 65
rect 29190 100 29230 105
rect 29190 65 29195 100
rect 29195 65 29225 100
rect 29225 65 29230 100
rect 29190 60 29230 65
rect 29360 100 29400 105
rect 29360 65 29365 100
rect 29365 65 29395 100
rect 29395 65 29400 100
rect 29360 60 29400 65
rect 29530 100 29570 105
rect 29530 65 29535 100
rect 29535 65 29565 100
rect 29565 65 29570 100
rect 29530 60 29570 65
rect 5335 -185 5385 -135
rect 5490 -190 5540 -140
rect 5845 -185 5895 -135
rect 5995 -190 6045 -140
rect 6335 -190 6385 -140
rect 6525 -185 6575 -135
rect 7210 -190 7260 -140
rect 8055 -190 8105 -140
rect 8190 -185 8240 -135
rect 8735 -185 8785 -135
rect 8870 -185 8920 -135
rect 9245 -185 9295 -135
rect 9380 -190 9430 -140
rect 9925 -190 9975 -140
rect 10060 -185 10110 -135
rect 10605 -185 10655 -135
rect 10740 -185 10790 -135
rect 11115 -185 11165 -135
rect 11250 -190 11300 -140
rect 11795 -185 11845 -135
rect 11930 -190 11980 -140
rect 12265 -190 12315 -140
rect 12475 -185 12525 -135
rect 13160 -190 13210 -140
rect 14005 -190 14055 -140
rect 14140 -185 14190 -135
rect 14685 -185 14735 -135
rect 14820 -185 14870 -135
rect 15195 -185 15245 -135
rect 15330 -190 15380 -140
rect 15875 -190 15925 -140
rect 16010 -185 16060 -135
rect 16555 -185 16605 -135
rect 16690 -185 16740 -135
rect 17065 -185 17115 -135
rect 17200 -190 17250 -140
rect 17745 -185 17795 -135
rect 17880 -190 17930 -140
rect 18215 -190 18265 -140
rect 18425 -185 18475 -135
rect 19110 -190 19160 -140
rect 19955 -190 20005 -140
rect 20635 -185 20685 -135
rect 21145 -185 21195 -135
rect 21280 -190 21330 -140
rect 21825 -190 21875 -135
rect 22300 -190 22350 -140
rect 22505 -185 22555 -135
rect 23190 -190 23240 -140
rect 24035 -190 24085 -140
rect 24170 -185 24220 -135
rect 24715 -185 24765 -135
rect 24850 -185 24900 -135
rect 25225 -185 25275 -135
rect 25360 -190 25410 -140
rect 25905 -190 25955 -140
rect 26040 -185 26090 -135
rect 26585 -185 26635 -135
rect 26720 -185 26770 -135
rect 27095 -185 27145 -135
rect 27605 -185 27655 -135
rect 27740 -190 27790 -140
rect 28285 -185 28335 -135
rect 28970 -190 29020 -140
rect 29815 -190 29865 -140
rect 30495 -185 30545 -135
rect 31005 -185 31055 -135
rect 31685 -190 31735 -140
rect 32365 -185 32415 -135
rect 32875 -185 32925 -135
rect 33555 -185 33605 -135
rect 34235 -185 34285 -135
rect 34920 -190 34970 -140
rect 35765 -190 35815 -140
rect 36445 -185 36495 -135
rect 36955 -185 37005 -135
rect 37635 -190 37685 -140
rect 38315 -185 38365 -135
rect 38825 -185 38875 -135
rect 39505 -185 39555 -135
rect 40185 -185 40235 -135
rect 40870 -190 40920 -140
rect 41715 -190 41765 -140
rect 42395 -185 42445 -135
rect 42905 -185 42955 -135
rect 43585 -190 43635 -140
rect 155 -440 195 -435
rect 155 -475 160 -440
rect 160 -475 190 -440
rect 190 -475 195 -440
rect 155 -480 195 -475
rect 325 -440 365 -435
rect 325 -475 330 -440
rect 330 -475 360 -440
rect 360 -475 365 -440
rect 325 -480 365 -475
rect 495 -440 535 -435
rect 495 -475 500 -440
rect 500 -475 530 -440
rect 530 -475 535 -440
rect 495 -480 535 -475
rect 665 -440 705 -435
rect 665 -475 670 -440
rect 670 -475 700 -440
rect 700 -475 705 -440
rect 665 -480 705 -475
rect 835 -440 875 -435
rect 835 -475 840 -440
rect 840 -475 870 -440
rect 870 -475 875 -440
rect 835 -480 875 -475
rect 1005 -440 1045 -435
rect 1005 -475 1010 -440
rect 1010 -475 1040 -440
rect 1040 -475 1045 -440
rect 1005 -480 1045 -475
rect 1175 -440 1215 -435
rect 1175 -475 1180 -440
rect 1180 -475 1210 -440
rect 1210 -475 1215 -440
rect 1175 -480 1215 -475
rect 1345 -440 1385 -435
rect 1345 -475 1350 -440
rect 1350 -475 1380 -440
rect 1380 -475 1385 -440
rect 1345 -480 1385 -475
rect 1515 -440 1555 -435
rect 1515 -475 1520 -440
rect 1520 -475 1550 -440
rect 1550 -475 1555 -440
rect 1515 -480 1555 -475
rect 1685 -440 1725 -435
rect 1685 -475 1690 -440
rect 1690 -475 1720 -440
rect 1720 -475 1725 -440
rect 1685 -480 1725 -475
rect 1855 -440 1895 -435
rect 1855 -475 1860 -440
rect 1860 -475 1890 -440
rect 1890 -475 1895 -440
rect 1855 -480 1895 -475
rect 2025 -440 2065 -435
rect 2025 -475 2030 -440
rect 2030 -475 2060 -440
rect 2060 -475 2065 -440
rect 2025 -480 2065 -475
rect 2195 -440 2235 -435
rect 2195 -475 2200 -440
rect 2200 -475 2230 -440
rect 2230 -475 2235 -440
rect 2195 -480 2235 -475
rect 2365 -440 2405 -435
rect 2365 -475 2370 -440
rect 2370 -475 2400 -440
rect 2400 -475 2405 -440
rect 2365 -480 2405 -475
rect 2535 -440 2575 -435
rect 2535 -475 2540 -440
rect 2540 -475 2570 -440
rect 2570 -475 2575 -440
rect 2535 -480 2575 -475
rect 2705 -440 2745 -435
rect 2705 -475 2710 -440
rect 2710 -475 2740 -440
rect 2740 -475 2745 -440
rect 2705 -480 2745 -475
rect 2875 -440 2915 -435
rect 2875 -475 2880 -440
rect 2880 -475 2910 -440
rect 2910 -475 2915 -440
rect 2875 -480 2915 -475
rect 3045 -440 3085 -435
rect 3045 -475 3050 -440
rect 3050 -475 3080 -440
rect 3080 -475 3085 -440
rect 3045 -480 3085 -475
rect 3215 -440 3255 -435
rect 3215 -475 3220 -440
rect 3220 -475 3250 -440
rect 3250 -475 3255 -440
rect 3215 -480 3255 -475
rect 3385 -440 3425 -435
rect 3385 -475 3390 -440
rect 3390 -475 3420 -440
rect 3420 -475 3425 -440
rect 3385 -480 3425 -475
rect 3555 -440 3595 -435
rect 3555 -475 3560 -440
rect 3560 -475 3590 -440
rect 3590 -475 3595 -440
rect 3555 -480 3595 -475
rect 3725 -440 3765 -435
rect 3725 -475 3730 -440
rect 3730 -475 3760 -440
rect 3760 -475 3765 -440
rect 3725 -480 3765 -475
rect 3895 -440 3935 -435
rect 3895 -475 3900 -440
rect 3900 -475 3930 -440
rect 3930 -475 3935 -440
rect 3895 -480 3935 -475
rect 4065 -440 4105 -435
rect 4065 -475 4070 -440
rect 4070 -475 4100 -440
rect 4100 -475 4105 -440
rect 4065 -480 4105 -475
rect 4235 -440 4275 -435
rect 4235 -475 4240 -440
rect 4240 -475 4270 -440
rect 4270 -475 4275 -440
rect 4235 -480 4275 -475
rect 4405 -440 4445 -435
rect 4405 -475 4410 -440
rect 4410 -475 4440 -440
rect 4440 -475 4445 -440
rect 4405 -480 4445 -475
rect 4575 -440 4615 -435
rect 4575 -475 4580 -440
rect 4580 -475 4610 -440
rect 4610 -475 4615 -440
rect 4575 -480 4615 -475
rect 4745 -440 4785 -435
rect 4745 -475 4750 -440
rect 4750 -475 4780 -440
rect 4780 -475 4785 -440
rect 4745 -480 4785 -475
rect 4915 -440 4955 -435
rect 4915 -475 4920 -440
rect 4920 -475 4950 -440
rect 4950 -475 4955 -440
rect 4915 -480 4955 -475
rect 5085 -440 5125 -435
rect 5085 -475 5090 -440
rect 5090 -475 5120 -440
rect 5120 -475 5125 -440
rect 5085 -480 5125 -475
rect 5255 -440 5295 -435
rect 5255 -475 5260 -440
rect 5260 -475 5290 -440
rect 5290 -475 5295 -440
rect 5255 -480 5295 -475
rect 5425 -440 5465 -435
rect 5425 -475 5430 -440
rect 5430 -475 5460 -440
rect 5460 -475 5465 -440
rect 5425 -480 5465 -475
rect 5595 -440 5635 -435
rect 5595 -475 5600 -440
rect 5600 -475 5630 -440
rect 5630 -475 5635 -440
rect 5595 -480 5635 -475
rect 5765 -440 5805 -435
rect 5765 -475 5770 -440
rect 5770 -475 5800 -440
rect 5800 -475 5805 -440
rect 5765 -480 5805 -475
rect 5935 -440 5975 -435
rect 5935 -475 5940 -440
rect 5940 -475 5970 -440
rect 5970 -475 5975 -440
rect 5935 -480 5975 -475
rect 6105 -440 6145 -435
rect 6105 -475 6110 -440
rect 6110 -475 6140 -440
rect 6140 -475 6145 -440
rect 6105 -480 6145 -475
rect 6275 -440 6315 -435
rect 6275 -475 6280 -440
rect 6280 -475 6310 -440
rect 6310 -475 6315 -440
rect 6275 -480 6315 -475
rect 6445 -440 6485 -435
rect 6445 -475 6450 -440
rect 6450 -475 6480 -440
rect 6480 -475 6485 -440
rect 6445 -480 6485 -475
rect 6615 -440 6655 -435
rect 6615 -475 6620 -440
rect 6620 -475 6650 -440
rect 6650 -475 6655 -440
rect 6615 -480 6655 -475
rect 6785 -440 6825 -435
rect 6785 -475 6790 -440
rect 6790 -475 6820 -440
rect 6820 -475 6825 -440
rect 6785 -480 6825 -475
rect 6955 -440 6995 -435
rect 6955 -475 6960 -440
rect 6960 -475 6990 -440
rect 6990 -475 6995 -440
rect 6955 -480 6995 -475
rect 7125 -440 7165 -435
rect 7125 -475 7130 -440
rect 7130 -475 7160 -440
rect 7160 -475 7165 -440
rect 7125 -480 7165 -475
rect 7295 -440 7335 -435
rect 7295 -475 7300 -440
rect 7300 -475 7330 -440
rect 7330 -475 7335 -440
rect 7295 -480 7335 -475
rect 7465 -440 7505 -435
rect 7465 -475 7470 -440
rect 7470 -475 7500 -440
rect 7500 -475 7505 -440
rect 7465 -480 7505 -475
rect 7635 -440 7675 -435
rect 7635 -475 7640 -440
rect 7640 -475 7670 -440
rect 7670 -475 7675 -440
rect 7635 -480 7675 -475
rect 7805 -440 7845 -435
rect 7805 -475 7810 -440
rect 7810 -475 7840 -440
rect 7840 -475 7845 -440
rect 7805 -480 7845 -475
rect 7975 -440 8015 -435
rect 7975 -475 7980 -440
rect 7980 -475 8010 -440
rect 8010 -475 8015 -440
rect 7975 -480 8015 -475
rect 8145 -440 8185 -435
rect 8145 -475 8150 -440
rect 8150 -475 8180 -440
rect 8180 -475 8185 -440
rect 8145 -480 8185 -475
rect 8315 -440 8355 -435
rect 8315 -475 8320 -440
rect 8320 -475 8350 -440
rect 8350 -475 8355 -440
rect 8315 -480 8355 -475
rect 8485 -440 8525 -435
rect 8485 -475 8490 -440
rect 8490 -475 8520 -440
rect 8520 -475 8525 -440
rect 8485 -480 8525 -475
rect 8655 -440 8695 -435
rect 8655 -475 8660 -440
rect 8660 -475 8690 -440
rect 8690 -475 8695 -440
rect 8655 -480 8695 -475
rect 8825 -440 8865 -435
rect 8825 -475 8830 -440
rect 8830 -475 8860 -440
rect 8860 -475 8865 -440
rect 8825 -480 8865 -475
rect 8995 -440 9035 -435
rect 8995 -475 9000 -440
rect 9000 -475 9030 -440
rect 9030 -475 9035 -440
rect 8995 -480 9035 -475
rect 9165 -440 9205 -435
rect 9165 -475 9170 -440
rect 9170 -475 9200 -440
rect 9200 -475 9205 -440
rect 9165 -480 9205 -475
rect 9335 -440 9375 -435
rect 9335 -475 9340 -440
rect 9340 -475 9370 -440
rect 9370 -475 9375 -440
rect 9335 -480 9375 -475
rect 9505 -440 9545 -435
rect 9505 -475 9510 -440
rect 9510 -475 9540 -440
rect 9540 -475 9545 -440
rect 9505 -480 9545 -475
rect 9675 -440 9715 -435
rect 9675 -475 9680 -440
rect 9680 -475 9710 -440
rect 9710 -475 9715 -440
rect 9675 -480 9715 -475
rect 9845 -440 9885 -435
rect 9845 -475 9850 -440
rect 9850 -475 9880 -440
rect 9880 -475 9885 -440
rect 9845 -480 9885 -475
rect 10015 -440 10055 -435
rect 10015 -475 10020 -440
rect 10020 -475 10050 -440
rect 10050 -475 10055 -440
rect 10015 -480 10055 -475
rect 10185 -440 10225 -435
rect 10185 -475 10190 -440
rect 10190 -475 10220 -440
rect 10220 -475 10225 -440
rect 10185 -480 10225 -475
rect 10355 -440 10395 -435
rect 10355 -475 10360 -440
rect 10360 -475 10390 -440
rect 10390 -475 10395 -440
rect 10355 -480 10395 -475
rect 10525 -440 10565 -435
rect 10525 -475 10530 -440
rect 10530 -475 10560 -440
rect 10560 -475 10565 -440
rect 10525 -480 10565 -475
rect 10695 -440 10735 -435
rect 10695 -475 10700 -440
rect 10700 -475 10730 -440
rect 10730 -475 10735 -440
rect 10695 -480 10735 -475
rect 10865 -440 10905 -435
rect 10865 -475 10870 -440
rect 10870 -475 10900 -440
rect 10900 -475 10905 -440
rect 10865 -480 10905 -475
rect 11035 -440 11075 -435
rect 11035 -475 11040 -440
rect 11040 -475 11070 -440
rect 11070 -475 11075 -440
rect 11035 -480 11075 -475
rect 11205 -440 11245 -435
rect 11205 -475 11210 -440
rect 11210 -475 11240 -440
rect 11240 -475 11245 -440
rect 11205 -480 11245 -475
rect 11375 -440 11415 -435
rect 11375 -475 11380 -440
rect 11380 -475 11410 -440
rect 11410 -475 11415 -440
rect 11375 -480 11415 -475
rect 11545 -440 11585 -435
rect 11545 -475 11550 -440
rect 11550 -475 11580 -440
rect 11580 -475 11585 -440
rect 11545 -480 11585 -475
rect 11715 -440 11755 -435
rect 11715 -475 11720 -440
rect 11720 -475 11750 -440
rect 11750 -475 11755 -440
rect 11715 -480 11755 -475
rect 11885 -440 11925 -435
rect 11885 -475 11890 -440
rect 11890 -475 11920 -440
rect 11920 -475 11925 -440
rect 11885 -480 11925 -475
rect 12055 -440 12095 -435
rect 12055 -475 12060 -440
rect 12060 -475 12090 -440
rect 12090 -475 12095 -440
rect 12055 -480 12095 -475
rect 12225 -440 12265 -435
rect 12225 -475 12230 -440
rect 12230 -475 12260 -440
rect 12260 -475 12265 -440
rect 12225 -480 12265 -475
rect 12395 -440 12435 -435
rect 12395 -475 12400 -440
rect 12400 -475 12430 -440
rect 12430 -475 12435 -440
rect 12395 -480 12435 -475
rect 12565 -440 12605 -435
rect 12565 -475 12570 -440
rect 12570 -475 12600 -440
rect 12600 -475 12605 -440
rect 12565 -480 12605 -475
rect 12735 -440 12775 -435
rect 12735 -475 12740 -440
rect 12740 -475 12770 -440
rect 12770 -475 12775 -440
rect 12735 -480 12775 -475
rect 12905 -440 12945 -435
rect 12905 -475 12910 -440
rect 12910 -475 12940 -440
rect 12940 -475 12945 -440
rect 12905 -480 12945 -475
rect 13075 -440 13115 -435
rect 13075 -475 13080 -440
rect 13080 -475 13110 -440
rect 13110 -475 13115 -440
rect 13075 -480 13115 -475
rect 13245 -440 13285 -435
rect 13245 -475 13250 -440
rect 13250 -475 13280 -440
rect 13280 -475 13285 -440
rect 13245 -480 13285 -475
rect 13415 -440 13455 -435
rect 13415 -475 13420 -440
rect 13420 -475 13450 -440
rect 13450 -475 13455 -440
rect 13415 -480 13455 -475
rect 13585 -440 13625 -435
rect 13585 -475 13590 -440
rect 13590 -475 13620 -440
rect 13620 -475 13625 -440
rect 13585 -480 13625 -475
rect 13755 -440 13795 -435
rect 13755 -475 13760 -440
rect 13760 -475 13790 -440
rect 13790 -475 13795 -440
rect 13755 -480 13795 -475
rect 13925 -440 13965 -435
rect 13925 -475 13930 -440
rect 13930 -475 13960 -440
rect 13960 -475 13965 -440
rect 13925 -480 13965 -475
rect 14095 -440 14135 -435
rect 14095 -475 14100 -440
rect 14100 -475 14130 -440
rect 14130 -475 14135 -440
rect 14095 -480 14135 -475
rect 14265 -440 14305 -435
rect 14265 -475 14270 -440
rect 14270 -475 14300 -440
rect 14300 -475 14305 -440
rect 14265 -480 14305 -475
rect 14435 -440 14475 -435
rect 14435 -475 14440 -440
rect 14440 -475 14470 -440
rect 14470 -475 14475 -440
rect 14435 -480 14475 -475
rect 14605 -440 14645 -435
rect 14605 -475 14610 -440
rect 14610 -475 14640 -440
rect 14640 -475 14645 -440
rect 14605 -480 14645 -475
rect 14775 -440 14815 -435
rect 14775 -475 14780 -440
rect 14780 -475 14810 -440
rect 14810 -475 14815 -440
rect 14775 -480 14815 -475
rect 14945 -440 14985 -435
rect 14945 -475 14950 -440
rect 14950 -475 14980 -440
rect 14980 -475 14985 -440
rect 14945 -480 14985 -475
rect 15115 -440 15155 -435
rect 15115 -475 15120 -440
rect 15120 -475 15150 -440
rect 15150 -475 15155 -440
rect 15115 -480 15155 -475
rect 15285 -440 15325 -435
rect 15285 -475 15290 -440
rect 15290 -475 15320 -440
rect 15320 -475 15325 -440
rect 15285 -480 15325 -475
rect 15455 -440 15495 -435
rect 15455 -475 15460 -440
rect 15460 -475 15490 -440
rect 15490 -475 15495 -440
rect 15455 -480 15495 -475
rect 15625 -440 15665 -435
rect 15625 -475 15630 -440
rect 15630 -475 15660 -440
rect 15660 -475 15665 -440
rect 15625 -480 15665 -475
rect 15795 -440 15835 -435
rect 15795 -475 15800 -440
rect 15800 -475 15830 -440
rect 15830 -475 15835 -440
rect 15795 -480 15835 -475
rect 15965 -440 16005 -435
rect 15965 -475 15970 -440
rect 15970 -475 16000 -440
rect 16000 -475 16005 -440
rect 15965 -480 16005 -475
rect 16135 -440 16175 -435
rect 16135 -475 16140 -440
rect 16140 -475 16170 -440
rect 16170 -475 16175 -440
rect 16135 -480 16175 -475
rect 16305 -440 16345 -435
rect 16305 -475 16310 -440
rect 16310 -475 16340 -440
rect 16340 -475 16345 -440
rect 16305 -480 16345 -475
rect 16475 -440 16515 -435
rect 16475 -475 16480 -440
rect 16480 -475 16510 -440
rect 16510 -475 16515 -440
rect 16475 -480 16515 -475
rect 16645 -440 16685 -435
rect 16645 -475 16650 -440
rect 16650 -475 16680 -440
rect 16680 -475 16685 -440
rect 16645 -480 16685 -475
rect 16815 -440 16855 -435
rect 16815 -475 16820 -440
rect 16820 -475 16850 -440
rect 16850 -475 16855 -440
rect 16815 -480 16855 -475
rect 16985 -440 17025 -435
rect 16985 -475 16990 -440
rect 16990 -475 17020 -440
rect 17020 -475 17025 -440
rect 16985 -480 17025 -475
rect 17155 -440 17195 -435
rect 17155 -475 17160 -440
rect 17160 -475 17190 -440
rect 17190 -475 17195 -440
rect 17155 -480 17195 -475
rect 17325 -440 17365 -435
rect 17325 -475 17330 -440
rect 17330 -475 17360 -440
rect 17360 -475 17365 -440
rect 17325 -480 17365 -475
rect 17495 -440 17535 -435
rect 17495 -475 17500 -440
rect 17500 -475 17530 -440
rect 17530 -475 17535 -440
rect 17495 -480 17535 -475
rect 17665 -440 17705 -435
rect 17665 -475 17670 -440
rect 17670 -475 17700 -440
rect 17700 -475 17705 -440
rect 17665 -480 17705 -475
rect 17835 -440 17875 -435
rect 17835 -475 17840 -440
rect 17840 -475 17870 -440
rect 17870 -475 17875 -440
rect 17835 -480 17875 -475
rect 18005 -440 18045 -435
rect 18005 -475 18010 -440
rect 18010 -475 18040 -440
rect 18040 -475 18045 -440
rect 18005 -480 18045 -475
rect 18175 -440 18215 -435
rect 18175 -475 18180 -440
rect 18180 -475 18210 -440
rect 18210 -475 18215 -440
rect 18175 -480 18215 -475
rect 18345 -440 18385 -435
rect 18345 -475 18350 -440
rect 18350 -475 18380 -440
rect 18380 -475 18385 -440
rect 18345 -480 18385 -475
rect 18515 -440 18555 -435
rect 18515 -475 18520 -440
rect 18520 -475 18550 -440
rect 18550 -475 18555 -440
rect 18515 -480 18555 -475
rect 18685 -440 18725 -435
rect 18685 -475 18690 -440
rect 18690 -475 18720 -440
rect 18720 -475 18725 -440
rect 18685 -480 18725 -475
rect 18855 -440 18895 -435
rect 18855 -475 18860 -440
rect 18860 -475 18890 -440
rect 18890 -475 18895 -440
rect 18855 -480 18895 -475
rect 19025 -440 19065 -435
rect 19025 -475 19030 -440
rect 19030 -475 19060 -440
rect 19060 -475 19065 -440
rect 19025 -480 19065 -475
rect 19195 -440 19235 -435
rect 19195 -475 19200 -440
rect 19200 -475 19230 -440
rect 19230 -475 19235 -440
rect 19195 -480 19235 -475
rect 19365 -440 19405 -435
rect 19365 -475 19370 -440
rect 19370 -475 19400 -440
rect 19400 -475 19405 -440
rect 19365 -480 19405 -475
rect 19535 -440 19575 -435
rect 19535 -475 19540 -440
rect 19540 -475 19570 -440
rect 19570 -475 19575 -440
rect 19535 -480 19575 -475
rect 19705 -440 19745 -435
rect 19705 -475 19710 -440
rect 19710 -475 19740 -440
rect 19740 -475 19745 -440
rect 19705 -480 19745 -475
rect 19875 -440 19915 -435
rect 19875 -475 19880 -440
rect 19880 -475 19910 -440
rect 19910 -475 19915 -440
rect 19875 -480 19915 -475
rect 20045 -440 20085 -435
rect 20045 -475 20050 -440
rect 20050 -475 20080 -440
rect 20080 -475 20085 -440
rect 20045 -480 20085 -475
rect 20215 -440 20255 -435
rect 20215 -475 20220 -440
rect 20220 -475 20250 -440
rect 20250 -475 20255 -440
rect 20215 -480 20255 -475
rect 20385 -440 20425 -435
rect 20385 -475 20390 -440
rect 20390 -475 20420 -440
rect 20420 -475 20425 -440
rect 20385 -480 20425 -475
rect 20555 -440 20595 -435
rect 20555 -475 20560 -440
rect 20560 -475 20590 -440
rect 20590 -475 20595 -440
rect 20555 -480 20595 -475
rect 20725 -440 20765 -435
rect 20725 -475 20730 -440
rect 20730 -475 20760 -440
rect 20760 -475 20765 -440
rect 20725 -480 20765 -475
rect 20895 -440 20935 -435
rect 20895 -475 20900 -440
rect 20900 -475 20930 -440
rect 20930 -475 20935 -440
rect 20895 -480 20935 -475
rect 21065 -440 21105 -435
rect 21065 -475 21070 -440
rect 21070 -475 21100 -440
rect 21100 -475 21105 -440
rect 21065 -480 21105 -475
rect 21235 -440 21275 -435
rect 21235 -475 21240 -440
rect 21240 -475 21270 -440
rect 21270 -475 21275 -440
rect 21235 -480 21275 -475
rect 21405 -440 21445 -435
rect 21405 -475 21410 -440
rect 21410 -475 21440 -440
rect 21440 -475 21445 -440
rect 21405 -480 21445 -475
rect 21575 -440 21615 -435
rect 21575 -475 21580 -440
rect 21580 -475 21610 -440
rect 21610 -475 21615 -440
rect 21575 -480 21615 -475
rect 21745 -440 21785 -435
rect 21745 -475 21750 -440
rect 21750 -475 21780 -440
rect 21780 -475 21785 -440
rect 21745 -480 21785 -475
rect 21915 -440 21955 -435
rect 21915 -475 21920 -440
rect 21920 -475 21950 -440
rect 21950 -475 21955 -440
rect 21915 -480 21955 -475
rect 22085 -440 22125 -435
rect 22085 -475 22090 -440
rect 22090 -475 22120 -440
rect 22120 -475 22125 -440
rect 22085 -480 22125 -475
rect 22255 -440 22295 -435
rect 22255 -475 22260 -440
rect 22260 -475 22290 -440
rect 22290 -475 22295 -440
rect 22255 -480 22295 -475
rect 22425 -440 22465 -435
rect 22425 -475 22430 -440
rect 22430 -475 22460 -440
rect 22460 -475 22465 -440
rect 22425 -480 22465 -475
rect 22595 -440 22635 -435
rect 22595 -475 22600 -440
rect 22600 -475 22630 -440
rect 22630 -475 22635 -440
rect 22595 -480 22635 -475
rect 22765 -440 22805 -435
rect 22765 -475 22770 -440
rect 22770 -475 22800 -440
rect 22800 -475 22805 -440
rect 22765 -480 22805 -475
rect 22935 -440 22975 -435
rect 22935 -475 22940 -440
rect 22940 -475 22970 -440
rect 22970 -475 22975 -440
rect 22935 -480 22975 -475
rect 23105 -440 23145 -435
rect 23105 -475 23110 -440
rect 23110 -475 23140 -440
rect 23140 -475 23145 -440
rect 23105 -480 23145 -475
rect 23275 -440 23315 -435
rect 23275 -475 23280 -440
rect 23280 -475 23310 -440
rect 23310 -475 23315 -440
rect 23275 -480 23315 -475
rect 23445 -440 23485 -435
rect 23445 -475 23450 -440
rect 23450 -475 23480 -440
rect 23480 -475 23485 -440
rect 23445 -480 23485 -475
rect 23615 -440 23655 -435
rect 23615 -475 23620 -440
rect 23620 -475 23650 -440
rect 23650 -475 23655 -440
rect 23615 -480 23655 -475
rect 23785 -440 23825 -435
rect 23785 -475 23790 -440
rect 23790 -475 23820 -440
rect 23820 -475 23825 -440
rect 23785 -480 23825 -475
rect 23955 -440 23995 -435
rect 23955 -475 23960 -440
rect 23960 -475 23990 -440
rect 23990 -475 23995 -440
rect 23955 -480 23995 -475
rect 24125 -440 24165 -435
rect 24125 -475 24130 -440
rect 24130 -475 24160 -440
rect 24160 -475 24165 -440
rect 24125 -480 24165 -475
rect 24295 -440 24335 -435
rect 24295 -475 24300 -440
rect 24300 -475 24330 -440
rect 24330 -475 24335 -440
rect 24295 -480 24335 -475
rect 24465 -440 24505 -435
rect 24465 -475 24470 -440
rect 24470 -475 24500 -440
rect 24500 -475 24505 -440
rect 24465 -480 24505 -475
rect 24635 -440 24675 -435
rect 24635 -475 24640 -440
rect 24640 -475 24670 -440
rect 24670 -475 24675 -440
rect 24635 -480 24675 -475
rect 24805 -440 24845 -435
rect 24805 -475 24810 -440
rect 24810 -475 24840 -440
rect 24840 -475 24845 -440
rect 24805 -480 24845 -475
rect 24975 -440 25015 -435
rect 24975 -475 24980 -440
rect 24980 -475 25010 -440
rect 25010 -475 25015 -440
rect 24975 -480 25015 -475
rect 25145 -440 25185 -435
rect 25145 -475 25150 -440
rect 25150 -475 25180 -440
rect 25180 -475 25185 -440
rect 25145 -480 25185 -475
rect 25315 -440 25355 -435
rect 25315 -475 25320 -440
rect 25320 -475 25350 -440
rect 25350 -475 25355 -440
rect 25315 -480 25355 -475
rect 25485 -440 25525 -435
rect 25485 -475 25490 -440
rect 25490 -475 25520 -440
rect 25520 -475 25525 -440
rect 25485 -480 25525 -475
rect 25655 -440 25695 -435
rect 25655 -475 25660 -440
rect 25660 -475 25690 -440
rect 25690 -475 25695 -440
rect 25655 -480 25695 -475
rect 25825 -440 25865 -435
rect 25825 -475 25830 -440
rect 25830 -475 25860 -440
rect 25860 -475 25865 -440
rect 25825 -480 25865 -475
rect 25995 -440 26035 -435
rect 25995 -475 26000 -440
rect 26000 -475 26030 -440
rect 26030 -475 26035 -440
rect 25995 -480 26035 -475
rect 26165 -440 26205 -435
rect 26165 -475 26170 -440
rect 26170 -475 26200 -440
rect 26200 -475 26205 -440
rect 26165 -480 26205 -475
rect 26335 -440 26375 -435
rect 26335 -475 26340 -440
rect 26340 -475 26370 -440
rect 26370 -475 26375 -440
rect 26335 -480 26375 -475
rect 26505 -440 26545 -435
rect 26505 -475 26510 -440
rect 26510 -475 26540 -440
rect 26540 -475 26545 -440
rect 26505 -480 26545 -475
rect 26675 -440 26715 -435
rect 26675 -475 26680 -440
rect 26680 -475 26710 -440
rect 26710 -475 26715 -440
rect 26675 -480 26715 -475
rect 26845 -440 26885 -435
rect 26845 -475 26850 -440
rect 26850 -475 26880 -440
rect 26880 -475 26885 -440
rect 26845 -480 26885 -475
rect 27015 -440 27055 -435
rect 27015 -475 27020 -440
rect 27020 -475 27050 -440
rect 27050 -475 27055 -440
rect 27015 -480 27055 -475
rect 27185 -440 27225 -435
rect 27185 -475 27190 -440
rect 27190 -475 27220 -440
rect 27220 -475 27225 -440
rect 27185 -480 27225 -475
rect 27355 -440 27395 -435
rect 27355 -475 27360 -440
rect 27360 -475 27390 -440
rect 27390 -475 27395 -440
rect 27355 -480 27395 -475
rect 27525 -440 27565 -435
rect 27525 -475 27530 -440
rect 27530 -475 27560 -440
rect 27560 -475 27565 -440
rect 27525 -480 27565 -475
rect 27695 -440 27735 -435
rect 27695 -475 27700 -440
rect 27700 -475 27730 -440
rect 27730 -475 27735 -440
rect 27695 -480 27735 -475
rect 27865 -440 27905 -435
rect 27865 -475 27870 -440
rect 27870 -475 27900 -440
rect 27900 -475 27905 -440
rect 27865 -480 27905 -475
rect 28035 -440 28075 -435
rect 28035 -475 28040 -440
rect 28040 -475 28070 -440
rect 28070 -475 28075 -440
rect 28035 -480 28075 -475
rect 28205 -440 28245 -435
rect 28205 -475 28210 -440
rect 28210 -475 28240 -440
rect 28240 -475 28245 -440
rect 28205 -480 28245 -475
rect 28375 -440 28415 -435
rect 28375 -475 28380 -440
rect 28380 -475 28410 -440
rect 28410 -475 28415 -440
rect 28375 -480 28415 -475
rect 28545 -440 28585 -435
rect 28545 -475 28550 -440
rect 28550 -475 28580 -440
rect 28580 -475 28585 -440
rect 28545 -480 28585 -475
rect 28715 -440 28755 -435
rect 28715 -475 28720 -440
rect 28720 -475 28750 -440
rect 28750 -475 28755 -440
rect 28715 -480 28755 -475
rect 28885 -440 28925 -435
rect 28885 -475 28890 -440
rect 28890 -475 28920 -440
rect 28920 -475 28925 -440
rect 28885 -480 28925 -475
rect 29055 -440 29095 -435
rect 29055 -475 29060 -440
rect 29060 -475 29090 -440
rect 29090 -475 29095 -440
rect 29055 -480 29095 -475
rect 29225 -440 29265 -435
rect 29225 -475 29230 -440
rect 29230 -475 29260 -440
rect 29260 -475 29265 -440
rect 29225 -480 29265 -475
rect 29395 -440 29435 -435
rect 29395 -475 29400 -440
rect 29400 -475 29430 -440
rect 29430 -475 29435 -440
rect 29395 -480 29435 -475
rect 29565 -440 29605 -435
rect 29565 -475 29570 -440
rect 29570 -475 29600 -440
rect 29600 -475 29605 -440
rect 29565 -480 29605 -475
rect 29735 -440 29775 -435
rect 29735 -475 29740 -440
rect 29740 -475 29770 -440
rect 29770 -475 29775 -440
rect 29735 -480 29775 -475
rect 29905 -440 29945 -435
rect 29905 -475 29910 -440
rect 29910 -475 29940 -440
rect 29940 -475 29945 -440
rect 29905 -480 29945 -475
rect 30075 -440 30115 -435
rect 30075 -475 30080 -440
rect 30080 -475 30110 -440
rect 30110 -475 30115 -440
rect 30075 -480 30115 -475
rect 30245 -440 30285 -435
rect 30245 -475 30250 -440
rect 30250 -475 30280 -440
rect 30280 -475 30285 -440
rect 30245 -480 30285 -475
rect 30415 -440 30455 -435
rect 30415 -475 30420 -440
rect 30420 -475 30450 -440
rect 30450 -475 30455 -440
rect 30415 -480 30455 -475
rect 30585 -440 30625 -435
rect 30585 -475 30590 -440
rect 30590 -475 30620 -440
rect 30620 -475 30625 -440
rect 30585 -480 30625 -475
rect 30755 -440 30795 -435
rect 30755 -475 30760 -440
rect 30760 -475 30790 -440
rect 30790 -475 30795 -440
rect 30755 -480 30795 -475
rect 30925 -440 30965 -435
rect 30925 -475 30930 -440
rect 30930 -475 30960 -440
rect 30960 -475 30965 -440
rect 30925 -480 30965 -475
rect 31095 -440 31135 -435
rect 31095 -475 31100 -440
rect 31100 -475 31130 -440
rect 31130 -475 31135 -440
rect 31095 -480 31135 -475
rect 31265 -440 31305 -435
rect 31265 -475 31270 -440
rect 31270 -475 31300 -440
rect 31300 -475 31305 -440
rect 31265 -480 31305 -475
rect 31435 -440 31475 -435
rect 31435 -475 31440 -440
rect 31440 -475 31470 -440
rect 31470 -475 31475 -440
rect 31435 -480 31475 -475
rect 31605 -440 31645 -435
rect 31605 -475 31610 -440
rect 31610 -475 31640 -440
rect 31640 -475 31645 -440
rect 31605 -480 31645 -475
rect 31775 -440 31815 -435
rect 31775 -475 31780 -440
rect 31780 -475 31810 -440
rect 31810 -475 31815 -440
rect 31775 -480 31815 -475
rect 31945 -440 31985 -435
rect 31945 -475 31950 -440
rect 31950 -475 31980 -440
rect 31980 -475 31985 -440
rect 31945 -480 31985 -475
rect 32115 -440 32155 -435
rect 32115 -475 32120 -440
rect 32120 -475 32150 -440
rect 32150 -475 32155 -440
rect 32115 -480 32155 -475
rect 32285 -440 32325 -435
rect 32285 -475 32290 -440
rect 32290 -475 32320 -440
rect 32320 -475 32325 -440
rect 32285 -480 32325 -475
rect 32455 -440 32495 -435
rect 32455 -475 32460 -440
rect 32460 -475 32490 -440
rect 32490 -475 32495 -440
rect 32455 -480 32495 -475
rect 32625 -440 32665 -435
rect 32625 -475 32630 -440
rect 32630 -475 32660 -440
rect 32660 -475 32665 -440
rect 32625 -480 32665 -475
rect 32795 -440 32835 -435
rect 32795 -475 32800 -440
rect 32800 -475 32830 -440
rect 32830 -475 32835 -440
rect 32795 -480 32835 -475
rect 32965 -440 33005 -435
rect 32965 -475 32970 -440
rect 32970 -475 33000 -440
rect 33000 -475 33005 -440
rect 32965 -480 33005 -475
rect 33135 -440 33175 -435
rect 33135 -475 33140 -440
rect 33140 -475 33170 -440
rect 33170 -475 33175 -440
rect 33135 -480 33175 -475
rect 33305 -440 33345 -435
rect 33305 -475 33310 -440
rect 33310 -475 33340 -440
rect 33340 -475 33345 -440
rect 33305 -480 33345 -475
rect 33475 -440 33515 -435
rect 33475 -475 33480 -440
rect 33480 -475 33510 -440
rect 33510 -475 33515 -440
rect 33475 -480 33515 -475
rect 33645 -440 33685 -435
rect 33645 -475 33650 -440
rect 33650 -475 33680 -440
rect 33680 -475 33685 -440
rect 33645 -480 33685 -475
rect 33815 -440 33855 -435
rect 33815 -475 33820 -440
rect 33820 -475 33850 -440
rect 33850 -475 33855 -440
rect 33815 -480 33855 -475
rect 33985 -440 34025 -435
rect 33985 -475 33990 -440
rect 33990 -475 34020 -440
rect 34020 -475 34025 -440
rect 33985 -480 34025 -475
rect 34155 -440 34195 -435
rect 34155 -475 34160 -440
rect 34160 -475 34190 -440
rect 34190 -475 34195 -440
rect 34155 -480 34195 -475
rect 34325 -440 34365 -435
rect 34325 -475 34330 -440
rect 34330 -475 34360 -440
rect 34360 -475 34365 -440
rect 34325 -480 34365 -475
rect 34495 -440 34535 -435
rect 34495 -475 34500 -440
rect 34500 -475 34530 -440
rect 34530 -475 34535 -440
rect 34495 -480 34535 -475
rect 34665 -440 34705 -435
rect 34665 -475 34670 -440
rect 34670 -475 34700 -440
rect 34700 -475 34705 -440
rect 34665 -480 34705 -475
rect 34835 -440 34875 -435
rect 34835 -475 34840 -440
rect 34840 -475 34870 -440
rect 34870 -475 34875 -440
rect 34835 -480 34875 -475
rect 35005 -440 35045 -435
rect 35005 -475 35010 -440
rect 35010 -475 35040 -440
rect 35040 -475 35045 -440
rect 35005 -480 35045 -475
rect 35175 -440 35215 -435
rect 35175 -475 35180 -440
rect 35180 -475 35210 -440
rect 35210 -475 35215 -440
rect 35175 -480 35215 -475
rect 35345 -440 35385 -435
rect 35345 -475 35350 -440
rect 35350 -475 35380 -440
rect 35380 -475 35385 -440
rect 35345 -480 35385 -475
rect 35515 -440 35555 -435
rect 35515 -475 35520 -440
rect 35520 -475 35550 -440
rect 35550 -475 35555 -440
rect 35515 -480 35555 -475
rect 35685 -440 35725 -435
rect 35685 -475 35690 -440
rect 35690 -475 35720 -440
rect 35720 -475 35725 -440
rect 35685 -480 35725 -475
rect 35855 -440 35895 -435
rect 35855 -475 35860 -440
rect 35860 -475 35890 -440
rect 35890 -475 35895 -440
rect 35855 -480 35895 -475
rect 36025 -440 36065 -435
rect 36025 -475 36030 -440
rect 36030 -475 36060 -440
rect 36060 -475 36065 -440
rect 36025 -480 36065 -475
rect 36195 -440 36235 -435
rect 36195 -475 36200 -440
rect 36200 -475 36230 -440
rect 36230 -475 36235 -440
rect 36195 -480 36235 -475
rect 36365 -440 36405 -435
rect 36365 -475 36370 -440
rect 36370 -475 36400 -440
rect 36400 -475 36405 -440
rect 36365 -480 36405 -475
rect 36535 -440 36575 -435
rect 36535 -475 36540 -440
rect 36540 -475 36570 -440
rect 36570 -475 36575 -440
rect 36535 -480 36575 -475
rect 36705 -440 36745 -435
rect 36705 -475 36710 -440
rect 36710 -475 36740 -440
rect 36740 -475 36745 -440
rect 36705 -480 36745 -475
rect 36875 -440 36915 -435
rect 36875 -475 36880 -440
rect 36880 -475 36910 -440
rect 36910 -475 36915 -440
rect 36875 -480 36915 -475
rect 37045 -440 37085 -435
rect 37045 -475 37050 -440
rect 37050 -475 37080 -440
rect 37080 -475 37085 -440
rect 37045 -480 37085 -475
rect 37215 -440 37255 -435
rect 37215 -475 37220 -440
rect 37220 -475 37250 -440
rect 37250 -475 37255 -440
rect 37215 -480 37255 -475
rect 37385 -440 37425 -435
rect 37385 -475 37390 -440
rect 37390 -475 37420 -440
rect 37420 -475 37425 -440
rect 37385 -480 37425 -475
rect 37555 -440 37595 -435
rect 37555 -475 37560 -440
rect 37560 -475 37590 -440
rect 37590 -475 37595 -440
rect 37555 -480 37595 -475
rect 37725 -440 37765 -435
rect 37725 -475 37730 -440
rect 37730 -475 37760 -440
rect 37760 -475 37765 -440
rect 37725 -480 37765 -475
rect 37895 -440 37935 -435
rect 37895 -475 37900 -440
rect 37900 -475 37930 -440
rect 37930 -475 37935 -440
rect 37895 -480 37935 -475
rect 38065 -440 38105 -435
rect 38065 -475 38070 -440
rect 38070 -475 38100 -440
rect 38100 -475 38105 -440
rect 38065 -480 38105 -475
rect 38235 -440 38275 -435
rect 38235 -475 38240 -440
rect 38240 -475 38270 -440
rect 38270 -475 38275 -440
rect 38235 -480 38275 -475
rect 38405 -440 38445 -435
rect 38405 -475 38410 -440
rect 38410 -475 38440 -440
rect 38440 -475 38445 -440
rect 38405 -480 38445 -475
rect 38575 -440 38615 -435
rect 38575 -475 38580 -440
rect 38580 -475 38610 -440
rect 38610 -475 38615 -440
rect 38575 -480 38615 -475
rect 38745 -440 38785 -435
rect 38745 -475 38750 -440
rect 38750 -475 38780 -440
rect 38780 -475 38785 -440
rect 38745 -480 38785 -475
rect 38915 -440 38955 -435
rect 38915 -475 38920 -440
rect 38920 -475 38950 -440
rect 38950 -475 38955 -440
rect 38915 -480 38955 -475
rect 39085 -440 39125 -435
rect 39085 -475 39090 -440
rect 39090 -475 39120 -440
rect 39120 -475 39125 -440
rect 39085 -480 39125 -475
rect 39255 -440 39295 -435
rect 39255 -475 39260 -440
rect 39260 -475 39290 -440
rect 39290 -475 39295 -440
rect 39255 -480 39295 -475
rect 39425 -440 39465 -435
rect 39425 -475 39430 -440
rect 39430 -475 39460 -440
rect 39460 -475 39465 -440
rect 39425 -480 39465 -475
rect 39595 -440 39635 -435
rect 39595 -475 39600 -440
rect 39600 -475 39630 -440
rect 39630 -475 39635 -440
rect 39595 -480 39635 -475
rect 39765 -440 39805 -435
rect 39765 -475 39770 -440
rect 39770 -475 39800 -440
rect 39800 -475 39805 -440
rect 39765 -480 39805 -475
rect 39935 -440 39975 -435
rect 39935 -475 39940 -440
rect 39940 -475 39970 -440
rect 39970 -475 39975 -440
rect 39935 -480 39975 -475
rect 40105 -440 40145 -435
rect 40105 -475 40110 -440
rect 40110 -475 40140 -440
rect 40140 -475 40145 -440
rect 40105 -480 40145 -475
rect 40275 -440 40315 -435
rect 40275 -475 40280 -440
rect 40280 -475 40310 -440
rect 40310 -475 40315 -440
rect 40275 -480 40315 -475
rect 40445 -440 40485 -435
rect 40445 -475 40450 -440
rect 40450 -475 40480 -440
rect 40480 -475 40485 -440
rect 40445 -480 40485 -475
rect 40615 -440 40655 -435
rect 40615 -475 40620 -440
rect 40620 -475 40650 -440
rect 40650 -475 40655 -440
rect 40615 -480 40655 -475
rect 40785 -440 40825 -435
rect 40785 -475 40790 -440
rect 40790 -475 40820 -440
rect 40820 -475 40825 -440
rect 40785 -480 40825 -475
rect 40955 -440 40995 -435
rect 40955 -475 40960 -440
rect 40960 -475 40990 -440
rect 40990 -475 40995 -440
rect 40955 -480 40995 -475
rect 41125 -440 41165 -435
rect 41125 -475 41130 -440
rect 41130 -475 41160 -440
rect 41160 -475 41165 -440
rect 41125 -480 41165 -475
rect 41295 -440 41335 -435
rect 41295 -475 41300 -440
rect 41300 -475 41330 -440
rect 41330 -475 41335 -440
rect 41295 -480 41335 -475
rect 41465 -440 41505 -435
rect 41465 -475 41470 -440
rect 41470 -475 41500 -440
rect 41500 -475 41505 -440
rect 41465 -480 41505 -475
rect 41635 -440 41675 -435
rect 41635 -475 41640 -440
rect 41640 -475 41670 -440
rect 41670 -475 41675 -440
rect 41635 -480 41675 -475
rect 41805 -440 41845 -435
rect 41805 -475 41810 -440
rect 41810 -475 41840 -440
rect 41840 -475 41845 -440
rect 41805 -480 41845 -475
rect 41975 -440 42015 -435
rect 41975 -475 41980 -440
rect 41980 -475 42010 -440
rect 42010 -475 42015 -440
rect 41975 -480 42015 -475
rect 42145 -440 42185 -435
rect 42145 -475 42150 -440
rect 42150 -475 42180 -440
rect 42180 -475 42185 -440
rect 42145 -480 42185 -475
rect 42315 -440 42355 -435
rect 42315 -475 42320 -440
rect 42320 -475 42350 -440
rect 42350 -475 42355 -440
rect 42315 -480 42355 -475
rect 42485 -440 42525 -435
rect 42485 -475 42490 -440
rect 42490 -475 42520 -440
rect 42520 -475 42525 -440
rect 42485 -480 42525 -475
rect 42655 -440 42695 -435
rect 42655 -475 42660 -440
rect 42660 -475 42690 -440
rect 42690 -475 42695 -440
rect 42655 -480 42695 -475
rect 42825 -440 42865 -435
rect 42825 -475 42830 -440
rect 42830 -475 42860 -440
rect 42860 -475 42865 -440
rect 42825 -480 42865 -475
rect 42995 -440 43035 -435
rect 42995 -475 43000 -440
rect 43000 -475 43030 -440
rect 43030 -475 43035 -440
rect 42995 -480 43035 -475
rect 43165 -440 43205 -435
rect 43165 -475 43170 -440
rect 43170 -475 43200 -440
rect 43200 -475 43205 -440
rect 43165 -480 43205 -475
rect 43335 -440 43375 -435
rect 43335 -475 43340 -440
rect 43340 -475 43370 -440
rect 43370 -475 43375 -440
rect 43335 -480 43375 -475
rect 43505 -440 43545 -435
rect 43505 -475 43510 -440
rect 43510 -475 43540 -440
rect 43540 -475 43545 -440
rect 43505 -480 43545 -475
rect 60 -760 120 -715
rect 740 -760 800 -715
rect 1420 -760 1480 -715
rect 2100 -760 2160 -715
rect 2780 -760 2840 -715
rect 3460 -760 3520 -715
rect 4140 -760 4200 -715
rect 4820 -760 4880 -715
rect 5500 -760 5560 -715
rect 6180 -760 6240 -715
rect 6860 -760 6920 -715
rect 7540 -760 7600 -715
rect 8220 -760 8280 -715
rect 8900 -760 8960 -715
rect 9580 -760 9640 -715
rect 10260 -760 10320 -715
rect 10940 -760 11000 -715
rect 11620 -760 11680 -715
rect 12300 -760 12360 -715
rect 12980 -760 13040 -715
rect 13660 -760 13720 -715
rect 14340 -760 14400 -715
rect 15020 -760 15080 -715
rect 15700 -760 15760 -715
rect 16380 -760 16440 -715
rect 17060 -760 17120 -715
rect 17740 -760 17800 -715
rect 18420 -760 18480 -715
rect 19100 -760 19160 -715
rect 19780 -760 19840 -715
rect 20460 -760 20520 -715
rect 21140 -760 21200 -715
rect 21820 -760 21880 -715
rect 22500 -760 22560 -715
rect 23180 -760 23240 -715
rect 23860 -760 23920 -715
rect 24540 -760 24600 -715
rect 25220 -760 25280 -715
rect 25900 -760 25960 -715
rect 26580 -760 26640 -715
rect 27260 -760 27320 -715
rect 27940 -760 28000 -715
rect 28620 -760 28680 -715
rect 29300 -760 29360 -715
rect 29980 -760 30040 -715
rect 30660 -760 30720 -715
rect 31340 -760 31400 -715
rect 32020 -760 32080 -715
rect 32700 -760 32760 -715
rect 33380 -760 33440 -715
rect 34060 -760 34120 -715
rect 34740 -760 34800 -715
rect 35420 -760 35480 -715
rect 36100 -760 36160 -715
rect 36780 -760 36840 -715
rect 37460 -760 37520 -715
rect 38140 -760 38200 -715
rect 38820 -760 38880 -715
rect 39500 -760 39560 -715
rect 40180 -760 40240 -715
rect 40860 -760 40920 -715
rect 41540 -760 41600 -715
rect 42220 -760 42280 -715
rect 42900 -760 42960 -715
<< metal4 >>
rect -284 370 -250 378
rect -284 335 -80 370
rect -284 200 -230 335
rect -100 330 -80 335
rect -100 290 180 330
rect -100 285 29670 290
rect -100 240 210 285
rect 270 240 550 285
rect 610 240 745 285
rect 805 240 1425 285
rect 1485 240 2105 285
rect 2165 240 2255 285
rect 2315 240 2935 285
rect 2995 240 3615 285
rect 3675 240 4295 285
rect 4355 240 4975 285
rect 5035 240 5655 285
rect 5715 240 6335 285
rect 6395 240 7015 285
rect 7075 240 7695 285
rect 7755 240 7845 285
rect 7905 240 8525 285
rect 8585 240 9205 285
rect 9265 240 9885 285
rect 9945 240 10565 285
rect 10625 240 11245 285
rect 11305 240 11925 285
rect 11985 240 12605 285
rect 12665 240 13285 285
rect 13345 240 13965 285
rect 14025 240 14645 285
rect 14705 240 15325 285
rect 15385 240 16005 285
rect 16065 240 16685 285
rect 16745 240 17365 285
rect 17425 240 18045 285
rect 18105 240 18725 285
rect 18785 240 19405 285
rect 19465 240 20085 285
rect 20145 240 20765 285
rect 20825 240 21445 285
rect 21505 240 22125 285
rect 22185 240 22805 285
rect 22865 240 23485 285
rect 23545 240 24165 285
rect 24225 240 24845 285
rect 24905 240 25525 285
rect 25585 240 26205 285
rect 26265 240 26885 285
rect 26945 240 27565 285
rect 27625 240 28245 285
rect 28305 240 28925 285
rect 28985 240 29605 285
rect 29665 240 29670 285
rect -100 235 29670 240
rect -100 205 180 235
rect -100 200 -80 205
rect -284 159 -80 200
rect -260 140 -80 159
rect 295 105 705 110
rect 295 60 305 105
rect 345 60 475 105
rect 515 60 645 105
rect 700 60 705 105
rect 295 55 705 60
rect 830 105 2245 110
rect 830 60 840 105
rect 880 60 1010 105
rect 1050 60 1180 105
rect 1220 60 1350 105
rect 1390 60 1520 105
rect 1560 60 1690 105
rect 1730 60 1860 105
rect 1900 60 2030 105
rect 2070 60 2185 105
rect 2240 60 2245 105
rect 830 55 2245 60
rect 2340 105 7835 110
rect 2340 60 2350 105
rect 2390 60 2520 105
rect 2560 60 2690 105
rect 2730 60 2860 105
rect 2900 60 3030 105
rect 3070 60 3200 105
rect 3240 60 3370 105
rect 3410 60 3540 105
rect 3580 60 3710 105
rect 3750 60 3880 105
rect 3920 60 4050 105
rect 4090 60 4220 105
rect 4260 60 4390 105
rect 4430 60 4560 105
rect 4600 60 4730 105
rect 4770 60 4900 105
rect 4940 60 5070 105
rect 5110 60 5240 105
rect 5280 60 5410 105
rect 5450 60 5580 105
rect 5620 60 5750 105
rect 5790 60 5920 105
rect 5960 60 6090 105
rect 6130 60 6260 105
rect 6300 60 6430 105
rect 6470 60 6600 105
rect 6640 60 6770 105
rect 6810 60 6940 105
rect 6980 60 7110 105
rect 7150 60 7280 105
rect 7320 60 7450 105
rect 7490 60 7620 105
rect 7660 60 7775 105
rect 7830 60 7835 105
rect 2340 55 7835 60
rect 7930 105 29600 110
rect 7930 60 7940 105
rect 7980 60 8110 105
rect 8150 60 8280 105
rect 8320 60 8450 105
rect 8490 60 8620 105
rect 8660 60 8790 105
rect 8830 60 8960 105
rect 9000 60 9130 105
rect 9170 60 9300 105
rect 9340 60 9470 105
rect 9510 60 9640 105
rect 9680 60 9810 105
rect 9850 60 9980 105
rect 10020 60 10150 105
rect 10190 60 10320 105
rect 10360 60 10490 105
rect 10530 60 10660 105
rect 10700 60 10830 105
rect 10870 60 11000 105
rect 11040 60 11170 105
rect 11210 60 11340 105
rect 11380 60 11510 105
rect 11550 60 11680 105
rect 11720 60 11850 105
rect 11890 60 12020 105
rect 12060 60 12190 105
rect 12230 60 12360 105
rect 12400 60 12530 105
rect 12570 60 12700 105
rect 12740 60 12870 105
rect 12910 60 13040 105
rect 13080 60 13210 105
rect 13250 60 13380 105
rect 13420 60 13550 105
rect 13590 60 13720 105
rect 13760 60 13890 105
rect 13930 60 14060 105
rect 14100 60 14230 105
rect 14270 60 14400 105
rect 14440 60 14570 105
rect 14610 60 14740 105
rect 14780 60 14910 105
rect 14950 60 15080 105
rect 15120 60 15250 105
rect 15290 60 15420 105
rect 15460 60 15590 105
rect 15630 60 15760 105
rect 15800 60 15930 105
rect 15970 60 16100 105
rect 16140 60 16270 105
rect 16310 60 16440 105
rect 16480 60 16610 105
rect 16650 60 16780 105
rect 16820 60 16950 105
rect 16990 60 17120 105
rect 17160 60 17290 105
rect 17330 60 17460 105
rect 17500 60 17630 105
rect 17670 60 17800 105
rect 17840 60 17970 105
rect 18010 60 18140 105
rect 18180 60 18310 105
rect 18350 60 18480 105
rect 18520 60 18650 105
rect 18690 60 18820 105
rect 18860 60 18990 105
rect 19030 60 19160 105
rect 19200 60 19330 105
rect 19370 60 19500 105
rect 19540 60 19670 105
rect 19710 60 19840 105
rect 19880 60 20010 105
rect 20050 60 20180 105
rect 20220 60 20350 105
rect 20390 60 20520 105
rect 20560 60 20690 105
rect 20730 60 20860 105
rect 20900 60 21030 105
rect 21070 60 21200 105
rect 21240 60 21370 105
rect 21410 60 21540 105
rect 21580 60 21710 105
rect 21750 60 21880 105
rect 21920 60 22050 105
rect 22090 60 22220 105
rect 22260 60 22390 105
rect 22430 60 22560 105
rect 22600 60 22730 105
rect 22770 60 22900 105
rect 22940 60 23070 105
rect 23110 60 23240 105
rect 23280 60 23410 105
rect 23450 60 23580 105
rect 23620 60 23750 105
rect 23790 60 23920 105
rect 23960 60 24090 105
rect 24130 60 24260 105
rect 24300 60 24430 105
rect 24470 60 24600 105
rect 24640 60 24770 105
rect 24810 60 24940 105
rect 24980 60 25110 105
rect 25150 60 25280 105
rect 25320 60 25450 105
rect 25490 60 25620 105
rect 25660 60 25790 105
rect 25830 60 25960 105
rect 26000 60 26130 105
rect 26170 60 26300 105
rect 26340 60 26470 105
rect 26510 60 26640 105
rect 26680 60 26810 105
rect 26850 60 26980 105
rect 27020 60 27150 105
rect 27190 60 27320 105
rect 27360 60 27490 105
rect 27530 60 27660 105
rect 27700 60 27830 105
rect 27870 60 28000 105
rect 28040 60 28170 105
rect 28210 60 28340 105
rect 28380 60 28510 105
rect 28550 60 28680 105
rect 28720 60 28850 105
rect 28890 60 29020 105
rect 29060 60 29190 105
rect 29230 60 29360 105
rect 29400 60 29530 105
rect 29570 60 29600 105
rect 7930 55 29600 60
rect -282 -110 175 -100
rect 39875 -110 40135 -105
rect -282 -135 43660 -110
rect -282 -185 65 -135
rect 115 -140 745 -135
rect 115 -185 215 -140
rect -282 -190 215 -185
rect 265 -190 555 -140
rect 605 -185 745 -140
rect 795 -140 2430 -135
rect 795 -185 1430 -140
rect 605 -190 1430 -185
rect 1480 -190 2275 -140
rect 2325 -185 2430 -140
rect 2480 -185 2955 -135
rect 3005 -185 3110 -135
rect 3160 -185 3465 -135
rect 3515 -140 4300 -135
rect 3515 -185 3620 -140
rect 2325 -190 3620 -185
rect 3670 -190 4145 -140
rect 4195 -185 4300 -140
rect 4350 -185 4825 -135
rect 4875 -185 4980 -135
rect 5030 -185 5335 -135
rect 5385 -140 5845 -135
rect 5385 -185 5490 -140
rect 4195 -190 5490 -185
rect 5540 -185 5845 -140
rect 5895 -140 6525 -135
rect 5895 -185 5995 -140
rect 5540 -190 5995 -185
rect 6045 -190 6335 -140
rect 6385 -185 6525 -140
rect 6575 -140 8190 -135
rect 6575 -185 7210 -140
rect 6385 -190 7210 -185
rect 7260 -190 8055 -140
rect 8105 -185 8190 -140
rect 8240 -185 8735 -135
rect 8785 -185 8870 -135
rect 8920 -185 9245 -135
rect 9295 -140 10060 -135
rect 9295 -185 9380 -140
rect 8105 -190 9380 -185
rect 9430 -190 9925 -140
rect 9975 -185 10060 -140
rect 10110 -185 10605 -135
rect 10655 -185 10740 -135
rect 10790 -185 11115 -135
rect 11165 -140 11795 -135
rect 11165 -185 11250 -140
rect 9975 -190 11250 -185
rect 11300 -185 11795 -140
rect 11845 -140 12475 -135
rect 11845 -185 11930 -140
rect 11300 -190 11930 -185
rect 11980 -190 12265 -140
rect 12315 -185 12475 -140
rect 12525 -140 14140 -135
rect 12525 -185 13160 -140
rect 12315 -190 13160 -185
rect 13210 -190 14005 -140
rect 14055 -185 14140 -140
rect 14190 -185 14685 -135
rect 14735 -185 14820 -135
rect 14870 -185 15195 -135
rect 15245 -140 16010 -135
rect 15245 -185 15330 -140
rect 14055 -190 15330 -185
rect 15380 -190 15875 -140
rect 15925 -185 16010 -140
rect 16060 -185 16555 -135
rect 16605 -185 16690 -135
rect 16740 -185 17065 -135
rect 17115 -140 17745 -135
rect 17115 -185 17200 -140
rect 15925 -190 17200 -185
rect 17250 -185 17745 -140
rect 17795 -140 18425 -135
rect 17795 -185 17880 -140
rect 17250 -190 17880 -185
rect 17930 -190 18215 -140
rect 18265 -185 18425 -140
rect 18475 -140 20635 -135
rect 18475 -185 19110 -140
rect 18265 -190 19110 -185
rect 19160 -190 19955 -140
rect 20005 -185 20635 -140
rect 20685 -185 21145 -135
rect 21195 -140 21825 -135
rect 21195 -185 21280 -140
rect 20005 -190 21280 -185
rect 21330 -190 21825 -140
rect 21875 -140 22505 -135
rect 21875 -190 22300 -140
rect 22350 -185 22505 -140
rect 22555 -140 24170 -135
rect 22555 -185 23190 -140
rect 22350 -190 23190 -185
rect 23240 -190 24035 -140
rect 24085 -185 24170 -140
rect 24220 -185 24715 -135
rect 24765 -185 24850 -135
rect 24900 -185 25225 -135
rect 25275 -140 26040 -135
rect 25275 -185 25360 -140
rect 24085 -190 25360 -185
rect 25410 -190 25905 -140
rect 25955 -185 26040 -140
rect 26090 -185 26585 -135
rect 26635 -185 26720 -135
rect 26770 -185 27095 -135
rect 27145 -185 27605 -135
rect 27655 -140 28285 -135
rect 27655 -185 27740 -140
rect 25955 -190 27740 -185
rect 27790 -185 28285 -140
rect 28335 -140 30495 -135
rect 28335 -185 28970 -140
rect 27790 -190 28970 -185
rect 29020 -190 29815 -140
rect 29865 -185 30495 -140
rect 30545 -185 31005 -135
rect 31055 -140 32365 -135
rect 31055 -185 31685 -140
rect 29865 -190 31685 -185
rect 31735 -185 32365 -140
rect 32415 -185 32875 -135
rect 32925 -185 33555 -135
rect 33605 -185 34235 -135
rect 34285 -140 36445 -135
rect 34285 -185 34920 -140
rect 31735 -190 34920 -185
rect 34970 -190 35765 -140
rect 35815 -185 36445 -140
rect 36495 -185 36955 -135
rect 37005 -140 38315 -135
rect 37005 -185 37635 -140
rect 35815 -190 37635 -185
rect 37685 -185 38315 -140
rect 38365 -185 38825 -135
rect 38875 -185 39505 -135
rect 39555 -185 40185 -135
rect 40235 -140 42395 -135
rect 40235 -185 40870 -140
rect 37685 -190 40870 -185
rect 40920 -190 41715 -140
rect 41765 -185 42395 -140
rect 42445 -185 42905 -135
rect 42955 -140 43660 -135
rect 42955 -185 43585 -140
rect 41765 -190 43585 -185
rect 43635 -190 43660 -140
rect -282 -215 43660 -190
rect -282 -225 175 -215
rect 39875 -220 40135 -215
rect -470 -410 180 -395
rect -470 -430 275 -410
rect -470 -435 43650 -430
rect -470 -480 155 -435
rect 195 -480 325 -435
rect 365 -480 495 -435
rect 535 -480 665 -435
rect 705 -480 835 -435
rect 875 -480 1005 -435
rect 1045 -480 1175 -435
rect 1215 -480 1345 -435
rect 1385 -480 1515 -435
rect 1555 -480 1685 -435
rect 1725 -480 1855 -435
rect 1895 -480 2025 -435
rect 2065 -480 2195 -435
rect 2235 -480 2365 -435
rect 2405 -480 2535 -435
rect 2575 -480 2705 -435
rect 2745 -480 2875 -435
rect 2915 -480 3045 -435
rect 3085 -480 3215 -435
rect 3255 -480 3385 -435
rect 3425 -480 3555 -435
rect 3595 -480 3725 -435
rect 3765 -480 3895 -435
rect 3935 -480 4065 -435
rect 4105 -480 4235 -435
rect 4275 -480 4405 -435
rect 4445 -480 4575 -435
rect 4615 -480 4745 -435
rect 4785 -480 4915 -435
rect 4955 -480 5085 -435
rect 5125 -480 5255 -435
rect 5295 -480 5425 -435
rect 5465 -480 5595 -435
rect 5635 -480 5765 -435
rect 5805 -480 5935 -435
rect 5975 -480 6105 -435
rect 6145 -480 6275 -435
rect 6315 -480 6445 -435
rect 6485 -480 6615 -435
rect 6655 -480 6785 -435
rect 6825 -480 6955 -435
rect 6995 -480 7125 -435
rect 7165 -480 7295 -435
rect 7335 -480 7465 -435
rect 7505 -480 7635 -435
rect 7675 -480 7805 -435
rect 7845 -480 7975 -435
rect 8015 -480 8145 -435
rect 8185 -480 8315 -435
rect 8355 -480 8485 -435
rect 8525 -480 8655 -435
rect 8695 -480 8825 -435
rect 8865 -480 8995 -435
rect 9035 -480 9165 -435
rect 9205 -480 9335 -435
rect 9375 -480 9505 -435
rect 9545 -480 9675 -435
rect 9715 -480 9845 -435
rect 9885 -480 10015 -435
rect 10055 -480 10185 -435
rect 10225 -480 10355 -435
rect 10395 -480 10525 -435
rect 10565 -480 10695 -435
rect 10735 -480 10865 -435
rect 10905 -480 11035 -435
rect 11075 -480 11205 -435
rect 11245 -480 11375 -435
rect 11415 -480 11545 -435
rect 11585 -480 11715 -435
rect 11755 -480 11885 -435
rect 11925 -480 12055 -435
rect 12095 -480 12225 -435
rect 12265 -480 12395 -435
rect 12435 -480 12565 -435
rect 12605 -480 12735 -435
rect 12775 -480 12905 -435
rect 12945 -480 13075 -435
rect 13115 -480 13245 -435
rect 13285 -480 13415 -435
rect 13455 -480 13585 -435
rect 13625 -480 13755 -435
rect 13795 -480 13925 -435
rect 13965 -480 14095 -435
rect 14135 -480 14265 -435
rect 14305 -480 14435 -435
rect 14475 -480 14605 -435
rect 14645 -480 14775 -435
rect 14815 -480 14945 -435
rect 14985 -480 15115 -435
rect 15155 -480 15285 -435
rect 15325 -480 15455 -435
rect 15495 -480 15625 -435
rect 15665 -480 15795 -435
rect 15835 -480 15965 -435
rect 16005 -480 16135 -435
rect 16175 -480 16305 -435
rect 16345 -480 16475 -435
rect 16515 -480 16645 -435
rect 16685 -480 16815 -435
rect 16855 -480 16985 -435
rect 17025 -480 17155 -435
rect 17195 -480 17325 -435
rect 17365 -480 17495 -435
rect 17535 -480 17665 -435
rect 17705 -480 17835 -435
rect 17875 -480 18005 -435
rect 18045 -480 18175 -435
rect 18215 -480 18345 -435
rect 18385 -480 18515 -435
rect 18555 -480 18685 -435
rect 18725 -480 18855 -435
rect 18895 -480 19025 -435
rect 19065 -480 19195 -435
rect 19235 -480 19365 -435
rect 19405 -480 19535 -435
rect 19575 -480 19705 -435
rect 19745 -480 19875 -435
rect 19915 -480 20045 -435
rect 20085 -480 20215 -435
rect 20255 -480 20385 -435
rect 20425 -480 20555 -435
rect 20595 -480 20725 -435
rect 20765 -480 20895 -435
rect 20935 -480 21065 -435
rect 21105 -480 21235 -435
rect 21275 -480 21405 -435
rect 21445 -480 21575 -435
rect 21615 -480 21745 -435
rect 21785 -480 21915 -435
rect 21955 -480 22085 -435
rect 22125 -480 22255 -435
rect 22295 -480 22425 -435
rect 22465 -480 22595 -435
rect 22635 -480 22765 -435
rect 22805 -480 22935 -435
rect 22975 -480 23105 -435
rect 23145 -480 23275 -435
rect 23315 -480 23445 -435
rect 23485 -480 23615 -435
rect 23655 -480 23785 -435
rect 23825 -480 23955 -435
rect 23995 -480 24125 -435
rect 24165 -480 24295 -435
rect 24335 -480 24465 -435
rect 24505 -480 24635 -435
rect 24675 -480 24805 -435
rect 24845 -480 24975 -435
rect 25015 -480 25145 -435
rect 25185 -480 25315 -435
rect 25355 -480 25485 -435
rect 25525 -480 25655 -435
rect 25695 -480 25825 -435
rect 25865 -480 25995 -435
rect 26035 -480 26165 -435
rect 26205 -480 26335 -435
rect 26375 -480 26505 -435
rect 26545 -480 26675 -435
rect 26715 -480 26845 -435
rect 26885 -480 27015 -435
rect 27055 -480 27185 -435
rect 27225 -480 27355 -435
rect 27395 -480 27525 -435
rect 27565 -480 27695 -435
rect 27735 -480 27865 -435
rect 27905 -480 28035 -435
rect 28075 -480 28205 -435
rect 28245 -480 28375 -435
rect 28415 -480 28545 -435
rect 28585 -480 28715 -435
rect 28755 -480 28885 -435
rect 28925 -480 29055 -435
rect 29095 -480 29225 -435
rect 29265 -480 29395 -435
rect 29435 -480 29565 -435
rect 29605 -480 29735 -435
rect 29775 -480 29905 -435
rect 29945 -480 30075 -435
rect 30115 -480 30245 -435
rect 30285 -480 30415 -435
rect 30455 -480 30585 -435
rect 30625 -480 30755 -435
rect 30795 -480 30925 -435
rect 30965 -480 31095 -435
rect 31135 -480 31265 -435
rect 31305 -480 31435 -435
rect 31475 -480 31605 -435
rect 31645 -480 31775 -435
rect 31815 -480 31945 -435
rect 31985 -480 32115 -435
rect 32155 -480 32285 -435
rect 32325 -480 32455 -435
rect 32495 -480 32625 -435
rect 32665 -480 32795 -435
rect 32835 -480 32965 -435
rect 33005 -480 33135 -435
rect 33175 -480 33305 -435
rect 33345 -480 33475 -435
rect 33515 -480 33645 -435
rect 33685 -480 33815 -435
rect 33855 -480 33985 -435
rect 34025 -480 34155 -435
rect 34195 -480 34325 -435
rect 34365 -480 34495 -435
rect 34535 -480 34665 -435
rect 34705 -480 34835 -435
rect 34875 -480 35005 -435
rect 35045 -480 35175 -435
rect 35215 -480 35345 -435
rect 35385 -480 35515 -435
rect 35555 -480 35685 -435
rect 35725 -480 35855 -435
rect 35895 -480 36025 -435
rect 36065 -480 36195 -435
rect 36235 -480 36365 -435
rect 36405 -480 36535 -435
rect 36575 -480 36705 -435
rect 36745 -480 36875 -435
rect 36915 -480 37045 -435
rect 37085 -480 37215 -435
rect 37255 -480 37385 -435
rect 37425 -480 37555 -435
rect 37595 -480 37725 -435
rect 37765 -480 37895 -435
rect 37935 -480 38065 -435
rect 38105 -480 38235 -435
rect 38275 -480 38405 -435
rect 38445 -480 38575 -435
rect 38615 -480 38745 -435
rect 38785 -480 38915 -435
rect 38955 -480 39085 -435
rect 39125 -480 39255 -435
rect 39295 -480 39425 -435
rect 39465 -480 39595 -435
rect 39635 -480 39765 -435
rect 39805 -480 39935 -435
rect 39975 -480 40105 -435
rect 40145 -480 40275 -435
rect 40315 -480 40445 -435
rect 40485 -480 40615 -435
rect 40655 -480 40785 -435
rect 40825 -480 40955 -435
rect 40995 -480 41125 -435
rect 41165 -480 41295 -435
rect 41335 -480 41465 -435
rect 41505 -480 41635 -435
rect 41675 -480 41805 -435
rect 41845 -480 41975 -435
rect 42015 -480 42145 -435
rect 42185 -480 42315 -435
rect 42355 -480 42485 -435
rect 42525 -480 42655 -435
rect 42695 -480 42825 -435
rect 42865 -480 42995 -435
rect 43035 -480 43165 -435
rect 43205 -480 43335 -435
rect 43375 -480 43505 -435
rect 43545 -480 43650 -435
rect -470 -485 43650 -480
rect -470 -505 275 -485
rect -470 -520 180 -505
rect -245 -670 -105 -660
rect -245 -700 -235 -670
rect -280 -775 -235 -700
rect -245 -805 -235 -775
rect -105 -710 195 -700
rect -105 -715 43660 -710
rect -105 -760 60 -715
rect 120 -760 740 -715
rect 800 -760 1420 -715
rect 1480 -760 2100 -715
rect 2160 -760 2780 -715
rect 2840 -760 3460 -715
rect 3520 -760 4140 -715
rect 4200 -760 4820 -715
rect 4880 -760 5500 -715
rect 5560 -760 6180 -715
rect 6240 -760 6860 -715
rect 6920 -760 7540 -715
rect 7600 -760 8220 -715
rect 8280 -760 8900 -715
rect 8960 -760 9580 -715
rect 9640 -760 10260 -715
rect 10320 -760 10940 -715
rect 11000 -760 11620 -715
rect 11680 -760 12300 -715
rect 12360 -760 12980 -715
rect 13040 -760 13660 -715
rect 13720 -760 14340 -715
rect 14400 -760 15020 -715
rect 15080 -760 15700 -715
rect 15760 -760 16380 -715
rect 16440 -760 17060 -715
rect 17120 -760 17740 -715
rect 17800 -760 18420 -715
rect 18480 -760 19100 -715
rect 19160 -760 19780 -715
rect 19840 -760 20460 -715
rect 20520 -760 21140 -715
rect 21200 -760 21820 -715
rect 21880 -760 22500 -715
rect 22560 -760 23180 -715
rect 23240 -760 23860 -715
rect 23920 -760 24540 -715
rect 24600 -760 25220 -715
rect 25280 -760 25900 -715
rect 25960 -760 26580 -715
rect 26640 -760 27260 -715
rect 27320 -760 27940 -715
rect 28000 -760 28620 -715
rect 28680 -760 29300 -715
rect 29360 -760 29980 -715
rect 30040 -760 30660 -715
rect 30720 -760 31340 -715
rect 31400 -760 32020 -715
rect 32080 -760 32700 -715
rect 32760 -760 33380 -715
rect 33440 -760 34060 -715
rect 34120 -760 34740 -715
rect 34800 -760 35420 -715
rect 35480 -760 36100 -715
rect 36160 -760 36780 -715
rect 36840 -760 37460 -715
rect 37520 -760 38140 -715
rect 38200 -760 38820 -715
rect 38880 -760 39500 -715
rect 39560 -760 40180 -715
rect 40240 -760 40860 -715
rect 40920 -760 41540 -715
rect 41600 -760 42220 -715
rect 42280 -760 42900 -715
rect 42960 -760 43660 -715
rect -105 -765 43660 -760
rect -105 -775 195 -765
rect -245 -815 -105 -805
<< via4 >>
rect -230 200 -100 335
rect -235 -805 -105 -670
<< metal5 >>
rect -280 378 -70 400
rect -284 335 -70 378
rect -284 200 -230 335
rect -100 200 -70 335
rect -284 159 -70 200
rect -280 -670 -70 159
rect -280 -805 -235 -670
rect -105 -805 -70 -670
rect -280 -910 -70 -805
<< labels >>
rlabel metal4 -376 -475 -376 -475 1 out
rlabel metal2 -410 25 -410 25 1 in
rlabel metal4 -15 276 -15 276 1 vdd!
rlabel metal4 -17 -186 -17 -186 1 gnd!
<< end >>
