magic
tech sky130A
timestamp 1647816202
<< locali >>
rect 4852 699 4944 707
rect 4852 625 4863 699
rect 4938 625 4944 699
rect 4852 616 4944 625
<< viali >>
rect 4863 625 4938 699
<< metal1 >>
rect 4852 706 4944 707
rect 5296 706 5397 710
rect 4852 699 5397 706
rect 4852 625 4863 699
rect 4938 625 5397 699
rect 4852 619 5397 625
rect 4852 616 4944 619
rect 5296 -143 5397 619
rect 2594 -145 5398 -143
rect 778 -147 5398 -145
rect -36 -251 5398 -147
rect -36 -252 2709 -251
rect -36 -314 40 -252
rect -76 -336 79 -314
rect -76 -455 -57 -336
rect 60 -455 79 -336
rect -76 -474 79 -455
<< via1 >>
rect -57 -455 60 -336
<< metal2 >>
rect -450 4360 -293 4383
rect -450 4256 -430 4360
rect -318 4256 -293 4360
rect -450 4239 -293 4256
rect -413 752 -333 4239
rect -191 2951 -32 2961
rect -191 2832 -174 2951
rect -50 2832 -32 2951
rect -191 2822 -32 2832
rect -144 2063 -69 2822
rect -144 2009 479 2063
rect -413 733 -320 752
rect -413 650 320 733
rect -413 648 235 650
rect -76 -336 79 -314
rect -76 -455 -57 -336
rect 60 -455 79 -336
rect -76 -474 79 -455
rect -38 -653 38 -474
<< via2 >>
rect -430 4256 -318 4360
rect -174 2832 -50 2951
<< metal3 >>
rect -450 4360 -293 4383
rect -450 4256 -430 4360
rect -318 4256 -293 4360
rect -450 4239 -293 4256
rect -191 2951 -32 2961
rect -191 2832 -174 2951
rect -50 2832 -32 2951
rect -191 2822 -32 2832
<< via3 >>
rect -430 4256 -318 4360
rect -174 2832 -50 2951
<< metal4 >>
rect -746 4517 342 4683
rect -736 3260 -610 4517
rect -450 4368 -293 4383
rect -453 4360 63 4368
rect -453 4256 -430 4360
rect -318 4256 63 4360
rect -453 4244 63 4256
rect -450 4239 -293 4244
rect -736 3094 377 3260
rect -736 -729 -610 3094
rect -191 2959 -32 2961
rect -198 2951 57 2959
rect -198 2832 -174 2951
rect -50 2832 57 2951
rect -198 2813 57 2832
rect 563 1476 707 1486
rect 563 1355 566 1476
rect 700 1355 707 1476
rect 563 1332 707 1355
rect -736 -895 367 -729
<< via4 >>
rect 566 1355 700 1476
<< metal5 >>
rect 185 3695 402 3949
rect 68 2350 404 2569
rect 69 1504 230 2350
rect 69 1476 732 1504
rect 69 1355 566 1476
rect 700 1355 732 1476
rect 69 1327 732 1355
rect 69 389 230 1327
rect 69 225 380 389
rect 163 -293 380 225
use tapered_buf  tapered_buf_1
timestamp 1647815768
transform 1 0 472 0 1 4762
box -470 -910 43675 404
use tapered_buf  tapered_buf_3
timestamp 1647815768
transform 1 0 447 0 1 -658
box -470 -910 43675 404
use tapered_buf  tapered_buf_0
timestamp 1647815768
transform 1 0 473 0 1 3342
box -470 -910 43675 404
use divider  divider_0
timestamp 1647816202
transform 1 0 489 0 1 235
box -490 -235 4690 2150
<< labels >>
rlabel space 44 3384 44 3384 1 mc2
rlabel space 30 -1142 30 -1142 1 out
rlabel metal4 -691 1606 -691 1606 1 gnd!
rlabel metal5 195 2465 195 2465 1 vdd!
rlabel space 24 4795 24 4795 1 clk
<< end >>
