magic
tech sky130A
timestamp 1647866489
<< locali >>
rect 4847 790 4958 799
rect -384 575 55 722
rect 4847 698 4859 790
rect 4949 698 4958 790
rect 4847 689 4958 698
<< viali >>
rect 4859 698 4949 790
<< metal1 >>
rect 4847 793 4958 799
rect 4847 790 5407 793
rect -480 730 -295 750
rect -480 568 -467 730
rect -308 568 -295 730
rect 4847 698 4859 790
rect 4949 698 5407 790
rect 4847 689 4958 698
rect -480 552 -295 568
rect 5301 -236 5407 698
rect -60 -316 29 -314
rect -60 -318 4956 -316
rect 5301 -318 5404 -236
rect -60 -402 5404 -318
rect -60 -707 29 -402
rect 2035 -404 5404 -402
rect 2035 -407 4956 -404
rect -143 -742 50 -707
rect -143 -873 -108 -742
rect 13 -873 50 -742
rect -143 -897 50 -873
<< via1 >>
rect -467 568 -308 730
rect -108 -873 13 -742
<< metal2 >>
rect -590 5259 -406 5277
rect -590 5126 -571 5259
rect -425 5126 -406 5259
rect -590 5110 -406 5126
rect -552 1658 -444 5110
rect -275 3858 -121 3870
rect -275 3743 -259 3858
rect -133 3743 -121 3858
rect -275 3729 -121 3743
rect -244 3039 -161 3729
rect -244 3037 252 3039
rect -244 2978 361 3037
rect -135 2976 361 2978
rect 300 2099 358 2976
rect -552 1568 7 1658
rect -86 794 4 1568
rect -86 791 258 794
rect -480 730 -295 750
rect -480 568 -467 730
rect -308 568 -295 730
rect -86 736 312 791
rect -86 725 258 736
rect -86 724 4 725
rect -480 552 -295 568
rect -143 -742 50 -707
rect -143 -873 -108 -742
rect 13 -873 50 -742
rect -143 -897 50 -873
<< via2 >>
rect -571 5126 -425 5259
rect -259 3743 -133 3858
rect -467 568 -308 730
<< metal3 >>
rect -590 5259 -406 5277
rect -590 5126 -571 5259
rect -425 5126 -406 5259
rect -590 5110 -406 5126
rect -275 3858 -121 3870
rect -275 3743 -259 3858
rect -133 3743 -121 3858
rect -275 3729 -121 3743
rect -480 730 -295 750
rect -480 568 -467 730
rect -308 568 -295 730
rect -480 552 -295 568
<< via3 >>
rect -571 5126 -425 5259
rect -259 3743 -133 3858
rect -467 568 -308 730
<< metal4 >>
rect -926 5386 308 5521
rect -924 4765 -768 5386
rect -590 5259 61 5293
rect -590 5126 -571 5259
rect -425 5126 61 5259
rect -590 5110 61 5126
rect -929 4173 -768 4765
rect -929 4164 308 4173
rect -926 4038 308 4164
rect -924 3845 -768 4038
rect -952 3373 -768 3845
rect -275 3858 63 3886
rect -275 3743 -259 3858
rect -133 3743 63 3858
rect -275 3729 63 3743
rect -924 713 -768 3373
rect 5673 1465 7697 1493
rect 4174 1421 7697 1465
rect 8466 1421 8575 3429
rect 4174 1403 8575 1421
rect 5673 1369 8575 1403
rect 5673 1343 7697 1369
rect -480 730 -295 750
rect -480 714 -467 730
rect -559 713 -467 714
rect -924 577 -467 713
rect -924 -959 -768 577
rect -559 573 -467 577
rect -480 568 -467 573
rect -308 568 -295 730
rect -480 552 -295 568
rect 8466 -612 8575 1369
rect -924 -1134 329 -959
rect -924 -1156 -768 -1134
<< metal5 >>
rect 186 4833 404 4838
rect 179 4404 414 4833
use tapered_buf  tapered_buf_1
timestamp 1647818295
transform 1 0 473 0 1 4272
box -470 -910 43675 401
use tapered_buf  tapered_buf_4
timestamp 1647818295
transform 1 0 473 0 1 5654
box -470 -910 43675 401
use divider  divider_0
timestamp 1647769399
transform 1 0 489 0 1 316
box -490 -235 4690 2150
use tapered_buf  tapered_buf_2
timestamp 1647818295
transform 1 0 434 0 1 -881
box -470 -910 43675 401
<< labels >>
rlabel space 40 -1345 40 -1345 1 up
rlabel metal4 8501 2091 8501 2091 1 vdd!
rlabel metal4 -877 1968 -877 1968 1 gnd!
rlabel metal4 48 3729 48 3729 1 ref
rlabel space 64 4302 64 4302 1 div
rlabel space 32 4313 32 4313 1 mc2
rlabel space 64 5650 64 5650 1 div
rlabel space 18 5671 18 5671 1 clk
<< end >>
