magic
tech sky130A
magscale 1 2
timestamp 1640983258
<< psubdiff >>
rect -3380 530 -3120 560
rect -3380 330 -3350 530
rect -3150 330 -3120 530
rect -3380 300 -3120 330
rect -2480 530 -2220 560
rect -2480 330 -2450 530
rect -2250 330 -2220 530
rect -2480 300 -2220 330
rect -1450 530 -1190 560
rect -1450 330 -1420 530
rect -1220 330 -1190 530
rect -1450 300 -1190 330
rect -420 530 -160 560
rect -420 330 -390 530
rect -190 330 -160 530
rect -420 300 -160 330
rect 610 530 870 560
rect 610 330 640 530
rect 840 330 870 530
rect 610 300 870 330
rect 1640 530 1900 560
rect 1640 330 1670 530
rect 1870 330 1900 530
rect 1640 300 1900 330
rect 2670 530 2930 560
rect 2670 330 2700 530
rect 2900 330 2930 530
rect 2670 300 2930 330
rect 4050 530 4310 560
rect 4050 330 4080 530
rect 4280 330 4310 530
rect 4050 300 4310 330
rect 5080 530 5340 560
rect 5080 330 5110 530
rect 5310 330 5340 530
rect 5080 300 5340 330
rect 6110 530 6370 560
rect 6110 330 6140 530
rect 6340 330 6370 530
rect 6110 300 6370 330
rect 7140 530 7400 560
rect 7140 330 7170 530
rect 7370 330 7400 530
rect 7140 300 7400 330
rect 8170 530 8430 560
rect 8170 330 8200 530
rect 8400 330 8430 530
rect 8170 300 8430 330
rect 9200 530 9460 560
rect 9200 330 9230 530
rect 9430 330 9460 530
rect 9200 300 9460 330
rect 10230 530 10490 560
rect 10230 330 10260 530
rect 10460 330 10490 530
rect 10230 300 10490 330
rect 11260 530 11520 560
rect 11260 330 11290 530
rect 11490 330 11520 530
rect 11260 300 11520 330
rect 11980 530 12240 560
rect 11980 330 12010 530
rect 12210 330 12240 530
rect 11980 300 12240 330
rect 11980 -710 12240 -680
rect -3380 -740 -3120 -710
rect -3380 -940 -3350 -740
rect -3150 -940 -3120 -740
rect 11980 -910 12010 -710
rect 12210 -910 12240 -710
rect 11980 -940 12240 -910
rect -3380 -970 -3120 -940
rect 11980 -1740 12240 -1710
rect -3380 -1770 -3120 -1740
rect -3380 -1970 -3350 -1770
rect -3150 -1970 -3120 -1770
rect 11980 -1940 12010 -1740
rect 12210 -1940 12240 -1740
rect 11980 -1970 12240 -1940
rect -3380 -2000 -3120 -1970
rect -3380 -2800 -3120 -2770
rect -3380 -3000 -3350 -2800
rect -3150 -3000 -3120 -2800
rect -3380 -3030 -3120 -3000
rect -3380 -3830 -3120 -3800
rect -3380 -4030 -3350 -3830
rect -3150 -4030 -3120 -3830
rect -3380 -4060 -3120 -4030
rect -3380 -4860 -3120 -4830
rect -3380 -5060 -3350 -4860
rect -3150 -5060 -3120 -4860
rect -3380 -5090 -3120 -5060
rect 11980 -2770 12240 -2740
rect 11980 -2970 12010 -2770
rect 12210 -2970 12240 -2770
rect 11980 -3000 12240 -2970
rect 11980 -3800 12240 -3770
rect 11980 -4000 12010 -3800
rect 12210 -4000 12240 -3800
rect 11980 -4030 12240 -4000
rect 11980 -4830 12240 -4800
rect 11980 -5030 12010 -4830
rect 12210 -5030 12240 -4830
rect 11980 -5060 12240 -5030
rect 11980 -5860 12240 -5830
rect -3380 -5890 -3120 -5860
rect -3380 -6090 -3350 -5890
rect -3150 -6090 -3120 -5890
rect 11980 -6060 12010 -5860
rect 12210 -6060 12240 -5860
rect 11980 -6090 12240 -6060
rect -3380 -6120 -3120 -6090
rect 11980 -6890 12240 -6860
rect -3380 -6920 -3120 -6890
rect -3380 -7120 -3350 -6920
rect -3150 -7120 -3120 -6920
rect 11980 -7090 12010 -6890
rect 12210 -7090 12240 -6890
rect 11980 -7120 12240 -7090
rect -3380 -7150 -3120 -7120
rect 11980 -8550 12240 -8520
rect -3380 -8580 -3120 -8550
rect -3380 -8780 -3350 -8580
rect -3150 -8780 -3120 -8580
rect 11980 -8750 12010 -8550
rect 12210 -8750 12240 -8550
rect 11980 -8780 12240 -8750
rect -3380 -8810 -3120 -8780
rect 11980 -9580 12240 -9550
rect -3380 -9610 -3120 -9580
rect -3380 -9810 -3350 -9610
rect -3150 -9810 -3120 -9610
rect 11980 -9780 12010 -9580
rect 12210 -9780 12240 -9580
rect 11980 -9810 12240 -9780
rect -3380 -9840 -3120 -9810
rect 11980 -10610 12240 -10580
rect -3380 -10640 -3120 -10610
rect -3380 -10840 -3350 -10640
rect -3150 -10840 -3120 -10640
rect 11980 -10810 12010 -10610
rect 12210 -10810 12240 -10610
rect 11980 -10840 12240 -10810
rect -3380 -10870 -3120 -10840
rect 11980 -11640 12240 -11610
rect -3380 -11670 -3120 -11640
rect -3380 -11870 -3350 -11670
rect -3150 -11870 -3120 -11670
rect 11980 -11840 12010 -11640
rect 12210 -11840 12240 -11640
rect 11980 -11870 12240 -11840
rect -3380 -11900 -3120 -11870
rect 11980 -12670 12240 -12640
rect -3380 -12700 -3120 -12670
rect -3380 -12900 -3350 -12700
rect -3150 -12900 -3120 -12700
rect 11980 -12870 12010 -12670
rect 12210 -12870 12240 -12670
rect 11980 -12900 12240 -12870
rect -3380 -12930 -3120 -12900
rect 11980 -13700 12240 -13670
rect -3380 -13730 -3120 -13700
rect -3380 -13930 -3350 -13730
rect -3150 -13930 -3120 -13730
rect 11980 -13900 12010 -13700
rect 12210 -13900 12240 -13700
rect 11980 -13930 12240 -13900
rect -3380 -13960 -3120 -13930
rect 11980 -15210 12240 -15180
rect -3380 -15240 -3120 -15210
rect -3380 -15440 -3350 -15240
rect -3150 -15440 -3120 -15240
rect 11980 -15410 12010 -15210
rect 12210 -15410 12240 -15210
rect 11980 -15440 12240 -15410
rect -3380 -15470 -3120 -15440
rect 11980 -16240 12240 -16210
rect -3380 -16270 -3120 -16240
rect -3380 -16470 -3350 -16270
rect -3150 -16470 -3120 -16270
rect 11980 -16440 12010 -16240
rect 12210 -16440 12240 -16240
rect 11980 -16470 12240 -16440
rect -3380 -16500 -3120 -16470
rect 11980 -17270 12240 -17240
rect -3380 -17300 -3120 -17270
rect -3380 -17500 -3350 -17300
rect -3150 -17500 -3120 -17300
rect 11980 -17470 12010 -17270
rect 12210 -17470 12240 -17270
rect 11980 -17500 12240 -17470
rect -3380 -17530 -3120 -17500
rect 11980 -18300 12240 -18270
rect -3380 -18330 -3120 -18300
rect -3380 -18530 -3350 -18330
rect -3150 -18530 -3120 -18330
rect 11980 -18500 12010 -18300
rect 12210 -18500 12240 -18300
rect 11980 -18530 12240 -18500
rect -3380 -18560 -3120 -18530
rect 11980 -19330 12240 -19300
rect -3380 -19360 -3120 -19330
rect -3380 -19560 -3350 -19360
rect -3150 -19560 -3120 -19360
rect 11980 -19530 12010 -19330
rect 12210 -19530 12240 -19330
rect 11980 -19560 12240 -19530
rect -3380 -19590 -3120 -19560
rect 11980 -20360 12240 -20330
rect -3380 -20390 -3120 -20360
rect -3380 -20590 -3350 -20390
rect -3150 -20590 -3120 -20390
rect 11980 -20560 12010 -20360
rect 12210 -20560 12240 -20360
rect 11980 -20590 12240 -20560
rect -3380 -20620 -3120 -20590
rect -3380 -21540 -3120 -21510
rect -3380 -21740 -3350 -21540
rect -3150 -21740 -3120 -21540
rect -3380 -21770 -3120 -21740
rect -2480 -21540 -2220 -21510
rect -2480 -21740 -2450 -21540
rect -2250 -21740 -2220 -21540
rect -2480 -21770 -2220 -21740
rect -1450 -21540 -1190 -21510
rect -1450 -21740 -1420 -21540
rect -1220 -21740 -1190 -21540
rect -1450 -21770 -1190 -21740
rect -420 -21540 -160 -21510
rect -420 -21740 -390 -21540
rect -190 -21740 -160 -21540
rect -420 -21770 -160 -21740
rect 610 -21540 870 -21510
rect 610 -21740 640 -21540
rect 840 -21740 870 -21540
rect 610 -21770 870 -21740
rect 1640 -21540 1900 -21510
rect 1640 -21740 1670 -21540
rect 1870 -21740 1900 -21540
rect 1640 -21770 1900 -21740
rect 2670 -21540 2930 -21510
rect 2670 -21740 2700 -21540
rect 2900 -21740 2930 -21540
rect 2670 -21770 2930 -21740
rect 3270 -21540 3530 -21510
rect 3270 -21740 3300 -21540
rect 3500 -21740 3530 -21540
rect 3270 -21770 3530 -21740
rect 4120 -21540 4380 -21510
rect 4120 -21740 4150 -21540
rect 4350 -21740 4380 -21540
rect 4120 -21770 4380 -21740
rect 4600 -21540 4860 -21510
rect 4600 -21740 4630 -21540
rect 4830 -21740 4860 -21540
rect 4600 -21770 4860 -21740
rect 5080 -21540 5340 -21510
rect 5080 -21740 5110 -21540
rect 5310 -21740 5340 -21540
rect 5080 -21770 5340 -21740
rect 6110 -21540 6370 -21510
rect 6110 -21740 6140 -21540
rect 6340 -21740 6370 -21540
rect 6110 -21770 6370 -21740
rect 7140 -21540 7400 -21510
rect 7140 -21740 7170 -21540
rect 7370 -21740 7400 -21540
rect 7140 -21770 7400 -21740
rect 8170 -21540 8430 -21510
rect 8170 -21740 8200 -21540
rect 8400 -21740 8430 -21540
rect 8170 -21770 8430 -21740
rect 9200 -21540 9460 -21510
rect 9200 -21740 9230 -21540
rect 9430 -21740 9460 -21540
rect 9200 -21770 9460 -21740
rect 10230 -21540 10490 -21510
rect 10230 -21740 10260 -21540
rect 10460 -21740 10490 -21540
rect 10230 -21770 10490 -21740
rect 11260 -21540 11520 -21510
rect 11260 -21740 11290 -21540
rect 11490 -21740 11520 -21540
rect 11260 -21770 11520 -21740
rect 11980 -21540 12240 -21510
rect 11980 -21740 12010 -21540
rect 12210 -21740 12240 -21540
rect 11980 -21770 12240 -21740
<< psubdiffcont >>
rect -3350 330 -3150 530
rect -2450 330 -2250 530
rect -1420 330 -1220 530
rect -390 330 -190 530
rect 640 330 840 530
rect 1670 330 1870 530
rect 2700 330 2900 530
rect 4080 330 4280 530
rect 5110 330 5310 530
rect 6140 330 6340 530
rect 7170 330 7370 530
rect 8200 330 8400 530
rect 9230 330 9430 530
rect 10260 330 10460 530
rect 11290 330 11490 530
rect 12010 330 12210 530
rect -3350 -940 -3150 -740
rect 12010 -910 12210 -710
rect -3350 -1970 -3150 -1770
rect 12010 -1940 12210 -1740
rect -3350 -3000 -3150 -2800
rect -3350 -4030 -3150 -3830
rect -3350 -5060 -3150 -4860
rect 12010 -2970 12210 -2770
rect 12010 -4000 12210 -3800
rect 12010 -5030 12210 -4830
rect -3350 -6090 -3150 -5890
rect 12010 -6060 12210 -5860
rect -3350 -7120 -3150 -6920
rect 12010 -7090 12210 -6890
rect -3350 -8780 -3150 -8580
rect 12010 -8750 12210 -8550
rect -3350 -9810 -3150 -9610
rect 12010 -9780 12210 -9580
rect -3350 -10840 -3150 -10640
rect 12010 -10810 12210 -10610
rect -3350 -11870 -3150 -11670
rect 12010 -11840 12210 -11640
rect -3350 -12900 -3150 -12700
rect 12010 -12870 12210 -12670
rect -3350 -13930 -3150 -13730
rect 12010 -13900 12210 -13700
rect -3350 -15440 -3150 -15240
rect 12010 -15410 12210 -15210
rect -3350 -16470 -3150 -16270
rect 12010 -16440 12210 -16240
rect -3350 -17500 -3150 -17300
rect 12010 -17470 12210 -17270
rect -3350 -18530 -3150 -18330
rect 12010 -18500 12210 -18300
rect -3350 -19560 -3150 -19360
rect 12010 -19530 12210 -19330
rect -3350 -20590 -3150 -20390
rect 12010 -20560 12210 -20360
rect -3350 -21740 -3150 -21540
rect -2450 -21740 -2250 -21540
rect -1420 -21740 -1220 -21540
rect -390 -21740 -190 -21540
rect 640 -21740 840 -21540
rect 1670 -21740 1870 -21540
rect 2700 -21740 2900 -21540
rect 3300 -21740 3500 -21540
rect 4150 -21740 4350 -21540
rect 4630 -21740 4830 -21540
rect 5110 -21740 5310 -21540
rect 6140 -21740 6340 -21540
rect 7170 -21740 7370 -21540
rect 8200 -21740 8400 -21540
rect 9230 -21740 9430 -21540
rect 10260 -21740 10460 -21540
rect 11290 -21740 11490 -21540
rect 12010 -21740 12210 -21540
<< xpolycontact >>
rect 4216 -2998 4286 -2566
rect 4216 -5230 4286 -4798
rect 4534 -2998 4604 -2566
rect 4534 -5230 4604 -4798
<< xpolyres >>
rect 4216 -4798 4286 -2998
rect 4534 -4798 4604 -2998
<< locali >>
rect -3600 530 12480 780
rect -3600 330 -3350 530
rect -3150 330 -2450 530
rect -2250 330 -1420 530
rect -1220 330 -390 530
rect -190 330 640 530
rect 840 330 1670 530
rect 1870 330 2700 530
rect 2900 330 4080 530
rect 4280 330 5110 530
rect 5310 330 6140 530
rect 6340 330 7170 530
rect 7370 330 8200 530
rect 8400 330 9230 530
rect 9430 330 10260 530
rect 10460 330 11290 530
rect 11490 330 12010 530
rect 12210 330 12480 530
rect -3600 60 12480 330
rect -3600 -740 -2880 60
rect -3600 -940 -3350 -740
rect -3150 -940 -2880 -740
rect -3600 -1770 -2880 -940
rect -3600 -1970 -3350 -1770
rect -3150 -1970 -2880 -1770
rect -3600 -2800 -2880 -1970
rect 11760 -710 12480 60
rect 11760 -910 12010 -710
rect 12210 -910 12480 -710
rect 11760 -1740 12480 -910
rect 11760 -1940 12010 -1740
rect 12210 -1940 12480 -1740
rect 4340 -2180 4670 -2160
rect 4340 -2380 4450 -2180
rect 4650 -2380 4670 -2180
rect 4340 -2400 4670 -2380
rect -3600 -3000 -3350 -2800
rect -3150 -3000 -2880 -2800
rect 11760 -2770 12480 -1940
rect 11760 -2970 12010 -2770
rect 12210 -2970 12480 -2770
rect -3600 -3830 -2880 -3000
rect -3600 -4030 -3350 -3830
rect -3150 -4030 -2880 -3830
rect -3600 -4860 -2880 -4030
rect 11760 -3800 12480 -2970
rect 11760 -4000 12010 -3800
rect 12210 -4000 12480 -3800
rect -3600 -5060 -3350 -4860
rect -3150 -5060 -2880 -4860
rect -3600 -5890 -2880 -5060
rect 11760 -4830 12480 -4000
rect 11760 -5030 12010 -4830
rect 12210 -5030 12480 -4830
rect -3600 -6090 -3350 -5890
rect -3150 -6090 -2880 -5890
rect -3600 -6920 -2880 -6090
rect -3600 -7120 -3350 -6920
rect -3150 -7120 -2880 -6920
rect -3600 -8580 -2880 -7120
rect -3600 -8780 -3350 -8580
rect -3150 -8780 -2880 -8580
rect -3600 -9610 -2880 -8780
rect -3600 -9810 -3350 -9610
rect -3150 -9810 -2880 -9610
rect -3600 -10640 -2880 -9810
rect -3600 -10840 -3350 -10640
rect -3150 -10840 -2880 -10640
rect -3600 -11670 -2880 -10840
rect -3600 -11870 -3350 -11670
rect -3150 -11870 -2880 -11670
rect -3600 -12700 -2880 -11870
rect -3600 -12900 -3350 -12700
rect -3150 -12900 -2880 -12700
rect -3600 -13730 -2880 -12900
rect -3600 -13930 -3350 -13730
rect -3150 -13930 -2880 -13730
rect -3600 -15240 -2880 -13930
rect -3600 -15440 -3350 -15240
rect -3150 -15440 -2880 -15240
rect -3600 -16270 -2880 -15440
rect -3600 -16470 -3350 -16270
rect -3150 -16470 -2880 -16270
rect -3600 -17300 -2880 -16470
rect -3600 -17500 -3350 -17300
rect -3150 -17500 -2880 -17300
rect -3600 -18330 -2880 -17500
rect -3600 -18530 -3350 -18330
rect -3150 -18530 -2880 -18330
rect -3600 -19360 -2880 -18530
rect -3600 -19560 -3350 -19360
rect -3150 -19560 -2880 -19360
rect -3600 -20390 -2880 -19560
rect -3600 -20590 -3350 -20390
rect -3150 -20590 -2880 -20390
rect -3600 -21290 -2880 -20590
rect 11760 -5860 12480 -5030
rect 11760 -6060 12010 -5860
rect 12210 -6060 12480 -5860
rect 11760 -6890 12480 -6060
rect 11760 -7090 12010 -6890
rect 12210 -7090 12480 -6890
rect 11760 -8550 12480 -7090
rect 11760 -8750 12010 -8550
rect 12210 -8750 12480 -8550
rect 11760 -9580 12480 -8750
rect 11760 -9780 12010 -9580
rect 12210 -9780 12480 -9580
rect 11760 -10610 12480 -9780
rect 11760 -10810 12010 -10610
rect 12210 -10810 12480 -10610
rect 11760 -11640 12480 -10810
rect 11760 -11840 12010 -11640
rect 12210 -11840 12480 -11640
rect 11760 -12670 12480 -11840
rect 11760 -12870 12010 -12670
rect 12210 -12870 12480 -12670
rect 11760 -13700 12480 -12870
rect 11760 -13900 12010 -13700
rect 12210 -13900 12480 -13700
rect 11760 -15210 12480 -13900
rect 11760 -15410 12010 -15210
rect 12210 -15410 12480 -15210
rect 11760 -16240 12480 -15410
rect 11760 -16440 12010 -16240
rect 12210 -16440 12480 -16240
rect 11760 -17270 12480 -16440
rect 11760 -17470 12010 -17270
rect 12210 -17470 12480 -17270
rect 11760 -18300 12480 -17470
rect 11760 -18500 12010 -18300
rect 12210 -18500 12480 -18300
rect 11760 -19330 12480 -18500
rect 11760 -19530 12010 -19330
rect 12210 -19530 12480 -19330
rect 11760 -20360 12480 -19530
rect 11760 -20560 12010 -20360
rect 12210 -20560 12480 -20360
rect 11760 -21290 12480 -20560
rect -3600 -21540 12480 -21290
rect -3600 -21740 -3350 -21540
rect -3150 -21740 -2450 -21540
rect -2250 -21740 -1420 -21540
rect -1220 -21740 -390 -21540
rect -190 -21740 640 -21540
rect 840 -21740 1670 -21540
rect 1870 -21740 2700 -21540
rect 2900 -21740 3300 -21540
rect 3500 -21740 4150 -21540
rect 4350 -21740 4630 -21540
rect 4830 -21740 5110 -21540
rect 5310 -21740 6140 -21540
rect 6340 -21740 7170 -21540
rect 7370 -21740 8200 -21540
rect 8400 -21740 9230 -21540
rect 9430 -21740 10260 -21540
rect 10460 -21740 11290 -21540
rect 11490 -21740 12010 -21540
rect 12210 -21740 12480 -21540
rect -3600 -22010 12480 -21740
<< viali >>
rect 4450 -2380 4650 -2180
rect 4232 -2981 4270 -2584
rect 4550 -2981 4588 -2584
rect 4232 -5212 4270 -4815
rect 4550 -5212 4588 -4815
rect 3300 -21740 3500 -21540
rect 4150 -21740 4350 -21540
rect 4630 -21740 4830 -21540
<< metal1 >>
rect 4420 -2180 4920 -2150
rect 4420 -2380 4450 -2180
rect 4650 -2380 4920 -2180
rect 4420 -2410 4920 -2380
rect 4226 -2580 4276 -2572
rect 4544 -2580 4594 -2572
rect 4226 -2584 4594 -2580
rect 4226 -2981 4232 -2584
rect 4270 -2981 4550 -2584
rect 4588 -2981 4594 -2584
rect 4226 -2990 4594 -2981
rect 4226 -2993 4276 -2990
rect 4544 -2993 4594 -2990
rect 4210 -4803 4240 -4800
rect 4210 -4810 4276 -4803
rect 3910 -4815 4276 -4810
rect 3910 -4950 4232 -4815
rect 3910 -5110 3950 -4950
rect 4110 -5110 4232 -4950
rect 3910 -5212 4232 -5110
rect 4270 -5212 4276 -4815
rect 3910 -5224 4276 -5212
rect 4544 -4810 4594 -4803
rect 4670 -4810 4920 -2410
rect 4544 -4815 4980 -4810
rect 4544 -5212 4550 -4815
rect 4588 -4960 4980 -4815
rect 4588 -5120 4680 -4960
rect 4840 -5120 4980 -4960
rect 4588 -5212 4980 -5120
rect 4544 -5224 4980 -5212
rect 3910 -5230 4240 -5224
rect 4580 -5230 4980 -5224
rect 3280 -21540 3520 -21520
rect 3280 -21740 3300 -21540
rect 3500 -21740 3520 -21540
rect 3280 -21760 3520 -21740
rect 4130 -21540 4370 -21520
rect 4130 -21740 4150 -21540
rect 4350 -21740 4370 -21540
rect 4130 -21760 4370 -21740
rect 4610 -21540 4850 -21520
rect 4610 -21740 4630 -21540
rect 4830 -21740 4850 -21540
rect 4610 -21760 4850 -21740
<< via1 >>
rect 3950 -5110 4110 -4950
rect 4680 -5120 4840 -4960
rect 3300 -21740 3500 -21540
rect 4150 -21740 4350 -21540
rect 4630 -21740 4830 -21540
<< metal2 >>
rect 3930 -4950 4130 -4930
rect 3930 -5110 3950 -4950
rect 4110 -5110 4130 -4950
rect 3930 -5130 4130 -5110
rect 4660 -4960 4860 -4940
rect 4660 -5120 4680 -4960
rect 4840 -5120 4860 -4960
rect 4660 -5140 4860 -5120
rect 3280 -21540 3520 -21520
rect 3280 -21740 3300 -21540
rect 3500 -21740 3520 -21540
rect 3280 -21760 3520 -21740
rect 4130 -21540 4370 -21520
rect 4130 -21740 4150 -21540
rect 4350 -21740 4370 -21540
rect 4130 -21760 4370 -21740
rect 4610 -21540 4850 -21520
rect 4610 -21740 4630 -21540
rect 4830 -21740 4850 -21540
rect 4610 -21760 4850 -21740
<< via2 >>
rect 3950 -5110 4110 -4950
rect 4680 -5120 4840 -4960
rect 3300 -21740 3500 -21540
rect 4150 -21740 4350 -21540
rect 4630 -21740 4830 -21540
<< metal3 >>
rect -2560 -6220 3600 -1030
rect 3930 -4950 4130 -4930
rect 3930 -5110 3950 -4950
rect 4110 -5110 4130 -4950
rect 3930 -5130 4130 -5110
rect 4660 -4960 4860 -4940
rect 4660 -5120 4680 -4960
rect 4840 -5120 4860 -4960
rect 4660 -5140 4860 -5120
rect 4960 -6220 11350 -970
rect -2560 -7520 11350 -6220
rect -2560 -7900 11180 -7520
rect -2560 -21120 10530 -7900
rect 140 -21130 920 -21120
rect 3190 -21540 4910 -21120
rect 3190 -21740 3300 -21540
rect 3500 -21740 4150 -21540
rect 4350 -21740 4630 -21540
rect 4830 -21740 4910 -21540
rect 3190 -21850 4910 -21740
<< via3 >>
rect 3950 -5110 4110 -4950
rect 4680 -5120 4840 -4960
<< mimcap >>
rect -2460 -1170 3540 -1130
rect -2460 -7090 -2420 -1170
rect 3500 -7090 3540 -1170
rect -2460 -7130 3540 -7090
rect 5290 -1170 11290 -1130
rect 5290 -7090 5330 -1170
rect 11250 -7090 11290 -1170
rect 5290 -7130 11290 -7090
rect 4470 -8010 10470 -7970
rect -2460 -8190 3540 -8150
rect -2460 -14110 -2420 -8190
rect 3500 -14110 3540 -8190
rect 4470 -13930 4510 -8010
rect 10430 -13930 10470 -8010
rect 4470 -13970 10470 -13930
rect -2460 -14150 3540 -14110
rect 4470 -14880 10470 -14840
rect -2460 -14980 3540 -14940
rect -2460 -20900 -2420 -14980
rect 3500 -20900 3540 -14980
rect 4470 -20800 4510 -14880
rect 10430 -20800 10470 -14880
rect 4470 -20840 10470 -20800
rect -2460 -20940 3540 -20900
<< mimcapcontact >>
rect -2420 -7090 3500 -1170
rect 5330 -7090 11250 -1170
rect -2420 -14110 3500 -8190
rect 4510 -13930 10430 -8010
rect -2420 -20900 3500 -14980
rect 4510 -20800 10430 -14880
<< metal4 >>
rect -2421 -1170 140 -1169
rect 920 -1170 3501 -1169
rect -2421 -7090 -2420 -1170
rect 3500 -4810 3501 -1170
rect 5329 -1170 7890 -1169
rect 8670 -1170 11251 -1169
rect 5329 -4810 5330 -1170
rect 3500 -4930 4070 -4810
rect 3500 -4950 4130 -4930
rect 4730 -4940 5330 -4810
rect 3500 -5110 3950 -4950
rect 4110 -5110 4130 -4950
rect 3500 -5130 4130 -5110
rect 4660 -4960 5330 -4940
rect 4660 -5120 4680 -4960
rect 4840 -5120 5330 -4960
rect 3500 -5230 4070 -5130
rect 4660 -5140 5330 -5120
rect 4730 -5230 5330 -5140
rect 3500 -7090 3501 -5230
rect -2421 -7091 3501 -7090
rect 5329 -7090 5330 -5230
rect 11250 -7090 11251 -1170
rect 5329 -7091 7890 -7090
rect 8670 -7091 11251 -7090
rect 140 -8189 920 -7091
rect 4509 -8010 7070 -8009
rect 7850 -8010 10431 -8009
rect -2421 -8190 3501 -8189
rect -2421 -14110 -2420 -8190
rect 3500 -14110 3501 -8190
rect 4509 -13930 4510 -8010
rect 10430 -13930 10431 -8010
rect 4509 -13931 10431 -13930
rect -2421 -14111 3501 -14110
rect 140 -14979 920 -14111
rect 7070 -14879 7850 -13931
rect 4509 -14880 10431 -14879
rect -2421 -14980 3501 -14979
rect -2421 -20900 -2420 -14980
rect 3500 -17580 3501 -14980
rect 4509 -17580 4510 -14880
rect 3500 -18450 4510 -17580
rect 3500 -20900 3501 -18450
rect 4509 -20800 4510 -18450
rect 10430 -20800 10431 -14880
rect 4509 -20801 7070 -20800
rect 7860 -20801 10431 -20800
rect -2421 -20901 140 -20900
rect 920 -20901 3501 -20900
<< labels >>
rlabel psubdiffcont 4660 -21680 4660 -21680 1 gnd!
rlabel psubdiffcont 4660 -21680 4660 -21680 1 gnd
rlabel locali 4370 -2280 4370 -2280 1 v
<< end >>
