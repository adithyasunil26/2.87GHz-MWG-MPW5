magic
tech sky130A
magscale 1 2
timestamp 1647903036
<< nwell >>
rect -70 170 59380 660
rect 70 -1610 87350 -940
<< pwell >>
rect 373 765 1515 1165
rect 5493 743 6635 1143
<< nmos >>
rect 550 0 580 100
rect 720 0 750 100
rect 890 0 920 100
rect 1060 0 1090 100
rect 1620 0 1650 100
rect 1790 0 1820 100
rect 1960 0 1990 100
rect 2130 0 2160 100
rect 2300 0 2330 100
rect 2470 0 2500 100
rect 2640 0 2670 100
rect 2810 0 2840 100
rect 2980 0 3010 100
rect 3150 0 3180 100
rect 3320 0 3350 100
rect 3490 0 3520 100
rect 3660 0 3690 100
rect 3830 0 3860 100
rect 4000 0 4030 100
rect 4170 0 4200 100
rect 4640 0 4670 100
rect 4810 0 4840 100
rect 4980 0 5010 100
rect 5150 0 5180 100
rect 5320 0 5350 100
rect 5490 0 5520 100
rect 5660 0 5690 100
rect 5830 0 5860 100
rect 6000 0 6030 100
rect 6170 0 6200 100
rect 6340 0 6370 100
rect 6510 0 6540 100
rect 6680 0 6710 100
rect 6850 0 6880 100
rect 7020 0 7050 100
rect 7190 0 7220 100
rect 7360 0 7390 100
rect 7530 0 7560 100
rect 7700 0 7730 100
rect 7870 0 7900 100
rect 8040 0 8070 100
rect 8210 0 8240 100
rect 8380 0 8410 100
rect 8550 0 8580 100
rect 8720 0 8750 100
rect 8890 0 8920 100
rect 9060 0 9090 100
rect 9230 0 9260 100
rect 9400 0 9430 100
rect 9570 0 9600 100
rect 9740 0 9770 100
rect 9910 0 9940 100
rect 10080 0 10110 100
rect 10250 0 10280 100
rect 10420 0 10450 100
rect 10590 0 10620 100
rect 10760 0 10790 100
rect 10930 0 10960 100
rect 11100 0 11130 100
rect 11270 0 11300 100
rect 11440 0 11470 100
rect 11610 0 11640 100
rect 11780 0 11810 100
rect 11950 0 11980 100
rect 12120 0 12150 100
rect 12290 0 12320 100
rect 12460 0 12490 100
rect 12630 0 12660 100
rect 12800 0 12830 100
rect 12970 0 13000 100
rect 13140 0 13170 100
rect 13310 0 13340 100
rect 13480 0 13510 100
rect 13650 0 13680 100
rect 13820 0 13850 100
rect 13990 0 14020 100
rect 14160 0 14190 100
rect 14330 0 14360 100
rect 14500 0 14530 100
rect 14670 0 14700 100
rect 14840 0 14870 100
rect 15010 0 15040 100
rect 15180 0 15210 100
rect 15350 0 15380 100
rect 15820 0 15850 100
rect 15990 0 16020 100
rect 16160 0 16190 100
rect 16330 0 16360 100
rect 16500 0 16530 100
rect 16670 0 16700 100
rect 16840 0 16870 100
rect 17010 0 17040 100
rect 17180 0 17210 100
rect 17350 0 17380 100
rect 17520 0 17550 100
rect 17690 0 17720 100
rect 17860 0 17890 100
rect 18030 0 18060 100
rect 18200 0 18230 100
rect 18370 0 18400 100
rect 18540 0 18570 100
rect 18710 0 18740 100
rect 18880 0 18910 100
rect 19050 0 19080 100
rect 19220 0 19250 100
rect 19390 0 19420 100
rect 19560 0 19590 100
rect 19730 0 19760 100
rect 19900 0 19930 100
rect 20070 0 20100 100
rect 20240 0 20270 100
rect 20410 0 20440 100
rect 20580 0 20610 100
rect 20750 0 20780 100
rect 20920 0 20950 100
rect 21090 0 21120 100
rect 21260 0 21290 100
rect 21430 0 21460 100
rect 21600 0 21630 100
rect 21770 0 21800 100
rect 21940 0 21970 100
rect 22110 0 22140 100
rect 22280 0 22310 100
rect 22450 0 22480 100
rect 22620 0 22650 100
rect 22790 0 22820 100
rect 22960 0 22990 100
rect 23130 0 23160 100
rect 23300 0 23330 100
rect 23470 0 23500 100
rect 23640 0 23670 100
rect 23810 0 23840 100
rect 23980 0 24010 100
rect 24150 0 24180 100
rect 24320 0 24350 100
rect 24490 0 24520 100
rect 24660 0 24690 100
rect 24830 0 24860 100
rect 25000 0 25030 100
rect 25170 0 25200 100
rect 25340 0 25370 100
rect 25510 0 25540 100
rect 25680 0 25710 100
rect 25850 0 25880 100
rect 26020 0 26050 100
rect 26190 0 26220 100
rect 26360 0 26390 100
rect 26530 0 26560 100
rect 26700 0 26730 100
rect 26870 0 26900 100
rect 27040 0 27070 100
rect 27210 0 27240 100
rect 27380 0 27410 100
rect 27550 0 27580 100
rect 27720 0 27750 100
rect 27890 0 27920 100
rect 28060 0 28090 100
rect 28230 0 28260 100
rect 28400 0 28430 100
rect 28570 0 28600 100
rect 28740 0 28770 100
rect 28910 0 28940 100
rect 29080 0 29110 100
rect 29250 0 29280 100
rect 29420 0 29450 100
rect 29590 0 29620 100
rect 29760 0 29790 100
rect 29930 0 29960 100
rect 30100 0 30130 100
rect 30270 0 30300 100
rect 30440 0 30470 100
rect 30610 0 30640 100
rect 30780 0 30810 100
rect 30950 0 30980 100
rect 31120 0 31150 100
rect 31290 0 31320 100
rect 31460 0 31490 100
rect 31630 0 31660 100
rect 31800 0 31830 100
rect 31970 0 32000 100
rect 32140 0 32170 100
rect 32310 0 32340 100
rect 32480 0 32510 100
rect 32650 0 32680 100
rect 32820 0 32850 100
rect 32990 0 33020 100
rect 33160 0 33190 100
rect 33330 0 33360 100
rect 33500 0 33530 100
rect 33670 0 33700 100
rect 33840 0 33870 100
rect 34010 0 34040 100
rect 34180 0 34210 100
rect 34350 0 34380 100
rect 34520 0 34550 100
rect 34690 0 34720 100
rect 34860 0 34890 100
rect 35030 0 35060 100
rect 35200 0 35230 100
rect 35370 0 35400 100
rect 35540 0 35570 100
rect 35710 0 35740 100
rect 35880 0 35910 100
rect 36050 0 36080 100
rect 36220 0 36250 100
rect 36390 0 36420 100
rect 36560 0 36590 100
rect 36730 0 36760 100
rect 36900 0 36930 100
rect 37070 0 37100 100
rect 37240 0 37270 100
rect 37410 0 37440 100
rect 37580 0 37610 100
rect 37750 0 37780 100
rect 37920 0 37950 100
rect 38090 0 38120 100
rect 38260 0 38290 100
rect 38430 0 38460 100
rect 38600 0 38630 100
rect 38770 0 38800 100
rect 38940 0 38970 100
rect 39110 0 39140 100
rect 39280 0 39310 100
rect 39450 0 39480 100
rect 39620 0 39650 100
rect 39790 0 39820 100
rect 39960 0 39990 100
rect 40130 0 40160 100
rect 40300 0 40330 100
rect 40470 0 40500 100
rect 40640 0 40670 100
rect 40810 0 40840 100
rect 40980 0 41010 100
rect 41150 0 41180 100
rect 41320 0 41350 100
rect 41490 0 41520 100
rect 41660 0 41690 100
rect 41830 0 41860 100
rect 42000 0 42030 100
rect 42170 0 42200 100
rect 42340 0 42370 100
rect 42510 0 42540 100
rect 42680 0 42710 100
rect 42850 0 42880 100
rect 43020 0 43050 100
rect 43190 0 43220 100
rect 43360 0 43390 100
rect 43530 0 43560 100
rect 43700 0 43730 100
rect 43870 0 43900 100
rect 44040 0 44070 100
rect 44210 0 44240 100
rect 44380 0 44410 100
rect 44550 0 44580 100
rect 44720 0 44750 100
rect 44890 0 44920 100
rect 45060 0 45090 100
rect 45230 0 45260 100
rect 45400 0 45430 100
rect 45570 0 45600 100
rect 45740 0 45770 100
rect 45910 0 45940 100
rect 46080 0 46110 100
rect 46250 0 46280 100
rect 46420 0 46450 100
rect 46590 0 46620 100
rect 46760 0 46790 100
rect 46930 0 46960 100
rect 47100 0 47130 100
rect 47270 0 47300 100
rect 47440 0 47470 100
rect 47610 0 47640 100
rect 47780 0 47810 100
rect 47950 0 47980 100
rect 48120 0 48150 100
rect 48290 0 48320 100
rect 48460 0 48490 100
rect 48630 0 48660 100
rect 48800 0 48830 100
rect 48970 0 49000 100
rect 49140 0 49170 100
rect 49310 0 49340 100
rect 49480 0 49510 100
rect 49650 0 49680 100
rect 49820 0 49850 100
rect 49990 0 50020 100
rect 50160 0 50190 100
rect 50330 0 50360 100
rect 50500 0 50530 100
rect 50670 0 50700 100
rect 50840 0 50870 100
rect 51010 0 51040 100
rect 51180 0 51210 100
rect 51350 0 51380 100
rect 51520 0 51550 100
rect 51690 0 51720 100
rect 51860 0 51890 100
rect 52030 0 52060 100
rect 52200 0 52230 100
rect 52370 0 52400 100
rect 52540 0 52570 100
rect 52710 0 52740 100
rect 52880 0 52910 100
rect 53050 0 53080 100
rect 53220 0 53250 100
rect 53390 0 53420 100
rect 53560 0 53590 100
rect 53730 0 53760 100
rect 53900 0 53930 100
rect 54070 0 54100 100
rect 54240 0 54270 100
rect 54410 0 54440 100
rect 54580 0 54610 100
rect 54750 0 54780 100
rect 54920 0 54950 100
rect 55090 0 55120 100
rect 55260 0 55290 100
rect 55430 0 55460 100
rect 55600 0 55630 100
rect 55770 0 55800 100
rect 55940 0 55970 100
rect 56110 0 56140 100
rect 56280 0 56310 100
rect 56450 0 56480 100
rect 56620 0 56650 100
rect 56790 0 56820 100
rect 56960 0 56990 100
rect 57130 0 57160 100
rect 57300 0 57330 100
rect 57470 0 57500 100
rect 57640 0 57670 100
rect 57810 0 57840 100
rect 57980 0 58010 100
rect 58150 0 58180 100
rect 58320 0 58350 100
rect 58490 0 58520 100
rect 58660 0 58690 100
rect 58830 0 58860 100
rect 59000 0 59030 100
rect 59170 0 59200 100
rect 130 -140 160 -40
rect 250 -850 280 -650
rect 420 -850 450 -650
rect 590 -850 620 -650
rect 760 -850 790 -650
rect 930 -850 960 -650
rect 1100 -850 1130 -650
rect 1270 -850 1300 -650
rect 1440 -850 1470 -650
rect 1610 -850 1640 -650
rect 1780 -850 1810 -650
rect 1950 -850 1980 -650
rect 2120 -850 2150 -650
rect 2290 -850 2320 -650
rect 2460 -850 2490 -650
rect 2630 -850 2660 -650
rect 2800 -850 2830 -650
rect 2970 -850 3000 -650
rect 3140 -850 3170 -650
rect 3310 -850 3340 -650
rect 3480 -850 3510 -650
rect 3650 -850 3680 -650
rect 3820 -850 3850 -650
rect 3990 -850 4020 -650
rect 4160 -850 4190 -650
rect 4330 -850 4360 -650
rect 4500 -850 4530 -650
rect 4670 -850 4700 -650
rect 4840 -850 4870 -650
rect 5010 -850 5040 -650
rect 5180 -850 5210 -650
rect 5350 -850 5380 -650
rect 5520 -850 5550 -650
rect 5690 -850 5720 -650
rect 5860 -850 5890 -650
rect 6030 -850 6060 -650
rect 6200 -850 6230 -650
rect 6370 -850 6400 -650
rect 6540 -850 6570 -650
rect 6710 -850 6740 -650
rect 6880 -850 6910 -650
rect 7050 -850 7080 -650
rect 7220 -850 7250 -650
rect 7390 -850 7420 -650
rect 7560 -850 7590 -650
rect 7730 -850 7760 -650
rect 7900 -850 7930 -650
rect 8070 -850 8100 -650
rect 8240 -850 8270 -650
rect 8410 -850 8440 -650
rect 8580 -850 8610 -650
rect 8750 -850 8780 -650
rect 8920 -850 8950 -650
rect 9090 -850 9120 -650
rect 9260 -850 9290 -650
rect 9430 -850 9460 -650
rect 9600 -850 9630 -650
rect 9770 -850 9800 -650
rect 9940 -850 9970 -650
rect 10110 -850 10140 -650
rect 10280 -850 10310 -650
rect 10450 -850 10480 -650
rect 10620 -850 10650 -650
rect 10790 -850 10820 -650
rect 10960 -850 10990 -650
rect 11130 -850 11160 -650
rect 11300 -850 11330 -650
rect 11470 -850 11500 -650
rect 11640 -850 11670 -650
rect 11810 -850 11840 -650
rect 11980 -850 12010 -650
rect 12150 -850 12180 -650
rect 12320 -850 12350 -650
rect 12490 -850 12520 -650
rect 12660 -850 12690 -650
rect 12830 -850 12860 -650
rect 13000 -850 13030 -650
rect 13170 -850 13200 -650
rect 13340 -850 13370 -650
rect 13510 -850 13540 -650
rect 13680 -850 13710 -650
rect 13850 -850 13880 -650
rect 14020 -850 14050 -650
rect 14190 -850 14220 -650
rect 14360 -850 14390 -650
rect 14530 -850 14560 -650
rect 14700 -850 14730 -650
rect 14870 -850 14900 -650
rect 15040 -850 15070 -650
rect 15210 -850 15240 -650
rect 15380 -850 15410 -650
rect 15550 -850 15580 -650
rect 15720 -850 15750 -650
rect 15890 -850 15920 -650
rect 16060 -850 16090 -650
rect 16230 -850 16260 -650
rect 16400 -850 16430 -650
rect 16570 -850 16600 -650
rect 16740 -850 16770 -650
rect 16910 -850 16940 -650
rect 17080 -850 17110 -650
rect 17250 -850 17280 -650
rect 17420 -850 17450 -650
rect 17590 -850 17620 -650
rect 17760 -850 17790 -650
rect 17930 -850 17960 -650
rect 18100 -850 18130 -650
rect 18270 -850 18300 -650
rect 18440 -850 18470 -650
rect 18610 -850 18640 -650
rect 18780 -850 18810 -650
rect 18950 -850 18980 -650
rect 19120 -850 19150 -650
rect 19290 -850 19320 -650
rect 19460 -850 19490 -650
rect 19630 -850 19660 -650
rect 19800 -850 19830 -650
rect 19970 -850 20000 -650
rect 20140 -850 20170 -650
rect 20310 -850 20340 -650
rect 20480 -850 20510 -650
rect 20650 -850 20680 -650
rect 20820 -850 20850 -650
rect 20990 -850 21020 -650
rect 21160 -850 21190 -650
rect 21330 -850 21360 -650
rect 21500 -850 21530 -650
rect 21670 -850 21700 -650
rect 21840 -850 21870 -650
rect 22010 -850 22040 -650
rect 22180 -850 22210 -650
rect 22350 -850 22380 -650
rect 22520 -850 22550 -650
rect 22690 -850 22720 -650
rect 22860 -850 22890 -650
rect 23030 -850 23060 -650
rect 23200 -850 23230 -650
rect 23370 -850 23400 -650
rect 23540 -850 23570 -650
rect 23710 -850 23740 -650
rect 23880 -850 23910 -650
rect 24050 -850 24080 -650
rect 24220 -850 24250 -650
rect 24390 -850 24420 -650
rect 24560 -850 24590 -650
rect 24730 -850 24760 -650
rect 24900 -850 24930 -650
rect 25070 -850 25100 -650
rect 25240 -850 25270 -650
rect 25410 -850 25440 -650
rect 25580 -850 25610 -650
rect 25750 -850 25780 -650
rect 25920 -850 25950 -650
rect 26090 -850 26120 -650
rect 26260 -850 26290 -650
rect 26430 -850 26460 -650
rect 26600 -850 26630 -650
rect 26770 -850 26800 -650
rect 26940 -850 26970 -650
rect 27110 -850 27140 -650
rect 27280 -850 27310 -650
rect 27450 -850 27480 -650
rect 27620 -850 27650 -650
rect 27790 -850 27820 -650
rect 27960 -850 27990 -650
rect 28130 -850 28160 -650
rect 28300 -850 28330 -650
rect 28470 -850 28500 -650
rect 28640 -850 28670 -650
rect 28810 -850 28840 -650
rect 28980 -850 29010 -650
rect 29150 -850 29180 -650
rect 29320 -850 29350 -650
rect 29490 -850 29520 -650
rect 29660 -850 29690 -650
rect 29830 -850 29860 -650
rect 30000 -850 30030 -650
rect 30170 -850 30200 -650
rect 30340 -850 30370 -650
rect 30510 -850 30540 -650
rect 30680 -850 30710 -650
rect 30850 -850 30880 -650
rect 31020 -850 31050 -650
rect 31190 -850 31220 -650
rect 31360 -850 31390 -650
rect 31530 -850 31560 -650
rect 31700 -850 31730 -650
rect 31870 -850 31900 -650
rect 32040 -850 32070 -650
rect 32210 -850 32240 -650
rect 32380 -850 32410 -650
rect 32550 -850 32580 -650
rect 32720 -850 32750 -650
rect 32890 -850 32920 -650
rect 33060 -850 33090 -650
rect 33230 -850 33260 -650
rect 33400 -850 33430 -650
rect 33570 -850 33600 -650
rect 33740 -850 33770 -650
rect 33910 -850 33940 -650
rect 34080 -850 34110 -650
rect 34250 -850 34280 -650
rect 34420 -850 34450 -650
rect 34590 -850 34620 -650
rect 34760 -850 34790 -650
rect 34930 -850 34960 -650
rect 35100 -850 35130 -650
rect 35270 -850 35300 -650
rect 35440 -850 35470 -650
rect 35610 -850 35640 -650
rect 35780 -850 35810 -650
rect 35950 -850 35980 -650
rect 36120 -850 36150 -650
rect 36290 -850 36320 -650
rect 36460 -850 36490 -650
rect 36630 -850 36660 -650
rect 36800 -850 36830 -650
rect 36970 -850 37000 -650
rect 37140 -850 37170 -650
rect 37310 -850 37340 -650
rect 37480 -850 37510 -650
rect 37650 -850 37680 -650
rect 37820 -850 37850 -650
rect 37990 -850 38020 -650
rect 38160 -850 38190 -650
rect 38330 -850 38360 -650
rect 38500 -850 38530 -650
rect 38670 -850 38700 -650
rect 38840 -850 38870 -650
rect 39010 -850 39040 -650
rect 39180 -850 39210 -650
rect 39350 -850 39380 -650
rect 39520 -850 39550 -650
rect 39690 -850 39720 -650
rect 39860 -850 39890 -650
rect 40030 -850 40060 -650
rect 40200 -850 40230 -650
rect 40370 -850 40400 -650
rect 40540 -850 40570 -650
rect 40710 -850 40740 -650
rect 40880 -850 40910 -650
rect 41050 -850 41080 -650
rect 41220 -850 41250 -650
rect 41390 -850 41420 -650
rect 41560 -850 41590 -650
rect 41730 -850 41760 -650
rect 41900 -850 41930 -650
rect 42070 -850 42100 -650
rect 42240 -850 42270 -650
rect 42410 -850 42440 -650
rect 42580 -850 42610 -650
rect 42750 -850 42780 -650
rect 42920 -850 42950 -650
rect 43090 -850 43120 -650
rect 43260 -850 43290 -650
rect 43430 -850 43460 -650
rect 43600 -850 43630 -650
rect 43770 -850 43800 -650
rect 43940 -850 43970 -650
rect 44110 -850 44140 -650
rect 44280 -850 44310 -650
rect 44450 -850 44480 -650
rect 44620 -850 44650 -650
rect 44790 -850 44820 -650
rect 44960 -850 44990 -650
rect 45130 -850 45160 -650
rect 45300 -850 45330 -650
rect 45470 -850 45500 -650
rect 45640 -850 45670 -650
rect 45810 -850 45840 -650
rect 45980 -850 46010 -650
rect 46150 -850 46180 -650
rect 46320 -850 46350 -650
rect 46490 -850 46520 -650
rect 46660 -850 46690 -650
rect 46830 -850 46860 -650
rect 47000 -850 47030 -650
rect 47170 -850 47200 -650
rect 47340 -850 47370 -650
rect 47510 -850 47540 -650
rect 47680 -850 47710 -650
rect 47850 -850 47880 -650
rect 48020 -850 48050 -650
rect 48190 -850 48220 -650
rect 48360 -850 48390 -650
rect 48530 -850 48560 -650
rect 48700 -850 48730 -650
rect 48870 -850 48900 -650
rect 49040 -850 49070 -650
rect 49210 -850 49240 -650
rect 49380 -850 49410 -650
rect 49550 -850 49580 -650
rect 49720 -850 49750 -650
rect 49890 -850 49920 -650
rect 50060 -850 50090 -650
rect 50230 -850 50260 -650
rect 50400 -850 50430 -650
rect 50570 -850 50600 -650
rect 50740 -850 50770 -650
rect 50910 -850 50940 -650
rect 51080 -850 51110 -650
rect 51250 -850 51280 -650
rect 51420 -850 51450 -650
rect 51590 -850 51620 -650
rect 51760 -850 51790 -650
rect 51930 -850 51960 -650
rect 52100 -850 52130 -650
rect 52270 -850 52300 -650
rect 52440 -850 52470 -650
rect 52610 -850 52640 -650
rect 52780 -850 52810 -650
rect 52950 -850 52980 -650
rect 53120 -850 53150 -650
rect 53290 -850 53320 -650
rect 53460 -850 53490 -650
rect 53630 -850 53660 -650
rect 53800 -850 53830 -650
rect 53970 -850 54000 -650
rect 54140 -850 54170 -650
rect 54310 -850 54340 -650
rect 54480 -850 54510 -650
rect 54650 -850 54680 -650
rect 54820 -850 54850 -650
rect 54990 -850 55020 -650
rect 55160 -850 55190 -650
rect 55330 -850 55360 -650
rect 55500 -850 55530 -650
rect 55670 -850 55700 -650
rect 55840 -850 55870 -650
rect 56010 -850 56040 -650
rect 56180 -850 56210 -650
rect 56350 -850 56380 -650
rect 56520 -850 56550 -650
rect 56690 -850 56720 -650
rect 56860 -850 56890 -650
rect 57030 -850 57060 -650
rect 57200 -850 57230 -650
rect 57370 -850 57400 -650
rect 57540 -850 57570 -650
rect 57710 -850 57740 -650
rect 57880 -850 57910 -650
rect 58050 -850 58080 -650
rect 58220 -850 58250 -650
rect 58390 -850 58420 -650
rect 58560 -850 58590 -650
rect 58730 -850 58760 -650
rect 58900 -850 58930 -650
rect 59070 -850 59100 -650
rect 59240 -850 59270 -650
rect 59410 -850 59440 -650
rect 59580 -850 59610 -650
rect 59750 -850 59780 -650
rect 59920 -850 59950 -650
rect 60090 -850 60120 -650
rect 60260 -850 60290 -650
rect 60430 -850 60460 -650
rect 60600 -850 60630 -650
rect 60770 -850 60800 -650
rect 60940 -850 60970 -650
rect 61110 -850 61140 -650
rect 61280 -850 61310 -650
rect 61450 -850 61480 -650
rect 61620 -850 61650 -650
rect 61790 -850 61820 -650
rect 61960 -850 61990 -650
rect 62130 -850 62160 -650
rect 62300 -850 62330 -650
rect 62470 -850 62500 -650
rect 62640 -850 62670 -650
rect 62810 -850 62840 -650
rect 62980 -850 63010 -650
rect 63150 -850 63180 -650
rect 63320 -850 63350 -650
rect 63490 -850 63520 -650
rect 63660 -850 63690 -650
rect 63830 -850 63860 -650
rect 64000 -850 64030 -650
rect 64170 -850 64200 -650
rect 64340 -850 64370 -650
rect 64510 -850 64540 -650
rect 64680 -850 64710 -650
rect 64850 -850 64880 -650
rect 65020 -850 65050 -650
rect 65190 -850 65220 -650
rect 65360 -850 65390 -650
rect 65530 -850 65560 -650
rect 65700 -850 65730 -650
rect 65870 -850 65900 -650
rect 66040 -850 66070 -650
rect 66210 -850 66240 -650
rect 66380 -850 66410 -650
rect 66550 -850 66580 -650
rect 66720 -850 66750 -650
rect 66890 -850 66920 -650
rect 67060 -850 67090 -650
rect 67230 -850 67260 -650
rect 67400 -850 67430 -650
rect 67570 -850 67600 -650
rect 67740 -850 67770 -650
rect 67910 -850 67940 -650
rect 68080 -850 68110 -650
rect 68250 -850 68280 -650
rect 68420 -850 68450 -650
rect 68590 -850 68620 -650
rect 68760 -850 68790 -650
rect 68930 -850 68960 -650
rect 69100 -850 69130 -650
rect 69270 -850 69300 -650
rect 69440 -850 69470 -650
rect 69610 -850 69640 -650
rect 69780 -850 69810 -650
rect 69950 -850 69980 -650
rect 70120 -850 70150 -650
rect 70290 -850 70320 -650
rect 70460 -850 70490 -650
rect 70630 -850 70660 -650
rect 70800 -850 70830 -650
rect 70970 -850 71000 -650
rect 71140 -850 71170 -650
rect 71310 -850 71340 -650
rect 71480 -850 71510 -650
rect 71650 -850 71680 -650
rect 71820 -850 71850 -650
rect 71990 -850 72020 -650
rect 72160 -850 72190 -650
rect 72330 -850 72360 -650
rect 72500 -850 72530 -650
rect 72670 -850 72700 -650
rect 72840 -850 72870 -650
rect 73010 -850 73040 -650
rect 73180 -850 73210 -650
rect 73350 -850 73380 -650
rect 73520 -850 73550 -650
rect 73690 -850 73720 -650
rect 73860 -850 73890 -650
rect 74030 -850 74060 -650
rect 74200 -850 74230 -650
rect 74370 -850 74400 -650
rect 74540 -850 74570 -650
rect 74710 -850 74740 -650
rect 74880 -850 74910 -650
rect 75050 -850 75080 -650
rect 75220 -850 75250 -650
rect 75390 -850 75420 -650
rect 75560 -850 75590 -650
rect 75730 -850 75760 -650
rect 75900 -850 75930 -650
rect 76070 -850 76100 -650
rect 76240 -850 76270 -650
rect 76410 -850 76440 -650
rect 76580 -850 76610 -650
rect 76750 -850 76780 -650
rect 76920 -850 76950 -650
rect 77090 -850 77120 -650
rect 77260 -850 77290 -650
rect 77430 -850 77460 -650
rect 77600 -850 77630 -650
rect 77770 -850 77800 -650
rect 77940 -850 77970 -650
rect 78110 -850 78140 -650
rect 78280 -850 78310 -650
rect 78450 -850 78480 -650
rect 78620 -850 78650 -650
rect 78790 -850 78820 -650
rect 78960 -850 78990 -650
rect 79130 -850 79160 -650
rect 79300 -850 79330 -650
rect 79470 -850 79500 -650
rect 79640 -850 79670 -650
rect 79810 -850 79840 -650
rect 79980 -850 80010 -650
rect 80150 -850 80180 -650
rect 80320 -850 80350 -650
rect 80490 -850 80520 -650
rect 80660 -850 80690 -650
rect 80830 -850 80860 -650
rect 81000 -850 81030 -650
rect 81170 -850 81200 -650
rect 81340 -850 81370 -650
rect 81510 -850 81540 -650
rect 81680 -850 81710 -650
rect 81850 -850 81880 -650
rect 82020 -850 82050 -650
rect 82190 -850 82220 -650
rect 82360 -850 82390 -650
rect 82530 -850 82560 -650
rect 82700 -850 82730 -650
rect 82870 -850 82900 -650
rect 83040 -850 83070 -650
rect 83210 -850 83240 -650
rect 83380 -850 83410 -650
rect 83550 -850 83580 -650
rect 83720 -850 83750 -650
rect 83890 -850 83920 -650
rect 84060 -850 84090 -650
rect 84230 -850 84260 -650
rect 84400 -850 84430 -650
rect 84570 -850 84600 -650
rect 84740 -850 84770 -650
rect 84910 -850 84940 -650
rect 85080 -850 85110 -650
rect 85250 -850 85280 -650
rect 85420 -850 85450 -650
rect 85590 -850 85620 -650
rect 85760 -850 85790 -650
rect 85930 -850 85960 -650
rect 86100 -850 86130 -650
rect 86270 -850 86300 -650
rect 86440 -850 86470 -650
rect 86610 -850 86640 -650
rect 86780 -850 86810 -650
rect 86950 -850 86980 -650
rect 87120 -850 87150 -650
<< pmos >>
rect 130 230 160 430
rect 550 230 580 430
rect 720 230 750 430
rect 890 230 920 430
rect 1060 230 1090 430
rect 1620 230 1650 430
rect 1790 230 1820 430
rect 1960 230 1990 430
rect 2130 230 2160 430
rect 2300 230 2330 430
rect 2470 230 2500 430
rect 2640 230 2670 430
rect 2810 230 2840 430
rect 2980 230 3010 430
rect 3150 230 3180 430
rect 3320 230 3350 430
rect 3490 230 3520 430
rect 3660 230 3690 430
rect 3830 230 3860 430
rect 4000 230 4030 430
rect 4170 230 4200 430
rect 4640 230 4670 430
rect 4810 230 4840 430
rect 4980 230 5010 430
rect 5150 230 5180 430
rect 5320 230 5350 430
rect 5490 230 5520 430
rect 5660 230 5690 430
rect 5830 230 5860 430
rect 6000 230 6030 430
rect 6170 230 6200 430
rect 6340 230 6370 430
rect 6510 230 6540 430
rect 6680 230 6710 430
rect 6850 230 6880 430
rect 7020 230 7050 430
rect 7190 230 7220 430
rect 7360 230 7390 430
rect 7530 230 7560 430
rect 7700 230 7730 430
rect 7870 230 7900 430
rect 8040 230 8070 430
rect 8210 230 8240 430
rect 8380 230 8410 430
rect 8550 230 8580 430
rect 8720 230 8750 430
rect 8890 230 8920 430
rect 9060 230 9090 430
rect 9230 230 9260 430
rect 9400 230 9430 430
rect 9570 230 9600 430
rect 9740 230 9770 430
rect 9910 230 9940 430
rect 10080 230 10110 430
rect 10250 230 10280 430
rect 10420 230 10450 430
rect 10590 230 10620 430
rect 10760 230 10790 430
rect 10930 230 10960 430
rect 11100 230 11130 430
rect 11270 230 11300 430
rect 11440 230 11470 430
rect 11610 230 11640 430
rect 11780 230 11810 430
rect 11950 230 11980 430
rect 12120 230 12150 430
rect 12290 230 12320 430
rect 12460 230 12490 430
rect 12630 230 12660 430
rect 12800 230 12830 430
rect 12970 230 13000 430
rect 13140 230 13170 430
rect 13310 230 13340 430
rect 13480 230 13510 430
rect 13650 230 13680 430
rect 13820 230 13850 430
rect 13990 230 14020 430
rect 14160 230 14190 430
rect 14330 230 14360 430
rect 14500 230 14530 430
rect 14670 230 14700 430
rect 14840 230 14870 430
rect 15010 230 15040 430
rect 15180 230 15210 430
rect 15350 230 15380 430
rect 15820 230 15850 430
rect 15990 230 16020 430
rect 16160 230 16190 430
rect 16330 230 16360 430
rect 16500 230 16530 430
rect 16670 230 16700 430
rect 16840 230 16870 430
rect 17010 230 17040 430
rect 17180 230 17210 430
rect 17350 230 17380 430
rect 17520 230 17550 430
rect 17690 230 17720 430
rect 17860 230 17890 430
rect 18030 230 18060 430
rect 18200 230 18230 430
rect 18370 230 18400 430
rect 18540 230 18570 430
rect 18710 230 18740 430
rect 18880 230 18910 430
rect 19050 230 19080 430
rect 19220 230 19250 430
rect 19390 230 19420 430
rect 19560 230 19590 430
rect 19730 230 19760 430
rect 19900 230 19930 430
rect 20070 230 20100 430
rect 20240 230 20270 430
rect 20410 230 20440 430
rect 20580 230 20610 430
rect 20750 230 20780 430
rect 20920 230 20950 430
rect 21090 230 21120 430
rect 21260 230 21290 430
rect 21430 230 21460 430
rect 21600 230 21630 430
rect 21770 230 21800 430
rect 21940 230 21970 430
rect 22110 230 22140 430
rect 22280 230 22310 430
rect 22450 230 22480 430
rect 22620 230 22650 430
rect 22790 230 22820 430
rect 22960 230 22990 430
rect 23130 230 23160 430
rect 23300 230 23330 430
rect 23470 230 23500 430
rect 23640 230 23670 430
rect 23810 230 23840 430
rect 23980 230 24010 430
rect 24150 230 24180 430
rect 24320 230 24350 430
rect 24490 230 24520 430
rect 24660 230 24690 430
rect 24830 230 24860 430
rect 25000 230 25030 430
rect 25170 230 25200 430
rect 25340 230 25370 430
rect 25510 230 25540 430
rect 25680 230 25710 430
rect 25850 230 25880 430
rect 26020 230 26050 430
rect 26190 230 26220 430
rect 26360 230 26390 430
rect 26530 230 26560 430
rect 26700 230 26730 430
rect 26870 230 26900 430
rect 27040 230 27070 430
rect 27210 230 27240 430
rect 27380 230 27410 430
rect 27550 230 27580 430
rect 27720 230 27750 430
rect 27890 230 27920 430
rect 28060 230 28090 430
rect 28230 230 28260 430
rect 28400 230 28430 430
rect 28570 230 28600 430
rect 28740 230 28770 430
rect 28910 230 28940 430
rect 29080 230 29110 430
rect 29250 230 29280 430
rect 29420 230 29450 430
rect 29590 230 29620 430
rect 29760 230 29790 430
rect 29930 230 29960 430
rect 30100 230 30130 430
rect 30270 230 30300 430
rect 30440 230 30470 430
rect 30610 230 30640 430
rect 30780 230 30810 430
rect 30950 230 30980 430
rect 31120 230 31150 430
rect 31290 230 31320 430
rect 31460 230 31490 430
rect 31630 230 31660 430
rect 31800 230 31830 430
rect 31970 230 32000 430
rect 32140 230 32170 430
rect 32310 230 32340 430
rect 32480 230 32510 430
rect 32650 230 32680 430
rect 32820 230 32850 430
rect 32990 230 33020 430
rect 33160 230 33190 430
rect 33330 230 33360 430
rect 33500 230 33530 430
rect 33670 230 33700 430
rect 33840 230 33870 430
rect 34010 230 34040 430
rect 34180 230 34210 430
rect 34350 230 34380 430
rect 34520 230 34550 430
rect 34690 230 34720 430
rect 34860 230 34890 430
rect 35030 230 35060 430
rect 35200 230 35230 430
rect 35370 230 35400 430
rect 35540 230 35570 430
rect 35710 230 35740 430
rect 35880 230 35910 430
rect 36050 230 36080 430
rect 36220 230 36250 430
rect 36390 230 36420 430
rect 36560 230 36590 430
rect 36730 230 36760 430
rect 36900 230 36930 430
rect 37070 230 37100 430
rect 37240 230 37270 430
rect 37410 230 37440 430
rect 37580 230 37610 430
rect 37750 230 37780 430
rect 37920 230 37950 430
rect 38090 230 38120 430
rect 38260 230 38290 430
rect 38430 230 38460 430
rect 38600 230 38630 430
rect 38770 230 38800 430
rect 38940 230 38970 430
rect 39110 230 39140 430
rect 39280 230 39310 430
rect 39450 230 39480 430
rect 39620 230 39650 430
rect 39790 230 39820 430
rect 39960 230 39990 430
rect 40130 230 40160 430
rect 40300 230 40330 430
rect 40470 230 40500 430
rect 40640 230 40670 430
rect 40810 230 40840 430
rect 40980 230 41010 430
rect 41150 230 41180 430
rect 41320 230 41350 430
rect 41490 230 41520 430
rect 41660 230 41690 430
rect 41830 230 41860 430
rect 42000 230 42030 430
rect 42170 230 42200 430
rect 42340 230 42370 430
rect 42510 230 42540 430
rect 42680 230 42710 430
rect 42850 230 42880 430
rect 43020 230 43050 430
rect 43190 230 43220 430
rect 43360 230 43390 430
rect 43530 230 43560 430
rect 43700 230 43730 430
rect 43870 230 43900 430
rect 44040 230 44070 430
rect 44210 230 44240 430
rect 44380 230 44410 430
rect 44550 230 44580 430
rect 44720 230 44750 430
rect 44890 230 44920 430
rect 45060 230 45090 430
rect 45230 230 45260 430
rect 45400 230 45430 430
rect 45570 230 45600 430
rect 45740 230 45770 430
rect 45910 230 45940 430
rect 46080 230 46110 430
rect 46250 230 46280 430
rect 46420 230 46450 430
rect 46590 230 46620 430
rect 46760 230 46790 430
rect 46930 230 46960 430
rect 47100 230 47130 430
rect 47270 230 47300 430
rect 47440 230 47470 430
rect 47610 230 47640 430
rect 47780 230 47810 430
rect 47950 230 47980 430
rect 48120 230 48150 430
rect 48290 230 48320 430
rect 48460 230 48490 430
rect 48630 230 48660 430
rect 48800 230 48830 430
rect 48970 230 49000 430
rect 49140 230 49170 430
rect 49310 230 49340 430
rect 49480 230 49510 430
rect 49650 230 49680 430
rect 49820 230 49850 430
rect 49990 230 50020 430
rect 50160 230 50190 430
rect 50330 230 50360 430
rect 50500 230 50530 430
rect 50670 230 50700 430
rect 50840 230 50870 430
rect 51010 230 51040 430
rect 51180 230 51210 430
rect 51350 230 51380 430
rect 51520 230 51550 430
rect 51690 230 51720 430
rect 51860 230 51890 430
rect 52030 230 52060 430
rect 52200 230 52230 430
rect 52370 230 52400 430
rect 52540 230 52570 430
rect 52710 230 52740 430
rect 52880 230 52910 430
rect 53050 230 53080 430
rect 53220 230 53250 430
rect 53390 230 53420 430
rect 53560 230 53590 430
rect 53730 230 53760 430
rect 53900 230 53930 430
rect 54070 230 54100 430
rect 54240 230 54270 430
rect 54410 230 54440 430
rect 54580 230 54610 430
rect 54750 230 54780 430
rect 54920 230 54950 430
rect 55090 230 55120 430
rect 55260 230 55290 430
rect 55430 230 55460 430
rect 55600 230 55630 430
rect 55770 230 55800 430
rect 55940 230 55970 430
rect 56110 230 56140 430
rect 56280 230 56310 430
rect 56450 230 56480 430
rect 56620 230 56650 430
rect 56790 230 56820 430
rect 56960 230 56990 430
rect 57130 230 57160 430
rect 57300 230 57330 430
rect 57470 230 57500 430
rect 57640 230 57670 430
rect 57810 230 57840 430
rect 57980 230 58010 430
rect 58150 230 58180 430
rect 58320 230 58350 430
rect 58490 230 58520 430
rect 58660 230 58690 430
rect 58830 230 58860 430
rect 59000 230 59030 430
rect 59170 230 59200 430
rect 250 -1380 280 -980
rect 420 -1380 450 -980
rect 590 -1380 620 -980
rect 760 -1380 790 -980
rect 930 -1380 960 -980
rect 1100 -1380 1130 -980
rect 1270 -1380 1300 -980
rect 1440 -1380 1470 -980
rect 1610 -1380 1640 -980
rect 1780 -1380 1810 -980
rect 1950 -1380 1980 -980
rect 2120 -1380 2150 -980
rect 2290 -1380 2320 -980
rect 2460 -1380 2490 -980
rect 2630 -1380 2660 -980
rect 2800 -1380 2830 -980
rect 2970 -1380 3000 -980
rect 3140 -1380 3170 -980
rect 3310 -1380 3340 -980
rect 3480 -1380 3510 -980
rect 3650 -1380 3680 -980
rect 3820 -1380 3850 -980
rect 3990 -1380 4020 -980
rect 4160 -1380 4190 -980
rect 4330 -1380 4360 -980
rect 4500 -1380 4530 -980
rect 4670 -1380 4700 -980
rect 4840 -1380 4870 -980
rect 5010 -1380 5040 -980
rect 5180 -1380 5210 -980
rect 5350 -1380 5380 -980
rect 5520 -1380 5550 -980
rect 5690 -1380 5720 -980
rect 5860 -1380 5890 -980
rect 6030 -1380 6060 -980
rect 6200 -1380 6230 -980
rect 6370 -1380 6400 -980
rect 6540 -1380 6570 -980
rect 6710 -1380 6740 -980
rect 6880 -1380 6910 -980
rect 7050 -1380 7080 -980
rect 7220 -1380 7250 -980
rect 7390 -1380 7420 -980
rect 7560 -1380 7590 -980
rect 7730 -1380 7760 -980
rect 7900 -1380 7930 -980
rect 8070 -1380 8100 -980
rect 8240 -1380 8270 -980
rect 8410 -1380 8440 -980
rect 8580 -1380 8610 -980
rect 8750 -1380 8780 -980
rect 8920 -1380 8950 -980
rect 9090 -1380 9120 -980
rect 9260 -1380 9290 -980
rect 9430 -1380 9460 -980
rect 9600 -1380 9630 -980
rect 9770 -1380 9800 -980
rect 9940 -1380 9970 -980
rect 10110 -1380 10140 -980
rect 10280 -1380 10310 -980
rect 10450 -1380 10480 -980
rect 10620 -1380 10650 -980
rect 10790 -1380 10820 -980
rect 10960 -1380 10990 -980
rect 11130 -1380 11160 -980
rect 11300 -1380 11330 -980
rect 11470 -1380 11500 -980
rect 11640 -1380 11670 -980
rect 11810 -1380 11840 -980
rect 11980 -1380 12010 -980
rect 12150 -1380 12180 -980
rect 12320 -1380 12350 -980
rect 12490 -1380 12520 -980
rect 12660 -1380 12690 -980
rect 12830 -1380 12860 -980
rect 13000 -1380 13030 -980
rect 13170 -1380 13200 -980
rect 13340 -1380 13370 -980
rect 13510 -1380 13540 -980
rect 13680 -1380 13710 -980
rect 13850 -1380 13880 -980
rect 14020 -1380 14050 -980
rect 14190 -1380 14220 -980
rect 14360 -1380 14390 -980
rect 14530 -1380 14560 -980
rect 14700 -1380 14730 -980
rect 14870 -1380 14900 -980
rect 15040 -1380 15070 -980
rect 15210 -1380 15240 -980
rect 15380 -1380 15410 -980
rect 15550 -1380 15580 -980
rect 15720 -1380 15750 -980
rect 15890 -1380 15920 -980
rect 16060 -1380 16090 -980
rect 16230 -1380 16260 -980
rect 16400 -1380 16430 -980
rect 16570 -1380 16600 -980
rect 16740 -1380 16770 -980
rect 16910 -1380 16940 -980
rect 17080 -1380 17110 -980
rect 17250 -1380 17280 -980
rect 17420 -1380 17450 -980
rect 17590 -1380 17620 -980
rect 17760 -1380 17790 -980
rect 17930 -1380 17960 -980
rect 18100 -1380 18130 -980
rect 18270 -1380 18300 -980
rect 18440 -1380 18470 -980
rect 18610 -1380 18640 -980
rect 18780 -1380 18810 -980
rect 18950 -1380 18980 -980
rect 19120 -1380 19150 -980
rect 19290 -1380 19320 -980
rect 19460 -1380 19490 -980
rect 19630 -1380 19660 -980
rect 19800 -1380 19830 -980
rect 19970 -1380 20000 -980
rect 20140 -1380 20170 -980
rect 20310 -1380 20340 -980
rect 20480 -1380 20510 -980
rect 20650 -1380 20680 -980
rect 20820 -1380 20850 -980
rect 20990 -1380 21020 -980
rect 21160 -1380 21190 -980
rect 21330 -1380 21360 -980
rect 21500 -1380 21530 -980
rect 21670 -1380 21700 -980
rect 21840 -1380 21870 -980
rect 22010 -1380 22040 -980
rect 22180 -1380 22210 -980
rect 22350 -1380 22380 -980
rect 22520 -1380 22550 -980
rect 22690 -1380 22720 -980
rect 22860 -1380 22890 -980
rect 23030 -1380 23060 -980
rect 23200 -1380 23230 -980
rect 23370 -1380 23400 -980
rect 23540 -1380 23570 -980
rect 23710 -1380 23740 -980
rect 23880 -1380 23910 -980
rect 24050 -1380 24080 -980
rect 24220 -1380 24250 -980
rect 24390 -1380 24420 -980
rect 24560 -1380 24590 -980
rect 24730 -1380 24760 -980
rect 24900 -1380 24930 -980
rect 25070 -1380 25100 -980
rect 25240 -1380 25270 -980
rect 25410 -1380 25440 -980
rect 25580 -1380 25610 -980
rect 25750 -1380 25780 -980
rect 25920 -1380 25950 -980
rect 26090 -1380 26120 -980
rect 26260 -1380 26290 -980
rect 26430 -1380 26460 -980
rect 26600 -1380 26630 -980
rect 26770 -1380 26800 -980
rect 26940 -1380 26970 -980
rect 27110 -1380 27140 -980
rect 27280 -1380 27310 -980
rect 27450 -1380 27480 -980
rect 27620 -1380 27650 -980
rect 27790 -1380 27820 -980
rect 27960 -1380 27990 -980
rect 28130 -1380 28160 -980
rect 28300 -1380 28330 -980
rect 28470 -1380 28500 -980
rect 28640 -1380 28670 -980
rect 28810 -1380 28840 -980
rect 28980 -1380 29010 -980
rect 29150 -1380 29180 -980
rect 29320 -1380 29350 -980
rect 29490 -1380 29520 -980
rect 29660 -1380 29690 -980
rect 29830 -1380 29860 -980
rect 30000 -1380 30030 -980
rect 30170 -1380 30200 -980
rect 30340 -1380 30370 -980
rect 30510 -1380 30540 -980
rect 30680 -1380 30710 -980
rect 30850 -1380 30880 -980
rect 31020 -1380 31050 -980
rect 31190 -1380 31220 -980
rect 31360 -1380 31390 -980
rect 31530 -1380 31560 -980
rect 31700 -1380 31730 -980
rect 31870 -1380 31900 -980
rect 32040 -1380 32070 -980
rect 32210 -1380 32240 -980
rect 32380 -1380 32410 -980
rect 32550 -1380 32580 -980
rect 32720 -1380 32750 -980
rect 32890 -1380 32920 -980
rect 33060 -1380 33090 -980
rect 33230 -1380 33260 -980
rect 33400 -1380 33430 -980
rect 33570 -1380 33600 -980
rect 33740 -1380 33770 -980
rect 33910 -1380 33940 -980
rect 34080 -1380 34110 -980
rect 34250 -1380 34280 -980
rect 34420 -1380 34450 -980
rect 34590 -1380 34620 -980
rect 34760 -1380 34790 -980
rect 34930 -1380 34960 -980
rect 35100 -1380 35130 -980
rect 35270 -1380 35300 -980
rect 35440 -1380 35470 -980
rect 35610 -1380 35640 -980
rect 35780 -1380 35810 -980
rect 35950 -1380 35980 -980
rect 36120 -1380 36150 -980
rect 36290 -1380 36320 -980
rect 36460 -1380 36490 -980
rect 36630 -1380 36660 -980
rect 36800 -1380 36830 -980
rect 36970 -1380 37000 -980
rect 37140 -1380 37170 -980
rect 37310 -1380 37340 -980
rect 37480 -1380 37510 -980
rect 37650 -1380 37680 -980
rect 37820 -1380 37850 -980
rect 37990 -1380 38020 -980
rect 38160 -1380 38190 -980
rect 38330 -1380 38360 -980
rect 38500 -1380 38530 -980
rect 38670 -1380 38700 -980
rect 38840 -1380 38870 -980
rect 39010 -1380 39040 -980
rect 39180 -1380 39210 -980
rect 39350 -1380 39380 -980
rect 39520 -1380 39550 -980
rect 39690 -1380 39720 -980
rect 39860 -1380 39890 -980
rect 40030 -1380 40060 -980
rect 40200 -1380 40230 -980
rect 40370 -1380 40400 -980
rect 40540 -1380 40570 -980
rect 40710 -1380 40740 -980
rect 40880 -1380 40910 -980
rect 41050 -1380 41080 -980
rect 41220 -1380 41250 -980
rect 41390 -1380 41420 -980
rect 41560 -1380 41590 -980
rect 41730 -1380 41760 -980
rect 41900 -1380 41930 -980
rect 42070 -1380 42100 -980
rect 42240 -1380 42270 -980
rect 42410 -1380 42440 -980
rect 42580 -1380 42610 -980
rect 42750 -1380 42780 -980
rect 42920 -1380 42950 -980
rect 43090 -1380 43120 -980
rect 43260 -1380 43290 -980
rect 43430 -1380 43460 -980
rect 43600 -1380 43630 -980
rect 43770 -1380 43800 -980
rect 43940 -1380 43970 -980
rect 44110 -1380 44140 -980
rect 44280 -1380 44310 -980
rect 44450 -1380 44480 -980
rect 44620 -1380 44650 -980
rect 44790 -1380 44820 -980
rect 44960 -1380 44990 -980
rect 45130 -1380 45160 -980
rect 45300 -1380 45330 -980
rect 45470 -1380 45500 -980
rect 45640 -1380 45670 -980
rect 45810 -1380 45840 -980
rect 45980 -1380 46010 -980
rect 46150 -1380 46180 -980
rect 46320 -1380 46350 -980
rect 46490 -1380 46520 -980
rect 46660 -1380 46690 -980
rect 46830 -1380 46860 -980
rect 47000 -1380 47030 -980
rect 47170 -1380 47200 -980
rect 47340 -1380 47370 -980
rect 47510 -1380 47540 -980
rect 47680 -1380 47710 -980
rect 47850 -1380 47880 -980
rect 48020 -1380 48050 -980
rect 48190 -1380 48220 -980
rect 48360 -1380 48390 -980
rect 48530 -1380 48560 -980
rect 48700 -1380 48730 -980
rect 48870 -1380 48900 -980
rect 49040 -1380 49070 -980
rect 49210 -1380 49240 -980
rect 49380 -1380 49410 -980
rect 49550 -1380 49580 -980
rect 49720 -1380 49750 -980
rect 49890 -1380 49920 -980
rect 50060 -1380 50090 -980
rect 50230 -1380 50260 -980
rect 50400 -1380 50430 -980
rect 50570 -1380 50600 -980
rect 50740 -1380 50770 -980
rect 50910 -1380 50940 -980
rect 51080 -1380 51110 -980
rect 51250 -1380 51280 -980
rect 51420 -1380 51450 -980
rect 51590 -1380 51620 -980
rect 51760 -1380 51790 -980
rect 51930 -1380 51960 -980
rect 52100 -1380 52130 -980
rect 52270 -1380 52300 -980
rect 52440 -1380 52470 -980
rect 52610 -1380 52640 -980
rect 52780 -1380 52810 -980
rect 52950 -1380 52980 -980
rect 53120 -1380 53150 -980
rect 53290 -1380 53320 -980
rect 53460 -1380 53490 -980
rect 53630 -1380 53660 -980
rect 53800 -1380 53830 -980
rect 53970 -1380 54000 -980
rect 54140 -1380 54170 -980
rect 54310 -1380 54340 -980
rect 54480 -1380 54510 -980
rect 54650 -1380 54680 -980
rect 54820 -1380 54850 -980
rect 54990 -1380 55020 -980
rect 55160 -1380 55190 -980
rect 55330 -1380 55360 -980
rect 55500 -1380 55530 -980
rect 55670 -1380 55700 -980
rect 55840 -1380 55870 -980
rect 56010 -1380 56040 -980
rect 56180 -1380 56210 -980
rect 56350 -1380 56380 -980
rect 56520 -1380 56550 -980
rect 56690 -1380 56720 -980
rect 56860 -1380 56890 -980
rect 57030 -1380 57060 -980
rect 57200 -1380 57230 -980
rect 57370 -1380 57400 -980
rect 57540 -1380 57570 -980
rect 57710 -1380 57740 -980
rect 57880 -1380 57910 -980
rect 58050 -1380 58080 -980
rect 58220 -1380 58250 -980
rect 58390 -1380 58420 -980
rect 58560 -1380 58590 -980
rect 58730 -1380 58760 -980
rect 58900 -1380 58930 -980
rect 59070 -1380 59100 -980
rect 59240 -1380 59270 -980
rect 59410 -1380 59440 -980
rect 59580 -1380 59610 -980
rect 59750 -1380 59780 -980
rect 59920 -1380 59950 -980
rect 60090 -1380 60120 -980
rect 60260 -1380 60290 -980
rect 60430 -1380 60460 -980
rect 60600 -1380 60630 -980
rect 60770 -1380 60800 -980
rect 60940 -1380 60970 -980
rect 61110 -1380 61140 -980
rect 61280 -1380 61310 -980
rect 61450 -1380 61480 -980
rect 61620 -1380 61650 -980
rect 61790 -1380 61820 -980
rect 61960 -1380 61990 -980
rect 62130 -1380 62160 -980
rect 62300 -1380 62330 -980
rect 62470 -1380 62500 -980
rect 62640 -1380 62670 -980
rect 62810 -1380 62840 -980
rect 62980 -1380 63010 -980
rect 63150 -1380 63180 -980
rect 63320 -1380 63350 -980
rect 63490 -1380 63520 -980
rect 63660 -1380 63690 -980
rect 63830 -1380 63860 -980
rect 64000 -1380 64030 -980
rect 64170 -1380 64200 -980
rect 64340 -1380 64370 -980
rect 64510 -1380 64540 -980
rect 64680 -1380 64710 -980
rect 64850 -1380 64880 -980
rect 65020 -1380 65050 -980
rect 65190 -1380 65220 -980
rect 65360 -1380 65390 -980
rect 65530 -1380 65560 -980
rect 65700 -1380 65730 -980
rect 65870 -1380 65900 -980
rect 66040 -1380 66070 -980
rect 66210 -1380 66240 -980
rect 66380 -1380 66410 -980
rect 66550 -1380 66580 -980
rect 66720 -1380 66750 -980
rect 66890 -1380 66920 -980
rect 67060 -1380 67090 -980
rect 67230 -1380 67260 -980
rect 67400 -1380 67430 -980
rect 67570 -1380 67600 -980
rect 67740 -1380 67770 -980
rect 67910 -1380 67940 -980
rect 68080 -1380 68110 -980
rect 68250 -1380 68280 -980
rect 68420 -1380 68450 -980
rect 68590 -1380 68620 -980
rect 68760 -1380 68790 -980
rect 68930 -1380 68960 -980
rect 69100 -1380 69130 -980
rect 69270 -1380 69300 -980
rect 69440 -1380 69470 -980
rect 69610 -1380 69640 -980
rect 69780 -1380 69810 -980
rect 69950 -1380 69980 -980
rect 70120 -1380 70150 -980
rect 70290 -1380 70320 -980
rect 70460 -1380 70490 -980
rect 70630 -1380 70660 -980
rect 70800 -1380 70830 -980
rect 70970 -1380 71000 -980
rect 71140 -1380 71170 -980
rect 71310 -1380 71340 -980
rect 71480 -1380 71510 -980
rect 71650 -1380 71680 -980
rect 71820 -1380 71850 -980
rect 71990 -1380 72020 -980
rect 72160 -1380 72190 -980
rect 72330 -1380 72360 -980
rect 72500 -1380 72530 -980
rect 72670 -1380 72700 -980
rect 72840 -1380 72870 -980
rect 73010 -1380 73040 -980
rect 73180 -1380 73210 -980
rect 73350 -1380 73380 -980
rect 73520 -1380 73550 -980
rect 73690 -1380 73720 -980
rect 73860 -1380 73890 -980
rect 74030 -1380 74060 -980
rect 74200 -1380 74230 -980
rect 74370 -1380 74400 -980
rect 74540 -1380 74570 -980
rect 74710 -1380 74740 -980
rect 74880 -1380 74910 -980
rect 75050 -1380 75080 -980
rect 75220 -1380 75250 -980
rect 75390 -1380 75420 -980
rect 75560 -1380 75590 -980
rect 75730 -1380 75760 -980
rect 75900 -1380 75930 -980
rect 76070 -1380 76100 -980
rect 76240 -1380 76270 -980
rect 76410 -1380 76440 -980
rect 76580 -1380 76610 -980
rect 76750 -1380 76780 -980
rect 76920 -1380 76950 -980
rect 77090 -1380 77120 -980
rect 77260 -1380 77290 -980
rect 77430 -1380 77460 -980
rect 77600 -1380 77630 -980
rect 77770 -1380 77800 -980
rect 77940 -1380 77970 -980
rect 78110 -1380 78140 -980
rect 78280 -1380 78310 -980
rect 78450 -1380 78480 -980
rect 78620 -1380 78650 -980
rect 78790 -1380 78820 -980
rect 78960 -1380 78990 -980
rect 79130 -1380 79160 -980
rect 79300 -1380 79330 -980
rect 79470 -1380 79500 -980
rect 79640 -1380 79670 -980
rect 79810 -1380 79840 -980
rect 79980 -1380 80010 -980
rect 80150 -1380 80180 -980
rect 80320 -1380 80350 -980
rect 80490 -1380 80520 -980
rect 80660 -1380 80690 -980
rect 80830 -1380 80860 -980
rect 81000 -1380 81030 -980
rect 81170 -1380 81200 -980
rect 81340 -1380 81370 -980
rect 81510 -1380 81540 -980
rect 81680 -1380 81710 -980
rect 81850 -1380 81880 -980
rect 82020 -1380 82050 -980
rect 82190 -1380 82220 -980
rect 82360 -1380 82390 -980
rect 82530 -1380 82560 -980
rect 82700 -1380 82730 -980
rect 82870 -1380 82900 -980
rect 83040 -1380 83070 -980
rect 83210 -1380 83240 -980
rect 83380 -1380 83410 -980
rect 83550 -1380 83580 -980
rect 83720 -1380 83750 -980
rect 83890 -1380 83920 -980
rect 84060 -1380 84090 -980
rect 84230 -1380 84260 -980
rect 84400 -1380 84430 -980
rect 84570 -1380 84600 -980
rect 84740 -1380 84770 -980
rect 84910 -1380 84940 -980
rect 85080 -1380 85110 -980
rect 85250 -1380 85280 -980
rect 85420 -1380 85450 -980
rect 85590 -1380 85620 -980
rect 85760 -1380 85790 -980
rect 85930 -1380 85960 -980
rect 86100 -1380 86130 -980
rect 86270 -1380 86300 -980
rect 86440 -1380 86470 -980
rect 86610 -1380 86640 -980
rect 86780 -1380 86810 -980
rect 86950 -1380 86980 -980
rect 87120 -1380 87150 -980
<< ndiff >>
rect 540 1007 580 1010
rect 531 995 634 1007
rect 531 935 543 995
rect 577 935 634 995
rect 531 923 634 935
rect 1254 995 1357 1007
rect 1254 935 1311 995
rect 1345 935 1357 995
rect 1254 923 1357 935
rect 540 910 580 923
rect 5651 973 5754 985
rect 5651 913 5663 973
rect 5697 913 5754 973
rect 5651 901 5754 913
rect 6374 973 6477 985
rect 6374 913 6431 973
rect 6465 913 6477 973
rect 6374 901 6477 913
rect 410 80 550 100
rect 410 20 450 80
rect 510 20 550 80
rect 410 0 550 20
rect 580 80 720 100
rect 580 20 620 80
rect 680 20 720 80
rect 580 0 720 20
rect 750 80 890 100
rect 750 20 790 80
rect 850 20 890 80
rect 750 0 890 20
rect 920 80 1060 100
rect 920 20 960 80
rect 1020 20 1060 80
rect 920 0 1060 20
rect 1090 80 1230 100
rect 1090 20 1130 80
rect 1190 20 1230 80
rect 1090 0 1230 20
rect 1480 80 1620 100
rect 1480 20 1520 80
rect 1580 20 1620 80
rect 1480 0 1620 20
rect 1650 80 1790 100
rect 1650 20 1690 80
rect 1750 20 1790 80
rect 1650 0 1790 20
rect 1820 80 1960 100
rect 1820 20 1860 80
rect 1920 20 1960 80
rect 1820 0 1960 20
rect 1990 80 2130 100
rect 1990 20 2030 80
rect 2090 20 2130 80
rect 1990 0 2130 20
rect 2160 80 2300 100
rect 2160 20 2200 80
rect 2260 20 2300 80
rect 2160 0 2300 20
rect 2330 80 2470 100
rect 2330 20 2370 80
rect 2430 20 2470 80
rect 2330 0 2470 20
rect 2500 80 2640 100
rect 2500 20 2540 80
rect 2600 20 2640 80
rect 2500 0 2640 20
rect 2670 80 2810 100
rect 2670 20 2710 80
rect 2770 20 2810 80
rect 2670 0 2810 20
rect 2840 80 2980 100
rect 2840 20 2880 80
rect 2940 20 2980 80
rect 2840 0 2980 20
rect 3010 80 3150 100
rect 3010 20 3050 80
rect 3110 20 3150 80
rect 3010 0 3150 20
rect 3180 80 3320 100
rect 3180 20 3220 80
rect 3280 20 3320 80
rect 3180 0 3320 20
rect 3350 80 3490 100
rect 3350 20 3390 80
rect 3450 20 3490 80
rect 3350 0 3490 20
rect 3520 80 3660 100
rect 3520 20 3560 80
rect 3620 20 3660 80
rect 3520 0 3660 20
rect 3690 80 3830 100
rect 3690 20 3730 80
rect 3790 20 3830 80
rect 3690 0 3830 20
rect 3860 80 4000 100
rect 3860 20 3900 80
rect 3960 20 4000 80
rect 3860 0 4000 20
rect 4030 80 4170 100
rect 4030 20 4070 80
rect 4130 20 4170 80
rect 4030 0 4170 20
rect 4200 80 4340 100
rect 4200 20 4240 80
rect 4300 20 4340 80
rect 4200 0 4340 20
rect 4500 80 4640 100
rect 4500 20 4540 80
rect 4600 20 4640 80
rect 4500 0 4640 20
rect 4670 80 4810 100
rect 4670 20 4710 80
rect 4770 20 4810 80
rect 4670 0 4810 20
rect 4840 80 4980 100
rect 4840 20 4880 80
rect 4940 20 4980 80
rect 4840 0 4980 20
rect 5010 80 5150 100
rect 5010 20 5050 80
rect 5110 20 5150 80
rect 5010 0 5150 20
rect 5180 80 5320 100
rect 5180 20 5220 80
rect 5280 20 5320 80
rect 5180 0 5320 20
rect 5350 80 5490 100
rect 5350 20 5390 80
rect 5450 20 5490 80
rect 5350 0 5490 20
rect 5520 80 5660 100
rect 5520 20 5560 80
rect 5620 20 5660 80
rect 5520 0 5660 20
rect 5690 80 5830 100
rect 5690 20 5730 80
rect 5790 20 5830 80
rect 5690 0 5830 20
rect 5860 80 6000 100
rect 5860 20 5900 80
rect 5960 20 6000 80
rect 5860 0 6000 20
rect 6030 80 6170 100
rect 6030 20 6070 80
rect 6130 20 6170 80
rect 6030 0 6170 20
rect 6200 80 6340 100
rect 6200 20 6240 80
rect 6300 20 6340 80
rect 6200 0 6340 20
rect 6370 80 6510 100
rect 6370 20 6410 80
rect 6470 20 6510 80
rect 6370 0 6510 20
rect 6540 80 6680 100
rect 6540 20 6580 80
rect 6640 20 6680 80
rect 6540 0 6680 20
rect 6710 80 6850 100
rect 6710 20 6750 80
rect 6810 20 6850 80
rect 6710 0 6850 20
rect 6880 80 7020 100
rect 6880 20 6920 80
rect 6980 20 7020 80
rect 6880 0 7020 20
rect 7050 80 7190 100
rect 7050 20 7090 80
rect 7150 20 7190 80
rect 7050 0 7190 20
rect 7220 80 7360 100
rect 7220 20 7260 80
rect 7320 20 7360 80
rect 7220 0 7360 20
rect 7390 80 7530 100
rect 7390 20 7430 80
rect 7490 20 7530 80
rect 7390 0 7530 20
rect 7560 80 7700 100
rect 7560 20 7600 80
rect 7660 20 7700 80
rect 7560 0 7700 20
rect 7730 80 7870 100
rect 7730 20 7770 80
rect 7830 20 7870 80
rect 7730 0 7870 20
rect 7900 80 8040 100
rect 7900 20 7940 80
rect 8000 20 8040 80
rect 7900 0 8040 20
rect 8070 80 8210 100
rect 8070 20 8110 80
rect 8170 20 8210 80
rect 8070 0 8210 20
rect 8240 80 8380 100
rect 8240 20 8280 80
rect 8340 20 8380 80
rect 8240 0 8380 20
rect 8410 80 8550 100
rect 8410 20 8450 80
rect 8510 20 8550 80
rect 8410 0 8550 20
rect 8580 80 8720 100
rect 8580 20 8620 80
rect 8680 20 8720 80
rect 8580 0 8720 20
rect 8750 80 8890 100
rect 8750 20 8790 80
rect 8850 20 8890 80
rect 8750 0 8890 20
rect 8920 80 9060 100
rect 8920 20 8960 80
rect 9020 20 9060 80
rect 8920 0 9060 20
rect 9090 80 9230 100
rect 9090 20 9130 80
rect 9190 20 9230 80
rect 9090 0 9230 20
rect 9260 80 9400 100
rect 9260 20 9300 80
rect 9360 20 9400 80
rect 9260 0 9400 20
rect 9430 80 9570 100
rect 9430 20 9470 80
rect 9530 20 9570 80
rect 9430 0 9570 20
rect 9600 80 9740 100
rect 9600 20 9640 80
rect 9700 20 9740 80
rect 9600 0 9740 20
rect 9770 80 9910 100
rect 9770 20 9810 80
rect 9870 20 9910 80
rect 9770 0 9910 20
rect 9940 80 10080 100
rect 9940 20 9980 80
rect 10040 20 10080 80
rect 9940 0 10080 20
rect 10110 80 10250 100
rect 10110 20 10150 80
rect 10210 20 10250 80
rect 10110 0 10250 20
rect 10280 80 10420 100
rect 10280 20 10320 80
rect 10380 20 10420 80
rect 10280 0 10420 20
rect 10450 80 10590 100
rect 10450 20 10490 80
rect 10550 20 10590 80
rect 10450 0 10590 20
rect 10620 80 10760 100
rect 10620 20 10660 80
rect 10720 20 10760 80
rect 10620 0 10760 20
rect 10790 80 10930 100
rect 10790 20 10830 80
rect 10890 20 10930 80
rect 10790 0 10930 20
rect 10960 80 11100 100
rect 10960 20 11000 80
rect 11060 20 11100 80
rect 10960 0 11100 20
rect 11130 80 11270 100
rect 11130 20 11170 80
rect 11230 20 11270 80
rect 11130 0 11270 20
rect 11300 80 11440 100
rect 11300 20 11340 80
rect 11400 20 11440 80
rect 11300 0 11440 20
rect 11470 80 11610 100
rect 11470 20 11510 80
rect 11570 20 11610 80
rect 11470 0 11610 20
rect 11640 80 11780 100
rect 11640 20 11680 80
rect 11740 20 11780 80
rect 11640 0 11780 20
rect 11810 80 11950 100
rect 11810 20 11850 80
rect 11910 20 11950 80
rect 11810 0 11950 20
rect 11980 80 12120 100
rect 11980 20 12020 80
rect 12080 20 12120 80
rect 11980 0 12120 20
rect 12150 80 12290 100
rect 12150 20 12190 80
rect 12250 20 12290 80
rect 12150 0 12290 20
rect 12320 80 12460 100
rect 12320 20 12360 80
rect 12420 20 12460 80
rect 12320 0 12460 20
rect 12490 80 12630 100
rect 12490 20 12530 80
rect 12590 20 12630 80
rect 12490 0 12630 20
rect 12660 80 12800 100
rect 12660 20 12700 80
rect 12760 20 12800 80
rect 12660 0 12800 20
rect 12830 80 12970 100
rect 12830 20 12870 80
rect 12930 20 12970 80
rect 12830 0 12970 20
rect 13000 80 13140 100
rect 13000 20 13040 80
rect 13100 20 13140 80
rect 13000 0 13140 20
rect 13170 80 13310 100
rect 13170 20 13210 80
rect 13270 20 13310 80
rect 13170 0 13310 20
rect 13340 80 13480 100
rect 13340 20 13380 80
rect 13440 20 13480 80
rect 13340 0 13480 20
rect 13510 80 13650 100
rect 13510 20 13550 80
rect 13610 20 13650 80
rect 13510 0 13650 20
rect 13680 80 13820 100
rect 13680 20 13720 80
rect 13780 20 13820 80
rect 13680 0 13820 20
rect 13850 80 13990 100
rect 13850 20 13890 80
rect 13950 20 13990 80
rect 13850 0 13990 20
rect 14020 80 14160 100
rect 14020 20 14060 80
rect 14120 20 14160 80
rect 14020 0 14160 20
rect 14190 80 14330 100
rect 14190 20 14230 80
rect 14290 20 14330 80
rect 14190 0 14330 20
rect 14360 80 14500 100
rect 14360 20 14400 80
rect 14460 20 14500 80
rect 14360 0 14500 20
rect 14530 80 14670 100
rect 14530 20 14570 80
rect 14630 20 14670 80
rect 14530 0 14670 20
rect 14700 80 14840 100
rect 14700 20 14740 80
rect 14800 20 14840 80
rect 14700 0 14840 20
rect 14870 80 15010 100
rect 14870 20 14910 80
rect 14970 20 15010 80
rect 14870 0 15010 20
rect 15040 80 15180 100
rect 15040 20 15080 80
rect 15140 20 15180 80
rect 15040 0 15180 20
rect 15210 80 15350 100
rect 15210 20 15250 80
rect 15310 20 15350 80
rect 15210 0 15350 20
rect 15380 80 15520 100
rect 15380 20 15420 80
rect 15480 20 15520 80
rect 15380 0 15520 20
rect 15680 80 15820 100
rect 15680 20 15720 80
rect 15780 20 15820 80
rect 15680 0 15820 20
rect 15850 80 15990 100
rect 15850 20 15890 80
rect 15950 20 15990 80
rect 15850 0 15990 20
rect 16020 80 16160 100
rect 16020 20 16060 80
rect 16120 20 16160 80
rect 16020 0 16160 20
rect 16190 80 16330 100
rect 16190 20 16230 80
rect 16290 20 16330 80
rect 16190 0 16330 20
rect 16360 80 16500 100
rect 16360 20 16400 80
rect 16460 20 16500 80
rect 16360 0 16500 20
rect 16530 80 16670 100
rect 16530 20 16570 80
rect 16630 20 16670 80
rect 16530 0 16670 20
rect 16700 80 16840 100
rect 16700 20 16740 80
rect 16800 20 16840 80
rect 16700 0 16840 20
rect 16870 80 17010 100
rect 16870 20 16910 80
rect 16970 20 17010 80
rect 16870 0 17010 20
rect 17040 80 17180 100
rect 17040 20 17080 80
rect 17140 20 17180 80
rect 17040 0 17180 20
rect 17210 80 17350 100
rect 17210 20 17250 80
rect 17310 20 17350 80
rect 17210 0 17350 20
rect 17380 80 17520 100
rect 17380 20 17420 80
rect 17480 20 17520 80
rect 17380 0 17520 20
rect 17550 80 17690 100
rect 17550 20 17590 80
rect 17650 20 17690 80
rect 17550 0 17690 20
rect 17720 80 17860 100
rect 17720 20 17760 80
rect 17820 20 17860 80
rect 17720 0 17860 20
rect 17890 80 18030 100
rect 17890 20 17930 80
rect 17990 20 18030 80
rect 17890 0 18030 20
rect 18060 80 18200 100
rect 18060 20 18100 80
rect 18160 20 18200 80
rect 18060 0 18200 20
rect 18230 80 18370 100
rect 18230 20 18270 80
rect 18330 20 18370 80
rect 18230 0 18370 20
rect 18400 80 18540 100
rect 18400 20 18440 80
rect 18500 20 18540 80
rect 18400 0 18540 20
rect 18570 80 18710 100
rect 18570 20 18610 80
rect 18670 20 18710 80
rect 18570 0 18710 20
rect 18740 80 18880 100
rect 18740 20 18780 80
rect 18840 20 18880 80
rect 18740 0 18880 20
rect 18910 80 19050 100
rect 18910 20 18950 80
rect 19010 20 19050 80
rect 18910 0 19050 20
rect 19080 80 19220 100
rect 19080 20 19120 80
rect 19180 20 19220 80
rect 19080 0 19220 20
rect 19250 80 19390 100
rect 19250 20 19290 80
rect 19350 20 19390 80
rect 19250 0 19390 20
rect 19420 80 19560 100
rect 19420 20 19460 80
rect 19520 20 19560 80
rect 19420 0 19560 20
rect 19590 80 19730 100
rect 19590 20 19630 80
rect 19690 20 19730 80
rect 19590 0 19730 20
rect 19760 80 19900 100
rect 19760 20 19800 80
rect 19860 20 19900 80
rect 19760 0 19900 20
rect 19930 80 20070 100
rect 19930 20 19970 80
rect 20030 20 20070 80
rect 19930 0 20070 20
rect 20100 80 20240 100
rect 20100 20 20140 80
rect 20200 20 20240 80
rect 20100 0 20240 20
rect 20270 80 20410 100
rect 20270 20 20310 80
rect 20370 20 20410 80
rect 20270 0 20410 20
rect 20440 80 20580 100
rect 20440 20 20480 80
rect 20540 20 20580 80
rect 20440 0 20580 20
rect 20610 80 20750 100
rect 20610 20 20650 80
rect 20710 20 20750 80
rect 20610 0 20750 20
rect 20780 80 20920 100
rect 20780 20 20820 80
rect 20880 20 20920 80
rect 20780 0 20920 20
rect 20950 80 21090 100
rect 20950 20 20990 80
rect 21050 20 21090 80
rect 20950 0 21090 20
rect 21120 80 21260 100
rect 21120 20 21160 80
rect 21220 20 21260 80
rect 21120 0 21260 20
rect 21290 80 21430 100
rect 21290 20 21330 80
rect 21390 20 21430 80
rect 21290 0 21430 20
rect 21460 80 21600 100
rect 21460 20 21500 80
rect 21560 20 21600 80
rect 21460 0 21600 20
rect 21630 80 21770 100
rect 21630 20 21670 80
rect 21730 20 21770 80
rect 21630 0 21770 20
rect 21800 80 21940 100
rect 21800 20 21840 80
rect 21900 20 21940 80
rect 21800 0 21940 20
rect 21970 80 22110 100
rect 21970 20 22010 80
rect 22070 20 22110 80
rect 21970 0 22110 20
rect 22140 80 22280 100
rect 22140 20 22180 80
rect 22240 20 22280 80
rect 22140 0 22280 20
rect 22310 80 22450 100
rect 22310 20 22350 80
rect 22410 20 22450 80
rect 22310 0 22450 20
rect 22480 80 22620 100
rect 22480 20 22520 80
rect 22580 20 22620 80
rect 22480 0 22620 20
rect 22650 80 22790 100
rect 22650 20 22690 80
rect 22750 20 22790 80
rect 22650 0 22790 20
rect 22820 80 22960 100
rect 22820 20 22860 80
rect 22920 20 22960 80
rect 22820 0 22960 20
rect 22990 80 23130 100
rect 22990 20 23030 80
rect 23090 20 23130 80
rect 22990 0 23130 20
rect 23160 80 23300 100
rect 23160 20 23200 80
rect 23260 20 23300 80
rect 23160 0 23300 20
rect 23330 80 23470 100
rect 23330 20 23370 80
rect 23430 20 23470 80
rect 23330 0 23470 20
rect 23500 80 23640 100
rect 23500 20 23540 80
rect 23600 20 23640 80
rect 23500 0 23640 20
rect 23670 80 23810 100
rect 23670 20 23710 80
rect 23770 20 23810 80
rect 23670 0 23810 20
rect 23840 80 23980 100
rect 23840 20 23880 80
rect 23940 20 23980 80
rect 23840 0 23980 20
rect 24010 80 24150 100
rect 24010 20 24050 80
rect 24110 20 24150 80
rect 24010 0 24150 20
rect 24180 80 24320 100
rect 24180 20 24220 80
rect 24280 20 24320 80
rect 24180 0 24320 20
rect 24350 80 24490 100
rect 24350 20 24390 80
rect 24450 20 24490 80
rect 24350 0 24490 20
rect 24520 80 24660 100
rect 24520 20 24560 80
rect 24620 20 24660 80
rect 24520 0 24660 20
rect 24690 80 24830 100
rect 24690 20 24730 80
rect 24790 20 24830 80
rect 24690 0 24830 20
rect 24860 80 25000 100
rect 24860 20 24900 80
rect 24960 20 25000 80
rect 24860 0 25000 20
rect 25030 80 25170 100
rect 25030 20 25070 80
rect 25130 20 25170 80
rect 25030 0 25170 20
rect 25200 80 25340 100
rect 25200 20 25240 80
rect 25300 20 25340 80
rect 25200 0 25340 20
rect 25370 80 25510 100
rect 25370 20 25410 80
rect 25470 20 25510 80
rect 25370 0 25510 20
rect 25540 80 25680 100
rect 25540 20 25580 80
rect 25640 20 25680 80
rect 25540 0 25680 20
rect 25710 80 25850 100
rect 25710 20 25750 80
rect 25810 20 25850 80
rect 25710 0 25850 20
rect 25880 80 26020 100
rect 25880 20 25920 80
rect 25980 20 26020 80
rect 25880 0 26020 20
rect 26050 80 26190 100
rect 26050 20 26090 80
rect 26150 20 26190 80
rect 26050 0 26190 20
rect 26220 80 26360 100
rect 26220 20 26260 80
rect 26320 20 26360 80
rect 26220 0 26360 20
rect 26390 80 26530 100
rect 26390 20 26430 80
rect 26490 20 26530 80
rect 26390 0 26530 20
rect 26560 80 26700 100
rect 26560 20 26600 80
rect 26660 20 26700 80
rect 26560 0 26700 20
rect 26730 80 26870 100
rect 26730 20 26770 80
rect 26830 20 26870 80
rect 26730 0 26870 20
rect 26900 80 27040 100
rect 26900 20 26940 80
rect 27000 20 27040 80
rect 26900 0 27040 20
rect 27070 80 27210 100
rect 27070 20 27110 80
rect 27170 20 27210 80
rect 27070 0 27210 20
rect 27240 80 27380 100
rect 27240 20 27280 80
rect 27340 20 27380 80
rect 27240 0 27380 20
rect 27410 80 27550 100
rect 27410 20 27450 80
rect 27510 20 27550 80
rect 27410 0 27550 20
rect 27580 80 27720 100
rect 27580 20 27620 80
rect 27680 20 27720 80
rect 27580 0 27720 20
rect 27750 80 27890 100
rect 27750 20 27790 80
rect 27850 20 27890 80
rect 27750 0 27890 20
rect 27920 80 28060 100
rect 27920 20 27960 80
rect 28020 20 28060 80
rect 27920 0 28060 20
rect 28090 80 28230 100
rect 28090 20 28130 80
rect 28190 20 28230 80
rect 28090 0 28230 20
rect 28260 80 28400 100
rect 28260 20 28300 80
rect 28360 20 28400 80
rect 28260 0 28400 20
rect 28430 80 28570 100
rect 28430 20 28470 80
rect 28530 20 28570 80
rect 28430 0 28570 20
rect 28600 80 28740 100
rect 28600 20 28640 80
rect 28700 20 28740 80
rect 28600 0 28740 20
rect 28770 80 28910 100
rect 28770 20 28810 80
rect 28870 20 28910 80
rect 28770 0 28910 20
rect 28940 80 29080 100
rect 28940 20 28980 80
rect 29040 20 29080 80
rect 28940 0 29080 20
rect 29110 80 29250 100
rect 29110 20 29150 80
rect 29210 20 29250 80
rect 29110 0 29250 20
rect 29280 80 29420 100
rect 29280 20 29320 80
rect 29380 20 29420 80
rect 29280 0 29420 20
rect 29450 80 29590 100
rect 29450 20 29490 80
rect 29550 20 29590 80
rect 29450 0 29590 20
rect 29620 80 29760 100
rect 29620 20 29660 80
rect 29720 20 29760 80
rect 29620 0 29760 20
rect 29790 80 29930 100
rect 29790 20 29830 80
rect 29890 20 29930 80
rect 29790 0 29930 20
rect 29960 80 30100 100
rect 29960 20 30000 80
rect 30060 20 30100 80
rect 29960 0 30100 20
rect 30130 80 30270 100
rect 30130 20 30170 80
rect 30230 20 30270 80
rect 30130 0 30270 20
rect 30300 80 30440 100
rect 30300 20 30340 80
rect 30400 20 30440 80
rect 30300 0 30440 20
rect 30470 80 30610 100
rect 30470 20 30510 80
rect 30570 20 30610 80
rect 30470 0 30610 20
rect 30640 80 30780 100
rect 30640 20 30680 80
rect 30740 20 30780 80
rect 30640 0 30780 20
rect 30810 80 30950 100
rect 30810 20 30850 80
rect 30910 20 30950 80
rect 30810 0 30950 20
rect 30980 80 31120 100
rect 30980 20 31020 80
rect 31080 20 31120 80
rect 30980 0 31120 20
rect 31150 80 31290 100
rect 31150 20 31190 80
rect 31250 20 31290 80
rect 31150 0 31290 20
rect 31320 80 31460 100
rect 31320 20 31360 80
rect 31420 20 31460 80
rect 31320 0 31460 20
rect 31490 80 31630 100
rect 31490 20 31530 80
rect 31590 20 31630 80
rect 31490 0 31630 20
rect 31660 80 31800 100
rect 31660 20 31700 80
rect 31760 20 31800 80
rect 31660 0 31800 20
rect 31830 80 31970 100
rect 31830 20 31870 80
rect 31930 20 31970 80
rect 31830 0 31970 20
rect 32000 80 32140 100
rect 32000 20 32040 80
rect 32100 20 32140 80
rect 32000 0 32140 20
rect 32170 80 32310 100
rect 32170 20 32210 80
rect 32270 20 32310 80
rect 32170 0 32310 20
rect 32340 80 32480 100
rect 32340 20 32380 80
rect 32440 20 32480 80
rect 32340 0 32480 20
rect 32510 80 32650 100
rect 32510 20 32550 80
rect 32610 20 32650 80
rect 32510 0 32650 20
rect 32680 80 32820 100
rect 32680 20 32720 80
rect 32780 20 32820 80
rect 32680 0 32820 20
rect 32850 80 32990 100
rect 32850 20 32890 80
rect 32950 20 32990 80
rect 32850 0 32990 20
rect 33020 80 33160 100
rect 33020 20 33060 80
rect 33120 20 33160 80
rect 33020 0 33160 20
rect 33190 80 33330 100
rect 33190 20 33230 80
rect 33290 20 33330 80
rect 33190 0 33330 20
rect 33360 80 33500 100
rect 33360 20 33400 80
rect 33460 20 33500 80
rect 33360 0 33500 20
rect 33530 80 33670 100
rect 33530 20 33570 80
rect 33630 20 33670 80
rect 33530 0 33670 20
rect 33700 80 33840 100
rect 33700 20 33740 80
rect 33800 20 33840 80
rect 33700 0 33840 20
rect 33870 80 34010 100
rect 33870 20 33910 80
rect 33970 20 34010 80
rect 33870 0 34010 20
rect 34040 80 34180 100
rect 34040 20 34080 80
rect 34140 20 34180 80
rect 34040 0 34180 20
rect 34210 80 34350 100
rect 34210 20 34250 80
rect 34310 20 34350 80
rect 34210 0 34350 20
rect 34380 80 34520 100
rect 34380 20 34420 80
rect 34480 20 34520 80
rect 34380 0 34520 20
rect 34550 80 34690 100
rect 34550 20 34590 80
rect 34650 20 34690 80
rect 34550 0 34690 20
rect 34720 80 34860 100
rect 34720 20 34760 80
rect 34820 20 34860 80
rect 34720 0 34860 20
rect 34890 80 35030 100
rect 34890 20 34930 80
rect 34990 20 35030 80
rect 34890 0 35030 20
rect 35060 80 35200 100
rect 35060 20 35100 80
rect 35160 20 35200 80
rect 35060 0 35200 20
rect 35230 80 35370 100
rect 35230 20 35270 80
rect 35330 20 35370 80
rect 35230 0 35370 20
rect 35400 80 35540 100
rect 35400 20 35440 80
rect 35500 20 35540 80
rect 35400 0 35540 20
rect 35570 80 35710 100
rect 35570 20 35610 80
rect 35670 20 35710 80
rect 35570 0 35710 20
rect 35740 80 35880 100
rect 35740 20 35780 80
rect 35840 20 35880 80
rect 35740 0 35880 20
rect 35910 80 36050 100
rect 35910 20 35950 80
rect 36010 20 36050 80
rect 35910 0 36050 20
rect 36080 80 36220 100
rect 36080 20 36120 80
rect 36180 20 36220 80
rect 36080 0 36220 20
rect 36250 80 36390 100
rect 36250 20 36290 80
rect 36350 20 36390 80
rect 36250 0 36390 20
rect 36420 80 36560 100
rect 36420 20 36460 80
rect 36520 20 36560 80
rect 36420 0 36560 20
rect 36590 80 36730 100
rect 36590 20 36630 80
rect 36690 20 36730 80
rect 36590 0 36730 20
rect 36760 80 36900 100
rect 36760 20 36800 80
rect 36860 20 36900 80
rect 36760 0 36900 20
rect 36930 80 37070 100
rect 36930 20 36970 80
rect 37030 20 37070 80
rect 36930 0 37070 20
rect 37100 80 37240 100
rect 37100 20 37140 80
rect 37200 20 37240 80
rect 37100 0 37240 20
rect 37270 80 37410 100
rect 37270 20 37310 80
rect 37370 20 37410 80
rect 37270 0 37410 20
rect 37440 80 37580 100
rect 37440 20 37480 80
rect 37540 20 37580 80
rect 37440 0 37580 20
rect 37610 80 37750 100
rect 37610 20 37650 80
rect 37710 20 37750 80
rect 37610 0 37750 20
rect 37780 80 37920 100
rect 37780 20 37820 80
rect 37880 20 37920 80
rect 37780 0 37920 20
rect 37950 80 38090 100
rect 37950 20 37990 80
rect 38050 20 38090 80
rect 37950 0 38090 20
rect 38120 80 38260 100
rect 38120 20 38160 80
rect 38220 20 38260 80
rect 38120 0 38260 20
rect 38290 80 38430 100
rect 38290 20 38330 80
rect 38390 20 38430 80
rect 38290 0 38430 20
rect 38460 80 38600 100
rect 38460 20 38500 80
rect 38560 20 38600 80
rect 38460 0 38600 20
rect 38630 80 38770 100
rect 38630 20 38670 80
rect 38730 20 38770 80
rect 38630 0 38770 20
rect 38800 80 38940 100
rect 38800 20 38840 80
rect 38900 20 38940 80
rect 38800 0 38940 20
rect 38970 80 39110 100
rect 38970 20 39010 80
rect 39070 20 39110 80
rect 38970 0 39110 20
rect 39140 80 39280 100
rect 39140 20 39180 80
rect 39240 20 39280 80
rect 39140 0 39280 20
rect 39310 80 39450 100
rect 39310 20 39350 80
rect 39410 20 39450 80
rect 39310 0 39450 20
rect 39480 80 39620 100
rect 39480 20 39520 80
rect 39580 20 39620 80
rect 39480 0 39620 20
rect 39650 80 39790 100
rect 39650 20 39690 80
rect 39750 20 39790 80
rect 39650 0 39790 20
rect 39820 80 39960 100
rect 39820 20 39860 80
rect 39920 20 39960 80
rect 39820 0 39960 20
rect 39990 80 40130 100
rect 39990 20 40030 80
rect 40090 20 40130 80
rect 39990 0 40130 20
rect 40160 80 40300 100
rect 40160 20 40200 80
rect 40260 20 40300 80
rect 40160 0 40300 20
rect 40330 80 40470 100
rect 40330 20 40370 80
rect 40430 20 40470 80
rect 40330 0 40470 20
rect 40500 80 40640 100
rect 40500 20 40540 80
rect 40600 20 40640 80
rect 40500 0 40640 20
rect 40670 80 40810 100
rect 40670 20 40710 80
rect 40770 20 40810 80
rect 40670 0 40810 20
rect 40840 80 40980 100
rect 40840 20 40880 80
rect 40940 20 40980 80
rect 40840 0 40980 20
rect 41010 80 41150 100
rect 41010 20 41050 80
rect 41110 20 41150 80
rect 41010 0 41150 20
rect 41180 80 41320 100
rect 41180 20 41220 80
rect 41280 20 41320 80
rect 41180 0 41320 20
rect 41350 80 41490 100
rect 41350 20 41390 80
rect 41450 20 41490 80
rect 41350 0 41490 20
rect 41520 80 41660 100
rect 41520 20 41560 80
rect 41620 20 41660 80
rect 41520 0 41660 20
rect 41690 80 41830 100
rect 41690 20 41730 80
rect 41790 20 41830 80
rect 41690 0 41830 20
rect 41860 80 42000 100
rect 41860 20 41900 80
rect 41960 20 42000 80
rect 41860 0 42000 20
rect 42030 80 42170 100
rect 42030 20 42070 80
rect 42130 20 42170 80
rect 42030 0 42170 20
rect 42200 80 42340 100
rect 42200 20 42240 80
rect 42300 20 42340 80
rect 42200 0 42340 20
rect 42370 80 42510 100
rect 42370 20 42410 80
rect 42470 20 42510 80
rect 42370 0 42510 20
rect 42540 80 42680 100
rect 42540 20 42580 80
rect 42640 20 42680 80
rect 42540 0 42680 20
rect 42710 80 42850 100
rect 42710 20 42750 80
rect 42810 20 42850 80
rect 42710 0 42850 20
rect 42880 80 43020 100
rect 42880 20 42920 80
rect 42980 20 43020 80
rect 42880 0 43020 20
rect 43050 80 43190 100
rect 43050 20 43090 80
rect 43150 20 43190 80
rect 43050 0 43190 20
rect 43220 80 43360 100
rect 43220 20 43260 80
rect 43320 20 43360 80
rect 43220 0 43360 20
rect 43390 80 43530 100
rect 43390 20 43430 80
rect 43490 20 43530 80
rect 43390 0 43530 20
rect 43560 80 43700 100
rect 43560 20 43600 80
rect 43660 20 43700 80
rect 43560 0 43700 20
rect 43730 80 43870 100
rect 43730 20 43770 80
rect 43830 20 43870 80
rect 43730 0 43870 20
rect 43900 80 44040 100
rect 43900 20 43940 80
rect 44000 20 44040 80
rect 43900 0 44040 20
rect 44070 80 44210 100
rect 44070 20 44110 80
rect 44170 20 44210 80
rect 44070 0 44210 20
rect 44240 80 44380 100
rect 44240 20 44280 80
rect 44340 20 44380 80
rect 44240 0 44380 20
rect 44410 80 44550 100
rect 44410 20 44450 80
rect 44510 20 44550 80
rect 44410 0 44550 20
rect 44580 80 44720 100
rect 44580 20 44620 80
rect 44680 20 44720 80
rect 44580 0 44720 20
rect 44750 80 44890 100
rect 44750 20 44790 80
rect 44850 20 44890 80
rect 44750 0 44890 20
rect 44920 80 45060 100
rect 44920 20 44960 80
rect 45020 20 45060 80
rect 44920 0 45060 20
rect 45090 80 45230 100
rect 45090 20 45130 80
rect 45190 20 45230 80
rect 45090 0 45230 20
rect 45260 80 45400 100
rect 45260 20 45300 80
rect 45360 20 45400 80
rect 45260 0 45400 20
rect 45430 80 45570 100
rect 45430 20 45470 80
rect 45530 20 45570 80
rect 45430 0 45570 20
rect 45600 80 45740 100
rect 45600 20 45640 80
rect 45700 20 45740 80
rect 45600 0 45740 20
rect 45770 80 45910 100
rect 45770 20 45810 80
rect 45870 20 45910 80
rect 45770 0 45910 20
rect 45940 80 46080 100
rect 45940 20 45980 80
rect 46040 20 46080 80
rect 45940 0 46080 20
rect 46110 80 46250 100
rect 46110 20 46150 80
rect 46210 20 46250 80
rect 46110 0 46250 20
rect 46280 80 46420 100
rect 46280 20 46320 80
rect 46380 20 46420 80
rect 46280 0 46420 20
rect 46450 80 46590 100
rect 46450 20 46490 80
rect 46550 20 46590 80
rect 46450 0 46590 20
rect 46620 80 46760 100
rect 46620 20 46660 80
rect 46720 20 46760 80
rect 46620 0 46760 20
rect 46790 80 46930 100
rect 46790 20 46830 80
rect 46890 20 46930 80
rect 46790 0 46930 20
rect 46960 80 47100 100
rect 46960 20 47000 80
rect 47060 20 47100 80
rect 46960 0 47100 20
rect 47130 80 47270 100
rect 47130 20 47170 80
rect 47230 20 47270 80
rect 47130 0 47270 20
rect 47300 80 47440 100
rect 47300 20 47340 80
rect 47400 20 47440 80
rect 47300 0 47440 20
rect 47470 80 47610 100
rect 47470 20 47510 80
rect 47570 20 47610 80
rect 47470 0 47610 20
rect 47640 80 47780 100
rect 47640 20 47680 80
rect 47740 20 47780 80
rect 47640 0 47780 20
rect 47810 80 47950 100
rect 47810 20 47850 80
rect 47910 20 47950 80
rect 47810 0 47950 20
rect 47980 80 48120 100
rect 47980 20 48020 80
rect 48080 20 48120 80
rect 47980 0 48120 20
rect 48150 80 48290 100
rect 48150 20 48190 80
rect 48250 20 48290 80
rect 48150 0 48290 20
rect 48320 80 48460 100
rect 48320 20 48360 80
rect 48420 20 48460 80
rect 48320 0 48460 20
rect 48490 80 48630 100
rect 48490 20 48530 80
rect 48590 20 48630 80
rect 48490 0 48630 20
rect 48660 80 48800 100
rect 48660 20 48700 80
rect 48760 20 48800 80
rect 48660 0 48800 20
rect 48830 80 48970 100
rect 48830 20 48870 80
rect 48930 20 48970 80
rect 48830 0 48970 20
rect 49000 80 49140 100
rect 49000 20 49040 80
rect 49100 20 49140 80
rect 49000 0 49140 20
rect 49170 80 49310 100
rect 49170 20 49210 80
rect 49270 20 49310 80
rect 49170 0 49310 20
rect 49340 80 49480 100
rect 49340 20 49380 80
rect 49440 20 49480 80
rect 49340 0 49480 20
rect 49510 80 49650 100
rect 49510 20 49550 80
rect 49610 20 49650 80
rect 49510 0 49650 20
rect 49680 80 49820 100
rect 49680 20 49720 80
rect 49780 20 49820 80
rect 49680 0 49820 20
rect 49850 80 49990 100
rect 49850 20 49890 80
rect 49950 20 49990 80
rect 49850 0 49990 20
rect 50020 80 50160 100
rect 50020 20 50060 80
rect 50120 20 50160 80
rect 50020 0 50160 20
rect 50190 80 50330 100
rect 50190 20 50230 80
rect 50290 20 50330 80
rect 50190 0 50330 20
rect 50360 80 50500 100
rect 50360 20 50400 80
rect 50460 20 50500 80
rect 50360 0 50500 20
rect 50530 80 50670 100
rect 50530 20 50570 80
rect 50630 20 50670 80
rect 50530 0 50670 20
rect 50700 80 50840 100
rect 50700 20 50740 80
rect 50800 20 50840 80
rect 50700 0 50840 20
rect 50870 80 51010 100
rect 50870 20 50910 80
rect 50970 20 51010 80
rect 50870 0 51010 20
rect 51040 80 51180 100
rect 51040 20 51080 80
rect 51140 20 51180 80
rect 51040 0 51180 20
rect 51210 80 51350 100
rect 51210 20 51250 80
rect 51310 20 51350 80
rect 51210 0 51350 20
rect 51380 80 51520 100
rect 51380 20 51420 80
rect 51480 20 51520 80
rect 51380 0 51520 20
rect 51550 80 51690 100
rect 51550 20 51590 80
rect 51650 20 51690 80
rect 51550 0 51690 20
rect 51720 80 51860 100
rect 51720 20 51760 80
rect 51820 20 51860 80
rect 51720 0 51860 20
rect 51890 80 52030 100
rect 51890 20 51930 80
rect 51990 20 52030 80
rect 51890 0 52030 20
rect 52060 80 52200 100
rect 52060 20 52100 80
rect 52160 20 52200 80
rect 52060 0 52200 20
rect 52230 80 52370 100
rect 52230 20 52270 80
rect 52330 20 52370 80
rect 52230 0 52370 20
rect 52400 80 52540 100
rect 52400 20 52440 80
rect 52500 20 52540 80
rect 52400 0 52540 20
rect 52570 80 52710 100
rect 52570 20 52610 80
rect 52670 20 52710 80
rect 52570 0 52710 20
rect 52740 80 52880 100
rect 52740 20 52780 80
rect 52840 20 52880 80
rect 52740 0 52880 20
rect 52910 80 53050 100
rect 52910 20 52950 80
rect 53010 20 53050 80
rect 52910 0 53050 20
rect 53080 80 53220 100
rect 53080 20 53120 80
rect 53180 20 53220 80
rect 53080 0 53220 20
rect 53250 80 53390 100
rect 53250 20 53290 80
rect 53350 20 53390 80
rect 53250 0 53390 20
rect 53420 80 53560 100
rect 53420 20 53460 80
rect 53520 20 53560 80
rect 53420 0 53560 20
rect 53590 80 53730 100
rect 53590 20 53630 80
rect 53690 20 53730 80
rect 53590 0 53730 20
rect 53760 80 53900 100
rect 53760 20 53800 80
rect 53860 20 53900 80
rect 53760 0 53900 20
rect 53930 80 54070 100
rect 53930 20 53970 80
rect 54030 20 54070 80
rect 53930 0 54070 20
rect 54100 80 54240 100
rect 54100 20 54140 80
rect 54200 20 54240 80
rect 54100 0 54240 20
rect 54270 80 54410 100
rect 54270 20 54310 80
rect 54370 20 54410 80
rect 54270 0 54410 20
rect 54440 80 54580 100
rect 54440 20 54480 80
rect 54540 20 54580 80
rect 54440 0 54580 20
rect 54610 80 54750 100
rect 54610 20 54650 80
rect 54710 20 54750 80
rect 54610 0 54750 20
rect 54780 80 54920 100
rect 54780 20 54820 80
rect 54880 20 54920 80
rect 54780 0 54920 20
rect 54950 80 55090 100
rect 54950 20 54990 80
rect 55050 20 55090 80
rect 54950 0 55090 20
rect 55120 80 55260 100
rect 55120 20 55160 80
rect 55220 20 55260 80
rect 55120 0 55260 20
rect 55290 80 55430 100
rect 55290 20 55330 80
rect 55390 20 55430 80
rect 55290 0 55430 20
rect 55460 80 55600 100
rect 55460 20 55500 80
rect 55560 20 55600 80
rect 55460 0 55600 20
rect 55630 80 55770 100
rect 55630 20 55670 80
rect 55730 20 55770 80
rect 55630 0 55770 20
rect 55800 80 55940 100
rect 55800 20 55840 80
rect 55900 20 55940 80
rect 55800 0 55940 20
rect 55970 80 56110 100
rect 55970 20 56010 80
rect 56070 20 56110 80
rect 55970 0 56110 20
rect 56140 80 56280 100
rect 56140 20 56180 80
rect 56240 20 56280 80
rect 56140 0 56280 20
rect 56310 80 56450 100
rect 56310 20 56350 80
rect 56410 20 56450 80
rect 56310 0 56450 20
rect 56480 80 56620 100
rect 56480 20 56520 80
rect 56580 20 56620 80
rect 56480 0 56620 20
rect 56650 80 56790 100
rect 56650 20 56690 80
rect 56750 20 56790 80
rect 56650 0 56790 20
rect 56820 80 56960 100
rect 56820 20 56860 80
rect 56920 20 56960 80
rect 56820 0 56960 20
rect 56990 80 57130 100
rect 56990 20 57030 80
rect 57090 20 57130 80
rect 56990 0 57130 20
rect 57160 80 57300 100
rect 57160 20 57200 80
rect 57260 20 57300 80
rect 57160 0 57300 20
rect 57330 80 57470 100
rect 57330 20 57370 80
rect 57430 20 57470 80
rect 57330 0 57470 20
rect 57500 80 57640 100
rect 57500 20 57540 80
rect 57600 20 57640 80
rect 57500 0 57640 20
rect 57670 80 57810 100
rect 57670 20 57710 80
rect 57770 20 57810 80
rect 57670 0 57810 20
rect 57840 80 57980 100
rect 57840 20 57880 80
rect 57940 20 57980 80
rect 57840 0 57980 20
rect 58010 80 58150 100
rect 58010 20 58050 80
rect 58110 20 58150 80
rect 58010 0 58150 20
rect 58180 80 58320 100
rect 58180 20 58220 80
rect 58280 20 58320 80
rect 58180 0 58320 20
rect 58350 80 58490 100
rect 58350 20 58390 80
rect 58450 20 58490 80
rect 58350 0 58490 20
rect 58520 80 58660 100
rect 58520 20 58560 80
rect 58620 20 58660 80
rect 58520 0 58660 20
rect 58690 80 58830 100
rect 58690 20 58730 80
rect 58790 20 58830 80
rect 58690 0 58830 20
rect 58860 80 59000 100
rect 58860 20 58900 80
rect 58960 20 59000 80
rect 58860 0 59000 20
rect 59030 80 59170 100
rect 59030 20 59070 80
rect 59130 20 59170 80
rect 59030 0 59170 20
rect 59200 80 59340 100
rect 59200 20 59240 80
rect 59300 20 59340 80
rect 59200 0 59340 20
rect -10 -60 130 -40
rect -10 -120 30 -60
rect 90 -120 130 -60
rect -10 -140 130 -120
rect 160 -60 300 -40
rect 160 -120 200 -60
rect 260 -120 300 -60
rect 160 -140 300 -120
rect 110 -670 250 -650
rect 110 -730 150 -670
rect 210 -730 250 -670
rect 110 -770 250 -730
rect 110 -830 150 -770
rect 210 -830 250 -770
rect 110 -850 250 -830
rect 280 -670 420 -650
rect 280 -730 320 -670
rect 380 -730 420 -670
rect 280 -770 420 -730
rect 280 -830 320 -770
rect 380 -830 420 -770
rect 280 -850 420 -830
rect 450 -670 590 -650
rect 450 -730 490 -670
rect 550 -730 590 -670
rect 450 -770 590 -730
rect 450 -830 490 -770
rect 550 -830 590 -770
rect 450 -850 590 -830
rect 620 -670 760 -650
rect 620 -730 660 -670
rect 720 -730 760 -670
rect 620 -770 760 -730
rect 620 -830 660 -770
rect 720 -830 760 -770
rect 620 -850 760 -830
rect 790 -670 930 -650
rect 790 -730 830 -670
rect 890 -730 930 -670
rect 790 -770 930 -730
rect 790 -830 830 -770
rect 890 -830 930 -770
rect 790 -850 930 -830
rect 960 -670 1100 -650
rect 960 -730 1000 -670
rect 1060 -730 1100 -670
rect 960 -770 1100 -730
rect 960 -830 1000 -770
rect 1060 -830 1100 -770
rect 960 -850 1100 -830
rect 1130 -670 1270 -650
rect 1130 -730 1170 -670
rect 1230 -730 1270 -670
rect 1130 -770 1270 -730
rect 1130 -830 1170 -770
rect 1230 -830 1270 -770
rect 1130 -850 1270 -830
rect 1300 -670 1440 -650
rect 1300 -730 1340 -670
rect 1400 -730 1440 -670
rect 1300 -770 1440 -730
rect 1300 -830 1340 -770
rect 1400 -830 1440 -770
rect 1300 -850 1440 -830
rect 1470 -670 1610 -650
rect 1470 -730 1510 -670
rect 1570 -730 1610 -670
rect 1470 -770 1610 -730
rect 1470 -830 1510 -770
rect 1570 -830 1610 -770
rect 1470 -850 1610 -830
rect 1640 -670 1780 -650
rect 1640 -730 1680 -670
rect 1740 -730 1780 -670
rect 1640 -770 1780 -730
rect 1640 -830 1680 -770
rect 1740 -830 1780 -770
rect 1640 -850 1780 -830
rect 1810 -670 1950 -650
rect 1810 -730 1850 -670
rect 1910 -730 1950 -670
rect 1810 -770 1950 -730
rect 1810 -830 1850 -770
rect 1910 -830 1950 -770
rect 1810 -850 1950 -830
rect 1980 -670 2120 -650
rect 1980 -730 2020 -670
rect 2080 -730 2120 -670
rect 1980 -770 2120 -730
rect 1980 -830 2020 -770
rect 2080 -830 2120 -770
rect 1980 -850 2120 -830
rect 2150 -670 2290 -650
rect 2150 -730 2190 -670
rect 2250 -730 2290 -670
rect 2150 -770 2290 -730
rect 2150 -830 2190 -770
rect 2250 -830 2290 -770
rect 2150 -850 2290 -830
rect 2320 -670 2460 -650
rect 2320 -730 2360 -670
rect 2420 -730 2460 -670
rect 2320 -770 2460 -730
rect 2320 -830 2360 -770
rect 2420 -830 2460 -770
rect 2320 -850 2460 -830
rect 2490 -670 2630 -650
rect 2490 -730 2530 -670
rect 2590 -730 2630 -670
rect 2490 -770 2630 -730
rect 2490 -830 2530 -770
rect 2590 -830 2630 -770
rect 2490 -850 2630 -830
rect 2660 -670 2800 -650
rect 2660 -730 2700 -670
rect 2760 -730 2800 -670
rect 2660 -770 2800 -730
rect 2660 -830 2700 -770
rect 2760 -830 2800 -770
rect 2660 -850 2800 -830
rect 2830 -670 2970 -650
rect 2830 -730 2870 -670
rect 2930 -730 2970 -670
rect 2830 -770 2970 -730
rect 2830 -830 2870 -770
rect 2930 -830 2970 -770
rect 2830 -850 2970 -830
rect 3000 -670 3140 -650
rect 3000 -730 3040 -670
rect 3100 -730 3140 -670
rect 3000 -770 3140 -730
rect 3000 -830 3040 -770
rect 3100 -830 3140 -770
rect 3000 -850 3140 -830
rect 3170 -670 3310 -650
rect 3170 -730 3210 -670
rect 3270 -730 3310 -670
rect 3170 -770 3310 -730
rect 3170 -830 3210 -770
rect 3270 -830 3310 -770
rect 3170 -850 3310 -830
rect 3340 -670 3480 -650
rect 3340 -730 3380 -670
rect 3440 -730 3480 -670
rect 3340 -770 3480 -730
rect 3340 -830 3380 -770
rect 3440 -830 3480 -770
rect 3340 -850 3480 -830
rect 3510 -670 3650 -650
rect 3510 -730 3550 -670
rect 3610 -730 3650 -670
rect 3510 -770 3650 -730
rect 3510 -830 3550 -770
rect 3610 -830 3650 -770
rect 3510 -850 3650 -830
rect 3680 -670 3820 -650
rect 3680 -730 3720 -670
rect 3780 -730 3820 -670
rect 3680 -770 3820 -730
rect 3680 -830 3720 -770
rect 3780 -830 3820 -770
rect 3680 -850 3820 -830
rect 3850 -670 3990 -650
rect 3850 -730 3890 -670
rect 3950 -730 3990 -670
rect 3850 -770 3990 -730
rect 3850 -830 3890 -770
rect 3950 -830 3990 -770
rect 3850 -850 3990 -830
rect 4020 -670 4160 -650
rect 4020 -730 4060 -670
rect 4120 -730 4160 -670
rect 4020 -770 4160 -730
rect 4020 -830 4060 -770
rect 4120 -830 4160 -770
rect 4020 -850 4160 -830
rect 4190 -670 4330 -650
rect 4190 -730 4230 -670
rect 4290 -730 4330 -670
rect 4190 -770 4330 -730
rect 4190 -830 4230 -770
rect 4290 -830 4330 -770
rect 4190 -850 4330 -830
rect 4360 -670 4500 -650
rect 4360 -730 4400 -670
rect 4460 -730 4500 -670
rect 4360 -770 4500 -730
rect 4360 -830 4400 -770
rect 4460 -830 4500 -770
rect 4360 -850 4500 -830
rect 4530 -670 4670 -650
rect 4530 -730 4570 -670
rect 4630 -730 4670 -670
rect 4530 -770 4670 -730
rect 4530 -830 4570 -770
rect 4630 -830 4670 -770
rect 4530 -850 4670 -830
rect 4700 -670 4840 -650
rect 4700 -730 4740 -670
rect 4800 -730 4840 -670
rect 4700 -770 4840 -730
rect 4700 -830 4740 -770
rect 4800 -830 4840 -770
rect 4700 -850 4840 -830
rect 4870 -670 5010 -650
rect 4870 -730 4910 -670
rect 4970 -730 5010 -670
rect 4870 -770 5010 -730
rect 4870 -830 4910 -770
rect 4970 -830 5010 -770
rect 4870 -850 5010 -830
rect 5040 -670 5180 -650
rect 5040 -730 5080 -670
rect 5140 -730 5180 -670
rect 5040 -770 5180 -730
rect 5040 -830 5080 -770
rect 5140 -830 5180 -770
rect 5040 -850 5180 -830
rect 5210 -670 5350 -650
rect 5210 -730 5250 -670
rect 5310 -730 5350 -670
rect 5210 -770 5350 -730
rect 5210 -830 5250 -770
rect 5310 -830 5350 -770
rect 5210 -850 5350 -830
rect 5380 -670 5520 -650
rect 5380 -730 5420 -670
rect 5480 -730 5520 -670
rect 5380 -770 5520 -730
rect 5380 -830 5420 -770
rect 5480 -830 5520 -770
rect 5380 -850 5520 -830
rect 5550 -670 5690 -650
rect 5550 -730 5590 -670
rect 5650 -730 5690 -670
rect 5550 -770 5690 -730
rect 5550 -830 5590 -770
rect 5650 -830 5690 -770
rect 5550 -850 5690 -830
rect 5720 -670 5860 -650
rect 5720 -730 5760 -670
rect 5820 -730 5860 -670
rect 5720 -770 5860 -730
rect 5720 -830 5760 -770
rect 5820 -830 5860 -770
rect 5720 -850 5860 -830
rect 5890 -670 6030 -650
rect 5890 -730 5930 -670
rect 5990 -730 6030 -670
rect 5890 -770 6030 -730
rect 5890 -830 5930 -770
rect 5990 -830 6030 -770
rect 5890 -850 6030 -830
rect 6060 -670 6200 -650
rect 6060 -730 6100 -670
rect 6160 -730 6200 -670
rect 6060 -770 6200 -730
rect 6060 -830 6100 -770
rect 6160 -830 6200 -770
rect 6060 -850 6200 -830
rect 6230 -670 6370 -650
rect 6230 -730 6270 -670
rect 6330 -730 6370 -670
rect 6230 -770 6370 -730
rect 6230 -830 6270 -770
rect 6330 -830 6370 -770
rect 6230 -850 6370 -830
rect 6400 -670 6540 -650
rect 6400 -730 6440 -670
rect 6500 -730 6540 -670
rect 6400 -770 6540 -730
rect 6400 -830 6440 -770
rect 6500 -830 6540 -770
rect 6400 -850 6540 -830
rect 6570 -670 6710 -650
rect 6570 -730 6610 -670
rect 6670 -730 6710 -670
rect 6570 -770 6710 -730
rect 6570 -830 6610 -770
rect 6670 -830 6710 -770
rect 6570 -850 6710 -830
rect 6740 -670 6880 -650
rect 6740 -730 6780 -670
rect 6840 -730 6880 -670
rect 6740 -770 6880 -730
rect 6740 -830 6780 -770
rect 6840 -830 6880 -770
rect 6740 -850 6880 -830
rect 6910 -670 7050 -650
rect 6910 -730 6950 -670
rect 7010 -730 7050 -670
rect 6910 -770 7050 -730
rect 6910 -830 6950 -770
rect 7010 -830 7050 -770
rect 6910 -850 7050 -830
rect 7080 -670 7220 -650
rect 7080 -730 7120 -670
rect 7180 -730 7220 -670
rect 7080 -770 7220 -730
rect 7080 -830 7120 -770
rect 7180 -830 7220 -770
rect 7080 -850 7220 -830
rect 7250 -670 7390 -650
rect 7250 -730 7290 -670
rect 7350 -730 7390 -670
rect 7250 -770 7390 -730
rect 7250 -830 7290 -770
rect 7350 -830 7390 -770
rect 7250 -850 7390 -830
rect 7420 -670 7560 -650
rect 7420 -730 7460 -670
rect 7520 -730 7560 -670
rect 7420 -770 7560 -730
rect 7420 -830 7460 -770
rect 7520 -830 7560 -770
rect 7420 -850 7560 -830
rect 7590 -670 7730 -650
rect 7590 -730 7630 -670
rect 7690 -730 7730 -670
rect 7590 -770 7730 -730
rect 7590 -830 7630 -770
rect 7690 -830 7730 -770
rect 7590 -850 7730 -830
rect 7760 -670 7900 -650
rect 7760 -730 7800 -670
rect 7860 -730 7900 -670
rect 7760 -770 7900 -730
rect 7760 -830 7800 -770
rect 7860 -830 7900 -770
rect 7760 -850 7900 -830
rect 7930 -670 8070 -650
rect 7930 -730 7970 -670
rect 8030 -730 8070 -670
rect 7930 -770 8070 -730
rect 7930 -830 7970 -770
rect 8030 -830 8070 -770
rect 7930 -850 8070 -830
rect 8100 -670 8240 -650
rect 8100 -730 8140 -670
rect 8200 -730 8240 -670
rect 8100 -770 8240 -730
rect 8100 -830 8140 -770
rect 8200 -830 8240 -770
rect 8100 -850 8240 -830
rect 8270 -670 8410 -650
rect 8270 -730 8310 -670
rect 8370 -730 8410 -670
rect 8270 -770 8410 -730
rect 8270 -830 8310 -770
rect 8370 -830 8410 -770
rect 8270 -850 8410 -830
rect 8440 -670 8580 -650
rect 8440 -730 8480 -670
rect 8540 -730 8580 -670
rect 8440 -770 8580 -730
rect 8440 -830 8480 -770
rect 8540 -830 8580 -770
rect 8440 -850 8580 -830
rect 8610 -670 8750 -650
rect 8610 -730 8650 -670
rect 8710 -730 8750 -670
rect 8610 -770 8750 -730
rect 8610 -830 8650 -770
rect 8710 -830 8750 -770
rect 8610 -850 8750 -830
rect 8780 -670 8920 -650
rect 8780 -730 8820 -670
rect 8880 -730 8920 -670
rect 8780 -770 8920 -730
rect 8780 -830 8820 -770
rect 8880 -830 8920 -770
rect 8780 -850 8920 -830
rect 8950 -670 9090 -650
rect 8950 -730 8990 -670
rect 9050 -730 9090 -670
rect 8950 -770 9090 -730
rect 8950 -830 8990 -770
rect 9050 -830 9090 -770
rect 8950 -850 9090 -830
rect 9120 -670 9260 -650
rect 9120 -730 9160 -670
rect 9220 -730 9260 -670
rect 9120 -770 9260 -730
rect 9120 -830 9160 -770
rect 9220 -830 9260 -770
rect 9120 -850 9260 -830
rect 9290 -670 9430 -650
rect 9290 -730 9330 -670
rect 9390 -730 9430 -670
rect 9290 -770 9430 -730
rect 9290 -830 9330 -770
rect 9390 -830 9430 -770
rect 9290 -850 9430 -830
rect 9460 -670 9600 -650
rect 9460 -730 9500 -670
rect 9560 -730 9600 -670
rect 9460 -770 9600 -730
rect 9460 -830 9500 -770
rect 9560 -830 9600 -770
rect 9460 -850 9600 -830
rect 9630 -670 9770 -650
rect 9630 -730 9670 -670
rect 9730 -730 9770 -670
rect 9630 -770 9770 -730
rect 9630 -830 9670 -770
rect 9730 -830 9770 -770
rect 9630 -850 9770 -830
rect 9800 -670 9940 -650
rect 9800 -730 9840 -670
rect 9900 -730 9940 -670
rect 9800 -770 9940 -730
rect 9800 -830 9840 -770
rect 9900 -830 9940 -770
rect 9800 -850 9940 -830
rect 9970 -670 10110 -650
rect 9970 -730 10010 -670
rect 10070 -730 10110 -670
rect 9970 -770 10110 -730
rect 9970 -830 10010 -770
rect 10070 -830 10110 -770
rect 9970 -850 10110 -830
rect 10140 -670 10280 -650
rect 10140 -730 10180 -670
rect 10240 -730 10280 -670
rect 10140 -770 10280 -730
rect 10140 -830 10180 -770
rect 10240 -830 10280 -770
rect 10140 -850 10280 -830
rect 10310 -670 10450 -650
rect 10310 -730 10350 -670
rect 10410 -730 10450 -670
rect 10310 -770 10450 -730
rect 10310 -830 10350 -770
rect 10410 -830 10450 -770
rect 10310 -850 10450 -830
rect 10480 -670 10620 -650
rect 10480 -730 10520 -670
rect 10580 -730 10620 -670
rect 10480 -770 10620 -730
rect 10480 -830 10520 -770
rect 10580 -830 10620 -770
rect 10480 -850 10620 -830
rect 10650 -670 10790 -650
rect 10650 -730 10690 -670
rect 10750 -730 10790 -670
rect 10650 -770 10790 -730
rect 10650 -830 10690 -770
rect 10750 -830 10790 -770
rect 10650 -850 10790 -830
rect 10820 -670 10960 -650
rect 10820 -730 10860 -670
rect 10920 -730 10960 -670
rect 10820 -770 10960 -730
rect 10820 -830 10860 -770
rect 10920 -830 10960 -770
rect 10820 -850 10960 -830
rect 10990 -670 11130 -650
rect 10990 -730 11030 -670
rect 11090 -730 11130 -670
rect 10990 -770 11130 -730
rect 10990 -830 11030 -770
rect 11090 -830 11130 -770
rect 10990 -850 11130 -830
rect 11160 -670 11300 -650
rect 11160 -730 11200 -670
rect 11260 -730 11300 -670
rect 11160 -770 11300 -730
rect 11160 -830 11200 -770
rect 11260 -830 11300 -770
rect 11160 -850 11300 -830
rect 11330 -670 11470 -650
rect 11330 -730 11370 -670
rect 11430 -730 11470 -670
rect 11330 -770 11470 -730
rect 11330 -830 11370 -770
rect 11430 -830 11470 -770
rect 11330 -850 11470 -830
rect 11500 -670 11640 -650
rect 11500 -730 11540 -670
rect 11600 -730 11640 -670
rect 11500 -770 11640 -730
rect 11500 -830 11540 -770
rect 11600 -830 11640 -770
rect 11500 -850 11640 -830
rect 11670 -670 11810 -650
rect 11670 -730 11710 -670
rect 11770 -730 11810 -670
rect 11670 -770 11810 -730
rect 11670 -830 11710 -770
rect 11770 -830 11810 -770
rect 11670 -850 11810 -830
rect 11840 -670 11980 -650
rect 11840 -730 11880 -670
rect 11940 -730 11980 -670
rect 11840 -770 11980 -730
rect 11840 -830 11880 -770
rect 11940 -830 11980 -770
rect 11840 -850 11980 -830
rect 12010 -670 12150 -650
rect 12010 -730 12050 -670
rect 12110 -730 12150 -670
rect 12010 -770 12150 -730
rect 12010 -830 12050 -770
rect 12110 -830 12150 -770
rect 12010 -850 12150 -830
rect 12180 -670 12320 -650
rect 12180 -730 12220 -670
rect 12280 -730 12320 -670
rect 12180 -770 12320 -730
rect 12180 -830 12220 -770
rect 12280 -830 12320 -770
rect 12180 -850 12320 -830
rect 12350 -670 12490 -650
rect 12350 -730 12390 -670
rect 12450 -730 12490 -670
rect 12350 -770 12490 -730
rect 12350 -830 12390 -770
rect 12450 -830 12490 -770
rect 12350 -850 12490 -830
rect 12520 -670 12660 -650
rect 12520 -730 12560 -670
rect 12620 -730 12660 -670
rect 12520 -770 12660 -730
rect 12520 -830 12560 -770
rect 12620 -830 12660 -770
rect 12520 -850 12660 -830
rect 12690 -670 12830 -650
rect 12690 -730 12730 -670
rect 12790 -730 12830 -670
rect 12690 -770 12830 -730
rect 12690 -830 12730 -770
rect 12790 -830 12830 -770
rect 12690 -850 12830 -830
rect 12860 -670 13000 -650
rect 12860 -730 12900 -670
rect 12960 -730 13000 -670
rect 12860 -770 13000 -730
rect 12860 -830 12900 -770
rect 12960 -830 13000 -770
rect 12860 -850 13000 -830
rect 13030 -670 13170 -650
rect 13030 -730 13070 -670
rect 13130 -730 13170 -670
rect 13030 -770 13170 -730
rect 13030 -830 13070 -770
rect 13130 -830 13170 -770
rect 13030 -850 13170 -830
rect 13200 -670 13340 -650
rect 13200 -730 13240 -670
rect 13300 -730 13340 -670
rect 13200 -770 13340 -730
rect 13200 -830 13240 -770
rect 13300 -830 13340 -770
rect 13200 -850 13340 -830
rect 13370 -670 13510 -650
rect 13370 -730 13410 -670
rect 13470 -730 13510 -670
rect 13370 -770 13510 -730
rect 13370 -830 13410 -770
rect 13470 -830 13510 -770
rect 13370 -850 13510 -830
rect 13540 -670 13680 -650
rect 13540 -730 13580 -670
rect 13640 -730 13680 -670
rect 13540 -770 13680 -730
rect 13540 -830 13580 -770
rect 13640 -830 13680 -770
rect 13540 -850 13680 -830
rect 13710 -670 13850 -650
rect 13710 -730 13750 -670
rect 13810 -730 13850 -670
rect 13710 -770 13850 -730
rect 13710 -830 13750 -770
rect 13810 -830 13850 -770
rect 13710 -850 13850 -830
rect 13880 -670 14020 -650
rect 13880 -730 13920 -670
rect 13980 -730 14020 -670
rect 13880 -770 14020 -730
rect 13880 -830 13920 -770
rect 13980 -830 14020 -770
rect 13880 -850 14020 -830
rect 14050 -670 14190 -650
rect 14050 -730 14090 -670
rect 14150 -730 14190 -670
rect 14050 -770 14190 -730
rect 14050 -830 14090 -770
rect 14150 -830 14190 -770
rect 14050 -850 14190 -830
rect 14220 -670 14360 -650
rect 14220 -730 14260 -670
rect 14320 -730 14360 -670
rect 14220 -770 14360 -730
rect 14220 -830 14260 -770
rect 14320 -830 14360 -770
rect 14220 -850 14360 -830
rect 14390 -670 14530 -650
rect 14390 -730 14430 -670
rect 14490 -730 14530 -670
rect 14390 -770 14530 -730
rect 14390 -830 14430 -770
rect 14490 -830 14530 -770
rect 14390 -850 14530 -830
rect 14560 -670 14700 -650
rect 14560 -730 14600 -670
rect 14660 -730 14700 -670
rect 14560 -770 14700 -730
rect 14560 -830 14600 -770
rect 14660 -830 14700 -770
rect 14560 -850 14700 -830
rect 14730 -670 14870 -650
rect 14730 -730 14770 -670
rect 14830 -730 14870 -670
rect 14730 -770 14870 -730
rect 14730 -830 14770 -770
rect 14830 -830 14870 -770
rect 14730 -850 14870 -830
rect 14900 -670 15040 -650
rect 14900 -730 14940 -670
rect 15000 -730 15040 -670
rect 14900 -770 15040 -730
rect 14900 -830 14940 -770
rect 15000 -830 15040 -770
rect 14900 -850 15040 -830
rect 15070 -670 15210 -650
rect 15070 -730 15110 -670
rect 15170 -730 15210 -670
rect 15070 -770 15210 -730
rect 15070 -830 15110 -770
rect 15170 -830 15210 -770
rect 15070 -850 15210 -830
rect 15240 -670 15380 -650
rect 15240 -730 15280 -670
rect 15340 -730 15380 -670
rect 15240 -770 15380 -730
rect 15240 -830 15280 -770
rect 15340 -830 15380 -770
rect 15240 -850 15380 -830
rect 15410 -670 15550 -650
rect 15410 -730 15450 -670
rect 15510 -730 15550 -670
rect 15410 -770 15550 -730
rect 15410 -830 15450 -770
rect 15510 -830 15550 -770
rect 15410 -850 15550 -830
rect 15580 -670 15720 -650
rect 15580 -730 15620 -670
rect 15680 -730 15720 -670
rect 15580 -770 15720 -730
rect 15580 -830 15620 -770
rect 15680 -830 15720 -770
rect 15580 -850 15720 -830
rect 15750 -670 15890 -650
rect 15750 -730 15790 -670
rect 15850 -730 15890 -670
rect 15750 -770 15890 -730
rect 15750 -830 15790 -770
rect 15850 -830 15890 -770
rect 15750 -850 15890 -830
rect 15920 -670 16060 -650
rect 15920 -730 15960 -670
rect 16020 -730 16060 -670
rect 15920 -770 16060 -730
rect 15920 -830 15960 -770
rect 16020 -830 16060 -770
rect 15920 -850 16060 -830
rect 16090 -670 16230 -650
rect 16090 -730 16130 -670
rect 16190 -730 16230 -670
rect 16090 -770 16230 -730
rect 16090 -830 16130 -770
rect 16190 -830 16230 -770
rect 16090 -850 16230 -830
rect 16260 -670 16400 -650
rect 16260 -730 16300 -670
rect 16360 -730 16400 -670
rect 16260 -770 16400 -730
rect 16260 -830 16300 -770
rect 16360 -830 16400 -770
rect 16260 -850 16400 -830
rect 16430 -670 16570 -650
rect 16430 -730 16470 -670
rect 16530 -730 16570 -670
rect 16430 -770 16570 -730
rect 16430 -830 16470 -770
rect 16530 -830 16570 -770
rect 16430 -850 16570 -830
rect 16600 -670 16740 -650
rect 16600 -730 16640 -670
rect 16700 -730 16740 -670
rect 16600 -770 16740 -730
rect 16600 -830 16640 -770
rect 16700 -830 16740 -770
rect 16600 -850 16740 -830
rect 16770 -670 16910 -650
rect 16770 -730 16810 -670
rect 16870 -730 16910 -670
rect 16770 -770 16910 -730
rect 16770 -830 16810 -770
rect 16870 -830 16910 -770
rect 16770 -850 16910 -830
rect 16940 -670 17080 -650
rect 16940 -730 16980 -670
rect 17040 -730 17080 -670
rect 16940 -770 17080 -730
rect 16940 -830 16980 -770
rect 17040 -830 17080 -770
rect 16940 -850 17080 -830
rect 17110 -670 17250 -650
rect 17110 -730 17150 -670
rect 17210 -730 17250 -670
rect 17110 -770 17250 -730
rect 17110 -830 17150 -770
rect 17210 -830 17250 -770
rect 17110 -850 17250 -830
rect 17280 -670 17420 -650
rect 17280 -730 17320 -670
rect 17380 -730 17420 -670
rect 17280 -770 17420 -730
rect 17280 -830 17320 -770
rect 17380 -830 17420 -770
rect 17280 -850 17420 -830
rect 17450 -670 17590 -650
rect 17450 -730 17490 -670
rect 17550 -730 17590 -670
rect 17450 -770 17590 -730
rect 17450 -830 17490 -770
rect 17550 -830 17590 -770
rect 17450 -850 17590 -830
rect 17620 -670 17760 -650
rect 17620 -730 17660 -670
rect 17720 -730 17760 -670
rect 17620 -770 17760 -730
rect 17620 -830 17660 -770
rect 17720 -830 17760 -770
rect 17620 -850 17760 -830
rect 17790 -670 17930 -650
rect 17790 -730 17830 -670
rect 17890 -730 17930 -670
rect 17790 -770 17930 -730
rect 17790 -830 17830 -770
rect 17890 -830 17930 -770
rect 17790 -850 17930 -830
rect 17960 -670 18100 -650
rect 17960 -730 18000 -670
rect 18060 -730 18100 -670
rect 17960 -770 18100 -730
rect 17960 -830 18000 -770
rect 18060 -830 18100 -770
rect 17960 -850 18100 -830
rect 18130 -670 18270 -650
rect 18130 -730 18170 -670
rect 18230 -730 18270 -670
rect 18130 -770 18270 -730
rect 18130 -830 18170 -770
rect 18230 -830 18270 -770
rect 18130 -850 18270 -830
rect 18300 -670 18440 -650
rect 18300 -730 18340 -670
rect 18400 -730 18440 -670
rect 18300 -770 18440 -730
rect 18300 -830 18340 -770
rect 18400 -830 18440 -770
rect 18300 -850 18440 -830
rect 18470 -670 18610 -650
rect 18470 -730 18510 -670
rect 18570 -730 18610 -670
rect 18470 -770 18610 -730
rect 18470 -830 18510 -770
rect 18570 -830 18610 -770
rect 18470 -850 18610 -830
rect 18640 -670 18780 -650
rect 18640 -730 18680 -670
rect 18740 -730 18780 -670
rect 18640 -770 18780 -730
rect 18640 -830 18680 -770
rect 18740 -830 18780 -770
rect 18640 -850 18780 -830
rect 18810 -670 18950 -650
rect 18810 -730 18850 -670
rect 18910 -730 18950 -670
rect 18810 -770 18950 -730
rect 18810 -830 18850 -770
rect 18910 -830 18950 -770
rect 18810 -850 18950 -830
rect 18980 -670 19120 -650
rect 18980 -730 19020 -670
rect 19080 -730 19120 -670
rect 18980 -770 19120 -730
rect 18980 -830 19020 -770
rect 19080 -830 19120 -770
rect 18980 -850 19120 -830
rect 19150 -670 19290 -650
rect 19150 -730 19190 -670
rect 19250 -730 19290 -670
rect 19150 -770 19290 -730
rect 19150 -830 19190 -770
rect 19250 -830 19290 -770
rect 19150 -850 19290 -830
rect 19320 -670 19460 -650
rect 19320 -730 19360 -670
rect 19420 -730 19460 -670
rect 19320 -770 19460 -730
rect 19320 -830 19360 -770
rect 19420 -830 19460 -770
rect 19320 -850 19460 -830
rect 19490 -670 19630 -650
rect 19490 -730 19530 -670
rect 19590 -730 19630 -670
rect 19490 -770 19630 -730
rect 19490 -830 19530 -770
rect 19590 -830 19630 -770
rect 19490 -850 19630 -830
rect 19660 -670 19800 -650
rect 19660 -730 19700 -670
rect 19760 -730 19800 -670
rect 19660 -770 19800 -730
rect 19660 -830 19700 -770
rect 19760 -830 19800 -770
rect 19660 -850 19800 -830
rect 19830 -670 19970 -650
rect 19830 -730 19870 -670
rect 19930 -730 19970 -670
rect 19830 -770 19970 -730
rect 19830 -830 19870 -770
rect 19930 -830 19970 -770
rect 19830 -850 19970 -830
rect 20000 -670 20140 -650
rect 20000 -730 20040 -670
rect 20100 -730 20140 -670
rect 20000 -770 20140 -730
rect 20000 -830 20040 -770
rect 20100 -830 20140 -770
rect 20000 -850 20140 -830
rect 20170 -670 20310 -650
rect 20170 -730 20210 -670
rect 20270 -730 20310 -670
rect 20170 -770 20310 -730
rect 20170 -830 20210 -770
rect 20270 -830 20310 -770
rect 20170 -850 20310 -830
rect 20340 -670 20480 -650
rect 20340 -730 20380 -670
rect 20440 -730 20480 -670
rect 20340 -770 20480 -730
rect 20340 -830 20380 -770
rect 20440 -830 20480 -770
rect 20340 -850 20480 -830
rect 20510 -670 20650 -650
rect 20510 -730 20550 -670
rect 20610 -730 20650 -670
rect 20510 -770 20650 -730
rect 20510 -830 20550 -770
rect 20610 -830 20650 -770
rect 20510 -850 20650 -830
rect 20680 -670 20820 -650
rect 20680 -730 20720 -670
rect 20780 -730 20820 -670
rect 20680 -770 20820 -730
rect 20680 -830 20720 -770
rect 20780 -830 20820 -770
rect 20680 -850 20820 -830
rect 20850 -670 20990 -650
rect 20850 -730 20890 -670
rect 20950 -730 20990 -670
rect 20850 -770 20990 -730
rect 20850 -830 20890 -770
rect 20950 -830 20990 -770
rect 20850 -850 20990 -830
rect 21020 -670 21160 -650
rect 21020 -730 21060 -670
rect 21120 -730 21160 -670
rect 21020 -770 21160 -730
rect 21020 -830 21060 -770
rect 21120 -830 21160 -770
rect 21020 -850 21160 -830
rect 21190 -670 21330 -650
rect 21190 -730 21230 -670
rect 21290 -730 21330 -670
rect 21190 -770 21330 -730
rect 21190 -830 21230 -770
rect 21290 -830 21330 -770
rect 21190 -850 21330 -830
rect 21360 -670 21500 -650
rect 21360 -730 21400 -670
rect 21460 -730 21500 -670
rect 21360 -770 21500 -730
rect 21360 -830 21400 -770
rect 21460 -830 21500 -770
rect 21360 -850 21500 -830
rect 21530 -670 21670 -650
rect 21530 -730 21570 -670
rect 21630 -730 21670 -670
rect 21530 -770 21670 -730
rect 21530 -830 21570 -770
rect 21630 -830 21670 -770
rect 21530 -850 21670 -830
rect 21700 -670 21840 -650
rect 21700 -730 21740 -670
rect 21800 -730 21840 -670
rect 21700 -770 21840 -730
rect 21700 -830 21740 -770
rect 21800 -830 21840 -770
rect 21700 -850 21840 -830
rect 21870 -670 22010 -650
rect 21870 -730 21910 -670
rect 21970 -730 22010 -670
rect 21870 -770 22010 -730
rect 21870 -830 21910 -770
rect 21970 -830 22010 -770
rect 21870 -850 22010 -830
rect 22040 -670 22180 -650
rect 22040 -730 22080 -670
rect 22140 -730 22180 -670
rect 22040 -770 22180 -730
rect 22040 -830 22080 -770
rect 22140 -830 22180 -770
rect 22040 -850 22180 -830
rect 22210 -670 22350 -650
rect 22210 -730 22250 -670
rect 22310 -730 22350 -670
rect 22210 -770 22350 -730
rect 22210 -830 22250 -770
rect 22310 -830 22350 -770
rect 22210 -850 22350 -830
rect 22380 -670 22520 -650
rect 22380 -730 22420 -670
rect 22480 -730 22520 -670
rect 22380 -770 22520 -730
rect 22380 -830 22420 -770
rect 22480 -830 22520 -770
rect 22380 -850 22520 -830
rect 22550 -670 22690 -650
rect 22550 -730 22590 -670
rect 22650 -730 22690 -670
rect 22550 -770 22690 -730
rect 22550 -830 22590 -770
rect 22650 -830 22690 -770
rect 22550 -850 22690 -830
rect 22720 -670 22860 -650
rect 22720 -730 22760 -670
rect 22820 -730 22860 -670
rect 22720 -770 22860 -730
rect 22720 -830 22760 -770
rect 22820 -830 22860 -770
rect 22720 -850 22860 -830
rect 22890 -670 23030 -650
rect 22890 -730 22930 -670
rect 22990 -730 23030 -670
rect 22890 -770 23030 -730
rect 22890 -830 22930 -770
rect 22990 -830 23030 -770
rect 22890 -850 23030 -830
rect 23060 -670 23200 -650
rect 23060 -730 23100 -670
rect 23160 -730 23200 -670
rect 23060 -770 23200 -730
rect 23060 -830 23100 -770
rect 23160 -830 23200 -770
rect 23060 -850 23200 -830
rect 23230 -670 23370 -650
rect 23230 -730 23270 -670
rect 23330 -730 23370 -670
rect 23230 -770 23370 -730
rect 23230 -830 23270 -770
rect 23330 -830 23370 -770
rect 23230 -850 23370 -830
rect 23400 -670 23540 -650
rect 23400 -730 23440 -670
rect 23500 -730 23540 -670
rect 23400 -770 23540 -730
rect 23400 -830 23440 -770
rect 23500 -830 23540 -770
rect 23400 -850 23540 -830
rect 23570 -670 23710 -650
rect 23570 -730 23610 -670
rect 23670 -730 23710 -670
rect 23570 -770 23710 -730
rect 23570 -830 23610 -770
rect 23670 -830 23710 -770
rect 23570 -850 23710 -830
rect 23740 -670 23880 -650
rect 23740 -730 23780 -670
rect 23840 -730 23880 -670
rect 23740 -770 23880 -730
rect 23740 -830 23780 -770
rect 23840 -830 23880 -770
rect 23740 -850 23880 -830
rect 23910 -670 24050 -650
rect 23910 -730 23950 -670
rect 24010 -730 24050 -670
rect 23910 -770 24050 -730
rect 23910 -830 23950 -770
rect 24010 -830 24050 -770
rect 23910 -850 24050 -830
rect 24080 -670 24220 -650
rect 24080 -730 24120 -670
rect 24180 -730 24220 -670
rect 24080 -770 24220 -730
rect 24080 -830 24120 -770
rect 24180 -830 24220 -770
rect 24080 -850 24220 -830
rect 24250 -670 24390 -650
rect 24250 -730 24290 -670
rect 24350 -730 24390 -670
rect 24250 -770 24390 -730
rect 24250 -830 24290 -770
rect 24350 -830 24390 -770
rect 24250 -850 24390 -830
rect 24420 -670 24560 -650
rect 24420 -730 24460 -670
rect 24520 -730 24560 -670
rect 24420 -770 24560 -730
rect 24420 -830 24460 -770
rect 24520 -830 24560 -770
rect 24420 -850 24560 -830
rect 24590 -670 24730 -650
rect 24590 -730 24630 -670
rect 24690 -730 24730 -670
rect 24590 -770 24730 -730
rect 24590 -830 24630 -770
rect 24690 -830 24730 -770
rect 24590 -850 24730 -830
rect 24760 -670 24900 -650
rect 24760 -730 24800 -670
rect 24860 -730 24900 -670
rect 24760 -770 24900 -730
rect 24760 -830 24800 -770
rect 24860 -830 24900 -770
rect 24760 -850 24900 -830
rect 24930 -670 25070 -650
rect 24930 -730 24970 -670
rect 25030 -730 25070 -670
rect 24930 -770 25070 -730
rect 24930 -830 24970 -770
rect 25030 -830 25070 -770
rect 24930 -850 25070 -830
rect 25100 -670 25240 -650
rect 25100 -730 25140 -670
rect 25200 -730 25240 -670
rect 25100 -770 25240 -730
rect 25100 -830 25140 -770
rect 25200 -830 25240 -770
rect 25100 -850 25240 -830
rect 25270 -670 25410 -650
rect 25270 -730 25310 -670
rect 25370 -730 25410 -670
rect 25270 -770 25410 -730
rect 25270 -830 25310 -770
rect 25370 -830 25410 -770
rect 25270 -850 25410 -830
rect 25440 -670 25580 -650
rect 25440 -730 25480 -670
rect 25540 -730 25580 -670
rect 25440 -770 25580 -730
rect 25440 -830 25480 -770
rect 25540 -830 25580 -770
rect 25440 -850 25580 -830
rect 25610 -670 25750 -650
rect 25610 -730 25650 -670
rect 25710 -730 25750 -670
rect 25610 -770 25750 -730
rect 25610 -830 25650 -770
rect 25710 -830 25750 -770
rect 25610 -850 25750 -830
rect 25780 -670 25920 -650
rect 25780 -730 25820 -670
rect 25880 -730 25920 -670
rect 25780 -770 25920 -730
rect 25780 -830 25820 -770
rect 25880 -830 25920 -770
rect 25780 -850 25920 -830
rect 25950 -670 26090 -650
rect 25950 -730 25990 -670
rect 26050 -730 26090 -670
rect 25950 -770 26090 -730
rect 25950 -830 25990 -770
rect 26050 -830 26090 -770
rect 25950 -850 26090 -830
rect 26120 -670 26260 -650
rect 26120 -730 26160 -670
rect 26220 -730 26260 -670
rect 26120 -770 26260 -730
rect 26120 -830 26160 -770
rect 26220 -830 26260 -770
rect 26120 -850 26260 -830
rect 26290 -670 26430 -650
rect 26290 -730 26330 -670
rect 26390 -730 26430 -670
rect 26290 -770 26430 -730
rect 26290 -830 26330 -770
rect 26390 -830 26430 -770
rect 26290 -850 26430 -830
rect 26460 -670 26600 -650
rect 26460 -730 26500 -670
rect 26560 -730 26600 -670
rect 26460 -770 26600 -730
rect 26460 -830 26500 -770
rect 26560 -830 26600 -770
rect 26460 -850 26600 -830
rect 26630 -670 26770 -650
rect 26630 -730 26670 -670
rect 26730 -730 26770 -670
rect 26630 -770 26770 -730
rect 26630 -830 26670 -770
rect 26730 -830 26770 -770
rect 26630 -850 26770 -830
rect 26800 -670 26940 -650
rect 26800 -730 26840 -670
rect 26900 -730 26940 -670
rect 26800 -770 26940 -730
rect 26800 -830 26840 -770
rect 26900 -830 26940 -770
rect 26800 -850 26940 -830
rect 26970 -670 27110 -650
rect 26970 -730 27010 -670
rect 27070 -730 27110 -670
rect 26970 -770 27110 -730
rect 26970 -830 27010 -770
rect 27070 -830 27110 -770
rect 26970 -850 27110 -830
rect 27140 -670 27280 -650
rect 27140 -730 27180 -670
rect 27240 -730 27280 -670
rect 27140 -770 27280 -730
rect 27140 -830 27180 -770
rect 27240 -830 27280 -770
rect 27140 -850 27280 -830
rect 27310 -670 27450 -650
rect 27310 -730 27350 -670
rect 27410 -730 27450 -670
rect 27310 -770 27450 -730
rect 27310 -830 27350 -770
rect 27410 -830 27450 -770
rect 27310 -850 27450 -830
rect 27480 -670 27620 -650
rect 27480 -730 27520 -670
rect 27580 -730 27620 -670
rect 27480 -770 27620 -730
rect 27480 -830 27520 -770
rect 27580 -830 27620 -770
rect 27480 -850 27620 -830
rect 27650 -670 27790 -650
rect 27650 -730 27690 -670
rect 27750 -730 27790 -670
rect 27650 -770 27790 -730
rect 27650 -830 27690 -770
rect 27750 -830 27790 -770
rect 27650 -850 27790 -830
rect 27820 -670 27960 -650
rect 27820 -730 27860 -670
rect 27920 -730 27960 -670
rect 27820 -770 27960 -730
rect 27820 -830 27860 -770
rect 27920 -830 27960 -770
rect 27820 -850 27960 -830
rect 27990 -670 28130 -650
rect 27990 -730 28030 -670
rect 28090 -730 28130 -670
rect 27990 -770 28130 -730
rect 27990 -830 28030 -770
rect 28090 -830 28130 -770
rect 27990 -850 28130 -830
rect 28160 -670 28300 -650
rect 28160 -730 28200 -670
rect 28260 -730 28300 -670
rect 28160 -770 28300 -730
rect 28160 -830 28200 -770
rect 28260 -830 28300 -770
rect 28160 -850 28300 -830
rect 28330 -670 28470 -650
rect 28330 -730 28370 -670
rect 28430 -730 28470 -670
rect 28330 -770 28470 -730
rect 28330 -830 28370 -770
rect 28430 -830 28470 -770
rect 28330 -850 28470 -830
rect 28500 -670 28640 -650
rect 28500 -730 28540 -670
rect 28600 -730 28640 -670
rect 28500 -770 28640 -730
rect 28500 -830 28540 -770
rect 28600 -830 28640 -770
rect 28500 -850 28640 -830
rect 28670 -670 28810 -650
rect 28670 -730 28710 -670
rect 28770 -730 28810 -670
rect 28670 -770 28810 -730
rect 28670 -830 28710 -770
rect 28770 -830 28810 -770
rect 28670 -850 28810 -830
rect 28840 -670 28980 -650
rect 28840 -730 28880 -670
rect 28940 -730 28980 -670
rect 28840 -770 28980 -730
rect 28840 -830 28880 -770
rect 28940 -830 28980 -770
rect 28840 -850 28980 -830
rect 29010 -670 29150 -650
rect 29010 -730 29050 -670
rect 29110 -730 29150 -670
rect 29010 -770 29150 -730
rect 29010 -830 29050 -770
rect 29110 -830 29150 -770
rect 29010 -850 29150 -830
rect 29180 -670 29320 -650
rect 29180 -730 29220 -670
rect 29280 -730 29320 -670
rect 29180 -770 29320 -730
rect 29180 -830 29220 -770
rect 29280 -830 29320 -770
rect 29180 -850 29320 -830
rect 29350 -670 29490 -650
rect 29350 -730 29390 -670
rect 29450 -730 29490 -670
rect 29350 -770 29490 -730
rect 29350 -830 29390 -770
rect 29450 -830 29490 -770
rect 29350 -850 29490 -830
rect 29520 -670 29660 -650
rect 29520 -730 29560 -670
rect 29620 -730 29660 -670
rect 29520 -770 29660 -730
rect 29520 -830 29560 -770
rect 29620 -830 29660 -770
rect 29520 -850 29660 -830
rect 29690 -670 29830 -650
rect 29690 -730 29730 -670
rect 29790 -730 29830 -670
rect 29690 -770 29830 -730
rect 29690 -830 29730 -770
rect 29790 -830 29830 -770
rect 29690 -850 29830 -830
rect 29860 -670 30000 -650
rect 29860 -730 29900 -670
rect 29960 -730 30000 -670
rect 29860 -770 30000 -730
rect 29860 -830 29900 -770
rect 29960 -830 30000 -770
rect 29860 -850 30000 -830
rect 30030 -670 30170 -650
rect 30030 -730 30070 -670
rect 30130 -730 30170 -670
rect 30030 -770 30170 -730
rect 30030 -830 30070 -770
rect 30130 -830 30170 -770
rect 30030 -850 30170 -830
rect 30200 -670 30340 -650
rect 30200 -730 30240 -670
rect 30300 -730 30340 -670
rect 30200 -770 30340 -730
rect 30200 -830 30240 -770
rect 30300 -830 30340 -770
rect 30200 -850 30340 -830
rect 30370 -670 30510 -650
rect 30370 -730 30410 -670
rect 30470 -730 30510 -670
rect 30370 -770 30510 -730
rect 30370 -830 30410 -770
rect 30470 -830 30510 -770
rect 30370 -850 30510 -830
rect 30540 -670 30680 -650
rect 30540 -730 30580 -670
rect 30640 -730 30680 -670
rect 30540 -770 30680 -730
rect 30540 -830 30580 -770
rect 30640 -830 30680 -770
rect 30540 -850 30680 -830
rect 30710 -670 30850 -650
rect 30710 -730 30750 -670
rect 30810 -730 30850 -670
rect 30710 -770 30850 -730
rect 30710 -830 30750 -770
rect 30810 -830 30850 -770
rect 30710 -850 30850 -830
rect 30880 -670 31020 -650
rect 30880 -730 30920 -670
rect 30980 -730 31020 -670
rect 30880 -770 31020 -730
rect 30880 -830 30920 -770
rect 30980 -830 31020 -770
rect 30880 -850 31020 -830
rect 31050 -670 31190 -650
rect 31050 -730 31090 -670
rect 31150 -730 31190 -670
rect 31050 -770 31190 -730
rect 31050 -830 31090 -770
rect 31150 -830 31190 -770
rect 31050 -850 31190 -830
rect 31220 -670 31360 -650
rect 31220 -730 31260 -670
rect 31320 -730 31360 -670
rect 31220 -770 31360 -730
rect 31220 -830 31260 -770
rect 31320 -830 31360 -770
rect 31220 -850 31360 -830
rect 31390 -670 31530 -650
rect 31390 -730 31430 -670
rect 31490 -730 31530 -670
rect 31390 -770 31530 -730
rect 31390 -830 31430 -770
rect 31490 -830 31530 -770
rect 31390 -850 31530 -830
rect 31560 -670 31700 -650
rect 31560 -730 31600 -670
rect 31660 -730 31700 -670
rect 31560 -770 31700 -730
rect 31560 -830 31600 -770
rect 31660 -830 31700 -770
rect 31560 -850 31700 -830
rect 31730 -670 31870 -650
rect 31730 -730 31770 -670
rect 31830 -730 31870 -670
rect 31730 -770 31870 -730
rect 31730 -830 31770 -770
rect 31830 -830 31870 -770
rect 31730 -850 31870 -830
rect 31900 -670 32040 -650
rect 31900 -730 31940 -670
rect 32000 -730 32040 -670
rect 31900 -770 32040 -730
rect 31900 -830 31940 -770
rect 32000 -830 32040 -770
rect 31900 -850 32040 -830
rect 32070 -670 32210 -650
rect 32070 -730 32110 -670
rect 32170 -730 32210 -670
rect 32070 -770 32210 -730
rect 32070 -830 32110 -770
rect 32170 -830 32210 -770
rect 32070 -850 32210 -830
rect 32240 -670 32380 -650
rect 32240 -730 32280 -670
rect 32340 -730 32380 -670
rect 32240 -770 32380 -730
rect 32240 -830 32280 -770
rect 32340 -830 32380 -770
rect 32240 -850 32380 -830
rect 32410 -670 32550 -650
rect 32410 -730 32450 -670
rect 32510 -730 32550 -670
rect 32410 -770 32550 -730
rect 32410 -830 32450 -770
rect 32510 -830 32550 -770
rect 32410 -850 32550 -830
rect 32580 -670 32720 -650
rect 32580 -730 32620 -670
rect 32680 -730 32720 -670
rect 32580 -770 32720 -730
rect 32580 -830 32620 -770
rect 32680 -830 32720 -770
rect 32580 -850 32720 -830
rect 32750 -670 32890 -650
rect 32750 -730 32790 -670
rect 32850 -730 32890 -670
rect 32750 -770 32890 -730
rect 32750 -830 32790 -770
rect 32850 -830 32890 -770
rect 32750 -850 32890 -830
rect 32920 -670 33060 -650
rect 32920 -730 32960 -670
rect 33020 -730 33060 -670
rect 32920 -770 33060 -730
rect 32920 -830 32960 -770
rect 33020 -830 33060 -770
rect 32920 -850 33060 -830
rect 33090 -670 33230 -650
rect 33090 -730 33130 -670
rect 33190 -730 33230 -670
rect 33090 -770 33230 -730
rect 33090 -830 33130 -770
rect 33190 -830 33230 -770
rect 33090 -850 33230 -830
rect 33260 -670 33400 -650
rect 33260 -730 33300 -670
rect 33360 -730 33400 -670
rect 33260 -770 33400 -730
rect 33260 -830 33300 -770
rect 33360 -830 33400 -770
rect 33260 -850 33400 -830
rect 33430 -670 33570 -650
rect 33430 -730 33470 -670
rect 33530 -730 33570 -670
rect 33430 -770 33570 -730
rect 33430 -830 33470 -770
rect 33530 -830 33570 -770
rect 33430 -850 33570 -830
rect 33600 -670 33740 -650
rect 33600 -730 33640 -670
rect 33700 -730 33740 -670
rect 33600 -770 33740 -730
rect 33600 -830 33640 -770
rect 33700 -830 33740 -770
rect 33600 -850 33740 -830
rect 33770 -670 33910 -650
rect 33770 -730 33810 -670
rect 33870 -730 33910 -670
rect 33770 -770 33910 -730
rect 33770 -830 33810 -770
rect 33870 -830 33910 -770
rect 33770 -850 33910 -830
rect 33940 -670 34080 -650
rect 33940 -730 33980 -670
rect 34040 -730 34080 -670
rect 33940 -770 34080 -730
rect 33940 -830 33980 -770
rect 34040 -830 34080 -770
rect 33940 -850 34080 -830
rect 34110 -670 34250 -650
rect 34110 -730 34150 -670
rect 34210 -730 34250 -670
rect 34110 -770 34250 -730
rect 34110 -830 34150 -770
rect 34210 -830 34250 -770
rect 34110 -850 34250 -830
rect 34280 -670 34420 -650
rect 34280 -730 34320 -670
rect 34380 -730 34420 -670
rect 34280 -770 34420 -730
rect 34280 -830 34320 -770
rect 34380 -830 34420 -770
rect 34280 -850 34420 -830
rect 34450 -670 34590 -650
rect 34450 -730 34490 -670
rect 34550 -730 34590 -670
rect 34450 -770 34590 -730
rect 34450 -830 34490 -770
rect 34550 -830 34590 -770
rect 34450 -850 34590 -830
rect 34620 -670 34760 -650
rect 34620 -730 34660 -670
rect 34720 -730 34760 -670
rect 34620 -770 34760 -730
rect 34620 -830 34660 -770
rect 34720 -830 34760 -770
rect 34620 -850 34760 -830
rect 34790 -670 34930 -650
rect 34790 -730 34830 -670
rect 34890 -730 34930 -670
rect 34790 -770 34930 -730
rect 34790 -830 34830 -770
rect 34890 -830 34930 -770
rect 34790 -850 34930 -830
rect 34960 -670 35100 -650
rect 34960 -730 35000 -670
rect 35060 -730 35100 -670
rect 34960 -770 35100 -730
rect 34960 -830 35000 -770
rect 35060 -830 35100 -770
rect 34960 -850 35100 -830
rect 35130 -670 35270 -650
rect 35130 -730 35170 -670
rect 35230 -730 35270 -670
rect 35130 -770 35270 -730
rect 35130 -830 35170 -770
rect 35230 -830 35270 -770
rect 35130 -850 35270 -830
rect 35300 -670 35440 -650
rect 35300 -730 35340 -670
rect 35400 -730 35440 -670
rect 35300 -770 35440 -730
rect 35300 -830 35340 -770
rect 35400 -830 35440 -770
rect 35300 -850 35440 -830
rect 35470 -670 35610 -650
rect 35470 -730 35510 -670
rect 35570 -730 35610 -670
rect 35470 -770 35610 -730
rect 35470 -830 35510 -770
rect 35570 -830 35610 -770
rect 35470 -850 35610 -830
rect 35640 -670 35780 -650
rect 35640 -730 35680 -670
rect 35740 -730 35780 -670
rect 35640 -770 35780 -730
rect 35640 -830 35680 -770
rect 35740 -830 35780 -770
rect 35640 -850 35780 -830
rect 35810 -670 35950 -650
rect 35810 -730 35850 -670
rect 35910 -730 35950 -670
rect 35810 -770 35950 -730
rect 35810 -830 35850 -770
rect 35910 -830 35950 -770
rect 35810 -850 35950 -830
rect 35980 -670 36120 -650
rect 35980 -730 36020 -670
rect 36080 -730 36120 -670
rect 35980 -770 36120 -730
rect 35980 -830 36020 -770
rect 36080 -830 36120 -770
rect 35980 -850 36120 -830
rect 36150 -670 36290 -650
rect 36150 -730 36190 -670
rect 36250 -730 36290 -670
rect 36150 -770 36290 -730
rect 36150 -830 36190 -770
rect 36250 -830 36290 -770
rect 36150 -850 36290 -830
rect 36320 -670 36460 -650
rect 36320 -730 36360 -670
rect 36420 -730 36460 -670
rect 36320 -770 36460 -730
rect 36320 -830 36360 -770
rect 36420 -830 36460 -770
rect 36320 -850 36460 -830
rect 36490 -670 36630 -650
rect 36490 -730 36530 -670
rect 36590 -730 36630 -670
rect 36490 -770 36630 -730
rect 36490 -830 36530 -770
rect 36590 -830 36630 -770
rect 36490 -850 36630 -830
rect 36660 -670 36800 -650
rect 36660 -730 36700 -670
rect 36760 -730 36800 -670
rect 36660 -770 36800 -730
rect 36660 -830 36700 -770
rect 36760 -830 36800 -770
rect 36660 -850 36800 -830
rect 36830 -670 36970 -650
rect 36830 -730 36870 -670
rect 36930 -730 36970 -670
rect 36830 -770 36970 -730
rect 36830 -830 36870 -770
rect 36930 -830 36970 -770
rect 36830 -850 36970 -830
rect 37000 -670 37140 -650
rect 37000 -730 37040 -670
rect 37100 -730 37140 -670
rect 37000 -770 37140 -730
rect 37000 -830 37040 -770
rect 37100 -830 37140 -770
rect 37000 -850 37140 -830
rect 37170 -670 37310 -650
rect 37170 -730 37210 -670
rect 37270 -730 37310 -670
rect 37170 -770 37310 -730
rect 37170 -830 37210 -770
rect 37270 -830 37310 -770
rect 37170 -850 37310 -830
rect 37340 -670 37480 -650
rect 37340 -730 37380 -670
rect 37440 -730 37480 -670
rect 37340 -770 37480 -730
rect 37340 -830 37380 -770
rect 37440 -830 37480 -770
rect 37340 -850 37480 -830
rect 37510 -670 37650 -650
rect 37510 -730 37550 -670
rect 37610 -730 37650 -670
rect 37510 -770 37650 -730
rect 37510 -830 37550 -770
rect 37610 -830 37650 -770
rect 37510 -850 37650 -830
rect 37680 -670 37820 -650
rect 37680 -730 37720 -670
rect 37780 -730 37820 -670
rect 37680 -770 37820 -730
rect 37680 -830 37720 -770
rect 37780 -830 37820 -770
rect 37680 -850 37820 -830
rect 37850 -670 37990 -650
rect 37850 -730 37890 -670
rect 37950 -730 37990 -670
rect 37850 -770 37990 -730
rect 37850 -830 37890 -770
rect 37950 -830 37990 -770
rect 37850 -850 37990 -830
rect 38020 -670 38160 -650
rect 38020 -730 38060 -670
rect 38120 -730 38160 -670
rect 38020 -770 38160 -730
rect 38020 -830 38060 -770
rect 38120 -830 38160 -770
rect 38020 -850 38160 -830
rect 38190 -670 38330 -650
rect 38190 -730 38230 -670
rect 38290 -730 38330 -670
rect 38190 -770 38330 -730
rect 38190 -830 38230 -770
rect 38290 -830 38330 -770
rect 38190 -850 38330 -830
rect 38360 -670 38500 -650
rect 38360 -730 38400 -670
rect 38460 -730 38500 -670
rect 38360 -770 38500 -730
rect 38360 -830 38400 -770
rect 38460 -830 38500 -770
rect 38360 -850 38500 -830
rect 38530 -670 38670 -650
rect 38530 -730 38570 -670
rect 38630 -730 38670 -670
rect 38530 -770 38670 -730
rect 38530 -830 38570 -770
rect 38630 -830 38670 -770
rect 38530 -850 38670 -830
rect 38700 -670 38840 -650
rect 38700 -730 38740 -670
rect 38800 -730 38840 -670
rect 38700 -770 38840 -730
rect 38700 -830 38740 -770
rect 38800 -830 38840 -770
rect 38700 -850 38840 -830
rect 38870 -670 39010 -650
rect 38870 -730 38910 -670
rect 38970 -730 39010 -670
rect 38870 -770 39010 -730
rect 38870 -830 38910 -770
rect 38970 -830 39010 -770
rect 38870 -850 39010 -830
rect 39040 -670 39180 -650
rect 39040 -730 39080 -670
rect 39140 -730 39180 -670
rect 39040 -770 39180 -730
rect 39040 -830 39080 -770
rect 39140 -830 39180 -770
rect 39040 -850 39180 -830
rect 39210 -670 39350 -650
rect 39210 -730 39250 -670
rect 39310 -730 39350 -670
rect 39210 -770 39350 -730
rect 39210 -830 39250 -770
rect 39310 -830 39350 -770
rect 39210 -850 39350 -830
rect 39380 -670 39520 -650
rect 39380 -730 39420 -670
rect 39480 -730 39520 -670
rect 39380 -770 39520 -730
rect 39380 -830 39420 -770
rect 39480 -830 39520 -770
rect 39380 -850 39520 -830
rect 39550 -670 39690 -650
rect 39550 -730 39590 -670
rect 39650 -730 39690 -670
rect 39550 -770 39690 -730
rect 39550 -830 39590 -770
rect 39650 -830 39690 -770
rect 39550 -850 39690 -830
rect 39720 -670 39860 -650
rect 39720 -730 39760 -670
rect 39820 -730 39860 -670
rect 39720 -770 39860 -730
rect 39720 -830 39760 -770
rect 39820 -830 39860 -770
rect 39720 -850 39860 -830
rect 39890 -670 40030 -650
rect 39890 -730 39930 -670
rect 39990 -730 40030 -670
rect 39890 -770 40030 -730
rect 39890 -830 39930 -770
rect 39990 -830 40030 -770
rect 39890 -850 40030 -830
rect 40060 -670 40200 -650
rect 40060 -730 40100 -670
rect 40160 -730 40200 -670
rect 40060 -770 40200 -730
rect 40060 -830 40100 -770
rect 40160 -830 40200 -770
rect 40060 -850 40200 -830
rect 40230 -670 40370 -650
rect 40230 -730 40270 -670
rect 40330 -730 40370 -670
rect 40230 -770 40370 -730
rect 40230 -830 40270 -770
rect 40330 -830 40370 -770
rect 40230 -850 40370 -830
rect 40400 -670 40540 -650
rect 40400 -730 40440 -670
rect 40500 -730 40540 -670
rect 40400 -770 40540 -730
rect 40400 -830 40440 -770
rect 40500 -830 40540 -770
rect 40400 -850 40540 -830
rect 40570 -670 40710 -650
rect 40570 -730 40610 -670
rect 40670 -730 40710 -670
rect 40570 -770 40710 -730
rect 40570 -830 40610 -770
rect 40670 -830 40710 -770
rect 40570 -850 40710 -830
rect 40740 -670 40880 -650
rect 40740 -730 40780 -670
rect 40840 -730 40880 -670
rect 40740 -770 40880 -730
rect 40740 -830 40780 -770
rect 40840 -830 40880 -770
rect 40740 -850 40880 -830
rect 40910 -670 41050 -650
rect 40910 -730 40950 -670
rect 41010 -730 41050 -670
rect 40910 -770 41050 -730
rect 40910 -830 40950 -770
rect 41010 -830 41050 -770
rect 40910 -850 41050 -830
rect 41080 -670 41220 -650
rect 41080 -730 41120 -670
rect 41180 -730 41220 -670
rect 41080 -770 41220 -730
rect 41080 -830 41120 -770
rect 41180 -830 41220 -770
rect 41080 -850 41220 -830
rect 41250 -670 41390 -650
rect 41250 -730 41290 -670
rect 41350 -730 41390 -670
rect 41250 -770 41390 -730
rect 41250 -830 41290 -770
rect 41350 -830 41390 -770
rect 41250 -850 41390 -830
rect 41420 -670 41560 -650
rect 41420 -730 41460 -670
rect 41520 -730 41560 -670
rect 41420 -770 41560 -730
rect 41420 -830 41460 -770
rect 41520 -830 41560 -770
rect 41420 -850 41560 -830
rect 41590 -670 41730 -650
rect 41590 -730 41630 -670
rect 41690 -730 41730 -670
rect 41590 -770 41730 -730
rect 41590 -830 41630 -770
rect 41690 -830 41730 -770
rect 41590 -850 41730 -830
rect 41760 -670 41900 -650
rect 41760 -730 41800 -670
rect 41860 -730 41900 -670
rect 41760 -770 41900 -730
rect 41760 -830 41800 -770
rect 41860 -830 41900 -770
rect 41760 -850 41900 -830
rect 41930 -670 42070 -650
rect 41930 -730 41970 -670
rect 42030 -730 42070 -670
rect 41930 -770 42070 -730
rect 41930 -830 41970 -770
rect 42030 -830 42070 -770
rect 41930 -850 42070 -830
rect 42100 -670 42240 -650
rect 42100 -730 42140 -670
rect 42200 -730 42240 -670
rect 42100 -770 42240 -730
rect 42100 -830 42140 -770
rect 42200 -830 42240 -770
rect 42100 -850 42240 -830
rect 42270 -670 42410 -650
rect 42270 -730 42310 -670
rect 42370 -730 42410 -670
rect 42270 -770 42410 -730
rect 42270 -830 42310 -770
rect 42370 -830 42410 -770
rect 42270 -850 42410 -830
rect 42440 -670 42580 -650
rect 42440 -730 42480 -670
rect 42540 -730 42580 -670
rect 42440 -770 42580 -730
rect 42440 -830 42480 -770
rect 42540 -830 42580 -770
rect 42440 -850 42580 -830
rect 42610 -670 42750 -650
rect 42610 -730 42650 -670
rect 42710 -730 42750 -670
rect 42610 -770 42750 -730
rect 42610 -830 42650 -770
rect 42710 -830 42750 -770
rect 42610 -850 42750 -830
rect 42780 -670 42920 -650
rect 42780 -730 42820 -670
rect 42880 -730 42920 -670
rect 42780 -770 42920 -730
rect 42780 -830 42820 -770
rect 42880 -830 42920 -770
rect 42780 -850 42920 -830
rect 42950 -670 43090 -650
rect 42950 -730 42990 -670
rect 43050 -730 43090 -670
rect 42950 -770 43090 -730
rect 42950 -830 42990 -770
rect 43050 -830 43090 -770
rect 42950 -850 43090 -830
rect 43120 -670 43260 -650
rect 43120 -730 43160 -670
rect 43220 -730 43260 -670
rect 43120 -770 43260 -730
rect 43120 -830 43160 -770
rect 43220 -830 43260 -770
rect 43120 -850 43260 -830
rect 43290 -670 43430 -650
rect 43290 -730 43330 -670
rect 43390 -730 43430 -670
rect 43290 -770 43430 -730
rect 43290 -830 43330 -770
rect 43390 -830 43430 -770
rect 43290 -850 43430 -830
rect 43460 -670 43600 -650
rect 43460 -730 43500 -670
rect 43560 -730 43600 -670
rect 43460 -770 43600 -730
rect 43460 -830 43500 -770
rect 43560 -830 43600 -770
rect 43460 -850 43600 -830
rect 43630 -670 43770 -650
rect 43630 -730 43670 -670
rect 43730 -730 43770 -670
rect 43630 -770 43770 -730
rect 43630 -830 43670 -770
rect 43730 -830 43770 -770
rect 43630 -850 43770 -830
rect 43800 -670 43940 -650
rect 43800 -730 43840 -670
rect 43900 -730 43940 -670
rect 43800 -770 43940 -730
rect 43800 -830 43840 -770
rect 43900 -830 43940 -770
rect 43800 -850 43940 -830
rect 43970 -670 44110 -650
rect 43970 -730 44010 -670
rect 44070 -730 44110 -670
rect 43970 -770 44110 -730
rect 43970 -830 44010 -770
rect 44070 -830 44110 -770
rect 43970 -850 44110 -830
rect 44140 -670 44280 -650
rect 44140 -730 44180 -670
rect 44240 -730 44280 -670
rect 44140 -770 44280 -730
rect 44140 -830 44180 -770
rect 44240 -830 44280 -770
rect 44140 -850 44280 -830
rect 44310 -670 44450 -650
rect 44310 -730 44350 -670
rect 44410 -730 44450 -670
rect 44310 -770 44450 -730
rect 44310 -830 44350 -770
rect 44410 -830 44450 -770
rect 44310 -850 44450 -830
rect 44480 -670 44620 -650
rect 44480 -730 44520 -670
rect 44580 -730 44620 -670
rect 44480 -770 44620 -730
rect 44480 -830 44520 -770
rect 44580 -830 44620 -770
rect 44480 -850 44620 -830
rect 44650 -670 44790 -650
rect 44650 -730 44690 -670
rect 44750 -730 44790 -670
rect 44650 -770 44790 -730
rect 44650 -830 44690 -770
rect 44750 -830 44790 -770
rect 44650 -850 44790 -830
rect 44820 -670 44960 -650
rect 44820 -730 44860 -670
rect 44920 -730 44960 -670
rect 44820 -770 44960 -730
rect 44820 -830 44860 -770
rect 44920 -830 44960 -770
rect 44820 -850 44960 -830
rect 44990 -670 45130 -650
rect 44990 -730 45030 -670
rect 45090 -730 45130 -670
rect 44990 -770 45130 -730
rect 44990 -830 45030 -770
rect 45090 -830 45130 -770
rect 44990 -850 45130 -830
rect 45160 -670 45300 -650
rect 45160 -730 45200 -670
rect 45260 -730 45300 -670
rect 45160 -770 45300 -730
rect 45160 -830 45200 -770
rect 45260 -830 45300 -770
rect 45160 -850 45300 -830
rect 45330 -670 45470 -650
rect 45330 -730 45370 -670
rect 45430 -730 45470 -670
rect 45330 -770 45470 -730
rect 45330 -830 45370 -770
rect 45430 -830 45470 -770
rect 45330 -850 45470 -830
rect 45500 -670 45640 -650
rect 45500 -730 45540 -670
rect 45600 -730 45640 -670
rect 45500 -770 45640 -730
rect 45500 -830 45540 -770
rect 45600 -830 45640 -770
rect 45500 -850 45640 -830
rect 45670 -670 45810 -650
rect 45670 -730 45710 -670
rect 45770 -730 45810 -670
rect 45670 -770 45810 -730
rect 45670 -830 45710 -770
rect 45770 -830 45810 -770
rect 45670 -850 45810 -830
rect 45840 -670 45980 -650
rect 45840 -730 45880 -670
rect 45940 -730 45980 -670
rect 45840 -770 45980 -730
rect 45840 -830 45880 -770
rect 45940 -830 45980 -770
rect 45840 -850 45980 -830
rect 46010 -670 46150 -650
rect 46010 -730 46050 -670
rect 46110 -730 46150 -670
rect 46010 -770 46150 -730
rect 46010 -830 46050 -770
rect 46110 -830 46150 -770
rect 46010 -850 46150 -830
rect 46180 -670 46320 -650
rect 46180 -730 46220 -670
rect 46280 -730 46320 -670
rect 46180 -770 46320 -730
rect 46180 -830 46220 -770
rect 46280 -830 46320 -770
rect 46180 -850 46320 -830
rect 46350 -670 46490 -650
rect 46350 -730 46390 -670
rect 46450 -730 46490 -670
rect 46350 -770 46490 -730
rect 46350 -830 46390 -770
rect 46450 -830 46490 -770
rect 46350 -850 46490 -830
rect 46520 -670 46660 -650
rect 46520 -730 46560 -670
rect 46620 -730 46660 -670
rect 46520 -770 46660 -730
rect 46520 -830 46560 -770
rect 46620 -830 46660 -770
rect 46520 -850 46660 -830
rect 46690 -670 46830 -650
rect 46690 -730 46730 -670
rect 46790 -730 46830 -670
rect 46690 -770 46830 -730
rect 46690 -830 46730 -770
rect 46790 -830 46830 -770
rect 46690 -850 46830 -830
rect 46860 -670 47000 -650
rect 46860 -730 46900 -670
rect 46960 -730 47000 -670
rect 46860 -770 47000 -730
rect 46860 -830 46900 -770
rect 46960 -830 47000 -770
rect 46860 -850 47000 -830
rect 47030 -670 47170 -650
rect 47030 -730 47070 -670
rect 47130 -730 47170 -670
rect 47030 -770 47170 -730
rect 47030 -830 47070 -770
rect 47130 -830 47170 -770
rect 47030 -850 47170 -830
rect 47200 -670 47340 -650
rect 47200 -730 47240 -670
rect 47300 -730 47340 -670
rect 47200 -770 47340 -730
rect 47200 -830 47240 -770
rect 47300 -830 47340 -770
rect 47200 -850 47340 -830
rect 47370 -670 47510 -650
rect 47370 -730 47410 -670
rect 47470 -730 47510 -670
rect 47370 -770 47510 -730
rect 47370 -830 47410 -770
rect 47470 -830 47510 -770
rect 47370 -850 47510 -830
rect 47540 -670 47680 -650
rect 47540 -730 47580 -670
rect 47640 -730 47680 -670
rect 47540 -770 47680 -730
rect 47540 -830 47580 -770
rect 47640 -830 47680 -770
rect 47540 -850 47680 -830
rect 47710 -670 47850 -650
rect 47710 -730 47750 -670
rect 47810 -730 47850 -670
rect 47710 -770 47850 -730
rect 47710 -830 47750 -770
rect 47810 -830 47850 -770
rect 47710 -850 47850 -830
rect 47880 -670 48020 -650
rect 47880 -730 47920 -670
rect 47980 -730 48020 -670
rect 47880 -770 48020 -730
rect 47880 -830 47920 -770
rect 47980 -830 48020 -770
rect 47880 -850 48020 -830
rect 48050 -670 48190 -650
rect 48050 -730 48090 -670
rect 48150 -730 48190 -670
rect 48050 -770 48190 -730
rect 48050 -830 48090 -770
rect 48150 -830 48190 -770
rect 48050 -850 48190 -830
rect 48220 -670 48360 -650
rect 48220 -730 48260 -670
rect 48320 -730 48360 -670
rect 48220 -770 48360 -730
rect 48220 -830 48260 -770
rect 48320 -830 48360 -770
rect 48220 -850 48360 -830
rect 48390 -670 48530 -650
rect 48390 -730 48430 -670
rect 48490 -730 48530 -670
rect 48390 -770 48530 -730
rect 48390 -830 48430 -770
rect 48490 -830 48530 -770
rect 48390 -850 48530 -830
rect 48560 -670 48700 -650
rect 48560 -730 48600 -670
rect 48660 -730 48700 -670
rect 48560 -770 48700 -730
rect 48560 -830 48600 -770
rect 48660 -830 48700 -770
rect 48560 -850 48700 -830
rect 48730 -670 48870 -650
rect 48730 -730 48770 -670
rect 48830 -730 48870 -670
rect 48730 -770 48870 -730
rect 48730 -830 48770 -770
rect 48830 -830 48870 -770
rect 48730 -850 48870 -830
rect 48900 -670 49040 -650
rect 48900 -730 48940 -670
rect 49000 -730 49040 -670
rect 48900 -770 49040 -730
rect 48900 -830 48940 -770
rect 49000 -830 49040 -770
rect 48900 -850 49040 -830
rect 49070 -670 49210 -650
rect 49070 -730 49110 -670
rect 49170 -730 49210 -670
rect 49070 -770 49210 -730
rect 49070 -830 49110 -770
rect 49170 -830 49210 -770
rect 49070 -850 49210 -830
rect 49240 -670 49380 -650
rect 49240 -730 49280 -670
rect 49340 -730 49380 -670
rect 49240 -770 49380 -730
rect 49240 -830 49280 -770
rect 49340 -830 49380 -770
rect 49240 -850 49380 -830
rect 49410 -670 49550 -650
rect 49410 -730 49450 -670
rect 49510 -730 49550 -670
rect 49410 -770 49550 -730
rect 49410 -830 49450 -770
rect 49510 -830 49550 -770
rect 49410 -850 49550 -830
rect 49580 -670 49720 -650
rect 49580 -730 49620 -670
rect 49680 -730 49720 -670
rect 49580 -770 49720 -730
rect 49580 -830 49620 -770
rect 49680 -830 49720 -770
rect 49580 -850 49720 -830
rect 49750 -670 49890 -650
rect 49750 -730 49790 -670
rect 49850 -730 49890 -670
rect 49750 -770 49890 -730
rect 49750 -830 49790 -770
rect 49850 -830 49890 -770
rect 49750 -850 49890 -830
rect 49920 -670 50060 -650
rect 49920 -730 49960 -670
rect 50020 -730 50060 -670
rect 49920 -770 50060 -730
rect 49920 -830 49960 -770
rect 50020 -830 50060 -770
rect 49920 -850 50060 -830
rect 50090 -670 50230 -650
rect 50090 -730 50130 -670
rect 50190 -730 50230 -670
rect 50090 -770 50230 -730
rect 50090 -830 50130 -770
rect 50190 -830 50230 -770
rect 50090 -850 50230 -830
rect 50260 -670 50400 -650
rect 50260 -730 50300 -670
rect 50360 -730 50400 -670
rect 50260 -770 50400 -730
rect 50260 -830 50300 -770
rect 50360 -830 50400 -770
rect 50260 -850 50400 -830
rect 50430 -670 50570 -650
rect 50430 -730 50470 -670
rect 50530 -730 50570 -670
rect 50430 -770 50570 -730
rect 50430 -830 50470 -770
rect 50530 -830 50570 -770
rect 50430 -850 50570 -830
rect 50600 -670 50740 -650
rect 50600 -730 50640 -670
rect 50700 -730 50740 -670
rect 50600 -770 50740 -730
rect 50600 -830 50640 -770
rect 50700 -830 50740 -770
rect 50600 -850 50740 -830
rect 50770 -670 50910 -650
rect 50770 -730 50810 -670
rect 50870 -730 50910 -670
rect 50770 -770 50910 -730
rect 50770 -830 50810 -770
rect 50870 -830 50910 -770
rect 50770 -850 50910 -830
rect 50940 -670 51080 -650
rect 50940 -730 50980 -670
rect 51040 -730 51080 -670
rect 50940 -770 51080 -730
rect 50940 -830 50980 -770
rect 51040 -830 51080 -770
rect 50940 -850 51080 -830
rect 51110 -670 51250 -650
rect 51110 -730 51150 -670
rect 51210 -730 51250 -670
rect 51110 -770 51250 -730
rect 51110 -830 51150 -770
rect 51210 -830 51250 -770
rect 51110 -850 51250 -830
rect 51280 -670 51420 -650
rect 51280 -730 51320 -670
rect 51380 -730 51420 -670
rect 51280 -770 51420 -730
rect 51280 -830 51320 -770
rect 51380 -830 51420 -770
rect 51280 -850 51420 -830
rect 51450 -670 51590 -650
rect 51450 -730 51490 -670
rect 51550 -730 51590 -670
rect 51450 -770 51590 -730
rect 51450 -830 51490 -770
rect 51550 -830 51590 -770
rect 51450 -850 51590 -830
rect 51620 -670 51760 -650
rect 51620 -730 51660 -670
rect 51720 -730 51760 -670
rect 51620 -770 51760 -730
rect 51620 -830 51660 -770
rect 51720 -830 51760 -770
rect 51620 -850 51760 -830
rect 51790 -670 51930 -650
rect 51790 -730 51830 -670
rect 51890 -730 51930 -670
rect 51790 -770 51930 -730
rect 51790 -830 51830 -770
rect 51890 -830 51930 -770
rect 51790 -850 51930 -830
rect 51960 -670 52100 -650
rect 51960 -730 52000 -670
rect 52060 -730 52100 -670
rect 51960 -770 52100 -730
rect 51960 -830 52000 -770
rect 52060 -830 52100 -770
rect 51960 -850 52100 -830
rect 52130 -670 52270 -650
rect 52130 -730 52170 -670
rect 52230 -730 52270 -670
rect 52130 -770 52270 -730
rect 52130 -830 52170 -770
rect 52230 -830 52270 -770
rect 52130 -850 52270 -830
rect 52300 -670 52440 -650
rect 52300 -730 52340 -670
rect 52400 -730 52440 -670
rect 52300 -770 52440 -730
rect 52300 -830 52340 -770
rect 52400 -830 52440 -770
rect 52300 -850 52440 -830
rect 52470 -670 52610 -650
rect 52470 -730 52510 -670
rect 52570 -730 52610 -670
rect 52470 -770 52610 -730
rect 52470 -830 52510 -770
rect 52570 -830 52610 -770
rect 52470 -850 52610 -830
rect 52640 -670 52780 -650
rect 52640 -730 52680 -670
rect 52740 -730 52780 -670
rect 52640 -770 52780 -730
rect 52640 -830 52680 -770
rect 52740 -830 52780 -770
rect 52640 -850 52780 -830
rect 52810 -670 52950 -650
rect 52810 -730 52850 -670
rect 52910 -730 52950 -670
rect 52810 -770 52950 -730
rect 52810 -830 52850 -770
rect 52910 -830 52950 -770
rect 52810 -850 52950 -830
rect 52980 -670 53120 -650
rect 52980 -730 53020 -670
rect 53080 -730 53120 -670
rect 52980 -770 53120 -730
rect 52980 -830 53020 -770
rect 53080 -830 53120 -770
rect 52980 -850 53120 -830
rect 53150 -670 53290 -650
rect 53150 -730 53190 -670
rect 53250 -730 53290 -670
rect 53150 -770 53290 -730
rect 53150 -830 53190 -770
rect 53250 -830 53290 -770
rect 53150 -850 53290 -830
rect 53320 -670 53460 -650
rect 53320 -730 53360 -670
rect 53420 -730 53460 -670
rect 53320 -770 53460 -730
rect 53320 -830 53360 -770
rect 53420 -830 53460 -770
rect 53320 -850 53460 -830
rect 53490 -670 53630 -650
rect 53490 -730 53530 -670
rect 53590 -730 53630 -670
rect 53490 -770 53630 -730
rect 53490 -830 53530 -770
rect 53590 -830 53630 -770
rect 53490 -850 53630 -830
rect 53660 -670 53800 -650
rect 53660 -730 53700 -670
rect 53760 -730 53800 -670
rect 53660 -770 53800 -730
rect 53660 -830 53700 -770
rect 53760 -830 53800 -770
rect 53660 -850 53800 -830
rect 53830 -670 53970 -650
rect 53830 -730 53870 -670
rect 53930 -730 53970 -670
rect 53830 -770 53970 -730
rect 53830 -830 53870 -770
rect 53930 -830 53970 -770
rect 53830 -850 53970 -830
rect 54000 -670 54140 -650
rect 54000 -730 54040 -670
rect 54100 -730 54140 -670
rect 54000 -770 54140 -730
rect 54000 -830 54040 -770
rect 54100 -830 54140 -770
rect 54000 -850 54140 -830
rect 54170 -670 54310 -650
rect 54170 -730 54210 -670
rect 54270 -730 54310 -670
rect 54170 -770 54310 -730
rect 54170 -830 54210 -770
rect 54270 -830 54310 -770
rect 54170 -850 54310 -830
rect 54340 -670 54480 -650
rect 54340 -730 54380 -670
rect 54440 -730 54480 -670
rect 54340 -770 54480 -730
rect 54340 -830 54380 -770
rect 54440 -830 54480 -770
rect 54340 -850 54480 -830
rect 54510 -670 54650 -650
rect 54510 -730 54550 -670
rect 54610 -730 54650 -670
rect 54510 -770 54650 -730
rect 54510 -830 54550 -770
rect 54610 -830 54650 -770
rect 54510 -850 54650 -830
rect 54680 -670 54820 -650
rect 54680 -730 54720 -670
rect 54780 -730 54820 -670
rect 54680 -770 54820 -730
rect 54680 -830 54720 -770
rect 54780 -830 54820 -770
rect 54680 -850 54820 -830
rect 54850 -670 54990 -650
rect 54850 -730 54890 -670
rect 54950 -730 54990 -670
rect 54850 -770 54990 -730
rect 54850 -830 54890 -770
rect 54950 -830 54990 -770
rect 54850 -850 54990 -830
rect 55020 -670 55160 -650
rect 55020 -730 55060 -670
rect 55120 -730 55160 -670
rect 55020 -770 55160 -730
rect 55020 -830 55060 -770
rect 55120 -830 55160 -770
rect 55020 -850 55160 -830
rect 55190 -670 55330 -650
rect 55190 -730 55230 -670
rect 55290 -730 55330 -670
rect 55190 -770 55330 -730
rect 55190 -830 55230 -770
rect 55290 -830 55330 -770
rect 55190 -850 55330 -830
rect 55360 -670 55500 -650
rect 55360 -730 55400 -670
rect 55460 -730 55500 -670
rect 55360 -770 55500 -730
rect 55360 -830 55400 -770
rect 55460 -830 55500 -770
rect 55360 -850 55500 -830
rect 55530 -670 55670 -650
rect 55530 -730 55570 -670
rect 55630 -730 55670 -670
rect 55530 -770 55670 -730
rect 55530 -830 55570 -770
rect 55630 -830 55670 -770
rect 55530 -850 55670 -830
rect 55700 -670 55840 -650
rect 55700 -730 55740 -670
rect 55800 -730 55840 -670
rect 55700 -770 55840 -730
rect 55700 -830 55740 -770
rect 55800 -830 55840 -770
rect 55700 -850 55840 -830
rect 55870 -670 56010 -650
rect 55870 -730 55910 -670
rect 55970 -730 56010 -670
rect 55870 -770 56010 -730
rect 55870 -830 55910 -770
rect 55970 -830 56010 -770
rect 55870 -850 56010 -830
rect 56040 -670 56180 -650
rect 56040 -730 56080 -670
rect 56140 -730 56180 -670
rect 56040 -770 56180 -730
rect 56040 -830 56080 -770
rect 56140 -830 56180 -770
rect 56040 -850 56180 -830
rect 56210 -670 56350 -650
rect 56210 -730 56250 -670
rect 56310 -730 56350 -670
rect 56210 -770 56350 -730
rect 56210 -830 56250 -770
rect 56310 -830 56350 -770
rect 56210 -850 56350 -830
rect 56380 -670 56520 -650
rect 56380 -730 56420 -670
rect 56480 -730 56520 -670
rect 56380 -770 56520 -730
rect 56380 -830 56420 -770
rect 56480 -830 56520 -770
rect 56380 -850 56520 -830
rect 56550 -670 56690 -650
rect 56550 -730 56590 -670
rect 56650 -730 56690 -670
rect 56550 -770 56690 -730
rect 56550 -830 56590 -770
rect 56650 -830 56690 -770
rect 56550 -850 56690 -830
rect 56720 -670 56860 -650
rect 56720 -730 56760 -670
rect 56820 -730 56860 -670
rect 56720 -770 56860 -730
rect 56720 -830 56760 -770
rect 56820 -830 56860 -770
rect 56720 -850 56860 -830
rect 56890 -670 57030 -650
rect 56890 -730 56930 -670
rect 56990 -730 57030 -670
rect 56890 -770 57030 -730
rect 56890 -830 56930 -770
rect 56990 -830 57030 -770
rect 56890 -850 57030 -830
rect 57060 -670 57200 -650
rect 57060 -730 57100 -670
rect 57160 -730 57200 -670
rect 57060 -770 57200 -730
rect 57060 -830 57100 -770
rect 57160 -830 57200 -770
rect 57060 -850 57200 -830
rect 57230 -670 57370 -650
rect 57230 -730 57270 -670
rect 57330 -730 57370 -670
rect 57230 -770 57370 -730
rect 57230 -830 57270 -770
rect 57330 -830 57370 -770
rect 57230 -850 57370 -830
rect 57400 -670 57540 -650
rect 57400 -730 57440 -670
rect 57500 -730 57540 -670
rect 57400 -770 57540 -730
rect 57400 -830 57440 -770
rect 57500 -830 57540 -770
rect 57400 -850 57540 -830
rect 57570 -670 57710 -650
rect 57570 -730 57610 -670
rect 57670 -730 57710 -670
rect 57570 -770 57710 -730
rect 57570 -830 57610 -770
rect 57670 -830 57710 -770
rect 57570 -850 57710 -830
rect 57740 -670 57880 -650
rect 57740 -730 57780 -670
rect 57840 -730 57880 -670
rect 57740 -770 57880 -730
rect 57740 -830 57780 -770
rect 57840 -830 57880 -770
rect 57740 -850 57880 -830
rect 57910 -670 58050 -650
rect 57910 -730 57950 -670
rect 58010 -730 58050 -670
rect 57910 -770 58050 -730
rect 57910 -830 57950 -770
rect 58010 -830 58050 -770
rect 57910 -850 58050 -830
rect 58080 -670 58220 -650
rect 58080 -730 58120 -670
rect 58180 -730 58220 -670
rect 58080 -770 58220 -730
rect 58080 -830 58120 -770
rect 58180 -830 58220 -770
rect 58080 -850 58220 -830
rect 58250 -670 58390 -650
rect 58250 -730 58290 -670
rect 58350 -730 58390 -670
rect 58250 -770 58390 -730
rect 58250 -830 58290 -770
rect 58350 -830 58390 -770
rect 58250 -850 58390 -830
rect 58420 -670 58560 -650
rect 58420 -730 58460 -670
rect 58520 -730 58560 -670
rect 58420 -770 58560 -730
rect 58420 -830 58460 -770
rect 58520 -830 58560 -770
rect 58420 -850 58560 -830
rect 58590 -670 58730 -650
rect 58590 -730 58630 -670
rect 58690 -730 58730 -670
rect 58590 -770 58730 -730
rect 58590 -830 58630 -770
rect 58690 -830 58730 -770
rect 58590 -850 58730 -830
rect 58760 -670 58900 -650
rect 58760 -730 58800 -670
rect 58860 -730 58900 -670
rect 58760 -770 58900 -730
rect 58760 -830 58800 -770
rect 58860 -830 58900 -770
rect 58760 -850 58900 -830
rect 58930 -670 59070 -650
rect 58930 -730 58970 -670
rect 59030 -730 59070 -670
rect 58930 -770 59070 -730
rect 58930 -830 58970 -770
rect 59030 -830 59070 -770
rect 58930 -850 59070 -830
rect 59100 -670 59240 -650
rect 59100 -730 59140 -670
rect 59200 -730 59240 -670
rect 59100 -770 59240 -730
rect 59100 -830 59140 -770
rect 59200 -830 59240 -770
rect 59100 -850 59240 -830
rect 59270 -670 59410 -650
rect 59270 -730 59310 -670
rect 59370 -730 59410 -670
rect 59270 -770 59410 -730
rect 59270 -830 59310 -770
rect 59370 -830 59410 -770
rect 59270 -850 59410 -830
rect 59440 -670 59580 -650
rect 59440 -730 59480 -670
rect 59540 -730 59580 -670
rect 59440 -770 59580 -730
rect 59440 -830 59480 -770
rect 59540 -830 59580 -770
rect 59440 -850 59580 -830
rect 59610 -670 59750 -650
rect 59610 -730 59650 -670
rect 59710 -730 59750 -670
rect 59610 -770 59750 -730
rect 59610 -830 59650 -770
rect 59710 -830 59750 -770
rect 59610 -850 59750 -830
rect 59780 -670 59920 -650
rect 59780 -730 59820 -670
rect 59880 -730 59920 -670
rect 59780 -770 59920 -730
rect 59780 -830 59820 -770
rect 59880 -830 59920 -770
rect 59780 -850 59920 -830
rect 59950 -670 60090 -650
rect 59950 -730 59990 -670
rect 60050 -730 60090 -670
rect 59950 -770 60090 -730
rect 59950 -830 59990 -770
rect 60050 -830 60090 -770
rect 59950 -850 60090 -830
rect 60120 -670 60260 -650
rect 60120 -730 60160 -670
rect 60220 -730 60260 -670
rect 60120 -770 60260 -730
rect 60120 -830 60160 -770
rect 60220 -830 60260 -770
rect 60120 -850 60260 -830
rect 60290 -670 60430 -650
rect 60290 -730 60330 -670
rect 60390 -730 60430 -670
rect 60290 -770 60430 -730
rect 60290 -830 60330 -770
rect 60390 -830 60430 -770
rect 60290 -850 60430 -830
rect 60460 -670 60600 -650
rect 60460 -730 60500 -670
rect 60560 -730 60600 -670
rect 60460 -770 60600 -730
rect 60460 -830 60500 -770
rect 60560 -830 60600 -770
rect 60460 -850 60600 -830
rect 60630 -670 60770 -650
rect 60630 -730 60670 -670
rect 60730 -730 60770 -670
rect 60630 -770 60770 -730
rect 60630 -830 60670 -770
rect 60730 -830 60770 -770
rect 60630 -850 60770 -830
rect 60800 -670 60940 -650
rect 60800 -730 60840 -670
rect 60900 -730 60940 -670
rect 60800 -770 60940 -730
rect 60800 -830 60840 -770
rect 60900 -830 60940 -770
rect 60800 -850 60940 -830
rect 60970 -670 61110 -650
rect 60970 -730 61010 -670
rect 61070 -730 61110 -670
rect 60970 -770 61110 -730
rect 60970 -830 61010 -770
rect 61070 -830 61110 -770
rect 60970 -850 61110 -830
rect 61140 -670 61280 -650
rect 61140 -730 61180 -670
rect 61240 -730 61280 -670
rect 61140 -770 61280 -730
rect 61140 -830 61180 -770
rect 61240 -830 61280 -770
rect 61140 -850 61280 -830
rect 61310 -670 61450 -650
rect 61310 -730 61350 -670
rect 61410 -730 61450 -670
rect 61310 -770 61450 -730
rect 61310 -830 61350 -770
rect 61410 -830 61450 -770
rect 61310 -850 61450 -830
rect 61480 -670 61620 -650
rect 61480 -730 61520 -670
rect 61580 -730 61620 -670
rect 61480 -770 61620 -730
rect 61480 -830 61520 -770
rect 61580 -830 61620 -770
rect 61480 -850 61620 -830
rect 61650 -670 61790 -650
rect 61650 -730 61690 -670
rect 61750 -730 61790 -670
rect 61650 -770 61790 -730
rect 61650 -830 61690 -770
rect 61750 -830 61790 -770
rect 61650 -850 61790 -830
rect 61820 -670 61960 -650
rect 61820 -730 61860 -670
rect 61920 -730 61960 -670
rect 61820 -770 61960 -730
rect 61820 -830 61860 -770
rect 61920 -830 61960 -770
rect 61820 -850 61960 -830
rect 61990 -670 62130 -650
rect 61990 -730 62030 -670
rect 62090 -730 62130 -670
rect 61990 -770 62130 -730
rect 61990 -830 62030 -770
rect 62090 -830 62130 -770
rect 61990 -850 62130 -830
rect 62160 -670 62300 -650
rect 62160 -730 62200 -670
rect 62260 -730 62300 -670
rect 62160 -770 62300 -730
rect 62160 -830 62200 -770
rect 62260 -830 62300 -770
rect 62160 -850 62300 -830
rect 62330 -670 62470 -650
rect 62330 -730 62370 -670
rect 62430 -730 62470 -670
rect 62330 -770 62470 -730
rect 62330 -830 62370 -770
rect 62430 -830 62470 -770
rect 62330 -850 62470 -830
rect 62500 -670 62640 -650
rect 62500 -730 62540 -670
rect 62600 -730 62640 -670
rect 62500 -770 62640 -730
rect 62500 -830 62540 -770
rect 62600 -830 62640 -770
rect 62500 -850 62640 -830
rect 62670 -670 62810 -650
rect 62670 -730 62710 -670
rect 62770 -730 62810 -670
rect 62670 -770 62810 -730
rect 62670 -830 62710 -770
rect 62770 -830 62810 -770
rect 62670 -850 62810 -830
rect 62840 -670 62980 -650
rect 62840 -730 62880 -670
rect 62940 -730 62980 -670
rect 62840 -770 62980 -730
rect 62840 -830 62880 -770
rect 62940 -830 62980 -770
rect 62840 -850 62980 -830
rect 63010 -670 63150 -650
rect 63010 -730 63050 -670
rect 63110 -730 63150 -670
rect 63010 -770 63150 -730
rect 63010 -830 63050 -770
rect 63110 -830 63150 -770
rect 63010 -850 63150 -830
rect 63180 -670 63320 -650
rect 63180 -730 63220 -670
rect 63280 -730 63320 -670
rect 63180 -770 63320 -730
rect 63180 -830 63220 -770
rect 63280 -830 63320 -770
rect 63180 -850 63320 -830
rect 63350 -670 63490 -650
rect 63350 -730 63390 -670
rect 63450 -730 63490 -670
rect 63350 -770 63490 -730
rect 63350 -830 63390 -770
rect 63450 -830 63490 -770
rect 63350 -850 63490 -830
rect 63520 -670 63660 -650
rect 63520 -730 63560 -670
rect 63620 -730 63660 -670
rect 63520 -770 63660 -730
rect 63520 -830 63560 -770
rect 63620 -830 63660 -770
rect 63520 -850 63660 -830
rect 63690 -670 63830 -650
rect 63690 -730 63730 -670
rect 63790 -730 63830 -670
rect 63690 -770 63830 -730
rect 63690 -830 63730 -770
rect 63790 -830 63830 -770
rect 63690 -850 63830 -830
rect 63860 -670 64000 -650
rect 63860 -730 63900 -670
rect 63960 -730 64000 -670
rect 63860 -770 64000 -730
rect 63860 -830 63900 -770
rect 63960 -830 64000 -770
rect 63860 -850 64000 -830
rect 64030 -670 64170 -650
rect 64030 -730 64070 -670
rect 64130 -730 64170 -670
rect 64030 -770 64170 -730
rect 64030 -830 64070 -770
rect 64130 -830 64170 -770
rect 64030 -850 64170 -830
rect 64200 -670 64340 -650
rect 64200 -730 64240 -670
rect 64300 -730 64340 -670
rect 64200 -770 64340 -730
rect 64200 -830 64240 -770
rect 64300 -830 64340 -770
rect 64200 -850 64340 -830
rect 64370 -670 64510 -650
rect 64370 -730 64410 -670
rect 64470 -730 64510 -670
rect 64370 -770 64510 -730
rect 64370 -830 64410 -770
rect 64470 -830 64510 -770
rect 64370 -850 64510 -830
rect 64540 -670 64680 -650
rect 64540 -730 64580 -670
rect 64640 -730 64680 -670
rect 64540 -770 64680 -730
rect 64540 -830 64580 -770
rect 64640 -830 64680 -770
rect 64540 -850 64680 -830
rect 64710 -670 64850 -650
rect 64710 -730 64750 -670
rect 64810 -730 64850 -670
rect 64710 -770 64850 -730
rect 64710 -830 64750 -770
rect 64810 -830 64850 -770
rect 64710 -850 64850 -830
rect 64880 -670 65020 -650
rect 64880 -730 64920 -670
rect 64980 -730 65020 -670
rect 64880 -770 65020 -730
rect 64880 -830 64920 -770
rect 64980 -830 65020 -770
rect 64880 -850 65020 -830
rect 65050 -670 65190 -650
rect 65050 -730 65090 -670
rect 65150 -730 65190 -670
rect 65050 -770 65190 -730
rect 65050 -830 65090 -770
rect 65150 -830 65190 -770
rect 65050 -850 65190 -830
rect 65220 -670 65360 -650
rect 65220 -730 65260 -670
rect 65320 -730 65360 -670
rect 65220 -770 65360 -730
rect 65220 -830 65260 -770
rect 65320 -830 65360 -770
rect 65220 -850 65360 -830
rect 65390 -670 65530 -650
rect 65390 -730 65430 -670
rect 65490 -730 65530 -670
rect 65390 -770 65530 -730
rect 65390 -830 65430 -770
rect 65490 -830 65530 -770
rect 65390 -850 65530 -830
rect 65560 -670 65700 -650
rect 65560 -730 65600 -670
rect 65660 -730 65700 -670
rect 65560 -770 65700 -730
rect 65560 -830 65600 -770
rect 65660 -830 65700 -770
rect 65560 -850 65700 -830
rect 65730 -670 65870 -650
rect 65730 -730 65770 -670
rect 65830 -730 65870 -670
rect 65730 -770 65870 -730
rect 65730 -830 65770 -770
rect 65830 -830 65870 -770
rect 65730 -850 65870 -830
rect 65900 -670 66040 -650
rect 65900 -730 65940 -670
rect 66000 -730 66040 -670
rect 65900 -770 66040 -730
rect 65900 -830 65940 -770
rect 66000 -830 66040 -770
rect 65900 -850 66040 -830
rect 66070 -670 66210 -650
rect 66070 -730 66110 -670
rect 66170 -730 66210 -670
rect 66070 -770 66210 -730
rect 66070 -830 66110 -770
rect 66170 -830 66210 -770
rect 66070 -850 66210 -830
rect 66240 -670 66380 -650
rect 66240 -730 66280 -670
rect 66340 -730 66380 -670
rect 66240 -770 66380 -730
rect 66240 -830 66280 -770
rect 66340 -830 66380 -770
rect 66240 -850 66380 -830
rect 66410 -670 66550 -650
rect 66410 -730 66450 -670
rect 66510 -730 66550 -670
rect 66410 -770 66550 -730
rect 66410 -830 66450 -770
rect 66510 -830 66550 -770
rect 66410 -850 66550 -830
rect 66580 -670 66720 -650
rect 66580 -730 66620 -670
rect 66680 -730 66720 -670
rect 66580 -770 66720 -730
rect 66580 -830 66620 -770
rect 66680 -830 66720 -770
rect 66580 -850 66720 -830
rect 66750 -670 66890 -650
rect 66750 -730 66790 -670
rect 66850 -730 66890 -670
rect 66750 -770 66890 -730
rect 66750 -830 66790 -770
rect 66850 -830 66890 -770
rect 66750 -850 66890 -830
rect 66920 -670 67060 -650
rect 66920 -730 66960 -670
rect 67020 -730 67060 -670
rect 66920 -770 67060 -730
rect 66920 -830 66960 -770
rect 67020 -830 67060 -770
rect 66920 -850 67060 -830
rect 67090 -670 67230 -650
rect 67090 -730 67130 -670
rect 67190 -730 67230 -670
rect 67090 -770 67230 -730
rect 67090 -830 67130 -770
rect 67190 -830 67230 -770
rect 67090 -850 67230 -830
rect 67260 -670 67400 -650
rect 67260 -730 67300 -670
rect 67360 -730 67400 -670
rect 67260 -770 67400 -730
rect 67260 -830 67300 -770
rect 67360 -830 67400 -770
rect 67260 -850 67400 -830
rect 67430 -670 67570 -650
rect 67430 -730 67470 -670
rect 67530 -730 67570 -670
rect 67430 -770 67570 -730
rect 67430 -830 67470 -770
rect 67530 -830 67570 -770
rect 67430 -850 67570 -830
rect 67600 -670 67740 -650
rect 67600 -730 67640 -670
rect 67700 -730 67740 -670
rect 67600 -770 67740 -730
rect 67600 -830 67640 -770
rect 67700 -830 67740 -770
rect 67600 -850 67740 -830
rect 67770 -670 67910 -650
rect 67770 -730 67810 -670
rect 67870 -730 67910 -670
rect 67770 -770 67910 -730
rect 67770 -830 67810 -770
rect 67870 -830 67910 -770
rect 67770 -850 67910 -830
rect 67940 -670 68080 -650
rect 67940 -730 67980 -670
rect 68040 -730 68080 -670
rect 67940 -770 68080 -730
rect 67940 -830 67980 -770
rect 68040 -830 68080 -770
rect 67940 -850 68080 -830
rect 68110 -670 68250 -650
rect 68110 -730 68150 -670
rect 68210 -730 68250 -670
rect 68110 -770 68250 -730
rect 68110 -830 68150 -770
rect 68210 -830 68250 -770
rect 68110 -850 68250 -830
rect 68280 -670 68420 -650
rect 68280 -730 68320 -670
rect 68380 -730 68420 -670
rect 68280 -770 68420 -730
rect 68280 -830 68320 -770
rect 68380 -830 68420 -770
rect 68280 -850 68420 -830
rect 68450 -670 68590 -650
rect 68450 -730 68490 -670
rect 68550 -730 68590 -670
rect 68450 -770 68590 -730
rect 68450 -830 68490 -770
rect 68550 -830 68590 -770
rect 68450 -850 68590 -830
rect 68620 -670 68760 -650
rect 68620 -730 68660 -670
rect 68720 -730 68760 -670
rect 68620 -770 68760 -730
rect 68620 -830 68660 -770
rect 68720 -830 68760 -770
rect 68620 -850 68760 -830
rect 68790 -670 68930 -650
rect 68790 -730 68830 -670
rect 68890 -730 68930 -670
rect 68790 -770 68930 -730
rect 68790 -830 68830 -770
rect 68890 -830 68930 -770
rect 68790 -850 68930 -830
rect 68960 -670 69100 -650
rect 68960 -730 69000 -670
rect 69060 -730 69100 -670
rect 68960 -770 69100 -730
rect 68960 -830 69000 -770
rect 69060 -830 69100 -770
rect 68960 -850 69100 -830
rect 69130 -670 69270 -650
rect 69130 -730 69170 -670
rect 69230 -730 69270 -670
rect 69130 -770 69270 -730
rect 69130 -830 69170 -770
rect 69230 -830 69270 -770
rect 69130 -850 69270 -830
rect 69300 -670 69440 -650
rect 69300 -730 69340 -670
rect 69400 -730 69440 -670
rect 69300 -770 69440 -730
rect 69300 -830 69340 -770
rect 69400 -830 69440 -770
rect 69300 -850 69440 -830
rect 69470 -670 69610 -650
rect 69470 -730 69510 -670
rect 69570 -730 69610 -670
rect 69470 -770 69610 -730
rect 69470 -830 69510 -770
rect 69570 -830 69610 -770
rect 69470 -850 69610 -830
rect 69640 -670 69780 -650
rect 69640 -730 69680 -670
rect 69740 -730 69780 -670
rect 69640 -770 69780 -730
rect 69640 -830 69680 -770
rect 69740 -830 69780 -770
rect 69640 -850 69780 -830
rect 69810 -670 69950 -650
rect 69810 -730 69850 -670
rect 69910 -730 69950 -670
rect 69810 -770 69950 -730
rect 69810 -830 69850 -770
rect 69910 -830 69950 -770
rect 69810 -850 69950 -830
rect 69980 -670 70120 -650
rect 69980 -730 70020 -670
rect 70080 -730 70120 -670
rect 69980 -770 70120 -730
rect 69980 -830 70020 -770
rect 70080 -830 70120 -770
rect 69980 -850 70120 -830
rect 70150 -670 70290 -650
rect 70150 -730 70190 -670
rect 70250 -730 70290 -670
rect 70150 -770 70290 -730
rect 70150 -830 70190 -770
rect 70250 -830 70290 -770
rect 70150 -850 70290 -830
rect 70320 -670 70460 -650
rect 70320 -730 70360 -670
rect 70420 -730 70460 -670
rect 70320 -770 70460 -730
rect 70320 -830 70360 -770
rect 70420 -830 70460 -770
rect 70320 -850 70460 -830
rect 70490 -670 70630 -650
rect 70490 -730 70530 -670
rect 70590 -730 70630 -670
rect 70490 -770 70630 -730
rect 70490 -830 70530 -770
rect 70590 -830 70630 -770
rect 70490 -850 70630 -830
rect 70660 -670 70800 -650
rect 70660 -730 70700 -670
rect 70760 -730 70800 -670
rect 70660 -770 70800 -730
rect 70660 -830 70700 -770
rect 70760 -830 70800 -770
rect 70660 -850 70800 -830
rect 70830 -670 70970 -650
rect 70830 -730 70870 -670
rect 70930 -730 70970 -670
rect 70830 -770 70970 -730
rect 70830 -830 70870 -770
rect 70930 -830 70970 -770
rect 70830 -850 70970 -830
rect 71000 -670 71140 -650
rect 71000 -730 71040 -670
rect 71100 -730 71140 -670
rect 71000 -770 71140 -730
rect 71000 -830 71040 -770
rect 71100 -830 71140 -770
rect 71000 -850 71140 -830
rect 71170 -670 71310 -650
rect 71170 -730 71210 -670
rect 71270 -730 71310 -670
rect 71170 -770 71310 -730
rect 71170 -830 71210 -770
rect 71270 -830 71310 -770
rect 71170 -850 71310 -830
rect 71340 -670 71480 -650
rect 71340 -730 71380 -670
rect 71440 -730 71480 -670
rect 71340 -770 71480 -730
rect 71340 -830 71380 -770
rect 71440 -830 71480 -770
rect 71340 -850 71480 -830
rect 71510 -670 71650 -650
rect 71510 -730 71550 -670
rect 71610 -730 71650 -670
rect 71510 -770 71650 -730
rect 71510 -830 71550 -770
rect 71610 -830 71650 -770
rect 71510 -850 71650 -830
rect 71680 -670 71820 -650
rect 71680 -730 71720 -670
rect 71780 -730 71820 -670
rect 71680 -770 71820 -730
rect 71680 -830 71720 -770
rect 71780 -830 71820 -770
rect 71680 -850 71820 -830
rect 71850 -670 71990 -650
rect 71850 -730 71890 -670
rect 71950 -730 71990 -670
rect 71850 -770 71990 -730
rect 71850 -830 71890 -770
rect 71950 -830 71990 -770
rect 71850 -850 71990 -830
rect 72020 -670 72160 -650
rect 72020 -730 72060 -670
rect 72120 -730 72160 -670
rect 72020 -770 72160 -730
rect 72020 -830 72060 -770
rect 72120 -830 72160 -770
rect 72020 -850 72160 -830
rect 72190 -670 72330 -650
rect 72190 -730 72230 -670
rect 72290 -730 72330 -670
rect 72190 -770 72330 -730
rect 72190 -830 72230 -770
rect 72290 -830 72330 -770
rect 72190 -850 72330 -830
rect 72360 -670 72500 -650
rect 72360 -730 72400 -670
rect 72460 -730 72500 -670
rect 72360 -770 72500 -730
rect 72360 -830 72400 -770
rect 72460 -830 72500 -770
rect 72360 -850 72500 -830
rect 72530 -670 72670 -650
rect 72530 -730 72570 -670
rect 72630 -730 72670 -670
rect 72530 -770 72670 -730
rect 72530 -830 72570 -770
rect 72630 -830 72670 -770
rect 72530 -850 72670 -830
rect 72700 -670 72840 -650
rect 72700 -730 72740 -670
rect 72800 -730 72840 -670
rect 72700 -770 72840 -730
rect 72700 -830 72740 -770
rect 72800 -830 72840 -770
rect 72700 -850 72840 -830
rect 72870 -670 73010 -650
rect 72870 -730 72910 -670
rect 72970 -730 73010 -670
rect 72870 -770 73010 -730
rect 72870 -830 72910 -770
rect 72970 -830 73010 -770
rect 72870 -850 73010 -830
rect 73040 -670 73180 -650
rect 73040 -730 73080 -670
rect 73140 -730 73180 -670
rect 73040 -770 73180 -730
rect 73040 -830 73080 -770
rect 73140 -830 73180 -770
rect 73040 -850 73180 -830
rect 73210 -670 73350 -650
rect 73210 -730 73250 -670
rect 73310 -730 73350 -670
rect 73210 -770 73350 -730
rect 73210 -830 73250 -770
rect 73310 -830 73350 -770
rect 73210 -850 73350 -830
rect 73380 -670 73520 -650
rect 73380 -730 73420 -670
rect 73480 -730 73520 -670
rect 73380 -770 73520 -730
rect 73380 -830 73420 -770
rect 73480 -830 73520 -770
rect 73380 -850 73520 -830
rect 73550 -670 73690 -650
rect 73550 -730 73590 -670
rect 73650 -730 73690 -670
rect 73550 -770 73690 -730
rect 73550 -830 73590 -770
rect 73650 -830 73690 -770
rect 73550 -850 73690 -830
rect 73720 -670 73860 -650
rect 73720 -730 73760 -670
rect 73820 -730 73860 -670
rect 73720 -770 73860 -730
rect 73720 -830 73760 -770
rect 73820 -830 73860 -770
rect 73720 -850 73860 -830
rect 73890 -670 74030 -650
rect 73890 -730 73930 -670
rect 73990 -730 74030 -670
rect 73890 -770 74030 -730
rect 73890 -830 73930 -770
rect 73990 -830 74030 -770
rect 73890 -850 74030 -830
rect 74060 -670 74200 -650
rect 74060 -730 74100 -670
rect 74160 -730 74200 -670
rect 74060 -770 74200 -730
rect 74060 -830 74100 -770
rect 74160 -830 74200 -770
rect 74060 -850 74200 -830
rect 74230 -670 74370 -650
rect 74230 -730 74270 -670
rect 74330 -730 74370 -670
rect 74230 -770 74370 -730
rect 74230 -830 74270 -770
rect 74330 -830 74370 -770
rect 74230 -850 74370 -830
rect 74400 -670 74540 -650
rect 74400 -730 74440 -670
rect 74500 -730 74540 -670
rect 74400 -770 74540 -730
rect 74400 -830 74440 -770
rect 74500 -830 74540 -770
rect 74400 -850 74540 -830
rect 74570 -670 74710 -650
rect 74570 -730 74610 -670
rect 74670 -730 74710 -670
rect 74570 -770 74710 -730
rect 74570 -830 74610 -770
rect 74670 -830 74710 -770
rect 74570 -850 74710 -830
rect 74740 -670 74880 -650
rect 74740 -730 74780 -670
rect 74840 -730 74880 -670
rect 74740 -770 74880 -730
rect 74740 -830 74780 -770
rect 74840 -830 74880 -770
rect 74740 -850 74880 -830
rect 74910 -670 75050 -650
rect 74910 -730 74950 -670
rect 75010 -730 75050 -670
rect 74910 -770 75050 -730
rect 74910 -830 74950 -770
rect 75010 -830 75050 -770
rect 74910 -850 75050 -830
rect 75080 -670 75220 -650
rect 75080 -730 75120 -670
rect 75180 -730 75220 -670
rect 75080 -770 75220 -730
rect 75080 -830 75120 -770
rect 75180 -830 75220 -770
rect 75080 -850 75220 -830
rect 75250 -670 75390 -650
rect 75250 -730 75290 -670
rect 75350 -730 75390 -670
rect 75250 -770 75390 -730
rect 75250 -830 75290 -770
rect 75350 -830 75390 -770
rect 75250 -850 75390 -830
rect 75420 -670 75560 -650
rect 75420 -730 75460 -670
rect 75520 -730 75560 -670
rect 75420 -770 75560 -730
rect 75420 -830 75460 -770
rect 75520 -830 75560 -770
rect 75420 -850 75560 -830
rect 75590 -670 75730 -650
rect 75590 -730 75630 -670
rect 75690 -730 75730 -670
rect 75590 -770 75730 -730
rect 75590 -830 75630 -770
rect 75690 -830 75730 -770
rect 75590 -850 75730 -830
rect 75760 -670 75900 -650
rect 75760 -730 75800 -670
rect 75860 -730 75900 -670
rect 75760 -770 75900 -730
rect 75760 -830 75800 -770
rect 75860 -830 75900 -770
rect 75760 -850 75900 -830
rect 75930 -670 76070 -650
rect 75930 -730 75970 -670
rect 76030 -730 76070 -670
rect 75930 -770 76070 -730
rect 75930 -830 75970 -770
rect 76030 -830 76070 -770
rect 75930 -850 76070 -830
rect 76100 -670 76240 -650
rect 76100 -730 76140 -670
rect 76200 -730 76240 -670
rect 76100 -770 76240 -730
rect 76100 -830 76140 -770
rect 76200 -830 76240 -770
rect 76100 -850 76240 -830
rect 76270 -670 76410 -650
rect 76270 -730 76310 -670
rect 76370 -730 76410 -670
rect 76270 -770 76410 -730
rect 76270 -830 76310 -770
rect 76370 -830 76410 -770
rect 76270 -850 76410 -830
rect 76440 -670 76580 -650
rect 76440 -730 76480 -670
rect 76540 -730 76580 -670
rect 76440 -770 76580 -730
rect 76440 -830 76480 -770
rect 76540 -830 76580 -770
rect 76440 -850 76580 -830
rect 76610 -670 76750 -650
rect 76610 -730 76650 -670
rect 76710 -730 76750 -670
rect 76610 -770 76750 -730
rect 76610 -830 76650 -770
rect 76710 -830 76750 -770
rect 76610 -850 76750 -830
rect 76780 -670 76920 -650
rect 76780 -730 76820 -670
rect 76880 -730 76920 -670
rect 76780 -770 76920 -730
rect 76780 -830 76820 -770
rect 76880 -830 76920 -770
rect 76780 -850 76920 -830
rect 76950 -670 77090 -650
rect 76950 -730 76990 -670
rect 77050 -730 77090 -670
rect 76950 -770 77090 -730
rect 76950 -830 76990 -770
rect 77050 -830 77090 -770
rect 76950 -850 77090 -830
rect 77120 -670 77260 -650
rect 77120 -730 77160 -670
rect 77220 -730 77260 -670
rect 77120 -770 77260 -730
rect 77120 -830 77160 -770
rect 77220 -830 77260 -770
rect 77120 -850 77260 -830
rect 77290 -670 77430 -650
rect 77290 -730 77330 -670
rect 77390 -730 77430 -670
rect 77290 -770 77430 -730
rect 77290 -830 77330 -770
rect 77390 -830 77430 -770
rect 77290 -850 77430 -830
rect 77460 -670 77600 -650
rect 77460 -730 77500 -670
rect 77560 -730 77600 -670
rect 77460 -770 77600 -730
rect 77460 -830 77500 -770
rect 77560 -830 77600 -770
rect 77460 -850 77600 -830
rect 77630 -670 77770 -650
rect 77630 -730 77670 -670
rect 77730 -730 77770 -670
rect 77630 -770 77770 -730
rect 77630 -830 77670 -770
rect 77730 -830 77770 -770
rect 77630 -850 77770 -830
rect 77800 -670 77940 -650
rect 77800 -730 77840 -670
rect 77900 -730 77940 -670
rect 77800 -770 77940 -730
rect 77800 -830 77840 -770
rect 77900 -830 77940 -770
rect 77800 -850 77940 -830
rect 77970 -670 78110 -650
rect 77970 -730 78010 -670
rect 78070 -730 78110 -670
rect 77970 -770 78110 -730
rect 77970 -830 78010 -770
rect 78070 -830 78110 -770
rect 77970 -850 78110 -830
rect 78140 -670 78280 -650
rect 78140 -730 78180 -670
rect 78240 -730 78280 -670
rect 78140 -770 78280 -730
rect 78140 -830 78180 -770
rect 78240 -830 78280 -770
rect 78140 -850 78280 -830
rect 78310 -670 78450 -650
rect 78310 -730 78350 -670
rect 78410 -730 78450 -670
rect 78310 -770 78450 -730
rect 78310 -830 78350 -770
rect 78410 -830 78450 -770
rect 78310 -850 78450 -830
rect 78480 -670 78620 -650
rect 78480 -730 78520 -670
rect 78580 -730 78620 -670
rect 78480 -770 78620 -730
rect 78480 -830 78520 -770
rect 78580 -830 78620 -770
rect 78480 -850 78620 -830
rect 78650 -670 78790 -650
rect 78650 -730 78690 -670
rect 78750 -730 78790 -670
rect 78650 -770 78790 -730
rect 78650 -830 78690 -770
rect 78750 -830 78790 -770
rect 78650 -850 78790 -830
rect 78820 -670 78960 -650
rect 78820 -730 78860 -670
rect 78920 -730 78960 -670
rect 78820 -770 78960 -730
rect 78820 -830 78860 -770
rect 78920 -830 78960 -770
rect 78820 -850 78960 -830
rect 78990 -670 79130 -650
rect 78990 -730 79030 -670
rect 79090 -730 79130 -670
rect 78990 -770 79130 -730
rect 78990 -830 79030 -770
rect 79090 -830 79130 -770
rect 78990 -850 79130 -830
rect 79160 -670 79300 -650
rect 79160 -730 79200 -670
rect 79260 -730 79300 -670
rect 79160 -770 79300 -730
rect 79160 -830 79200 -770
rect 79260 -830 79300 -770
rect 79160 -850 79300 -830
rect 79330 -670 79470 -650
rect 79330 -730 79370 -670
rect 79430 -730 79470 -670
rect 79330 -770 79470 -730
rect 79330 -830 79370 -770
rect 79430 -830 79470 -770
rect 79330 -850 79470 -830
rect 79500 -670 79640 -650
rect 79500 -730 79540 -670
rect 79600 -730 79640 -670
rect 79500 -770 79640 -730
rect 79500 -830 79540 -770
rect 79600 -830 79640 -770
rect 79500 -850 79640 -830
rect 79670 -670 79810 -650
rect 79670 -730 79710 -670
rect 79770 -730 79810 -670
rect 79670 -770 79810 -730
rect 79670 -830 79710 -770
rect 79770 -830 79810 -770
rect 79670 -850 79810 -830
rect 79840 -670 79980 -650
rect 79840 -730 79880 -670
rect 79940 -730 79980 -670
rect 79840 -770 79980 -730
rect 79840 -830 79880 -770
rect 79940 -830 79980 -770
rect 79840 -850 79980 -830
rect 80010 -670 80150 -650
rect 80010 -730 80050 -670
rect 80110 -730 80150 -670
rect 80010 -770 80150 -730
rect 80010 -830 80050 -770
rect 80110 -830 80150 -770
rect 80010 -850 80150 -830
rect 80180 -670 80320 -650
rect 80180 -730 80220 -670
rect 80280 -730 80320 -670
rect 80180 -770 80320 -730
rect 80180 -830 80220 -770
rect 80280 -830 80320 -770
rect 80180 -850 80320 -830
rect 80350 -670 80490 -650
rect 80350 -730 80390 -670
rect 80450 -730 80490 -670
rect 80350 -770 80490 -730
rect 80350 -830 80390 -770
rect 80450 -830 80490 -770
rect 80350 -850 80490 -830
rect 80520 -670 80660 -650
rect 80520 -730 80560 -670
rect 80620 -730 80660 -670
rect 80520 -770 80660 -730
rect 80520 -830 80560 -770
rect 80620 -830 80660 -770
rect 80520 -850 80660 -830
rect 80690 -670 80830 -650
rect 80690 -730 80730 -670
rect 80790 -730 80830 -670
rect 80690 -770 80830 -730
rect 80690 -830 80730 -770
rect 80790 -830 80830 -770
rect 80690 -850 80830 -830
rect 80860 -670 81000 -650
rect 80860 -730 80900 -670
rect 80960 -730 81000 -670
rect 80860 -770 81000 -730
rect 80860 -830 80900 -770
rect 80960 -830 81000 -770
rect 80860 -850 81000 -830
rect 81030 -670 81170 -650
rect 81030 -730 81070 -670
rect 81130 -730 81170 -670
rect 81030 -770 81170 -730
rect 81030 -830 81070 -770
rect 81130 -830 81170 -770
rect 81030 -850 81170 -830
rect 81200 -670 81340 -650
rect 81200 -730 81240 -670
rect 81300 -730 81340 -670
rect 81200 -770 81340 -730
rect 81200 -830 81240 -770
rect 81300 -830 81340 -770
rect 81200 -850 81340 -830
rect 81370 -670 81510 -650
rect 81370 -730 81410 -670
rect 81470 -730 81510 -670
rect 81370 -770 81510 -730
rect 81370 -830 81410 -770
rect 81470 -830 81510 -770
rect 81370 -850 81510 -830
rect 81540 -670 81680 -650
rect 81540 -730 81580 -670
rect 81640 -730 81680 -670
rect 81540 -770 81680 -730
rect 81540 -830 81580 -770
rect 81640 -830 81680 -770
rect 81540 -850 81680 -830
rect 81710 -670 81850 -650
rect 81710 -730 81750 -670
rect 81810 -730 81850 -670
rect 81710 -770 81850 -730
rect 81710 -830 81750 -770
rect 81810 -830 81850 -770
rect 81710 -850 81850 -830
rect 81880 -670 82020 -650
rect 81880 -730 81920 -670
rect 81980 -730 82020 -670
rect 81880 -770 82020 -730
rect 81880 -830 81920 -770
rect 81980 -830 82020 -770
rect 81880 -850 82020 -830
rect 82050 -670 82190 -650
rect 82050 -730 82090 -670
rect 82150 -730 82190 -670
rect 82050 -770 82190 -730
rect 82050 -830 82090 -770
rect 82150 -830 82190 -770
rect 82050 -850 82190 -830
rect 82220 -670 82360 -650
rect 82220 -730 82260 -670
rect 82320 -730 82360 -670
rect 82220 -770 82360 -730
rect 82220 -830 82260 -770
rect 82320 -830 82360 -770
rect 82220 -850 82360 -830
rect 82390 -670 82530 -650
rect 82390 -730 82430 -670
rect 82490 -730 82530 -670
rect 82390 -770 82530 -730
rect 82390 -830 82430 -770
rect 82490 -830 82530 -770
rect 82390 -850 82530 -830
rect 82560 -670 82700 -650
rect 82560 -730 82600 -670
rect 82660 -730 82700 -670
rect 82560 -770 82700 -730
rect 82560 -830 82600 -770
rect 82660 -830 82700 -770
rect 82560 -850 82700 -830
rect 82730 -670 82870 -650
rect 82730 -730 82770 -670
rect 82830 -730 82870 -670
rect 82730 -770 82870 -730
rect 82730 -830 82770 -770
rect 82830 -830 82870 -770
rect 82730 -850 82870 -830
rect 82900 -670 83040 -650
rect 82900 -730 82940 -670
rect 83000 -730 83040 -670
rect 82900 -770 83040 -730
rect 82900 -830 82940 -770
rect 83000 -830 83040 -770
rect 82900 -850 83040 -830
rect 83070 -670 83210 -650
rect 83070 -730 83110 -670
rect 83170 -730 83210 -670
rect 83070 -770 83210 -730
rect 83070 -830 83110 -770
rect 83170 -830 83210 -770
rect 83070 -850 83210 -830
rect 83240 -670 83380 -650
rect 83240 -730 83280 -670
rect 83340 -730 83380 -670
rect 83240 -770 83380 -730
rect 83240 -830 83280 -770
rect 83340 -830 83380 -770
rect 83240 -850 83380 -830
rect 83410 -670 83550 -650
rect 83410 -730 83450 -670
rect 83510 -730 83550 -670
rect 83410 -770 83550 -730
rect 83410 -830 83450 -770
rect 83510 -830 83550 -770
rect 83410 -850 83550 -830
rect 83580 -670 83720 -650
rect 83580 -730 83620 -670
rect 83680 -730 83720 -670
rect 83580 -770 83720 -730
rect 83580 -830 83620 -770
rect 83680 -830 83720 -770
rect 83580 -850 83720 -830
rect 83750 -670 83890 -650
rect 83750 -730 83790 -670
rect 83850 -730 83890 -670
rect 83750 -770 83890 -730
rect 83750 -830 83790 -770
rect 83850 -830 83890 -770
rect 83750 -850 83890 -830
rect 83920 -670 84060 -650
rect 83920 -730 83960 -670
rect 84020 -730 84060 -670
rect 83920 -770 84060 -730
rect 83920 -830 83960 -770
rect 84020 -830 84060 -770
rect 83920 -850 84060 -830
rect 84090 -670 84230 -650
rect 84090 -730 84130 -670
rect 84190 -730 84230 -670
rect 84090 -770 84230 -730
rect 84090 -830 84130 -770
rect 84190 -830 84230 -770
rect 84090 -850 84230 -830
rect 84260 -670 84400 -650
rect 84260 -730 84300 -670
rect 84360 -730 84400 -670
rect 84260 -770 84400 -730
rect 84260 -830 84300 -770
rect 84360 -830 84400 -770
rect 84260 -850 84400 -830
rect 84430 -670 84570 -650
rect 84430 -730 84470 -670
rect 84530 -730 84570 -670
rect 84430 -770 84570 -730
rect 84430 -830 84470 -770
rect 84530 -830 84570 -770
rect 84430 -850 84570 -830
rect 84600 -670 84740 -650
rect 84600 -730 84640 -670
rect 84700 -730 84740 -670
rect 84600 -770 84740 -730
rect 84600 -830 84640 -770
rect 84700 -830 84740 -770
rect 84600 -850 84740 -830
rect 84770 -670 84910 -650
rect 84770 -730 84810 -670
rect 84870 -730 84910 -670
rect 84770 -770 84910 -730
rect 84770 -830 84810 -770
rect 84870 -830 84910 -770
rect 84770 -850 84910 -830
rect 84940 -670 85080 -650
rect 84940 -730 84980 -670
rect 85040 -730 85080 -670
rect 84940 -770 85080 -730
rect 84940 -830 84980 -770
rect 85040 -830 85080 -770
rect 84940 -850 85080 -830
rect 85110 -670 85250 -650
rect 85110 -730 85150 -670
rect 85210 -730 85250 -670
rect 85110 -770 85250 -730
rect 85110 -830 85150 -770
rect 85210 -830 85250 -770
rect 85110 -850 85250 -830
rect 85280 -670 85420 -650
rect 85280 -730 85320 -670
rect 85380 -730 85420 -670
rect 85280 -770 85420 -730
rect 85280 -830 85320 -770
rect 85380 -830 85420 -770
rect 85280 -850 85420 -830
rect 85450 -670 85590 -650
rect 85450 -730 85490 -670
rect 85550 -730 85590 -670
rect 85450 -770 85590 -730
rect 85450 -830 85490 -770
rect 85550 -830 85590 -770
rect 85450 -850 85590 -830
rect 85620 -670 85760 -650
rect 85620 -730 85660 -670
rect 85720 -730 85760 -670
rect 85620 -770 85760 -730
rect 85620 -830 85660 -770
rect 85720 -830 85760 -770
rect 85620 -850 85760 -830
rect 85790 -670 85930 -650
rect 85790 -730 85830 -670
rect 85890 -730 85930 -670
rect 85790 -770 85930 -730
rect 85790 -830 85830 -770
rect 85890 -830 85930 -770
rect 85790 -850 85930 -830
rect 85960 -670 86100 -650
rect 85960 -730 86000 -670
rect 86060 -730 86100 -670
rect 85960 -770 86100 -730
rect 85960 -830 86000 -770
rect 86060 -830 86100 -770
rect 85960 -850 86100 -830
rect 86130 -670 86270 -650
rect 86130 -730 86170 -670
rect 86230 -730 86270 -670
rect 86130 -770 86270 -730
rect 86130 -830 86170 -770
rect 86230 -830 86270 -770
rect 86130 -850 86270 -830
rect 86300 -670 86440 -650
rect 86300 -730 86340 -670
rect 86400 -730 86440 -670
rect 86300 -770 86440 -730
rect 86300 -830 86340 -770
rect 86400 -830 86440 -770
rect 86300 -850 86440 -830
rect 86470 -670 86610 -650
rect 86470 -730 86510 -670
rect 86570 -730 86610 -670
rect 86470 -770 86610 -730
rect 86470 -830 86510 -770
rect 86570 -830 86610 -770
rect 86470 -850 86610 -830
rect 86640 -670 86780 -650
rect 86640 -730 86680 -670
rect 86740 -730 86780 -670
rect 86640 -770 86780 -730
rect 86640 -830 86680 -770
rect 86740 -830 86780 -770
rect 86640 -850 86780 -830
rect 86810 -670 86950 -650
rect 86810 -730 86850 -670
rect 86910 -730 86950 -670
rect 86810 -770 86950 -730
rect 86810 -830 86850 -770
rect 86910 -830 86950 -770
rect 86810 -850 86950 -830
rect 86980 -670 87120 -650
rect 86980 -730 87020 -670
rect 87080 -730 87120 -670
rect 86980 -770 87120 -730
rect 86980 -830 87020 -770
rect 87080 -830 87120 -770
rect 86980 -850 87120 -830
rect 87150 -670 87290 -650
rect 87150 -730 87190 -670
rect 87250 -730 87290 -670
rect 87150 -770 87290 -730
rect 87150 -830 87190 -770
rect 87250 -830 87290 -770
rect 87150 -850 87290 -830
<< pdiff >>
rect -10 410 130 430
rect -10 350 30 410
rect 90 350 130 410
rect -10 310 130 350
rect -10 250 30 310
rect 90 250 130 310
rect -10 230 130 250
rect 160 410 300 430
rect 160 350 200 410
rect 260 350 300 410
rect 160 310 300 350
rect 160 250 200 310
rect 260 250 300 310
rect 160 230 300 250
rect 410 410 550 430
rect 410 350 450 410
rect 510 350 550 410
rect 410 310 550 350
rect 410 250 450 310
rect 510 250 550 310
rect 410 230 550 250
rect 580 410 720 430
rect 580 350 620 410
rect 680 350 720 410
rect 580 310 720 350
rect 580 250 620 310
rect 680 250 720 310
rect 580 230 720 250
rect 750 410 890 430
rect 750 350 790 410
rect 850 350 890 410
rect 750 310 890 350
rect 750 250 790 310
rect 850 250 890 310
rect 750 230 890 250
rect 920 410 1060 430
rect 920 350 960 410
rect 1020 350 1060 410
rect 920 310 1060 350
rect 920 250 960 310
rect 1020 250 1060 310
rect 920 230 1060 250
rect 1090 410 1230 430
rect 1090 350 1130 410
rect 1190 350 1230 410
rect 1090 310 1230 350
rect 1090 250 1130 310
rect 1190 250 1230 310
rect 1090 230 1230 250
rect 1480 410 1620 430
rect 1480 350 1520 410
rect 1580 350 1620 410
rect 1480 310 1620 350
rect 1480 250 1520 310
rect 1580 250 1620 310
rect 1480 230 1620 250
rect 1650 410 1790 430
rect 1650 350 1690 410
rect 1750 350 1790 410
rect 1650 310 1790 350
rect 1650 250 1690 310
rect 1750 250 1790 310
rect 1650 230 1790 250
rect 1820 410 1960 430
rect 1820 350 1860 410
rect 1920 350 1960 410
rect 1820 310 1960 350
rect 1820 250 1860 310
rect 1920 250 1960 310
rect 1820 230 1960 250
rect 1990 410 2130 430
rect 1990 350 2030 410
rect 2090 350 2130 410
rect 1990 310 2130 350
rect 1990 250 2030 310
rect 2090 250 2130 310
rect 1990 230 2130 250
rect 2160 410 2300 430
rect 2160 350 2200 410
rect 2260 350 2300 410
rect 2160 310 2300 350
rect 2160 250 2200 310
rect 2260 250 2300 310
rect 2160 230 2300 250
rect 2330 410 2470 430
rect 2330 350 2370 410
rect 2430 350 2470 410
rect 2330 310 2470 350
rect 2330 250 2370 310
rect 2430 250 2470 310
rect 2330 230 2470 250
rect 2500 410 2640 430
rect 2500 350 2540 410
rect 2600 350 2640 410
rect 2500 310 2640 350
rect 2500 250 2540 310
rect 2600 250 2640 310
rect 2500 230 2640 250
rect 2670 410 2810 430
rect 2670 350 2710 410
rect 2770 350 2810 410
rect 2670 310 2810 350
rect 2670 250 2710 310
rect 2770 250 2810 310
rect 2670 230 2810 250
rect 2840 410 2980 430
rect 2840 350 2880 410
rect 2940 350 2980 410
rect 2840 310 2980 350
rect 2840 250 2880 310
rect 2940 250 2980 310
rect 2840 230 2980 250
rect 3010 410 3150 430
rect 3010 350 3050 410
rect 3110 350 3150 410
rect 3010 310 3150 350
rect 3010 250 3050 310
rect 3110 250 3150 310
rect 3010 230 3150 250
rect 3180 410 3320 430
rect 3180 350 3220 410
rect 3280 350 3320 410
rect 3180 310 3320 350
rect 3180 250 3220 310
rect 3280 250 3320 310
rect 3180 230 3320 250
rect 3350 410 3490 430
rect 3350 350 3390 410
rect 3450 350 3490 410
rect 3350 310 3490 350
rect 3350 250 3390 310
rect 3450 250 3490 310
rect 3350 230 3490 250
rect 3520 410 3660 430
rect 3520 350 3560 410
rect 3620 350 3660 410
rect 3520 310 3660 350
rect 3520 250 3560 310
rect 3620 250 3660 310
rect 3520 230 3660 250
rect 3690 410 3830 430
rect 3690 350 3730 410
rect 3790 350 3830 410
rect 3690 310 3830 350
rect 3690 250 3730 310
rect 3790 250 3830 310
rect 3690 230 3830 250
rect 3860 410 4000 430
rect 3860 350 3900 410
rect 3960 350 4000 410
rect 3860 310 4000 350
rect 3860 250 3900 310
rect 3960 250 4000 310
rect 3860 230 4000 250
rect 4030 410 4170 430
rect 4030 350 4070 410
rect 4130 350 4170 410
rect 4030 310 4170 350
rect 4030 250 4070 310
rect 4130 250 4170 310
rect 4030 230 4170 250
rect 4200 410 4340 430
rect 4200 350 4240 410
rect 4300 350 4340 410
rect 4200 310 4340 350
rect 4200 250 4240 310
rect 4300 250 4340 310
rect 4200 230 4340 250
rect 4500 410 4640 430
rect 4500 350 4540 410
rect 4600 350 4640 410
rect 4500 310 4640 350
rect 4500 250 4540 310
rect 4600 250 4640 310
rect 4500 230 4640 250
rect 4670 410 4810 430
rect 4670 350 4710 410
rect 4770 350 4810 410
rect 4670 310 4810 350
rect 4670 250 4710 310
rect 4770 250 4810 310
rect 4670 230 4810 250
rect 4840 410 4980 430
rect 4840 350 4880 410
rect 4940 350 4980 410
rect 4840 310 4980 350
rect 4840 250 4880 310
rect 4940 250 4980 310
rect 4840 230 4980 250
rect 5010 410 5150 430
rect 5010 350 5050 410
rect 5110 350 5150 410
rect 5010 310 5150 350
rect 5010 250 5050 310
rect 5110 250 5150 310
rect 5010 230 5150 250
rect 5180 410 5320 430
rect 5180 350 5220 410
rect 5280 350 5320 410
rect 5180 310 5320 350
rect 5180 250 5220 310
rect 5280 250 5320 310
rect 5180 230 5320 250
rect 5350 410 5490 430
rect 5350 350 5390 410
rect 5450 350 5490 410
rect 5350 310 5490 350
rect 5350 250 5390 310
rect 5450 250 5490 310
rect 5350 230 5490 250
rect 5520 410 5660 430
rect 5520 350 5560 410
rect 5620 350 5660 410
rect 5520 310 5660 350
rect 5520 250 5560 310
rect 5620 250 5660 310
rect 5520 230 5660 250
rect 5690 410 5830 430
rect 5690 350 5730 410
rect 5790 350 5830 410
rect 5690 310 5830 350
rect 5690 250 5730 310
rect 5790 250 5830 310
rect 5690 230 5830 250
rect 5860 410 6000 430
rect 5860 350 5900 410
rect 5960 350 6000 410
rect 5860 310 6000 350
rect 5860 250 5900 310
rect 5960 250 6000 310
rect 5860 230 6000 250
rect 6030 410 6170 430
rect 6030 350 6070 410
rect 6130 350 6170 410
rect 6030 310 6170 350
rect 6030 250 6070 310
rect 6130 250 6170 310
rect 6030 230 6170 250
rect 6200 410 6340 430
rect 6200 350 6240 410
rect 6300 350 6340 410
rect 6200 310 6340 350
rect 6200 250 6240 310
rect 6300 250 6340 310
rect 6200 230 6340 250
rect 6370 410 6510 430
rect 6370 350 6410 410
rect 6470 350 6510 410
rect 6370 310 6510 350
rect 6370 250 6410 310
rect 6470 250 6510 310
rect 6370 230 6510 250
rect 6540 410 6680 430
rect 6540 350 6580 410
rect 6640 350 6680 410
rect 6540 310 6680 350
rect 6540 250 6580 310
rect 6640 250 6680 310
rect 6540 230 6680 250
rect 6710 410 6850 430
rect 6710 350 6750 410
rect 6810 350 6850 410
rect 6710 310 6850 350
rect 6710 250 6750 310
rect 6810 250 6850 310
rect 6710 230 6850 250
rect 6880 410 7020 430
rect 6880 350 6920 410
rect 6980 350 7020 410
rect 6880 310 7020 350
rect 6880 250 6920 310
rect 6980 250 7020 310
rect 6880 230 7020 250
rect 7050 410 7190 430
rect 7050 350 7090 410
rect 7150 350 7190 410
rect 7050 310 7190 350
rect 7050 250 7090 310
rect 7150 250 7190 310
rect 7050 230 7190 250
rect 7220 410 7360 430
rect 7220 350 7260 410
rect 7320 350 7360 410
rect 7220 310 7360 350
rect 7220 250 7260 310
rect 7320 250 7360 310
rect 7220 230 7360 250
rect 7390 410 7530 430
rect 7390 350 7430 410
rect 7490 350 7530 410
rect 7390 310 7530 350
rect 7390 250 7430 310
rect 7490 250 7530 310
rect 7390 230 7530 250
rect 7560 410 7700 430
rect 7560 350 7600 410
rect 7660 350 7700 410
rect 7560 310 7700 350
rect 7560 250 7600 310
rect 7660 250 7700 310
rect 7560 230 7700 250
rect 7730 410 7870 430
rect 7730 350 7770 410
rect 7830 350 7870 410
rect 7730 310 7870 350
rect 7730 250 7770 310
rect 7830 250 7870 310
rect 7730 230 7870 250
rect 7900 410 8040 430
rect 7900 350 7940 410
rect 8000 350 8040 410
rect 7900 310 8040 350
rect 7900 250 7940 310
rect 8000 250 8040 310
rect 7900 230 8040 250
rect 8070 410 8210 430
rect 8070 350 8110 410
rect 8170 350 8210 410
rect 8070 310 8210 350
rect 8070 250 8110 310
rect 8170 250 8210 310
rect 8070 230 8210 250
rect 8240 410 8380 430
rect 8240 350 8280 410
rect 8340 350 8380 410
rect 8240 310 8380 350
rect 8240 250 8280 310
rect 8340 250 8380 310
rect 8240 230 8380 250
rect 8410 410 8550 430
rect 8410 350 8450 410
rect 8510 350 8550 410
rect 8410 310 8550 350
rect 8410 250 8450 310
rect 8510 250 8550 310
rect 8410 230 8550 250
rect 8580 410 8720 430
rect 8580 350 8620 410
rect 8680 350 8720 410
rect 8580 310 8720 350
rect 8580 250 8620 310
rect 8680 250 8720 310
rect 8580 230 8720 250
rect 8750 410 8890 430
rect 8750 350 8790 410
rect 8850 350 8890 410
rect 8750 310 8890 350
rect 8750 250 8790 310
rect 8850 250 8890 310
rect 8750 230 8890 250
rect 8920 410 9060 430
rect 8920 350 8960 410
rect 9020 350 9060 410
rect 8920 310 9060 350
rect 8920 250 8960 310
rect 9020 250 9060 310
rect 8920 230 9060 250
rect 9090 410 9230 430
rect 9090 350 9130 410
rect 9190 350 9230 410
rect 9090 310 9230 350
rect 9090 250 9130 310
rect 9190 250 9230 310
rect 9090 230 9230 250
rect 9260 410 9400 430
rect 9260 350 9300 410
rect 9360 350 9400 410
rect 9260 310 9400 350
rect 9260 250 9300 310
rect 9360 250 9400 310
rect 9260 230 9400 250
rect 9430 410 9570 430
rect 9430 350 9470 410
rect 9530 350 9570 410
rect 9430 310 9570 350
rect 9430 250 9470 310
rect 9530 250 9570 310
rect 9430 230 9570 250
rect 9600 410 9740 430
rect 9600 350 9640 410
rect 9700 350 9740 410
rect 9600 310 9740 350
rect 9600 250 9640 310
rect 9700 250 9740 310
rect 9600 230 9740 250
rect 9770 410 9910 430
rect 9770 350 9810 410
rect 9870 350 9910 410
rect 9770 310 9910 350
rect 9770 250 9810 310
rect 9870 250 9910 310
rect 9770 230 9910 250
rect 9940 410 10080 430
rect 9940 350 9980 410
rect 10040 350 10080 410
rect 9940 310 10080 350
rect 9940 250 9980 310
rect 10040 250 10080 310
rect 9940 230 10080 250
rect 10110 410 10250 430
rect 10110 350 10150 410
rect 10210 350 10250 410
rect 10110 310 10250 350
rect 10110 250 10150 310
rect 10210 250 10250 310
rect 10110 230 10250 250
rect 10280 410 10420 430
rect 10280 350 10320 410
rect 10380 350 10420 410
rect 10280 310 10420 350
rect 10280 250 10320 310
rect 10380 250 10420 310
rect 10280 230 10420 250
rect 10450 410 10590 430
rect 10450 350 10490 410
rect 10550 350 10590 410
rect 10450 310 10590 350
rect 10450 250 10490 310
rect 10550 250 10590 310
rect 10450 230 10590 250
rect 10620 410 10760 430
rect 10620 350 10660 410
rect 10720 350 10760 410
rect 10620 310 10760 350
rect 10620 250 10660 310
rect 10720 250 10760 310
rect 10620 230 10760 250
rect 10790 410 10930 430
rect 10790 350 10830 410
rect 10890 350 10930 410
rect 10790 310 10930 350
rect 10790 250 10830 310
rect 10890 250 10930 310
rect 10790 230 10930 250
rect 10960 410 11100 430
rect 10960 350 11000 410
rect 11060 350 11100 410
rect 10960 310 11100 350
rect 10960 250 11000 310
rect 11060 250 11100 310
rect 10960 230 11100 250
rect 11130 410 11270 430
rect 11130 350 11170 410
rect 11230 350 11270 410
rect 11130 310 11270 350
rect 11130 250 11170 310
rect 11230 250 11270 310
rect 11130 230 11270 250
rect 11300 410 11440 430
rect 11300 350 11340 410
rect 11400 350 11440 410
rect 11300 310 11440 350
rect 11300 250 11340 310
rect 11400 250 11440 310
rect 11300 230 11440 250
rect 11470 410 11610 430
rect 11470 350 11510 410
rect 11570 350 11610 410
rect 11470 310 11610 350
rect 11470 250 11510 310
rect 11570 250 11610 310
rect 11470 230 11610 250
rect 11640 410 11780 430
rect 11640 350 11680 410
rect 11740 350 11780 410
rect 11640 310 11780 350
rect 11640 250 11680 310
rect 11740 250 11780 310
rect 11640 230 11780 250
rect 11810 410 11950 430
rect 11810 350 11850 410
rect 11910 350 11950 410
rect 11810 310 11950 350
rect 11810 250 11850 310
rect 11910 250 11950 310
rect 11810 230 11950 250
rect 11980 410 12120 430
rect 11980 350 12020 410
rect 12080 350 12120 410
rect 11980 310 12120 350
rect 11980 250 12020 310
rect 12080 250 12120 310
rect 11980 230 12120 250
rect 12150 410 12290 430
rect 12150 350 12190 410
rect 12250 350 12290 410
rect 12150 310 12290 350
rect 12150 250 12190 310
rect 12250 250 12290 310
rect 12150 230 12290 250
rect 12320 410 12460 430
rect 12320 350 12360 410
rect 12420 350 12460 410
rect 12320 310 12460 350
rect 12320 250 12360 310
rect 12420 250 12460 310
rect 12320 230 12460 250
rect 12490 410 12630 430
rect 12490 350 12530 410
rect 12590 350 12630 410
rect 12490 310 12630 350
rect 12490 250 12530 310
rect 12590 250 12630 310
rect 12490 230 12630 250
rect 12660 410 12800 430
rect 12660 350 12700 410
rect 12760 350 12800 410
rect 12660 310 12800 350
rect 12660 250 12700 310
rect 12760 250 12800 310
rect 12660 230 12800 250
rect 12830 410 12970 430
rect 12830 350 12870 410
rect 12930 350 12970 410
rect 12830 310 12970 350
rect 12830 250 12870 310
rect 12930 250 12970 310
rect 12830 230 12970 250
rect 13000 410 13140 430
rect 13000 350 13040 410
rect 13100 350 13140 410
rect 13000 310 13140 350
rect 13000 250 13040 310
rect 13100 250 13140 310
rect 13000 230 13140 250
rect 13170 410 13310 430
rect 13170 350 13210 410
rect 13270 350 13310 410
rect 13170 310 13310 350
rect 13170 250 13210 310
rect 13270 250 13310 310
rect 13170 230 13310 250
rect 13340 410 13480 430
rect 13340 350 13380 410
rect 13440 350 13480 410
rect 13340 310 13480 350
rect 13340 250 13380 310
rect 13440 250 13480 310
rect 13340 230 13480 250
rect 13510 410 13650 430
rect 13510 350 13550 410
rect 13610 350 13650 410
rect 13510 310 13650 350
rect 13510 250 13550 310
rect 13610 250 13650 310
rect 13510 230 13650 250
rect 13680 410 13820 430
rect 13680 350 13720 410
rect 13780 350 13820 410
rect 13680 310 13820 350
rect 13680 250 13720 310
rect 13780 250 13820 310
rect 13680 230 13820 250
rect 13850 410 13990 430
rect 13850 350 13890 410
rect 13950 350 13990 410
rect 13850 310 13990 350
rect 13850 250 13890 310
rect 13950 250 13990 310
rect 13850 230 13990 250
rect 14020 410 14160 430
rect 14020 350 14060 410
rect 14120 350 14160 410
rect 14020 310 14160 350
rect 14020 250 14060 310
rect 14120 250 14160 310
rect 14020 230 14160 250
rect 14190 410 14330 430
rect 14190 350 14230 410
rect 14290 350 14330 410
rect 14190 310 14330 350
rect 14190 250 14230 310
rect 14290 250 14330 310
rect 14190 230 14330 250
rect 14360 410 14500 430
rect 14360 350 14400 410
rect 14460 350 14500 410
rect 14360 310 14500 350
rect 14360 250 14400 310
rect 14460 250 14500 310
rect 14360 230 14500 250
rect 14530 410 14670 430
rect 14530 350 14570 410
rect 14630 350 14670 410
rect 14530 310 14670 350
rect 14530 250 14570 310
rect 14630 250 14670 310
rect 14530 230 14670 250
rect 14700 410 14840 430
rect 14700 350 14740 410
rect 14800 350 14840 410
rect 14700 310 14840 350
rect 14700 250 14740 310
rect 14800 250 14840 310
rect 14700 230 14840 250
rect 14870 410 15010 430
rect 14870 350 14910 410
rect 14970 350 15010 410
rect 14870 310 15010 350
rect 14870 250 14910 310
rect 14970 250 15010 310
rect 14870 230 15010 250
rect 15040 410 15180 430
rect 15040 350 15080 410
rect 15140 350 15180 410
rect 15040 310 15180 350
rect 15040 250 15080 310
rect 15140 250 15180 310
rect 15040 230 15180 250
rect 15210 410 15350 430
rect 15210 350 15250 410
rect 15310 350 15350 410
rect 15210 310 15350 350
rect 15210 250 15250 310
rect 15310 250 15350 310
rect 15210 230 15350 250
rect 15380 410 15520 430
rect 15380 350 15420 410
rect 15480 350 15520 410
rect 15380 310 15520 350
rect 15380 250 15420 310
rect 15480 250 15520 310
rect 15380 230 15520 250
rect 15680 410 15820 430
rect 15680 350 15720 410
rect 15780 350 15820 410
rect 15680 310 15820 350
rect 15680 250 15720 310
rect 15780 250 15820 310
rect 15680 230 15820 250
rect 15850 410 15990 430
rect 15850 350 15890 410
rect 15950 350 15990 410
rect 15850 310 15990 350
rect 15850 250 15890 310
rect 15950 250 15990 310
rect 15850 230 15990 250
rect 16020 410 16160 430
rect 16020 350 16060 410
rect 16120 350 16160 410
rect 16020 310 16160 350
rect 16020 250 16060 310
rect 16120 250 16160 310
rect 16020 230 16160 250
rect 16190 410 16330 430
rect 16190 350 16230 410
rect 16290 350 16330 410
rect 16190 310 16330 350
rect 16190 250 16230 310
rect 16290 250 16330 310
rect 16190 230 16330 250
rect 16360 410 16500 430
rect 16360 350 16400 410
rect 16460 350 16500 410
rect 16360 310 16500 350
rect 16360 250 16400 310
rect 16460 250 16500 310
rect 16360 230 16500 250
rect 16530 410 16670 430
rect 16530 350 16570 410
rect 16630 350 16670 410
rect 16530 310 16670 350
rect 16530 250 16570 310
rect 16630 250 16670 310
rect 16530 230 16670 250
rect 16700 410 16840 430
rect 16700 350 16740 410
rect 16800 350 16840 410
rect 16700 310 16840 350
rect 16700 250 16740 310
rect 16800 250 16840 310
rect 16700 230 16840 250
rect 16870 410 17010 430
rect 16870 350 16910 410
rect 16970 350 17010 410
rect 16870 310 17010 350
rect 16870 250 16910 310
rect 16970 250 17010 310
rect 16870 230 17010 250
rect 17040 410 17180 430
rect 17040 350 17080 410
rect 17140 350 17180 410
rect 17040 310 17180 350
rect 17040 250 17080 310
rect 17140 250 17180 310
rect 17040 230 17180 250
rect 17210 410 17350 430
rect 17210 350 17250 410
rect 17310 350 17350 410
rect 17210 310 17350 350
rect 17210 250 17250 310
rect 17310 250 17350 310
rect 17210 230 17350 250
rect 17380 410 17520 430
rect 17380 350 17420 410
rect 17480 350 17520 410
rect 17380 310 17520 350
rect 17380 250 17420 310
rect 17480 250 17520 310
rect 17380 230 17520 250
rect 17550 410 17690 430
rect 17550 350 17590 410
rect 17650 350 17690 410
rect 17550 310 17690 350
rect 17550 250 17590 310
rect 17650 250 17690 310
rect 17550 230 17690 250
rect 17720 410 17860 430
rect 17720 350 17760 410
rect 17820 350 17860 410
rect 17720 310 17860 350
rect 17720 250 17760 310
rect 17820 250 17860 310
rect 17720 230 17860 250
rect 17890 410 18030 430
rect 17890 350 17930 410
rect 17990 350 18030 410
rect 17890 310 18030 350
rect 17890 250 17930 310
rect 17990 250 18030 310
rect 17890 230 18030 250
rect 18060 410 18200 430
rect 18060 350 18100 410
rect 18160 350 18200 410
rect 18060 310 18200 350
rect 18060 250 18100 310
rect 18160 250 18200 310
rect 18060 230 18200 250
rect 18230 410 18370 430
rect 18230 350 18270 410
rect 18330 350 18370 410
rect 18230 310 18370 350
rect 18230 250 18270 310
rect 18330 250 18370 310
rect 18230 230 18370 250
rect 18400 410 18540 430
rect 18400 350 18440 410
rect 18500 350 18540 410
rect 18400 310 18540 350
rect 18400 250 18440 310
rect 18500 250 18540 310
rect 18400 230 18540 250
rect 18570 410 18710 430
rect 18570 350 18610 410
rect 18670 350 18710 410
rect 18570 310 18710 350
rect 18570 250 18610 310
rect 18670 250 18710 310
rect 18570 230 18710 250
rect 18740 410 18880 430
rect 18740 350 18780 410
rect 18840 350 18880 410
rect 18740 310 18880 350
rect 18740 250 18780 310
rect 18840 250 18880 310
rect 18740 230 18880 250
rect 18910 410 19050 430
rect 18910 350 18950 410
rect 19010 350 19050 410
rect 18910 310 19050 350
rect 18910 250 18950 310
rect 19010 250 19050 310
rect 18910 230 19050 250
rect 19080 410 19220 430
rect 19080 350 19120 410
rect 19180 350 19220 410
rect 19080 310 19220 350
rect 19080 250 19120 310
rect 19180 250 19220 310
rect 19080 230 19220 250
rect 19250 410 19390 430
rect 19250 350 19290 410
rect 19350 350 19390 410
rect 19250 310 19390 350
rect 19250 250 19290 310
rect 19350 250 19390 310
rect 19250 230 19390 250
rect 19420 410 19560 430
rect 19420 350 19460 410
rect 19520 350 19560 410
rect 19420 310 19560 350
rect 19420 250 19460 310
rect 19520 250 19560 310
rect 19420 230 19560 250
rect 19590 410 19730 430
rect 19590 350 19630 410
rect 19690 350 19730 410
rect 19590 310 19730 350
rect 19590 250 19630 310
rect 19690 250 19730 310
rect 19590 230 19730 250
rect 19760 410 19900 430
rect 19760 350 19800 410
rect 19860 350 19900 410
rect 19760 310 19900 350
rect 19760 250 19800 310
rect 19860 250 19900 310
rect 19760 230 19900 250
rect 19930 410 20070 430
rect 19930 350 19970 410
rect 20030 350 20070 410
rect 19930 310 20070 350
rect 19930 250 19970 310
rect 20030 250 20070 310
rect 19930 230 20070 250
rect 20100 410 20240 430
rect 20100 350 20140 410
rect 20200 350 20240 410
rect 20100 310 20240 350
rect 20100 250 20140 310
rect 20200 250 20240 310
rect 20100 230 20240 250
rect 20270 410 20410 430
rect 20270 350 20310 410
rect 20370 350 20410 410
rect 20270 310 20410 350
rect 20270 250 20310 310
rect 20370 250 20410 310
rect 20270 230 20410 250
rect 20440 410 20580 430
rect 20440 350 20480 410
rect 20540 350 20580 410
rect 20440 310 20580 350
rect 20440 250 20480 310
rect 20540 250 20580 310
rect 20440 230 20580 250
rect 20610 410 20750 430
rect 20610 350 20650 410
rect 20710 350 20750 410
rect 20610 310 20750 350
rect 20610 250 20650 310
rect 20710 250 20750 310
rect 20610 230 20750 250
rect 20780 410 20920 430
rect 20780 350 20820 410
rect 20880 350 20920 410
rect 20780 310 20920 350
rect 20780 250 20820 310
rect 20880 250 20920 310
rect 20780 230 20920 250
rect 20950 410 21090 430
rect 20950 350 20990 410
rect 21050 350 21090 410
rect 20950 310 21090 350
rect 20950 250 20990 310
rect 21050 250 21090 310
rect 20950 230 21090 250
rect 21120 410 21260 430
rect 21120 350 21160 410
rect 21220 350 21260 410
rect 21120 310 21260 350
rect 21120 250 21160 310
rect 21220 250 21260 310
rect 21120 230 21260 250
rect 21290 410 21430 430
rect 21290 350 21330 410
rect 21390 350 21430 410
rect 21290 310 21430 350
rect 21290 250 21330 310
rect 21390 250 21430 310
rect 21290 230 21430 250
rect 21460 410 21600 430
rect 21460 350 21500 410
rect 21560 350 21600 410
rect 21460 310 21600 350
rect 21460 250 21500 310
rect 21560 250 21600 310
rect 21460 230 21600 250
rect 21630 410 21770 430
rect 21630 350 21670 410
rect 21730 350 21770 410
rect 21630 310 21770 350
rect 21630 250 21670 310
rect 21730 250 21770 310
rect 21630 230 21770 250
rect 21800 410 21940 430
rect 21800 350 21840 410
rect 21900 350 21940 410
rect 21800 310 21940 350
rect 21800 250 21840 310
rect 21900 250 21940 310
rect 21800 230 21940 250
rect 21970 410 22110 430
rect 21970 350 22010 410
rect 22070 350 22110 410
rect 21970 310 22110 350
rect 21970 250 22010 310
rect 22070 250 22110 310
rect 21970 230 22110 250
rect 22140 410 22280 430
rect 22140 350 22180 410
rect 22240 350 22280 410
rect 22140 310 22280 350
rect 22140 250 22180 310
rect 22240 250 22280 310
rect 22140 230 22280 250
rect 22310 410 22450 430
rect 22310 350 22350 410
rect 22410 350 22450 410
rect 22310 310 22450 350
rect 22310 250 22350 310
rect 22410 250 22450 310
rect 22310 230 22450 250
rect 22480 410 22620 430
rect 22480 350 22520 410
rect 22580 350 22620 410
rect 22480 310 22620 350
rect 22480 250 22520 310
rect 22580 250 22620 310
rect 22480 230 22620 250
rect 22650 410 22790 430
rect 22650 350 22690 410
rect 22750 350 22790 410
rect 22650 310 22790 350
rect 22650 250 22690 310
rect 22750 250 22790 310
rect 22650 230 22790 250
rect 22820 410 22960 430
rect 22820 350 22860 410
rect 22920 350 22960 410
rect 22820 310 22960 350
rect 22820 250 22860 310
rect 22920 250 22960 310
rect 22820 230 22960 250
rect 22990 410 23130 430
rect 22990 350 23030 410
rect 23090 350 23130 410
rect 22990 310 23130 350
rect 22990 250 23030 310
rect 23090 250 23130 310
rect 22990 230 23130 250
rect 23160 410 23300 430
rect 23160 350 23200 410
rect 23260 350 23300 410
rect 23160 310 23300 350
rect 23160 250 23200 310
rect 23260 250 23300 310
rect 23160 230 23300 250
rect 23330 410 23470 430
rect 23330 350 23370 410
rect 23430 350 23470 410
rect 23330 310 23470 350
rect 23330 250 23370 310
rect 23430 250 23470 310
rect 23330 230 23470 250
rect 23500 410 23640 430
rect 23500 350 23540 410
rect 23600 350 23640 410
rect 23500 310 23640 350
rect 23500 250 23540 310
rect 23600 250 23640 310
rect 23500 230 23640 250
rect 23670 410 23810 430
rect 23670 350 23710 410
rect 23770 350 23810 410
rect 23670 310 23810 350
rect 23670 250 23710 310
rect 23770 250 23810 310
rect 23670 230 23810 250
rect 23840 410 23980 430
rect 23840 350 23880 410
rect 23940 350 23980 410
rect 23840 310 23980 350
rect 23840 250 23880 310
rect 23940 250 23980 310
rect 23840 230 23980 250
rect 24010 410 24150 430
rect 24010 350 24050 410
rect 24110 350 24150 410
rect 24010 310 24150 350
rect 24010 250 24050 310
rect 24110 250 24150 310
rect 24010 230 24150 250
rect 24180 410 24320 430
rect 24180 350 24220 410
rect 24280 350 24320 410
rect 24180 310 24320 350
rect 24180 250 24220 310
rect 24280 250 24320 310
rect 24180 230 24320 250
rect 24350 410 24490 430
rect 24350 350 24390 410
rect 24450 350 24490 410
rect 24350 310 24490 350
rect 24350 250 24390 310
rect 24450 250 24490 310
rect 24350 230 24490 250
rect 24520 410 24660 430
rect 24520 350 24560 410
rect 24620 350 24660 410
rect 24520 310 24660 350
rect 24520 250 24560 310
rect 24620 250 24660 310
rect 24520 230 24660 250
rect 24690 410 24830 430
rect 24690 350 24730 410
rect 24790 350 24830 410
rect 24690 310 24830 350
rect 24690 250 24730 310
rect 24790 250 24830 310
rect 24690 230 24830 250
rect 24860 410 25000 430
rect 24860 350 24900 410
rect 24960 350 25000 410
rect 24860 310 25000 350
rect 24860 250 24900 310
rect 24960 250 25000 310
rect 24860 230 25000 250
rect 25030 410 25170 430
rect 25030 350 25070 410
rect 25130 350 25170 410
rect 25030 310 25170 350
rect 25030 250 25070 310
rect 25130 250 25170 310
rect 25030 230 25170 250
rect 25200 410 25340 430
rect 25200 350 25240 410
rect 25300 350 25340 410
rect 25200 310 25340 350
rect 25200 250 25240 310
rect 25300 250 25340 310
rect 25200 230 25340 250
rect 25370 410 25510 430
rect 25370 350 25410 410
rect 25470 350 25510 410
rect 25370 310 25510 350
rect 25370 250 25410 310
rect 25470 250 25510 310
rect 25370 230 25510 250
rect 25540 410 25680 430
rect 25540 350 25580 410
rect 25640 350 25680 410
rect 25540 310 25680 350
rect 25540 250 25580 310
rect 25640 250 25680 310
rect 25540 230 25680 250
rect 25710 410 25850 430
rect 25710 350 25750 410
rect 25810 350 25850 410
rect 25710 310 25850 350
rect 25710 250 25750 310
rect 25810 250 25850 310
rect 25710 230 25850 250
rect 25880 410 26020 430
rect 25880 350 25920 410
rect 25980 350 26020 410
rect 25880 310 26020 350
rect 25880 250 25920 310
rect 25980 250 26020 310
rect 25880 230 26020 250
rect 26050 410 26190 430
rect 26050 350 26090 410
rect 26150 350 26190 410
rect 26050 310 26190 350
rect 26050 250 26090 310
rect 26150 250 26190 310
rect 26050 230 26190 250
rect 26220 410 26360 430
rect 26220 350 26260 410
rect 26320 350 26360 410
rect 26220 310 26360 350
rect 26220 250 26260 310
rect 26320 250 26360 310
rect 26220 230 26360 250
rect 26390 410 26530 430
rect 26390 350 26430 410
rect 26490 350 26530 410
rect 26390 310 26530 350
rect 26390 250 26430 310
rect 26490 250 26530 310
rect 26390 230 26530 250
rect 26560 410 26700 430
rect 26560 350 26600 410
rect 26660 350 26700 410
rect 26560 310 26700 350
rect 26560 250 26600 310
rect 26660 250 26700 310
rect 26560 230 26700 250
rect 26730 410 26870 430
rect 26730 350 26770 410
rect 26830 350 26870 410
rect 26730 310 26870 350
rect 26730 250 26770 310
rect 26830 250 26870 310
rect 26730 230 26870 250
rect 26900 410 27040 430
rect 26900 350 26940 410
rect 27000 350 27040 410
rect 26900 310 27040 350
rect 26900 250 26940 310
rect 27000 250 27040 310
rect 26900 230 27040 250
rect 27070 410 27210 430
rect 27070 350 27110 410
rect 27170 350 27210 410
rect 27070 310 27210 350
rect 27070 250 27110 310
rect 27170 250 27210 310
rect 27070 230 27210 250
rect 27240 410 27380 430
rect 27240 350 27280 410
rect 27340 350 27380 410
rect 27240 310 27380 350
rect 27240 250 27280 310
rect 27340 250 27380 310
rect 27240 230 27380 250
rect 27410 410 27550 430
rect 27410 350 27450 410
rect 27510 350 27550 410
rect 27410 310 27550 350
rect 27410 250 27450 310
rect 27510 250 27550 310
rect 27410 230 27550 250
rect 27580 410 27720 430
rect 27580 350 27620 410
rect 27680 350 27720 410
rect 27580 310 27720 350
rect 27580 250 27620 310
rect 27680 250 27720 310
rect 27580 230 27720 250
rect 27750 410 27890 430
rect 27750 350 27790 410
rect 27850 350 27890 410
rect 27750 310 27890 350
rect 27750 250 27790 310
rect 27850 250 27890 310
rect 27750 230 27890 250
rect 27920 410 28060 430
rect 27920 350 27960 410
rect 28020 350 28060 410
rect 27920 310 28060 350
rect 27920 250 27960 310
rect 28020 250 28060 310
rect 27920 230 28060 250
rect 28090 410 28230 430
rect 28090 350 28130 410
rect 28190 350 28230 410
rect 28090 310 28230 350
rect 28090 250 28130 310
rect 28190 250 28230 310
rect 28090 230 28230 250
rect 28260 410 28400 430
rect 28260 350 28300 410
rect 28360 350 28400 410
rect 28260 310 28400 350
rect 28260 250 28300 310
rect 28360 250 28400 310
rect 28260 230 28400 250
rect 28430 410 28570 430
rect 28430 350 28470 410
rect 28530 350 28570 410
rect 28430 310 28570 350
rect 28430 250 28470 310
rect 28530 250 28570 310
rect 28430 230 28570 250
rect 28600 410 28740 430
rect 28600 350 28640 410
rect 28700 350 28740 410
rect 28600 310 28740 350
rect 28600 250 28640 310
rect 28700 250 28740 310
rect 28600 230 28740 250
rect 28770 410 28910 430
rect 28770 350 28810 410
rect 28870 350 28910 410
rect 28770 310 28910 350
rect 28770 250 28810 310
rect 28870 250 28910 310
rect 28770 230 28910 250
rect 28940 410 29080 430
rect 28940 350 28980 410
rect 29040 350 29080 410
rect 28940 310 29080 350
rect 28940 250 28980 310
rect 29040 250 29080 310
rect 28940 230 29080 250
rect 29110 410 29250 430
rect 29110 350 29150 410
rect 29210 350 29250 410
rect 29110 310 29250 350
rect 29110 250 29150 310
rect 29210 250 29250 310
rect 29110 230 29250 250
rect 29280 410 29420 430
rect 29280 350 29320 410
rect 29380 350 29420 410
rect 29280 310 29420 350
rect 29280 250 29320 310
rect 29380 250 29420 310
rect 29280 230 29420 250
rect 29450 410 29590 430
rect 29450 350 29490 410
rect 29550 350 29590 410
rect 29450 310 29590 350
rect 29450 250 29490 310
rect 29550 250 29590 310
rect 29450 230 29590 250
rect 29620 410 29760 430
rect 29620 350 29660 410
rect 29720 350 29760 410
rect 29620 310 29760 350
rect 29620 250 29660 310
rect 29720 250 29760 310
rect 29620 230 29760 250
rect 29790 410 29930 430
rect 29790 350 29830 410
rect 29890 350 29930 410
rect 29790 310 29930 350
rect 29790 250 29830 310
rect 29890 250 29930 310
rect 29790 230 29930 250
rect 29960 410 30100 430
rect 29960 350 30000 410
rect 30060 350 30100 410
rect 29960 310 30100 350
rect 29960 250 30000 310
rect 30060 250 30100 310
rect 29960 230 30100 250
rect 30130 410 30270 430
rect 30130 350 30170 410
rect 30230 350 30270 410
rect 30130 310 30270 350
rect 30130 250 30170 310
rect 30230 250 30270 310
rect 30130 230 30270 250
rect 30300 410 30440 430
rect 30300 350 30340 410
rect 30400 350 30440 410
rect 30300 310 30440 350
rect 30300 250 30340 310
rect 30400 250 30440 310
rect 30300 230 30440 250
rect 30470 410 30610 430
rect 30470 350 30510 410
rect 30570 350 30610 410
rect 30470 310 30610 350
rect 30470 250 30510 310
rect 30570 250 30610 310
rect 30470 230 30610 250
rect 30640 410 30780 430
rect 30640 350 30680 410
rect 30740 350 30780 410
rect 30640 310 30780 350
rect 30640 250 30680 310
rect 30740 250 30780 310
rect 30640 230 30780 250
rect 30810 410 30950 430
rect 30810 350 30850 410
rect 30910 350 30950 410
rect 30810 310 30950 350
rect 30810 250 30850 310
rect 30910 250 30950 310
rect 30810 230 30950 250
rect 30980 410 31120 430
rect 30980 350 31020 410
rect 31080 350 31120 410
rect 30980 310 31120 350
rect 30980 250 31020 310
rect 31080 250 31120 310
rect 30980 230 31120 250
rect 31150 410 31290 430
rect 31150 350 31190 410
rect 31250 350 31290 410
rect 31150 310 31290 350
rect 31150 250 31190 310
rect 31250 250 31290 310
rect 31150 230 31290 250
rect 31320 410 31460 430
rect 31320 350 31360 410
rect 31420 350 31460 410
rect 31320 310 31460 350
rect 31320 250 31360 310
rect 31420 250 31460 310
rect 31320 230 31460 250
rect 31490 410 31630 430
rect 31490 350 31530 410
rect 31590 350 31630 410
rect 31490 310 31630 350
rect 31490 250 31530 310
rect 31590 250 31630 310
rect 31490 230 31630 250
rect 31660 410 31800 430
rect 31660 350 31700 410
rect 31760 350 31800 410
rect 31660 310 31800 350
rect 31660 250 31700 310
rect 31760 250 31800 310
rect 31660 230 31800 250
rect 31830 410 31970 430
rect 31830 350 31870 410
rect 31930 350 31970 410
rect 31830 310 31970 350
rect 31830 250 31870 310
rect 31930 250 31970 310
rect 31830 230 31970 250
rect 32000 410 32140 430
rect 32000 350 32040 410
rect 32100 350 32140 410
rect 32000 310 32140 350
rect 32000 250 32040 310
rect 32100 250 32140 310
rect 32000 230 32140 250
rect 32170 410 32310 430
rect 32170 350 32210 410
rect 32270 350 32310 410
rect 32170 310 32310 350
rect 32170 250 32210 310
rect 32270 250 32310 310
rect 32170 230 32310 250
rect 32340 410 32480 430
rect 32340 350 32380 410
rect 32440 350 32480 410
rect 32340 310 32480 350
rect 32340 250 32380 310
rect 32440 250 32480 310
rect 32340 230 32480 250
rect 32510 410 32650 430
rect 32510 350 32550 410
rect 32610 350 32650 410
rect 32510 310 32650 350
rect 32510 250 32550 310
rect 32610 250 32650 310
rect 32510 230 32650 250
rect 32680 410 32820 430
rect 32680 350 32720 410
rect 32780 350 32820 410
rect 32680 310 32820 350
rect 32680 250 32720 310
rect 32780 250 32820 310
rect 32680 230 32820 250
rect 32850 410 32990 430
rect 32850 350 32890 410
rect 32950 350 32990 410
rect 32850 310 32990 350
rect 32850 250 32890 310
rect 32950 250 32990 310
rect 32850 230 32990 250
rect 33020 410 33160 430
rect 33020 350 33060 410
rect 33120 350 33160 410
rect 33020 310 33160 350
rect 33020 250 33060 310
rect 33120 250 33160 310
rect 33020 230 33160 250
rect 33190 410 33330 430
rect 33190 350 33230 410
rect 33290 350 33330 410
rect 33190 310 33330 350
rect 33190 250 33230 310
rect 33290 250 33330 310
rect 33190 230 33330 250
rect 33360 410 33500 430
rect 33360 350 33400 410
rect 33460 350 33500 410
rect 33360 310 33500 350
rect 33360 250 33400 310
rect 33460 250 33500 310
rect 33360 230 33500 250
rect 33530 410 33670 430
rect 33530 350 33570 410
rect 33630 350 33670 410
rect 33530 310 33670 350
rect 33530 250 33570 310
rect 33630 250 33670 310
rect 33530 230 33670 250
rect 33700 410 33840 430
rect 33700 350 33740 410
rect 33800 350 33840 410
rect 33700 310 33840 350
rect 33700 250 33740 310
rect 33800 250 33840 310
rect 33700 230 33840 250
rect 33870 410 34010 430
rect 33870 350 33910 410
rect 33970 350 34010 410
rect 33870 310 34010 350
rect 33870 250 33910 310
rect 33970 250 34010 310
rect 33870 230 34010 250
rect 34040 410 34180 430
rect 34040 350 34080 410
rect 34140 350 34180 410
rect 34040 310 34180 350
rect 34040 250 34080 310
rect 34140 250 34180 310
rect 34040 230 34180 250
rect 34210 410 34350 430
rect 34210 350 34250 410
rect 34310 350 34350 410
rect 34210 310 34350 350
rect 34210 250 34250 310
rect 34310 250 34350 310
rect 34210 230 34350 250
rect 34380 410 34520 430
rect 34380 350 34420 410
rect 34480 350 34520 410
rect 34380 310 34520 350
rect 34380 250 34420 310
rect 34480 250 34520 310
rect 34380 230 34520 250
rect 34550 410 34690 430
rect 34550 350 34590 410
rect 34650 350 34690 410
rect 34550 310 34690 350
rect 34550 250 34590 310
rect 34650 250 34690 310
rect 34550 230 34690 250
rect 34720 410 34860 430
rect 34720 350 34760 410
rect 34820 350 34860 410
rect 34720 310 34860 350
rect 34720 250 34760 310
rect 34820 250 34860 310
rect 34720 230 34860 250
rect 34890 410 35030 430
rect 34890 350 34930 410
rect 34990 350 35030 410
rect 34890 310 35030 350
rect 34890 250 34930 310
rect 34990 250 35030 310
rect 34890 230 35030 250
rect 35060 410 35200 430
rect 35060 350 35100 410
rect 35160 350 35200 410
rect 35060 310 35200 350
rect 35060 250 35100 310
rect 35160 250 35200 310
rect 35060 230 35200 250
rect 35230 410 35370 430
rect 35230 350 35270 410
rect 35330 350 35370 410
rect 35230 310 35370 350
rect 35230 250 35270 310
rect 35330 250 35370 310
rect 35230 230 35370 250
rect 35400 410 35540 430
rect 35400 350 35440 410
rect 35500 350 35540 410
rect 35400 310 35540 350
rect 35400 250 35440 310
rect 35500 250 35540 310
rect 35400 230 35540 250
rect 35570 410 35710 430
rect 35570 350 35610 410
rect 35670 350 35710 410
rect 35570 310 35710 350
rect 35570 250 35610 310
rect 35670 250 35710 310
rect 35570 230 35710 250
rect 35740 410 35880 430
rect 35740 350 35780 410
rect 35840 350 35880 410
rect 35740 310 35880 350
rect 35740 250 35780 310
rect 35840 250 35880 310
rect 35740 230 35880 250
rect 35910 410 36050 430
rect 35910 350 35950 410
rect 36010 350 36050 410
rect 35910 310 36050 350
rect 35910 250 35950 310
rect 36010 250 36050 310
rect 35910 230 36050 250
rect 36080 410 36220 430
rect 36080 350 36120 410
rect 36180 350 36220 410
rect 36080 310 36220 350
rect 36080 250 36120 310
rect 36180 250 36220 310
rect 36080 230 36220 250
rect 36250 410 36390 430
rect 36250 350 36290 410
rect 36350 350 36390 410
rect 36250 310 36390 350
rect 36250 250 36290 310
rect 36350 250 36390 310
rect 36250 230 36390 250
rect 36420 410 36560 430
rect 36420 350 36460 410
rect 36520 350 36560 410
rect 36420 310 36560 350
rect 36420 250 36460 310
rect 36520 250 36560 310
rect 36420 230 36560 250
rect 36590 410 36730 430
rect 36590 350 36630 410
rect 36690 350 36730 410
rect 36590 310 36730 350
rect 36590 250 36630 310
rect 36690 250 36730 310
rect 36590 230 36730 250
rect 36760 410 36900 430
rect 36760 350 36800 410
rect 36860 350 36900 410
rect 36760 310 36900 350
rect 36760 250 36800 310
rect 36860 250 36900 310
rect 36760 230 36900 250
rect 36930 410 37070 430
rect 36930 350 36970 410
rect 37030 350 37070 410
rect 36930 310 37070 350
rect 36930 250 36970 310
rect 37030 250 37070 310
rect 36930 230 37070 250
rect 37100 410 37240 430
rect 37100 350 37140 410
rect 37200 350 37240 410
rect 37100 310 37240 350
rect 37100 250 37140 310
rect 37200 250 37240 310
rect 37100 230 37240 250
rect 37270 410 37410 430
rect 37270 350 37310 410
rect 37370 350 37410 410
rect 37270 310 37410 350
rect 37270 250 37310 310
rect 37370 250 37410 310
rect 37270 230 37410 250
rect 37440 410 37580 430
rect 37440 350 37480 410
rect 37540 350 37580 410
rect 37440 310 37580 350
rect 37440 250 37480 310
rect 37540 250 37580 310
rect 37440 230 37580 250
rect 37610 410 37750 430
rect 37610 350 37650 410
rect 37710 350 37750 410
rect 37610 310 37750 350
rect 37610 250 37650 310
rect 37710 250 37750 310
rect 37610 230 37750 250
rect 37780 410 37920 430
rect 37780 350 37820 410
rect 37880 350 37920 410
rect 37780 310 37920 350
rect 37780 250 37820 310
rect 37880 250 37920 310
rect 37780 230 37920 250
rect 37950 410 38090 430
rect 37950 350 37990 410
rect 38050 350 38090 410
rect 37950 310 38090 350
rect 37950 250 37990 310
rect 38050 250 38090 310
rect 37950 230 38090 250
rect 38120 410 38260 430
rect 38120 350 38160 410
rect 38220 350 38260 410
rect 38120 310 38260 350
rect 38120 250 38160 310
rect 38220 250 38260 310
rect 38120 230 38260 250
rect 38290 410 38430 430
rect 38290 350 38330 410
rect 38390 350 38430 410
rect 38290 310 38430 350
rect 38290 250 38330 310
rect 38390 250 38430 310
rect 38290 230 38430 250
rect 38460 410 38600 430
rect 38460 350 38500 410
rect 38560 350 38600 410
rect 38460 310 38600 350
rect 38460 250 38500 310
rect 38560 250 38600 310
rect 38460 230 38600 250
rect 38630 410 38770 430
rect 38630 350 38670 410
rect 38730 350 38770 410
rect 38630 310 38770 350
rect 38630 250 38670 310
rect 38730 250 38770 310
rect 38630 230 38770 250
rect 38800 410 38940 430
rect 38800 350 38840 410
rect 38900 350 38940 410
rect 38800 310 38940 350
rect 38800 250 38840 310
rect 38900 250 38940 310
rect 38800 230 38940 250
rect 38970 410 39110 430
rect 38970 350 39010 410
rect 39070 350 39110 410
rect 38970 310 39110 350
rect 38970 250 39010 310
rect 39070 250 39110 310
rect 38970 230 39110 250
rect 39140 410 39280 430
rect 39140 350 39180 410
rect 39240 350 39280 410
rect 39140 310 39280 350
rect 39140 250 39180 310
rect 39240 250 39280 310
rect 39140 230 39280 250
rect 39310 410 39450 430
rect 39310 350 39350 410
rect 39410 350 39450 410
rect 39310 310 39450 350
rect 39310 250 39350 310
rect 39410 250 39450 310
rect 39310 230 39450 250
rect 39480 410 39620 430
rect 39480 350 39520 410
rect 39580 350 39620 410
rect 39480 310 39620 350
rect 39480 250 39520 310
rect 39580 250 39620 310
rect 39480 230 39620 250
rect 39650 410 39790 430
rect 39650 350 39690 410
rect 39750 350 39790 410
rect 39650 310 39790 350
rect 39650 250 39690 310
rect 39750 250 39790 310
rect 39650 230 39790 250
rect 39820 410 39960 430
rect 39820 350 39860 410
rect 39920 350 39960 410
rect 39820 310 39960 350
rect 39820 250 39860 310
rect 39920 250 39960 310
rect 39820 230 39960 250
rect 39990 410 40130 430
rect 39990 350 40030 410
rect 40090 350 40130 410
rect 39990 310 40130 350
rect 39990 250 40030 310
rect 40090 250 40130 310
rect 39990 230 40130 250
rect 40160 410 40300 430
rect 40160 350 40200 410
rect 40260 350 40300 410
rect 40160 310 40300 350
rect 40160 250 40200 310
rect 40260 250 40300 310
rect 40160 230 40300 250
rect 40330 410 40470 430
rect 40330 350 40370 410
rect 40430 350 40470 410
rect 40330 310 40470 350
rect 40330 250 40370 310
rect 40430 250 40470 310
rect 40330 230 40470 250
rect 40500 410 40640 430
rect 40500 350 40540 410
rect 40600 350 40640 410
rect 40500 310 40640 350
rect 40500 250 40540 310
rect 40600 250 40640 310
rect 40500 230 40640 250
rect 40670 410 40810 430
rect 40670 350 40710 410
rect 40770 350 40810 410
rect 40670 310 40810 350
rect 40670 250 40710 310
rect 40770 250 40810 310
rect 40670 230 40810 250
rect 40840 410 40980 430
rect 40840 350 40880 410
rect 40940 350 40980 410
rect 40840 310 40980 350
rect 40840 250 40880 310
rect 40940 250 40980 310
rect 40840 230 40980 250
rect 41010 410 41150 430
rect 41010 350 41050 410
rect 41110 350 41150 410
rect 41010 310 41150 350
rect 41010 250 41050 310
rect 41110 250 41150 310
rect 41010 230 41150 250
rect 41180 410 41320 430
rect 41180 350 41220 410
rect 41280 350 41320 410
rect 41180 310 41320 350
rect 41180 250 41220 310
rect 41280 250 41320 310
rect 41180 230 41320 250
rect 41350 410 41490 430
rect 41350 350 41390 410
rect 41450 350 41490 410
rect 41350 310 41490 350
rect 41350 250 41390 310
rect 41450 250 41490 310
rect 41350 230 41490 250
rect 41520 410 41660 430
rect 41520 350 41560 410
rect 41620 350 41660 410
rect 41520 310 41660 350
rect 41520 250 41560 310
rect 41620 250 41660 310
rect 41520 230 41660 250
rect 41690 410 41830 430
rect 41690 350 41730 410
rect 41790 350 41830 410
rect 41690 310 41830 350
rect 41690 250 41730 310
rect 41790 250 41830 310
rect 41690 230 41830 250
rect 41860 410 42000 430
rect 41860 350 41900 410
rect 41960 350 42000 410
rect 41860 310 42000 350
rect 41860 250 41900 310
rect 41960 250 42000 310
rect 41860 230 42000 250
rect 42030 410 42170 430
rect 42030 350 42070 410
rect 42130 350 42170 410
rect 42030 310 42170 350
rect 42030 250 42070 310
rect 42130 250 42170 310
rect 42030 230 42170 250
rect 42200 410 42340 430
rect 42200 350 42240 410
rect 42300 350 42340 410
rect 42200 310 42340 350
rect 42200 250 42240 310
rect 42300 250 42340 310
rect 42200 230 42340 250
rect 42370 410 42510 430
rect 42370 350 42410 410
rect 42470 350 42510 410
rect 42370 310 42510 350
rect 42370 250 42410 310
rect 42470 250 42510 310
rect 42370 230 42510 250
rect 42540 410 42680 430
rect 42540 350 42580 410
rect 42640 350 42680 410
rect 42540 310 42680 350
rect 42540 250 42580 310
rect 42640 250 42680 310
rect 42540 230 42680 250
rect 42710 410 42850 430
rect 42710 350 42750 410
rect 42810 350 42850 410
rect 42710 310 42850 350
rect 42710 250 42750 310
rect 42810 250 42850 310
rect 42710 230 42850 250
rect 42880 410 43020 430
rect 42880 350 42920 410
rect 42980 350 43020 410
rect 42880 310 43020 350
rect 42880 250 42920 310
rect 42980 250 43020 310
rect 42880 230 43020 250
rect 43050 410 43190 430
rect 43050 350 43090 410
rect 43150 350 43190 410
rect 43050 310 43190 350
rect 43050 250 43090 310
rect 43150 250 43190 310
rect 43050 230 43190 250
rect 43220 410 43360 430
rect 43220 350 43260 410
rect 43320 350 43360 410
rect 43220 310 43360 350
rect 43220 250 43260 310
rect 43320 250 43360 310
rect 43220 230 43360 250
rect 43390 410 43530 430
rect 43390 350 43430 410
rect 43490 350 43530 410
rect 43390 310 43530 350
rect 43390 250 43430 310
rect 43490 250 43530 310
rect 43390 230 43530 250
rect 43560 410 43700 430
rect 43560 350 43600 410
rect 43660 350 43700 410
rect 43560 310 43700 350
rect 43560 250 43600 310
rect 43660 250 43700 310
rect 43560 230 43700 250
rect 43730 410 43870 430
rect 43730 350 43770 410
rect 43830 350 43870 410
rect 43730 310 43870 350
rect 43730 250 43770 310
rect 43830 250 43870 310
rect 43730 230 43870 250
rect 43900 410 44040 430
rect 43900 350 43940 410
rect 44000 350 44040 410
rect 43900 310 44040 350
rect 43900 250 43940 310
rect 44000 250 44040 310
rect 43900 230 44040 250
rect 44070 410 44210 430
rect 44070 350 44110 410
rect 44170 350 44210 410
rect 44070 310 44210 350
rect 44070 250 44110 310
rect 44170 250 44210 310
rect 44070 230 44210 250
rect 44240 410 44380 430
rect 44240 350 44280 410
rect 44340 350 44380 410
rect 44240 310 44380 350
rect 44240 250 44280 310
rect 44340 250 44380 310
rect 44240 230 44380 250
rect 44410 410 44550 430
rect 44410 350 44450 410
rect 44510 350 44550 410
rect 44410 310 44550 350
rect 44410 250 44450 310
rect 44510 250 44550 310
rect 44410 230 44550 250
rect 44580 410 44720 430
rect 44580 350 44620 410
rect 44680 350 44720 410
rect 44580 310 44720 350
rect 44580 250 44620 310
rect 44680 250 44720 310
rect 44580 230 44720 250
rect 44750 410 44890 430
rect 44750 350 44790 410
rect 44850 350 44890 410
rect 44750 310 44890 350
rect 44750 250 44790 310
rect 44850 250 44890 310
rect 44750 230 44890 250
rect 44920 410 45060 430
rect 44920 350 44960 410
rect 45020 350 45060 410
rect 44920 310 45060 350
rect 44920 250 44960 310
rect 45020 250 45060 310
rect 44920 230 45060 250
rect 45090 410 45230 430
rect 45090 350 45130 410
rect 45190 350 45230 410
rect 45090 310 45230 350
rect 45090 250 45130 310
rect 45190 250 45230 310
rect 45090 230 45230 250
rect 45260 410 45400 430
rect 45260 350 45300 410
rect 45360 350 45400 410
rect 45260 310 45400 350
rect 45260 250 45300 310
rect 45360 250 45400 310
rect 45260 230 45400 250
rect 45430 410 45570 430
rect 45430 350 45470 410
rect 45530 350 45570 410
rect 45430 310 45570 350
rect 45430 250 45470 310
rect 45530 250 45570 310
rect 45430 230 45570 250
rect 45600 410 45740 430
rect 45600 350 45640 410
rect 45700 350 45740 410
rect 45600 310 45740 350
rect 45600 250 45640 310
rect 45700 250 45740 310
rect 45600 230 45740 250
rect 45770 410 45910 430
rect 45770 350 45810 410
rect 45870 350 45910 410
rect 45770 310 45910 350
rect 45770 250 45810 310
rect 45870 250 45910 310
rect 45770 230 45910 250
rect 45940 410 46080 430
rect 45940 350 45980 410
rect 46040 350 46080 410
rect 45940 310 46080 350
rect 45940 250 45980 310
rect 46040 250 46080 310
rect 45940 230 46080 250
rect 46110 410 46250 430
rect 46110 350 46150 410
rect 46210 350 46250 410
rect 46110 310 46250 350
rect 46110 250 46150 310
rect 46210 250 46250 310
rect 46110 230 46250 250
rect 46280 410 46420 430
rect 46280 350 46320 410
rect 46380 350 46420 410
rect 46280 310 46420 350
rect 46280 250 46320 310
rect 46380 250 46420 310
rect 46280 230 46420 250
rect 46450 410 46590 430
rect 46450 350 46490 410
rect 46550 350 46590 410
rect 46450 310 46590 350
rect 46450 250 46490 310
rect 46550 250 46590 310
rect 46450 230 46590 250
rect 46620 410 46760 430
rect 46620 350 46660 410
rect 46720 350 46760 410
rect 46620 310 46760 350
rect 46620 250 46660 310
rect 46720 250 46760 310
rect 46620 230 46760 250
rect 46790 410 46930 430
rect 46790 350 46830 410
rect 46890 350 46930 410
rect 46790 310 46930 350
rect 46790 250 46830 310
rect 46890 250 46930 310
rect 46790 230 46930 250
rect 46960 410 47100 430
rect 46960 350 47000 410
rect 47060 350 47100 410
rect 46960 310 47100 350
rect 46960 250 47000 310
rect 47060 250 47100 310
rect 46960 230 47100 250
rect 47130 410 47270 430
rect 47130 350 47170 410
rect 47230 350 47270 410
rect 47130 310 47270 350
rect 47130 250 47170 310
rect 47230 250 47270 310
rect 47130 230 47270 250
rect 47300 410 47440 430
rect 47300 350 47340 410
rect 47400 350 47440 410
rect 47300 310 47440 350
rect 47300 250 47340 310
rect 47400 250 47440 310
rect 47300 230 47440 250
rect 47470 410 47610 430
rect 47470 350 47510 410
rect 47570 350 47610 410
rect 47470 310 47610 350
rect 47470 250 47510 310
rect 47570 250 47610 310
rect 47470 230 47610 250
rect 47640 410 47780 430
rect 47640 350 47680 410
rect 47740 350 47780 410
rect 47640 310 47780 350
rect 47640 250 47680 310
rect 47740 250 47780 310
rect 47640 230 47780 250
rect 47810 410 47950 430
rect 47810 350 47850 410
rect 47910 350 47950 410
rect 47810 310 47950 350
rect 47810 250 47850 310
rect 47910 250 47950 310
rect 47810 230 47950 250
rect 47980 410 48120 430
rect 47980 350 48020 410
rect 48080 350 48120 410
rect 47980 310 48120 350
rect 47980 250 48020 310
rect 48080 250 48120 310
rect 47980 230 48120 250
rect 48150 410 48290 430
rect 48150 350 48190 410
rect 48250 350 48290 410
rect 48150 310 48290 350
rect 48150 250 48190 310
rect 48250 250 48290 310
rect 48150 230 48290 250
rect 48320 410 48460 430
rect 48320 350 48360 410
rect 48420 350 48460 410
rect 48320 310 48460 350
rect 48320 250 48360 310
rect 48420 250 48460 310
rect 48320 230 48460 250
rect 48490 410 48630 430
rect 48490 350 48530 410
rect 48590 350 48630 410
rect 48490 310 48630 350
rect 48490 250 48530 310
rect 48590 250 48630 310
rect 48490 230 48630 250
rect 48660 410 48800 430
rect 48660 350 48700 410
rect 48760 350 48800 410
rect 48660 310 48800 350
rect 48660 250 48700 310
rect 48760 250 48800 310
rect 48660 230 48800 250
rect 48830 410 48970 430
rect 48830 350 48870 410
rect 48930 350 48970 410
rect 48830 310 48970 350
rect 48830 250 48870 310
rect 48930 250 48970 310
rect 48830 230 48970 250
rect 49000 410 49140 430
rect 49000 350 49040 410
rect 49100 350 49140 410
rect 49000 310 49140 350
rect 49000 250 49040 310
rect 49100 250 49140 310
rect 49000 230 49140 250
rect 49170 410 49310 430
rect 49170 350 49210 410
rect 49270 350 49310 410
rect 49170 310 49310 350
rect 49170 250 49210 310
rect 49270 250 49310 310
rect 49170 230 49310 250
rect 49340 410 49480 430
rect 49340 350 49380 410
rect 49440 350 49480 410
rect 49340 310 49480 350
rect 49340 250 49380 310
rect 49440 250 49480 310
rect 49340 230 49480 250
rect 49510 410 49650 430
rect 49510 350 49550 410
rect 49610 350 49650 410
rect 49510 310 49650 350
rect 49510 250 49550 310
rect 49610 250 49650 310
rect 49510 230 49650 250
rect 49680 410 49820 430
rect 49680 350 49720 410
rect 49780 350 49820 410
rect 49680 310 49820 350
rect 49680 250 49720 310
rect 49780 250 49820 310
rect 49680 230 49820 250
rect 49850 410 49990 430
rect 49850 350 49890 410
rect 49950 350 49990 410
rect 49850 310 49990 350
rect 49850 250 49890 310
rect 49950 250 49990 310
rect 49850 230 49990 250
rect 50020 410 50160 430
rect 50020 350 50060 410
rect 50120 350 50160 410
rect 50020 310 50160 350
rect 50020 250 50060 310
rect 50120 250 50160 310
rect 50020 230 50160 250
rect 50190 410 50330 430
rect 50190 350 50230 410
rect 50290 350 50330 410
rect 50190 310 50330 350
rect 50190 250 50230 310
rect 50290 250 50330 310
rect 50190 230 50330 250
rect 50360 410 50500 430
rect 50360 350 50400 410
rect 50460 350 50500 410
rect 50360 310 50500 350
rect 50360 250 50400 310
rect 50460 250 50500 310
rect 50360 230 50500 250
rect 50530 410 50670 430
rect 50530 350 50570 410
rect 50630 350 50670 410
rect 50530 310 50670 350
rect 50530 250 50570 310
rect 50630 250 50670 310
rect 50530 230 50670 250
rect 50700 410 50840 430
rect 50700 350 50740 410
rect 50800 350 50840 410
rect 50700 310 50840 350
rect 50700 250 50740 310
rect 50800 250 50840 310
rect 50700 230 50840 250
rect 50870 410 51010 430
rect 50870 350 50910 410
rect 50970 350 51010 410
rect 50870 310 51010 350
rect 50870 250 50910 310
rect 50970 250 51010 310
rect 50870 230 51010 250
rect 51040 410 51180 430
rect 51040 350 51080 410
rect 51140 350 51180 410
rect 51040 310 51180 350
rect 51040 250 51080 310
rect 51140 250 51180 310
rect 51040 230 51180 250
rect 51210 410 51350 430
rect 51210 350 51250 410
rect 51310 350 51350 410
rect 51210 310 51350 350
rect 51210 250 51250 310
rect 51310 250 51350 310
rect 51210 230 51350 250
rect 51380 410 51520 430
rect 51380 350 51420 410
rect 51480 350 51520 410
rect 51380 310 51520 350
rect 51380 250 51420 310
rect 51480 250 51520 310
rect 51380 230 51520 250
rect 51550 410 51690 430
rect 51550 350 51590 410
rect 51650 350 51690 410
rect 51550 310 51690 350
rect 51550 250 51590 310
rect 51650 250 51690 310
rect 51550 230 51690 250
rect 51720 410 51860 430
rect 51720 350 51760 410
rect 51820 350 51860 410
rect 51720 310 51860 350
rect 51720 250 51760 310
rect 51820 250 51860 310
rect 51720 230 51860 250
rect 51890 410 52030 430
rect 51890 350 51930 410
rect 51990 350 52030 410
rect 51890 310 52030 350
rect 51890 250 51930 310
rect 51990 250 52030 310
rect 51890 230 52030 250
rect 52060 410 52200 430
rect 52060 350 52100 410
rect 52160 350 52200 410
rect 52060 310 52200 350
rect 52060 250 52100 310
rect 52160 250 52200 310
rect 52060 230 52200 250
rect 52230 410 52370 430
rect 52230 350 52270 410
rect 52330 350 52370 410
rect 52230 310 52370 350
rect 52230 250 52270 310
rect 52330 250 52370 310
rect 52230 230 52370 250
rect 52400 410 52540 430
rect 52400 350 52440 410
rect 52500 350 52540 410
rect 52400 310 52540 350
rect 52400 250 52440 310
rect 52500 250 52540 310
rect 52400 230 52540 250
rect 52570 410 52710 430
rect 52570 350 52610 410
rect 52670 350 52710 410
rect 52570 310 52710 350
rect 52570 250 52610 310
rect 52670 250 52710 310
rect 52570 230 52710 250
rect 52740 410 52880 430
rect 52740 350 52780 410
rect 52840 350 52880 410
rect 52740 310 52880 350
rect 52740 250 52780 310
rect 52840 250 52880 310
rect 52740 230 52880 250
rect 52910 410 53050 430
rect 52910 350 52950 410
rect 53010 350 53050 410
rect 52910 310 53050 350
rect 52910 250 52950 310
rect 53010 250 53050 310
rect 52910 230 53050 250
rect 53080 410 53220 430
rect 53080 350 53120 410
rect 53180 350 53220 410
rect 53080 310 53220 350
rect 53080 250 53120 310
rect 53180 250 53220 310
rect 53080 230 53220 250
rect 53250 410 53390 430
rect 53250 350 53290 410
rect 53350 350 53390 410
rect 53250 310 53390 350
rect 53250 250 53290 310
rect 53350 250 53390 310
rect 53250 230 53390 250
rect 53420 410 53560 430
rect 53420 350 53460 410
rect 53520 350 53560 410
rect 53420 310 53560 350
rect 53420 250 53460 310
rect 53520 250 53560 310
rect 53420 230 53560 250
rect 53590 410 53730 430
rect 53590 350 53630 410
rect 53690 350 53730 410
rect 53590 310 53730 350
rect 53590 250 53630 310
rect 53690 250 53730 310
rect 53590 230 53730 250
rect 53760 410 53900 430
rect 53760 350 53800 410
rect 53860 350 53900 410
rect 53760 310 53900 350
rect 53760 250 53800 310
rect 53860 250 53900 310
rect 53760 230 53900 250
rect 53930 410 54070 430
rect 53930 350 53970 410
rect 54030 350 54070 410
rect 53930 310 54070 350
rect 53930 250 53970 310
rect 54030 250 54070 310
rect 53930 230 54070 250
rect 54100 410 54240 430
rect 54100 350 54140 410
rect 54200 350 54240 410
rect 54100 310 54240 350
rect 54100 250 54140 310
rect 54200 250 54240 310
rect 54100 230 54240 250
rect 54270 410 54410 430
rect 54270 350 54310 410
rect 54370 350 54410 410
rect 54270 310 54410 350
rect 54270 250 54310 310
rect 54370 250 54410 310
rect 54270 230 54410 250
rect 54440 410 54580 430
rect 54440 350 54480 410
rect 54540 350 54580 410
rect 54440 310 54580 350
rect 54440 250 54480 310
rect 54540 250 54580 310
rect 54440 230 54580 250
rect 54610 410 54750 430
rect 54610 350 54650 410
rect 54710 350 54750 410
rect 54610 310 54750 350
rect 54610 250 54650 310
rect 54710 250 54750 310
rect 54610 230 54750 250
rect 54780 410 54920 430
rect 54780 350 54820 410
rect 54880 350 54920 410
rect 54780 310 54920 350
rect 54780 250 54820 310
rect 54880 250 54920 310
rect 54780 230 54920 250
rect 54950 410 55090 430
rect 54950 350 54990 410
rect 55050 350 55090 410
rect 54950 310 55090 350
rect 54950 250 54990 310
rect 55050 250 55090 310
rect 54950 230 55090 250
rect 55120 410 55260 430
rect 55120 350 55160 410
rect 55220 350 55260 410
rect 55120 310 55260 350
rect 55120 250 55160 310
rect 55220 250 55260 310
rect 55120 230 55260 250
rect 55290 410 55430 430
rect 55290 350 55330 410
rect 55390 350 55430 410
rect 55290 310 55430 350
rect 55290 250 55330 310
rect 55390 250 55430 310
rect 55290 230 55430 250
rect 55460 410 55600 430
rect 55460 350 55500 410
rect 55560 350 55600 410
rect 55460 310 55600 350
rect 55460 250 55500 310
rect 55560 250 55600 310
rect 55460 230 55600 250
rect 55630 410 55770 430
rect 55630 350 55670 410
rect 55730 350 55770 410
rect 55630 310 55770 350
rect 55630 250 55670 310
rect 55730 250 55770 310
rect 55630 230 55770 250
rect 55800 410 55940 430
rect 55800 350 55840 410
rect 55900 350 55940 410
rect 55800 310 55940 350
rect 55800 250 55840 310
rect 55900 250 55940 310
rect 55800 230 55940 250
rect 55970 410 56110 430
rect 55970 350 56010 410
rect 56070 350 56110 410
rect 55970 310 56110 350
rect 55970 250 56010 310
rect 56070 250 56110 310
rect 55970 230 56110 250
rect 56140 410 56280 430
rect 56140 350 56180 410
rect 56240 350 56280 410
rect 56140 310 56280 350
rect 56140 250 56180 310
rect 56240 250 56280 310
rect 56140 230 56280 250
rect 56310 410 56450 430
rect 56310 350 56350 410
rect 56410 350 56450 410
rect 56310 310 56450 350
rect 56310 250 56350 310
rect 56410 250 56450 310
rect 56310 230 56450 250
rect 56480 410 56620 430
rect 56480 350 56520 410
rect 56580 350 56620 410
rect 56480 310 56620 350
rect 56480 250 56520 310
rect 56580 250 56620 310
rect 56480 230 56620 250
rect 56650 410 56790 430
rect 56650 350 56690 410
rect 56750 350 56790 410
rect 56650 310 56790 350
rect 56650 250 56690 310
rect 56750 250 56790 310
rect 56650 230 56790 250
rect 56820 410 56960 430
rect 56820 350 56860 410
rect 56920 350 56960 410
rect 56820 310 56960 350
rect 56820 250 56860 310
rect 56920 250 56960 310
rect 56820 230 56960 250
rect 56990 410 57130 430
rect 56990 350 57030 410
rect 57090 350 57130 410
rect 56990 310 57130 350
rect 56990 250 57030 310
rect 57090 250 57130 310
rect 56990 230 57130 250
rect 57160 410 57300 430
rect 57160 350 57200 410
rect 57260 350 57300 410
rect 57160 310 57300 350
rect 57160 250 57200 310
rect 57260 250 57300 310
rect 57160 230 57300 250
rect 57330 410 57470 430
rect 57330 350 57370 410
rect 57430 350 57470 410
rect 57330 310 57470 350
rect 57330 250 57370 310
rect 57430 250 57470 310
rect 57330 230 57470 250
rect 57500 410 57640 430
rect 57500 350 57540 410
rect 57600 350 57640 410
rect 57500 310 57640 350
rect 57500 250 57540 310
rect 57600 250 57640 310
rect 57500 230 57640 250
rect 57670 410 57810 430
rect 57670 350 57710 410
rect 57770 350 57810 410
rect 57670 310 57810 350
rect 57670 250 57710 310
rect 57770 250 57810 310
rect 57670 230 57810 250
rect 57840 410 57980 430
rect 57840 350 57880 410
rect 57940 350 57980 410
rect 57840 310 57980 350
rect 57840 250 57880 310
rect 57940 250 57980 310
rect 57840 230 57980 250
rect 58010 410 58150 430
rect 58010 350 58050 410
rect 58110 350 58150 410
rect 58010 310 58150 350
rect 58010 250 58050 310
rect 58110 250 58150 310
rect 58010 230 58150 250
rect 58180 410 58320 430
rect 58180 350 58220 410
rect 58280 350 58320 410
rect 58180 310 58320 350
rect 58180 250 58220 310
rect 58280 250 58320 310
rect 58180 230 58320 250
rect 58350 410 58490 430
rect 58350 350 58390 410
rect 58450 350 58490 410
rect 58350 310 58490 350
rect 58350 250 58390 310
rect 58450 250 58490 310
rect 58350 230 58490 250
rect 58520 410 58660 430
rect 58520 350 58560 410
rect 58620 350 58660 410
rect 58520 310 58660 350
rect 58520 250 58560 310
rect 58620 250 58660 310
rect 58520 230 58660 250
rect 58690 410 58830 430
rect 58690 350 58730 410
rect 58790 350 58830 410
rect 58690 310 58830 350
rect 58690 250 58730 310
rect 58790 250 58830 310
rect 58690 230 58830 250
rect 58860 410 59000 430
rect 58860 350 58900 410
rect 58960 350 59000 410
rect 58860 310 59000 350
rect 58860 250 58900 310
rect 58960 250 59000 310
rect 58860 230 59000 250
rect 59030 410 59170 430
rect 59030 350 59070 410
rect 59130 350 59170 410
rect 59030 310 59170 350
rect 59030 250 59070 310
rect 59130 250 59170 310
rect 59030 230 59170 250
rect 59200 410 59340 430
rect 59200 350 59240 410
rect 59300 350 59340 410
rect 59200 310 59340 350
rect 59200 250 59240 310
rect 59300 250 59340 310
rect 59200 230 59340 250
rect 110 -1000 250 -980
rect 110 -1060 150 -1000
rect 210 -1060 250 -1000
rect 110 -1100 250 -1060
rect 110 -1160 150 -1100
rect 210 -1160 250 -1100
rect 110 -1200 250 -1160
rect 110 -1260 150 -1200
rect 210 -1260 250 -1200
rect 110 -1300 250 -1260
rect 110 -1360 150 -1300
rect 210 -1360 250 -1300
rect 110 -1380 250 -1360
rect 280 -1000 420 -980
rect 280 -1060 320 -1000
rect 380 -1060 420 -1000
rect 280 -1100 420 -1060
rect 280 -1160 320 -1100
rect 380 -1160 420 -1100
rect 280 -1200 420 -1160
rect 280 -1260 320 -1200
rect 380 -1260 420 -1200
rect 280 -1300 420 -1260
rect 280 -1360 320 -1300
rect 380 -1360 420 -1300
rect 280 -1380 420 -1360
rect 450 -1000 590 -980
rect 450 -1060 490 -1000
rect 550 -1060 590 -1000
rect 450 -1100 590 -1060
rect 450 -1160 490 -1100
rect 550 -1160 590 -1100
rect 450 -1200 590 -1160
rect 450 -1260 490 -1200
rect 550 -1260 590 -1200
rect 450 -1300 590 -1260
rect 450 -1360 490 -1300
rect 550 -1360 590 -1300
rect 450 -1380 590 -1360
rect 620 -1000 760 -980
rect 620 -1060 660 -1000
rect 720 -1060 760 -1000
rect 620 -1100 760 -1060
rect 620 -1160 660 -1100
rect 720 -1160 760 -1100
rect 620 -1200 760 -1160
rect 620 -1260 660 -1200
rect 720 -1260 760 -1200
rect 620 -1300 760 -1260
rect 620 -1360 660 -1300
rect 720 -1360 760 -1300
rect 620 -1380 760 -1360
rect 790 -1000 930 -980
rect 790 -1060 830 -1000
rect 890 -1060 930 -1000
rect 790 -1100 930 -1060
rect 790 -1160 830 -1100
rect 890 -1160 930 -1100
rect 790 -1200 930 -1160
rect 790 -1260 830 -1200
rect 890 -1260 930 -1200
rect 790 -1300 930 -1260
rect 790 -1360 830 -1300
rect 890 -1360 930 -1300
rect 790 -1380 930 -1360
rect 960 -1000 1100 -980
rect 960 -1060 1000 -1000
rect 1060 -1060 1100 -1000
rect 960 -1100 1100 -1060
rect 960 -1160 1000 -1100
rect 1060 -1160 1100 -1100
rect 960 -1200 1100 -1160
rect 960 -1260 1000 -1200
rect 1060 -1260 1100 -1200
rect 960 -1300 1100 -1260
rect 960 -1360 1000 -1300
rect 1060 -1360 1100 -1300
rect 960 -1380 1100 -1360
rect 1130 -1000 1270 -980
rect 1130 -1060 1170 -1000
rect 1230 -1060 1270 -1000
rect 1130 -1100 1270 -1060
rect 1130 -1160 1170 -1100
rect 1230 -1160 1270 -1100
rect 1130 -1200 1270 -1160
rect 1130 -1260 1170 -1200
rect 1230 -1260 1270 -1200
rect 1130 -1300 1270 -1260
rect 1130 -1360 1170 -1300
rect 1230 -1360 1270 -1300
rect 1130 -1380 1270 -1360
rect 1300 -1000 1440 -980
rect 1300 -1060 1340 -1000
rect 1400 -1060 1440 -1000
rect 1300 -1100 1440 -1060
rect 1300 -1160 1340 -1100
rect 1400 -1160 1440 -1100
rect 1300 -1200 1440 -1160
rect 1300 -1260 1340 -1200
rect 1400 -1260 1440 -1200
rect 1300 -1300 1440 -1260
rect 1300 -1360 1340 -1300
rect 1400 -1360 1440 -1300
rect 1300 -1380 1440 -1360
rect 1470 -1000 1610 -980
rect 1470 -1060 1510 -1000
rect 1570 -1060 1610 -1000
rect 1470 -1100 1610 -1060
rect 1470 -1160 1510 -1100
rect 1570 -1160 1610 -1100
rect 1470 -1200 1610 -1160
rect 1470 -1260 1510 -1200
rect 1570 -1260 1610 -1200
rect 1470 -1300 1610 -1260
rect 1470 -1360 1510 -1300
rect 1570 -1360 1610 -1300
rect 1470 -1380 1610 -1360
rect 1640 -1000 1780 -980
rect 1640 -1060 1680 -1000
rect 1740 -1060 1780 -1000
rect 1640 -1100 1780 -1060
rect 1640 -1160 1680 -1100
rect 1740 -1160 1780 -1100
rect 1640 -1200 1780 -1160
rect 1640 -1260 1680 -1200
rect 1740 -1260 1780 -1200
rect 1640 -1300 1780 -1260
rect 1640 -1360 1680 -1300
rect 1740 -1360 1780 -1300
rect 1640 -1380 1780 -1360
rect 1810 -1000 1950 -980
rect 1810 -1060 1850 -1000
rect 1910 -1060 1950 -1000
rect 1810 -1100 1950 -1060
rect 1810 -1160 1850 -1100
rect 1910 -1160 1950 -1100
rect 1810 -1200 1950 -1160
rect 1810 -1260 1850 -1200
rect 1910 -1260 1950 -1200
rect 1810 -1300 1950 -1260
rect 1810 -1360 1850 -1300
rect 1910 -1360 1950 -1300
rect 1810 -1380 1950 -1360
rect 1980 -1000 2120 -980
rect 1980 -1060 2020 -1000
rect 2080 -1060 2120 -1000
rect 1980 -1100 2120 -1060
rect 1980 -1160 2020 -1100
rect 2080 -1160 2120 -1100
rect 1980 -1200 2120 -1160
rect 1980 -1260 2020 -1200
rect 2080 -1260 2120 -1200
rect 1980 -1300 2120 -1260
rect 1980 -1360 2020 -1300
rect 2080 -1360 2120 -1300
rect 1980 -1380 2120 -1360
rect 2150 -1000 2290 -980
rect 2150 -1060 2190 -1000
rect 2250 -1060 2290 -1000
rect 2150 -1100 2290 -1060
rect 2150 -1160 2190 -1100
rect 2250 -1160 2290 -1100
rect 2150 -1200 2290 -1160
rect 2150 -1260 2190 -1200
rect 2250 -1260 2290 -1200
rect 2150 -1300 2290 -1260
rect 2150 -1360 2190 -1300
rect 2250 -1360 2290 -1300
rect 2150 -1380 2290 -1360
rect 2320 -1000 2460 -980
rect 2320 -1060 2360 -1000
rect 2420 -1060 2460 -1000
rect 2320 -1100 2460 -1060
rect 2320 -1160 2360 -1100
rect 2420 -1160 2460 -1100
rect 2320 -1200 2460 -1160
rect 2320 -1260 2360 -1200
rect 2420 -1260 2460 -1200
rect 2320 -1300 2460 -1260
rect 2320 -1360 2360 -1300
rect 2420 -1360 2460 -1300
rect 2320 -1380 2460 -1360
rect 2490 -1000 2630 -980
rect 2490 -1060 2530 -1000
rect 2590 -1060 2630 -1000
rect 2490 -1100 2630 -1060
rect 2490 -1160 2530 -1100
rect 2590 -1160 2630 -1100
rect 2490 -1200 2630 -1160
rect 2490 -1260 2530 -1200
rect 2590 -1260 2630 -1200
rect 2490 -1300 2630 -1260
rect 2490 -1360 2530 -1300
rect 2590 -1360 2630 -1300
rect 2490 -1380 2630 -1360
rect 2660 -1000 2800 -980
rect 2660 -1060 2700 -1000
rect 2760 -1060 2800 -1000
rect 2660 -1100 2800 -1060
rect 2660 -1160 2700 -1100
rect 2760 -1160 2800 -1100
rect 2660 -1200 2800 -1160
rect 2660 -1260 2700 -1200
rect 2760 -1260 2800 -1200
rect 2660 -1300 2800 -1260
rect 2660 -1360 2700 -1300
rect 2760 -1360 2800 -1300
rect 2660 -1380 2800 -1360
rect 2830 -1000 2970 -980
rect 2830 -1060 2870 -1000
rect 2930 -1060 2970 -1000
rect 2830 -1100 2970 -1060
rect 2830 -1160 2870 -1100
rect 2930 -1160 2970 -1100
rect 2830 -1200 2970 -1160
rect 2830 -1260 2870 -1200
rect 2930 -1260 2970 -1200
rect 2830 -1300 2970 -1260
rect 2830 -1360 2870 -1300
rect 2930 -1360 2970 -1300
rect 2830 -1380 2970 -1360
rect 3000 -1000 3140 -980
rect 3000 -1060 3040 -1000
rect 3100 -1060 3140 -1000
rect 3000 -1100 3140 -1060
rect 3000 -1160 3040 -1100
rect 3100 -1160 3140 -1100
rect 3000 -1200 3140 -1160
rect 3000 -1260 3040 -1200
rect 3100 -1260 3140 -1200
rect 3000 -1300 3140 -1260
rect 3000 -1360 3040 -1300
rect 3100 -1360 3140 -1300
rect 3000 -1380 3140 -1360
rect 3170 -1000 3310 -980
rect 3170 -1060 3210 -1000
rect 3270 -1060 3310 -1000
rect 3170 -1100 3310 -1060
rect 3170 -1160 3210 -1100
rect 3270 -1160 3310 -1100
rect 3170 -1200 3310 -1160
rect 3170 -1260 3210 -1200
rect 3270 -1260 3310 -1200
rect 3170 -1300 3310 -1260
rect 3170 -1360 3210 -1300
rect 3270 -1360 3310 -1300
rect 3170 -1380 3310 -1360
rect 3340 -1000 3480 -980
rect 3340 -1060 3380 -1000
rect 3440 -1060 3480 -1000
rect 3340 -1100 3480 -1060
rect 3340 -1160 3380 -1100
rect 3440 -1160 3480 -1100
rect 3340 -1200 3480 -1160
rect 3340 -1260 3380 -1200
rect 3440 -1260 3480 -1200
rect 3340 -1300 3480 -1260
rect 3340 -1360 3380 -1300
rect 3440 -1360 3480 -1300
rect 3340 -1380 3480 -1360
rect 3510 -1000 3650 -980
rect 3510 -1060 3550 -1000
rect 3610 -1060 3650 -1000
rect 3510 -1100 3650 -1060
rect 3510 -1160 3550 -1100
rect 3610 -1160 3650 -1100
rect 3510 -1200 3650 -1160
rect 3510 -1260 3550 -1200
rect 3610 -1260 3650 -1200
rect 3510 -1300 3650 -1260
rect 3510 -1360 3550 -1300
rect 3610 -1360 3650 -1300
rect 3510 -1380 3650 -1360
rect 3680 -1000 3820 -980
rect 3680 -1060 3720 -1000
rect 3780 -1060 3820 -1000
rect 3680 -1100 3820 -1060
rect 3680 -1160 3720 -1100
rect 3780 -1160 3820 -1100
rect 3680 -1200 3820 -1160
rect 3680 -1260 3720 -1200
rect 3780 -1260 3820 -1200
rect 3680 -1300 3820 -1260
rect 3680 -1360 3720 -1300
rect 3780 -1360 3820 -1300
rect 3680 -1380 3820 -1360
rect 3850 -1000 3990 -980
rect 3850 -1060 3890 -1000
rect 3950 -1060 3990 -1000
rect 3850 -1100 3990 -1060
rect 3850 -1160 3890 -1100
rect 3950 -1160 3990 -1100
rect 3850 -1200 3990 -1160
rect 3850 -1260 3890 -1200
rect 3950 -1260 3990 -1200
rect 3850 -1300 3990 -1260
rect 3850 -1360 3890 -1300
rect 3950 -1360 3990 -1300
rect 3850 -1380 3990 -1360
rect 4020 -1000 4160 -980
rect 4020 -1060 4060 -1000
rect 4120 -1060 4160 -1000
rect 4020 -1100 4160 -1060
rect 4020 -1160 4060 -1100
rect 4120 -1160 4160 -1100
rect 4020 -1200 4160 -1160
rect 4020 -1260 4060 -1200
rect 4120 -1260 4160 -1200
rect 4020 -1300 4160 -1260
rect 4020 -1360 4060 -1300
rect 4120 -1360 4160 -1300
rect 4020 -1380 4160 -1360
rect 4190 -1000 4330 -980
rect 4190 -1060 4230 -1000
rect 4290 -1060 4330 -1000
rect 4190 -1100 4330 -1060
rect 4190 -1160 4230 -1100
rect 4290 -1160 4330 -1100
rect 4190 -1200 4330 -1160
rect 4190 -1260 4230 -1200
rect 4290 -1260 4330 -1200
rect 4190 -1300 4330 -1260
rect 4190 -1360 4230 -1300
rect 4290 -1360 4330 -1300
rect 4190 -1380 4330 -1360
rect 4360 -1000 4500 -980
rect 4360 -1060 4400 -1000
rect 4460 -1060 4500 -1000
rect 4360 -1100 4500 -1060
rect 4360 -1160 4400 -1100
rect 4460 -1160 4500 -1100
rect 4360 -1200 4500 -1160
rect 4360 -1260 4400 -1200
rect 4460 -1260 4500 -1200
rect 4360 -1300 4500 -1260
rect 4360 -1360 4400 -1300
rect 4460 -1360 4500 -1300
rect 4360 -1380 4500 -1360
rect 4530 -1000 4670 -980
rect 4530 -1060 4570 -1000
rect 4630 -1060 4670 -1000
rect 4530 -1100 4670 -1060
rect 4530 -1160 4570 -1100
rect 4630 -1160 4670 -1100
rect 4530 -1200 4670 -1160
rect 4530 -1260 4570 -1200
rect 4630 -1260 4670 -1200
rect 4530 -1300 4670 -1260
rect 4530 -1360 4570 -1300
rect 4630 -1360 4670 -1300
rect 4530 -1380 4670 -1360
rect 4700 -1000 4840 -980
rect 4700 -1060 4740 -1000
rect 4800 -1060 4840 -1000
rect 4700 -1100 4840 -1060
rect 4700 -1160 4740 -1100
rect 4800 -1160 4840 -1100
rect 4700 -1200 4840 -1160
rect 4700 -1260 4740 -1200
rect 4800 -1260 4840 -1200
rect 4700 -1300 4840 -1260
rect 4700 -1360 4740 -1300
rect 4800 -1360 4840 -1300
rect 4700 -1380 4840 -1360
rect 4870 -1000 5010 -980
rect 4870 -1060 4910 -1000
rect 4970 -1060 5010 -1000
rect 4870 -1100 5010 -1060
rect 4870 -1160 4910 -1100
rect 4970 -1160 5010 -1100
rect 4870 -1200 5010 -1160
rect 4870 -1260 4910 -1200
rect 4970 -1260 5010 -1200
rect 4870 -1300 5010 -1260
rect 4870 -1360 4910 -1300
rect 4970 -1360 5010 -1300
rect 4870 -1380 5010 -1360
rect 5040 -1000 5180 -980
rect 5040 -1060 5080 -1000
rect 5140 -1060 5180 -1000
rect 5040 -1100 5180 -1060
rect 5040 -1160 5080 -1100
rect 5140 -1160 5180 -1100
rect 5040 -1200 5180 -1160
rect 5040 -1260 5080 -1200
rect 5140 -1260 5180 -1200
rect 5040 -1300 5180 -1260
rect 5040 -1360 5080 -1300
rect 5140 -1360 5180 -1300
rect 5040 -1380 5180 -1360
rect 5210 -1000 5350 -980
rect 5210 -1060 5250 -1000
rect 5310 -1060 5350 -1000
rect 5210 -1100 5350 -1060
rect 5210 -1160 5250 -1100
rect 5310 -1160 5350 -1100
rect 5210 -1200 5350 -1160
rect 5210 -1260 5250 -1200
rect 5310 -1260 5350 -1200
rect 5210 -1300 5350 -1260
rect 5210 -1360 5250 -1300
rect 5310 -1360 5350 -1300
rect 5210 -1380 5350 -1360
rect 5380 -1000 5520 -980
rect 5380 -1060 5420 -1000
rect 5480 -1060 5520 -1000
rect 5380 -1100 5520 -1060
rect 5380 -1160 5420 -1100
rect 5480 -1160 5520 -1100
rect 5380 -1200 5520 -1160
rect 5380 -1260 5420 -1200
rect 5480 -1260 5520 -1200
rect 5380 -1300 5520 -1260
rect 5380 -1360 5420 -1300
rect 5480 -1360 5520 -1300
rect 5380 -1380 5520 -1360
rect 5550 -1000 5690 -980
rect 5550 -1060 5590 -1000
rect 5650 -1060 5690 -1000
rect 5550 -1100 5690 -1060
rect 5550 -1160 5590 -1100
rect 5650 -1160 5690 -1100
rect 5550 -1200 5690 -1160
rect 5550 -1260 5590 -1200
rect 5650 -1260 5690 -1200
rect 5550 -1300 5690 -1260
rect 5550 -1360 5590 -1300
rect 5650 -1360 5690 -1300
rect 5550 -1380 5690 -1360
rect 5720 -1000 5860 -980
rect 5720 -1060 5760 -1000
rect 5820 -1060 5860 -1000
rect 5720 -1100 5860 -1060
rect 5720 -1160 5760 -1100
rect 5820 -1160 5860 -1100
rect 5720 -1200 5860 -1160
rect 5720 -1260 5760 -1200
rect 5820 -1260 5860 -1200
rect 5720 -1300 5860 -1260
rect 5720 -1360 5760 -1300
rect 5820 -1360 5860 -1300
rect 5720 -1380 5860 -1360
rect 5890 -1000 6030 -980
rect 5890 -1060 5930 -1000
rect 5990 -1060 6030 -1000
rect 5890 -1100 6030 -1060
rect 5890 -1160 5930 -1100
rect 5990 -1160 6030 -1100
rect 5890 -1200 6030 -1160
rect 5890 -1260 5930 -1200
rect 5990 -1260 6030 -1200
rect 5890 -1300 6030 -1260
rect 5890 -1360 5930 -1300
rect 5990 -1360 6030 -1300
rect 5890 -1380 6030 -1360
rect 6060 -1000 6200 -980
rect 6060 -1060 6100 -1000
rect 6160 -1060 6200 -1000
rect 6060 -1100 6200 -1060
rect 6060 -1160 6100 -1100
rect 6160 -1160 6200 -1100
rect 6060 -1200 6200 -1160
rect 6060 -1260 6100 -1200
rect 6160 -1260 6200 -1200
rect 6060 -1300 6200 -1260
rect 6060 -1360 6100 -1300
rect 6160 -1360 6200 -1300
rect 6060 -1380 6200 -1360
rect 6230 -1000 6370 -980
rect 6230 -1060 6270 -1000
rect 6330 -1060 6370 -1000
rect 6230 -1100 6370 -1060
rect 6230 -1160 6270 -1100
rect 6330 -1160 6370 -1100
rect 6230 -1200 6370 -1160
rect 6230 -1260 6270 -1200
rect 6330 -1260 6370 -1200
rect 6230 -1300 6370 -1260
rect 6230 -1360 6270 -1300
rect 6330 -1360 6370 -1300
rect 6230 -1380 6370 -1360
rect 6400 -1000 6540 -980
rect 6400 -1060 6440 -1000
rect 6500 -1060 6540 -1000
rect 6400 -1100 6540 -1060
rect 6400 -1160 6440 -1100
rect 6500 -1160 6540 -1100
rect 6400 -1200 6540 -1160
rect 6400 -1260 6440 -1200
rect 6500 -1260 6540 -1200
rect 6400 -1300 6540 -1260
rect 6400 -1360 6440 -1300
rect 6500 -1360 6540 -1300
rect 6400 -1380 6540 -1360
rect 6570 -1000 6710 -980
rect 6570 -1060 6610 -1000
rect 6670 -1060 6710 -1000
rect 6570 -1100 6710 -1060
rect 6570 -1160 6610 -1100
rect 6670 -1160 6710 -1100
rect 6570 -1200 6710 -1160
rect 6570 -1260 6610 -1200
rect 6670 -1260 6710 -1200
rect 6570 -1300 6710 -1260
rect 6570 -1360 6610 -1300
rect 6670 -1360 6710 -1300
rect 6570 -1380 6710 -1360
rect 6740 -1000 6880 -980
rect 6740 -1060 6780 -1000
rect 6840 -1060 6880 -1000
rect 6740 -1100 6880 -1060
rect 6740 -1160 6780 -1100
rect 6840 -1160 6880 -1100
rect 6740 -1200 6880 -1160
rect 6740 -1260 6780 -1200
rect 6840 -1260 6880 -1200
rect 6740 -1300 6880 -1260
rect 6740 -1360 6780 -1300
rect 6840 -1360 6880 -1300
rect 6740 -1380 6880 -1360
rect 6910 -1000 7050 -980
rect 6910 -1060 6950 -1000
rect 7010 -1060 7050 -1000
rect 6910 -1100 7050 -1060
rect 6910 -1160 6950 -1100
rect 7010 -1160 7050 -1100
rect 6910 -1200 7050 -1160
rect 6910 -1260 6950 -1200
rect 7010 -1260 7050 -1200
rect 6910 -1300 7050 -1260
rect 6910 -1360 6950 -1300
rect 7010 -1360 7050 -1300
rect 6910 -1380 7050 -1360
rect 7080 -1000 7220 -980
rect 7080 -1060 7120 -1000
rect 7180 -1060 7220 -1000
rect 7080 -1100 7220 -1060
rect 7080 -1160 7120 -1100
rect 7180 -1160 7220 -1100
rect 7080 -1200 7220 -1160
rect 7080 -1260 7120 -1200
rect 7180 -1260 7220 -1200
rect 7080 -1300 7220 -1260
rect 7080 -1360 7120 -1300
rect 7180 -1360 7220 -1300
rect 7080 -1380 7220 -1360
rect 7250 -1000 7390 -980
rect 7250 -1060 7290 -1000
rect 7350 -1060 7390 -1000
rect 7250 -1100 7390 -1060
rect 7250 -1160 7290 -1100
rect 7350 -1160 7390 -1100
rect 7250 -1200 7390 -1160
rect 7250 -1260 7290 -1200
rect 7350 -1260 7390 -1200
rect 7250 -1300 7390 -1260
rect 7250 -1360 7290 -1300
rect 7350 -1360 7390 -1300
rect 7250 -1380 7390 -1360
rect 7420 -1000 7560 -980
rect 7420 -1060 7460 -1000
rect 7520 -1060 7560 -1000
rect 7420 -1100 7560 -1060
rect 7420 -1160 7460 -1100
rect 7520 -1160 7560 -1100
rect 7420 -1200 7560 -1160
rect 7420 -1260 7460 -1200
rect 7520 -1260 7560 -1200
rect 7420 -1300 7560 -1260
rect 7420 -1360 7460 -1300
rect 7520 -1360 7560 -1300
rect 7420 -1380 7560 -1360
rect 7590 -1000 7730 -980
rect 7590 -1060 7630 -1000
rect 7690 -1060 7730 -1000
rect 7590 -1100 7730 -1060
rect 7590 -1160 7630 -1100
rect 7690 -1160 7730 -1100
rect 7590 -1200 7730 -1160
rect 7590 -1260 7630 -1200
rect 7690 -1260 7730 -1200
rect 7590 -1300 7730 -1260
rect 7590 -1360 7630 -1300
rect 7690 -1360 7730 -1300
rect 7590 -1380 7730 -1360
rect 7760 -1000 7900 -980
rect 7760 -1060 7800 -1000
rect 7860 -1060 7900 -1000
rect 7760 -1100 7900 -1060
rect 7760 -1160 7800 -1100
rect 7860 -1160 7900 -1100
rect 7760 -1200 7900 -1160
rect 7760 -1260 7800 -1200
rect 7860 -1260 7900 -1200
rect 7760 -1300 7900 -1260
rect 7760 -1360 7800 -1300
rect 7860 -1360 7900 -1300
rect 7760 -1380 7900 -1360
rect 7930 -1000 8070 -980
rect 7930 -1060 7970 -1000
rect 8030 -1060 8070 -1000
rect 7930 -1100 8070 -1060
rect 7930 -1160 7970 -1100
rect 8030 -1160 8070 -1100
rect 7930 -1200 8070 -1160
rect 7930 -1260 7970 -1200
rect 8030 -1260 8070 -1200
rect 7930 -1300 8070 -1260
rect 7930 -1360 7970 -1300
rect 8030 -1360 8070 -1300
rect 7930 -1380 8070 -1360
rect 8100 -1000 8240 -980
rect 8100 -1060 8140 -1000
rect 8200 -1060 8240 -1000
rect 8100 -1100 8240 -1060
rect 8100 -1160 8140 -1100
rect 8200 -1160 8240 -1100
rect 8100 -1200 8240 -1160
rect 8100 -1260 8140 -1200
rect 8200 -1260 8240 -1200
rect 8100 -1300 8240 -1260
rect 8100 -1360 8140 -1300
rect 8200 -1360 8240 -1300
rect 8100 -1380 8240 -1360
rect 8270 -1000 8410 -980
rect 8270 -1060 8310 -1000
rect 8370 -1060 8410 -1000
rect 8270 -1100 8410 -1060
rect 8270 -1160 8310 -1100
rect 8370 -1160 8410 -1100
rect 8270 -1200 8410 -1160
rect 8270 -1260 8310 -1200
rect 8370 -1260 8410 -1200
rect 8270 -1300 8410 -1260
rect 8270 -1360 8310 -1300
rect 8370 -1360 8410 -1300
rect 8270 -1380 8410 -1360
rect 8440 -1000 8580 -980
rect 8440 -1060 8480 -1000
rect 8540 -1060 8580 -1000
rect 8440 -1100 8580 -1060
rect 8440 -1160 8480 -1100
rect 8540 -1160 8580 -1100
rect 8440 -1200 8580 -1160
rect 8440 -1260 8480 -1200
rect 8540 -1260 8580 -1200
rect 8440 -1300 8580 -1260
rect 8440 -1360 8480 -1300
rect 8540 -1360 8580 -1300
rect 8440 -1380 8580 -1360
rect 8610 -1000 8750 -980
rect 8610 -1060 8650 -1000
rect 8710 -1060 8750 -1000
rect 8610 -1100 8750 -1060
rect 8610 -1160 8650 -1100
rect 8710 -1160 8750 -1100
rect 8610 -1200 8750 -1160
rect 8610 -1260 8650 -1200
rect 8710 -1260 8750 -1200
rect 8610 -1300 8750 -1260
rect 8610 -1360 8650 -1300
rect 8710 -1360 8750 -1300
rect 8610 -1380 8750 -1360
rect 8780 -1000 8920 -980
rect 8780 -1060 8820 -1000
rect 8880 -1060 8920 -1000
rect 8780 -1100 8920 -1060
rect 8780 -1160 8820 -1100
rect 8880 -1160 8920 -1100
rect 8780 -1200 8920 -1160
rect 8780 -1260 8820 -1200
rect 8880 -1260 8920 -1200
rect 8780 -1300 8920 -1260
rect 8780 -1360 8820 -1300
rect 8880 -1360 8920 -1300
rect 8780 -1380 8920 -1360
rect 8950 -1000 9090 -980
rect 8950 -1060 8990 -1000
rect 9050 -1060 9090 -1000
rect 8950 -1100 9090 -1060
rect 8950 -1160 8990 -1100
rect 9050 -1160 9090 -1100
rect 8950 -1200 9090 -1160
rect 8950 -1260 8990 -1200
rect 9050 -1260 9090 -1200
rect 8950 -1300 9090 -1260
rect 8950 -1360 8990 -1300
rect 9050 -1360 9090 -1300
rect 8950 -1380 9090 -1360
rect 9120 -1000 9260 -980
rect 9120 -1060 9160 -1000
rect 9220 -1060 9260 -1000
rect 9120 -1100 9260 -1060
rect 9120 -1160 9160 -1100
rect 9220 -1160 9260 -1100
rect 9120 -1200 9260 -1160
rect 9120 -1260 9160 -1200
rect 9220 -1260 9260 -1200
rect 9120 -1300 9260 -1260
rect 9120 -1360 9160 -1300
rect 9220 -1360 9260 -1300
rect 9120 -1380 9260 -1360
rect 9290 -1000 9430 -980
rect 9290 -1060 9330 -1000
rect 9390 -1060 9430 -1000
rect 9290 -1100 9430 -1060
rect 9290 -1160 9330 -1100
rect 9390 -1160 9430 -1100
rect 9290 -1200 9430 -1160
rect 9290 -1260 9330 -1200
rect 9390 -1260 9430 -1200
rect 9290 -1300 9430 -1260
rect 9290 -1360 9330 -1300
rect 9390 -1360 9430 -1300
rect 9290 -1380 9430 -1360
rect 9460 -1000 9600 -980
rect 9460 -1060 9500 -1000
rect 9560 -1060 9600 -1000
rect 9460 -1100 9600 -1060
rect 9460 -1160 9500 -1100
rect 9560 -1160 9600 -1100
rect 9460 -1200 9600 -1160
rect 9460 -1260 9500 -1200
rect 9560 -1260 9600 -1200
rect 9460 -1300 9600 -1260
rect 9460 -1360 9500 -1300
rect 9560 -1360 9600 -1300
rect 9460 -1380 9600 -1360
rect 9630 -1000 9770 -980
rect 9630 -1060 9670 -1000
rect 9730 -1060 9770 -1000
rect 9630 -1100 9770 -1060
rect 9630 -1160 9670 -1100
rect 9730 -1160 9770 -1100
rect 9630 -1200 9770 -1160
rect 9630 -1260 9670 -1200
rect 9730 -1260 9770 -1200
rect 9630 -1300 9770 -1260
rect 9630 -1360 9670 -1300
rect 9730 -1360 9770 -1300
rect 9630 -1380 9770 -1360
rect 9800 -1000 9940 -980
rect 9800 -1060 9840 -1000
rect 9900 -1060 9940 -1000
rect 9800 -1100 9940 -1060
rect 9800 -1160 9840 -1100
rect 9900 -1160 9940 -1100
rect 9800 -1200 9940 -1160
rect 9800 -1260 9840 -1200
rect 9900 -1260 9940 -1200
rect 9800 -1300 9940 -1260
rect 9800 -1360 9840 -1300
rect 9900 -1360 9940 -1300
rect 9800 -1380 9940 -1360
rect 9970 -1000 10110 -980
rect 9970 -1060 10010 -1000
rect 10070 -1060 10110 -1000
rect 9970 -1100 10110 -1060
rect 9970 -1160 10010 -1100
rect 10070 -1160 10110 -1100
rect 9970 -1200 10110 -1160
rect 9970 -1260 10010 -1200
rect 10070 -1260 10110 -1200
rect 9970 -1300 10110 -1260
rect 9970 -1360 10010 -1300
rect 10070 -1360 10110 -1300
rect 9970 -1380 10110 -1360
rect 10140 -1000 10280 -980
rect 10140 -1060 10180 -1000
rect 10240 -1060 10280 -1000
rect 10140 -1100 10280 -1060
rect 10140 -1160 10180 -1100
rect 10240 -1160 10280 -1100
rect 10140 -1200 10280 -1160
rect 10140 -1260 10180 -1200
rect 10240 -1260 10280 -1200
rect 10140 -1300 10280 -1260
rect 10140 -1360 10180 -1300
rect 10240 -1360 10280 -1300
rect 10140 -1380 10280 -1360
rect 10310 -1000 10450 -980
rect 10310 -1060 10350 -1000
rect 10410 -1060 10450 -1000
rect 10310 -1100 10450 -1060
rect 10310 -1160 10350 -1100
rect 10410 -1160 10450 -1100
rect 10310 -1200 10450 -1160
rect 10310 -1260 10350 -1200
rect 10410 -1260 10450 -1200
rect 10310 -1300 10450 -1260
rect 10310 -1360 10350 -1300
rect 10410 -1360 10450 -1300
rect 10310 -1380 10450 -1360
rect 10480 -1000 10620 -980
rect 10480 -1060 10520 -1000
rect 10580 -1060 10620 -1000
rect 10480 -1100 10620 -1060
rect 10480 -1160 10520 -1100
rect 10580 -1160 10620 -1100
rect 10480 -1200 10620 -1160
rect 10480 -1260 10520 -1200
rect 10580 -1260 10620 -1200
rect 10480 -1300 10620 -1260
rect 10480 -1360 10520 -1300
rect 10580 -1360 10620 -1300
rect 10480 -1380 10620 -1360
rect 10650 -1000 10790 -980
rect 10650 -1060 10690 -1000
rect 10750 -1060 10790 -1000
rect 10650 -1100 10790 -1060
rect 10650 -1160 10690 -1100
rect 10750 -1160 10790 -1100
rect 10650 -1200 10790 -1160
rect 10650 -1260 10690 -1200
rect 10750 -1260 10790 -1200
rect 10650 -1300 10790 -1260
rect 10650 -1360 10690 -1300
rect 10750 -1360 10790 -1300
rect 10650 -1380 10790 -1360
rect 10820 -1000 10960 -980
rect 10820 -1060 10860 -1000
rect 10920 -1060 10960 -1000
rect 10820 -1100 10960 -1060
rect 10820 -1160 10860 -1100
rect 10920 -1160 10960 -1100
rect 10820 -1200 10960 -1160
rect 10820 -1260 10860 -1200
rect 10920 -1260 10960 -1200
rect 10820 -1300 10960 -1260
rect 10820 -1360 10860 -1300
rect 10920 -1360 10960 -1300
rect 10820 -1380 10960 -1360
rect 10990 -1000 11130 -980
rect 10990 -1060 11030 -1000
rect 11090 -1060 11130 -1000
rect 10990 -1100 11130 -1060
rect 10990 -1160 11030 -1100
rect 11090 -1160 11130 -1100
rect 10990 -1200 11130 -1160
rect 10990 -1260 11030 -1200
rect 11090 -1260 11130 -1200
rect 10990 -1300 11130 -1260
rect 10990 -1360 11030 -1300
rect 11090 -1360 11130 -1300
rect 10990 -1380 11130 -1360
rect 11160 -1000 11300 -980
rect 11160 -1060 11200 -1000
rect 11260 -1060 11300 -1000
rect 11160 -1100 11300 -1060
rect 11160 -1160 11200 -1100
rect 11260 -1160 11300 -1100
rect 11160 -1200 11300 -1160
rect 11160 -1260 11200 -1200
rect 11260 -1260 11300 -1200
rect 11160 -1300 11300 -1260
rect 11160 -1360 11200 -1300
rect 11260 -1360 11300 -1300
rect 11160 -1380 11300 -1360
rect 11330 -1000 11470 -980
rect 11330 -1060 11370 -1000
rect 11430 -1060 11470 -1000
rect 11330 -1100 11470 -1060
rect 11330 -1160 11370 -1100
rect 11430 -1160 11470 -1100
rect 11330 -1200 11470 -1160
rect 11330 -1260 11370 -1200
rect 11430 -1260 11470 -1200
rect 11330 -1300 11470 -1260
rect 11330 -1360 11370 -1300
rect 11430 -1360 11470 -1300
rect 11330 -1380 11470 -1360
rect 11500 -1000 11640 -980
rect 11500 -1060 11540 -1000
rect 11600 -1060 11640 -1000
rect 11500 -1100 11640 -1060
rect 11500 -1160 11540 -1100
rect 11600 -1160 11640 -1100
rect 11500 -1200 11640 -1160
rect 11500 -1260 11540 -1200
rect 11600 -1260 11640 -1200
rect 11500 -1300 11640 -1260
rect 11500 -1360 11540 -1300
rect 11600 -1360 11640 -1300
rect 11500 -1380 11640 -1360
rect 11670 -1000 11810 -980
rect 11670 -1060 11710 -1000
rect 11770 -1060 11810 -1000
rect 11670 -1100 11810 -1060
rect 11670 -1160 11710 -1100
rect 11770 -1160 11810 -1100
rect 11670 -1200 11810 -1160
rect 11670 -1260 11710 -1200
rect 11770 -1260 11810 -1200
rect 11670 -1300 11810 -1260
rect 11670 -1360 11710 -1300
rect 11770 -1360 11810 -1300
rect 11670 -1380 11810 -1360
rect 11840 -1000 11980 -980
rect 11840 -1060 11880 -1000
rect 11940 -1060 11980 -1000
rect 11840 -1100 11980 -1060
rect 11840 -1160 11880 -1100
rect 11940 -1160 11980 -1100
rect 11840 -1200 11980 -1160
rect 11840 -1260 11880 -1200
rect 11940 -1260 11980 -1200
rect 11840 -1300 11980 -1260
rect 11840 -1360 11880 -1300
rect 11940 -1360 11980 -1300
rect 11840 -1380 11980 -1360
rect 12010 -1000 12150 -980
rect 12010 -1060 12050 -1000
rect 12110 -1060 12150 -1000
rect 12010 -1100 12150 -1060
rect 12010 -1160 12050 -1100
rect 12110 -1160 12150 -1100
rect 12010 -1200 12150 -1160
rect 12010 -1260 12050 -1200
rect 12110 -1260 12150 -1200
rect 12010 -1300 12150 -1260
rect 12010 -1360 12050 -1300
rect 12110 -1360 12150 -1300
rect 12010 -1380 12150 -1360
rect 12180 -1000 12320 -980
rect 12180 -1060 12220 -1000
rect 12280 -1060 12320 -1000
rect 12180 -1100 12320 -1060
rect 12180 -1160 12220 -1100
rect 12280 -1160 12320 -1100
rect 12180 -1200 12320 -1160
rect 12180 -1260 12220 -1200
rect 12280 -1260 12320 -1200
rect 12180 -1300 12320 -1260
rect 12180 -1360 12220 -1300
rect 12280 -1360 12320 -1300
rect 12180 -1380 12320 -1360
rect 12350 -1000 12490 -980
rect 12350 -1060 12390 -1000
rect 12450 -1060 12490 -1000
rect 12350 -1100 12490 -1060
rect 12350 -1160 12390 -1100
rect 12450 -1160 12490 -1100
rect 12350 -1200 12490 -1160
rect 12350 -1260 12390 -1200
rect 12450 -1260 12490 -1200
rect 12350 -1300 12490 -1260
rect 12350 -1360 12390 -1300
rect 12450 -1360 12490 -1300
rect 12350 -1380 12490 -1360
rect 12520 -1000 12660 -980
rect 12520 -1060 12560 -1000
rect 12620 -1060 12660 -1000
rect 12520 -1100 12660 -1060
rect 12520 -1160 12560 -1100
rect 12620 -1160 12660 -1100
rect 12520 -1200 12660 -1160
rect 12520 -1260 12560 -1200
rect 12620 -1260 12660 -1200
rect 12520 -1300 12660 -1260
rect 12520 -1360 12560 -1300
rect 12620 -1360 12660 -1300
rect 12520 -1380 12660 -1360
rect 12690 -1000 12830 -980
rect 12690 -1060 12730 -1000
rect 12790 -1060 12830 -1000
rect 12690 -1100 12830 -1060
rect 12690 -1160 12730 -1100
rect 12790 -1160 12830 -1100
rect 12690 -1200 12830 -1160
rect 12690 -1260 12730 -1200
rect 12790 -1260 12830 -1200
rect 12690 -1300 12830 -1260
rect 12690 -1360 12730 -1300
rect 12790 -1360 12830 -1300
rect 12690 -1380 12830 -1360
rect 12860 -1000 13000 -980
rect 12860 -1060 12900 -1000
rect 12960 -1060 13000 -1000
rect 12860 -1100 13000 -1060
rect 12860 -1160 12900 -1100
rect 12960 -1160 13000 -1100
rect 12860 -1200 13000 -1160
rect 12860 -1260 12900 -1200
rect 12960 -1260 13000 -1200
rect 12860 -1300 13000 -1260
rect 12860 -1360 12900 -1300
rect 12960 -1360 13000 -1300
rect 12860 -1380 13000 -1360
rect 13030 -1000 13170 -980
rect 13030 -1060 13070 -1000
rect 13130 -1060 13170 -1000
rect 13030 -1100 13170 -1060
rect 13030 -1160 13070 -1100
rect 13130 -1160 13170 -1100
rect 13030 -1200 13170 -1160
rect 13030 -1260 13070 -1200
rect 13130 -1260 13170 -1200
rect 13030 -1300 13170 -1260
rect 13030 -1360 13070 -1300
rect 13130 -1360 13170 -1300
rect 13030 -1380 13170 -1360
rect 13200 -1000 13340 -980
rect 13200 -1060 13240 -1000
rect 13300 -1060 13340 -1000
rect 13200 -1100 13340 -1060
rect 13200 -1160 13240 -1100
rect 13300 -1160 13340 -1100
rect 13200 -1200 13340 -1160
rect 13200 -1260 13240 -1200
rect 13300 -1260 13340 -1200
rect 13200 -1300 13340 -1260
rect 13200 -1360 13240 -1300
rect 13300 -1360 13340 -1300
rect 13200 -1380 13340 -1360
rect 13370 -1000 13510 -980
rect 13370 -1060 13410 -1000
rect 13470 -1060 13510 -1000
rect 13370 -1100 13510 -1060
rect 13370 -1160 13410 -1100
rect 13470 -1160 13510 -1100
rect 13370 -1200 13510 -1160
rect 13370 -1260 13410 -1200
rect 13470 -1260 13510 -1200
rect 13370 -1300 13510 -1260
rect 13370 -1360 13410 -1300
rect 13470 -1360 13510 -1300
rect 13370 -1380 13510 -1360
rect 13540 -1000 13680 -980
rect 13540 -1060 13580 -1000
rect 13640 -1060 13680 -1000
rect 13540 -1100 13680 -1060
rect 13540 -1160 13580 -1100
rect 13640 -1160 13680 -1100
rect 13540 -1200 13680 -1160
rect 13540 -1260 13580 -1200
rect 13640 -1260 13680 -1200
rect 13540 -1300 13680 -1260
rect 13540 -1360 13580 -1300
rect 13640 -1360 13680 -1300
rect 13540 -1380 13680 -1360
rect 13710 -1000 13850 -980
rect 13710 -1060 13750 -1000
rect 13810 -1060 13850 -1000
rect 13710 -1100 13850 -1060
rect 13710 -1160 13750 -1100
rect 13810 -1160 13850 -1100
rect 13710 -1200 13850 -1160
rect 13710 -1260 13750 -1200
rect 13810 -1260 13850 -1200
rect 13710 -1300 13850 -1260
rect 13710 -1360 13750 -1300
rect 13810 -1360 13850 -1300
rect 13710 -1380 13850 -1360
rect 13880 -1000 14020 -980
rect 13880 -1060 13920 -1000
rect 13980 -1060 14020 -1000
rect 13880 -1100 14020 -1060
rect 13880 -1160 13920 -1100
rect 13980 -1160 14020 -1100
rect 13880 -1200 14020 -1160
rect 13880 -1260 13920 -1200
rect 13980 -1260 14020 -1200
rect 13880 -1300 14020 -1260
rect 13880 -1360 13920 -1300
rect 13980 -1360 14020 -1300
rect 13880 -1380 14020 -1360
rect 14050 -1000 14190 -980
rect 14050 -1060 14090 -1000
rect 14150 -1060 14190 -1000
rect 14050 -1100 14190 -1060
rect 14050 -1160 14090 -1100
rect 14150 -1160 14190 -1100
rect 14050 -1200 14190 -1160
rect 14050 -1260 14090 -1200
rect 14150 -1260 14190 -1200
rect 14050 -1300 14190 -1260
rect 14050 -1360 14090 -1300
rect 14150 -1360 14190 -1300
rect 14050 -1380 14190 -1360
rect 14220 -1000 14360 -980
rect 14220 -1060 14260 -1000
rect 14320 -1060 14360 -1000
rect 14220 -1100 14360 -1060
rect 14220 -1160 14260 -1100
rect 14320 -1160 14360 -1100
rect 14220 -1200 14360 -1160
rect 14220 -1260 14260 -1200
rect 14320 -1260 14360 -1200
rect 14220 -1300 14360 -1260
rect 14220 -1360 14260 -1300
rect 14320 -1360 14360 -1300
rect 14220 -1380 14360 -1360
rect 14390 -1000 14530 -980
rect 14390 -1060 14430 -1000
rect 14490 -1060 14530 -1000
rect 14390 -1100 14530 -1060
rect 14390 -1160 14430 -1100
rect 14490 -1160 14530 -1100
rect 14390 -1200 14530 -1160
rect 14390 -1260 14430 -1200
rect 14490 -1260 14530 -1200
rect 14390 -1300 14530 -1260
rect 14390 -1360 14430 -1300
rect 14490 -1360 14530 -1300
rect 14390 -1380 14530 -1360
rect 14560 -1000 14700 -980
rect 14560 -1060 14600 -1000
rect 14660 -1060 14700 -1000
rect 14560 -1100 14700 -1060
rect 14560 -1160 14600 -1100
rect 14660 -1160 14700 -1100
rect 14560 -1200 14700 -1160
rect 14560 -1260 14600 -1200
rect 14660 -1260 14700 -1200
rect 14560 -1300 14700 -1260
rect 14560 -1360 14600 -1300
rect 14660 -1360 14700 -1300
rect 14560 -1380 14700 -1360
rect 14730 -1000 14870 -980
rect 14730 -1060 14770 -1000
rect 14830 -1060 14870 -1000
rect 14730 -1100 14870 -1060
rect 14730 -1160 14770 -1100
rect 14830 -1160 14870 -1100
rect 14730 -1200 14870 -1160
rect 14730 -1260 14770 -1200
rect 14830 -1260 14870 -1200
rect 14730 -1300 14870 -1260
rect 14730 -1360 14770 -1300
rect 14830 -1360 14870 -1300
rect 14730 -1380 14870 -1360
rect 14900 -1000 15040 -980
rect 14900 -1060 14940 -1000
rect 15000 -1060 15040 -1000
rect 14900 -1100 15040 -1060
rect 14900 -1160 14940 -1100
rect 15000 -1160 15040 -1100
rect 14900 -1200 15040 -1160
rect 14900 -1260 14940 -1200
rect 15000 -1260 15040 -1200
rect 14900 -1300 15040 -1260
rect 14900 -1360 14940 -1300
rect 15000 -1360 15040 -1300
rect 14900 -1380 15040 -1360
rect 15070 -1000 15210 -980
rect 15070 -1060 15110 -1000
rect 15170 -1060 15210 -1000
rect 15070 -1100 15210 -1060
rect 15070 -1160 15110 -1100
rect 15170 -1160 15210 -1100
rect 15070 -1200 15210 -1160
rect 15070 -1260 15110 -1200
rect 15170 -1260 15210 -1200
rect 15070 -1300 15210 -1260
rect 15070 -1360 15110 -1300
rect 15170 -1360 15210 -1300
rect 15070 -1380 15210 -1360
rect 15240 -1000 15380 -980
rect 15240 -1060 15280 -1000
rect 15340 -1060 15380 -1000
rect 15240 -1100 15380 -1060
rect 15240 -1160 15280 -1100
rect 15340 -1160 15380 -1100
rect 15240 -1200 15380 -1160
rect 15240 -1260 15280 -1200
rect 15340 -1260 15380 -1200
rect 15240 -1300 15380 -1260
rect 15240 -1360 15280 -1300
rect 15340 -1360 15380 -1300
rect 15240 -1380 15380 -1360
rect 15410 -1000 15550 -980
rect 15410 -1060 15450 -1000
rect 15510 -1060 15550 -1000
rect 15410 -1100 15550 -1060
rect 15410 -1160 15450 -1100
rect 15510 -1160 15550 -1100
rect 15410 -1200 15550 -1160
rect 15410 -1260 15450 -1200
rect 15510 -1260 15550 -1200
rect 15410 -1300 15550 -1260
rect 15410 -1360 15450 -1300
rect 15510 -1360 15550 -1300
rect 15410 -1380 15550 -1360
rect 15580 -1000 15720 -980
rect 15580 -1060 15620 -1000
rect 15680 -1060 15720 -1000
rect 15580 -1100 15720 -1060
rect 15580 -1160 15620 -1100
rect 15680 -1160 15720 -1100
rect 15580 -1200 15720 -1160
rect 15580 -1260 15620 -1200
rect 15680 -1260 15720 -1200
rect 15580 -1300 15720 -1260
rect 15580 -1360 15620 -1300
rect 15680 -1360 15720 -1300
rect 15580 -1380 15720 -1360
rect 15750 -1000 15890 -980
rect 15750 -1060 15790 -1000
rect 15850 -1060 15890 -1000
rect 15750 -1100 15890 -1060
rect 15750 -1160 15790 -1100
rect 15850 -1160 15890 -1100
rect 15750 -1200 15890 -1160
rect 15750 -1260 15790 -1200
rect 15850 -1260 15890 -1200
rect 15750 -1300 15890 -1260
rect 15750 -1360 15790 -1300
rect 15850 -1360 15890 -1300
rect 15750 -1380 15890 -1360
rect 15920 -1000 16060 -980
rect 15920 -1060 15960 -1000
rect 16020 -1060 16060 -1000
rect 15920 -1100 16060 -1060
rect 15920 -1160 15960 -1100
rect 16020 -1160 16060 -1100
rect 15920 -1200 16060 -1160
rect 15920 -1260 15960 -1200
rect 16020 -1260 16060 -1200
rect 15920 -1300 16060 -1260
rect 15920 -1360 15960 -1300
rect 16020 -1360 16060 -1300
rect 15920 -1380 16060 -1360
rect 16090 -1000 16230 -980
rect 16090 -1060 16130 -1000
rect 16190 -1060 16230 -1000
rect 16090 -1100 16230 -1060
rect 16090 -1160 16130 -1100
rect 16190 -1160 16230 -1100
rect 16090 -1200 16230 -1160
rect 16090 -1260 16130 -1200
rect 16190 -1260 16230 -1200
rect 16090 -1300 16230 -1260
rect 16090 -1360 16130 -1300
rect 16190 -1360 16230 -1300
rect 16090 -1380 16230 -1360
rect 16260 -1000 16400 -980
rect 16260 -1060 16300 -1000
rect 16360 -1060 16400 -1000
rect 16260 -1100 16400 -1060
rect 16260 -1160 16300 -1100
rect 16360 -1160 16400 -1100
rect 16260 -1200 16400 -1160
rect 16260 -1260 16300 -1200
rect 16360 -1260 16400 -1200
rect 16260 -1300 16400 -1260
rect 16260 -1360 16300 -1300
rect 16360 -1360 16400 -1300
rect 16260 -1380 16400 -1360
rect 16430 -1000 16570 -980
rect 16430 -1060 16470 -1000
rect 16530 -1060 16570 -1000
rect 16430 -1100 16570 -1060
rect 16430 -1160 16470 -1100
rect 16530 -1160 16570 -1100
rect 16430 -1200 16570 -1160
rect 16430 -1260 16470 -1200
rect 16530 -1260 16570 -1200
rect 16430 -1300 16570 -1260
rect 16430 -1360 16470 -1300
rect 16530 -1360 16570 -1300
rect 16430 -1380 16570 -1360
rect 16600 -1000 16740 -980
rect 16600 -1060 16640 -1000
rect 16700 -1060 16740 -1000
rect 16600 -1100 16740 -1060
rect 16600 -1160 16640 -1100
rect 16700 -1160 16740 -1100
rect 16600 -1200 16740 -1160
rect 16600 -1260 16640 -1200
rect 16700 -1260 16740 -1200
rect 16600 -1300 16740 -1260
rect 16600 -1360 16640 -1300
rect 16700 -1360 16740 -1300
rect 16600 -1380 16740 -1360
rect 16770 -1000 16910 -980
rect 16770 -1060 16810 -1000
rect 16870 -1060 16910 -1000
rect 16770 -1100 16910 -1060
rect 16770 -1160 16810 -1100
rect 16870 -1160 16910 -1100
rect 16770 -1200 16910 -1160
rect 16770 -1260 16810 -1200
rect 16870 -1260 16910 -1200
rect 16770 -1300 16910 -1260
rect 16770 -1360 16810 -1300
rect 16870 -1360 16910 -1300
rect 16770 -1380 16910 -1360
rect 16940 -1000 17080 -980
rect 16940 -1060 16980 -1000
rect 17040 -1060 17080 -1000
rect 16940 -1100 17080 -1060
rect 16940 -1160 16980 -1100
rect 17040 -1160 17080 -1100
rect 16940 -1200 17080 -1160
rect 16940 -1260 16980 -1200
rect 17040 -1260 17080 -1200
rect 16940 -1300 17080 -1260
rect 16940 -1360 16980 -1300
rect 17040 -1360 17080 -1300
rect 16940 -1380 17080 -1360
rect 17110 -1000 17250 -980
rect 17110 -1060 17150 -1000
rect 17210 -1060 17250 -1000
rect 17110 -1100 17250 -1060
rect 17110 -1160 17150 -1100
rect 17210 -1160 17250 -1100
rect 17110 -1200 17250 -1160
rect 17110 -1260 17150 -1200
rect 17210 -1260 17250 -1200
rect 17110 -1300 17250 -1260
rect 17110 -1360 17150 -1300
rect 17210 -1360 17250 -1300
rect 17110 -1380 17250 -1360
rect 17280 -1000 17420 -980
rect 17280 -1060 17320 -1000
rect 17380 -1060 17420 -1000
rect 17280 -1100 17420 -1060
rect 17280 -1160 17320 -1100
rect 17380 -1160 17420 -1100
rect 17280 -1200 17420 -1160
rect 17280 -1260 17320 -1200
rect 17380 -1260 17420 -1200
rect 17280 -1300 17420 -1260
rect 17280 -1360 17320 -1300
rect 17380 -1360 17420 -1300
rect 17280 -1380 17420 -1360
rect 17450 -1000 17590 -980
rect 17450 -1060 17490 -1000
rect 17550 -1060 17590 -1000
rect 17450 -1100 17590 -1060
rect 17450 -1160 17490 -1100
rect 17550 -1160 17590 -1100
rect 17450 -1200 17590 -1160
rect 17450 -1260 17490 -1200
rect 17550 -1260 17590 -1200
rect 17450 -1300 17590 -1260
rect 17450 -1360 17490 -1300
rect 17550 -1360 17590 -1300
rect 17450 -1380 17590 -1360
rect 17620 -1000 17760 -980
rect 17620 -1060 17660 -1000
rect 17720 -1060 17760 -1000
rect 17620 -1100 17760 -1060
rect 17620 -1160 17660 -1100
rect 17720 -1160 17760 -1100
rect 17620 -1200 17760 -1160
rect 17620 -1260 17660 -1200
rect 17720 -1260 17760 -1200
rect 17620 -1300 17760 -1260
rect 17620 -1360 17660 -1300
rect 17720 -1360 17760 -1300
rect 17620 -1380 17760 -1360
rect 17790 -1000 17930 -980
rect 17790 -1060 17830 -1000
rect 17890 -1060 17930 -1000
rect 17790 -1100 17930 -1060
rect 17790 -1160 17830 -1100
rect 17890 -1160 17930 -1100
rect 17790 -1200 17930 -1160
rect 17790 -1260 17830 -1200
rect 17890 -1260 17930 -1200
rect 17790 -1300 17930 -1260
rect 17790 -1360 17830 -1300
rect 17890 -1360 17930 -1300
rect 17790 -1380 17930 -1360
rect 17960 -1000 18100 -980
rect 17960 -1060 18000 -1000
rect 18060 -1060 18100 -1000
rect 17960 -1100 18100 -1060
rect 17960 -1160 18000 -1100
rect 18060 -1160 18100 -1100
rect 17960 -1200 18100 -1160
rect 17960 -1260 18000 -1200
rect 18060 -1260 18100 -1200
rect 17960 -1300 18100 -1260
rect 17960 -1360 18000 -1300
rect 18060 -1360 18100 -1300
rect 17960 -1380 18100 -1360
rect 18130 -1000 18270 -980
rect 18130 -1060 18170 -1000
rect 18230 -1060 18270 -1000
rect 18130 -1100 18270 -1060
rect 18130 -1160 18170 -1100
rect 18230 -1160 18270 -1100
rect 18130 -1200 18270 -1160
rect 18130 -1260 18170 -1200
rect 18230 -1260 18270 -1200
rect 18130 -1300 18270 -1260
rect 18130 -1360 18170 -1300
rect 18230 -1360 18270 -1300
rect 18130 -1380 18270 -1360
rect 18300 -1000 18440 -980
rect 18300 -1060 18340 -1000
rect 18400 -1060 18440 -1000
rect 18300 -1100 18440 -1060
rect 18300 -1160 18340 -1100
rect 18400 -1160 18440 -1100
rect 18300 -1200 18440 -1160
rect 18300 -1260 18340 -1200
rect 18400 -1260 18440 -1200
rect 18300 -1300 18440 -1260
rect 18300 -1360 18340 -1300
rect 18400 -1360 18440 -1300
rect 18300 -1380 18440 -1360
rect 18470 -1000 18610 -980
rect 18470 -1060 18510 -1000
rect 18570 -1060 18610 -1000
rect 18470 -1100 18610 -1060
rect 18470 -1160 18510 -1100
rect 18570 -1160 18610 -1100
rect 18470 -1200 18610 -1160
rect 18470 -1260 18510 -1200
rect 18570 -1260 18610 -1200
rect 18470 -1300 18610 -1260
rect 18470 -1360 18510 -1300
rect 18570 -1360 18610 -1300
rect 18470 -1380 18610 -1360
rect 18640 -1000 18780 -980
rect 18640 -1060 18680 -1000
rect 18740 -1060 18780 -1000
rect 18640 -1100 18780 -1060
rect 18640 -1160 18680 -1100
rect 18740 -1160 18780 -1100
rect 18640 -1200 18780 -1160
rect 18640 -1260 18680 -1200
rect 18740 -1260 18780 -1200
rect 18640 -1300 18780 -1260
rect 18640 -1360 18680 -1300
rect 18740 -1360 18780 -1300
rect 18640 -1380 18780 -1360
rect 18810 -1000 18950 -980
rect 18810 -1060 18850 -1000
rect 18910 -1060 18950 -1000
rect 18810 -1100 18950 -1060
rect 18810 -1160 18850 -1100
rect 18910 -1160 18950 -1100
rect 18810 -1200 18950 -1160
rect 18810 -1260 18850 -1200
rect 18910 -1260 18950 -1200
rect 18810 -1300 18950 -1260
rect 18810 -1360 18850 -1300
rect 18910 -1360 18950 -1300
rect 18810 -1380 18950 -1360
rect 18980 -1000 19120 -980
rect 18980 -1060 19020 -1000
rect 19080 -1060 19120 -1000
rect 18980 -1100 19120 -1060
rect 18980 -1160 19020 -1100
rect 19080 -1160 19120 -1100
rect 18980 -1200 19120 -1160
rect 18980 -1260 19020 -1200
rect 19080 -1260 19120 -1200
rect 18980 -1300 19120 -1260
rect 18980 -1360 19020 -1300
rect 19080 -1360 19120 -1300
rect 18980 -1380 19120 -1360
rect 19150 -1000 19290 -980
rect 19150 -1060 19190 -1000
rect 19250 -1060 19290 -1000
rect 19150 -1100 19290 -1060
rect 19150 -1160 19190 -1100
rect 19250 -1160 19290 -1100
rect 19150 -1200 19290 -1160
rect 19150 -1260 19190 -1200
rect 19250 -1260 19290 -1200
rect 19150 -1300 19290 -1260
rect 19150 -1360 19190 -1300
rect 19250 -1360 19290 -1300
rect 19150 -1380 19290 -1360
rect 19320 -1000 19460 -980
rect 19320 -1060 19360 -1000
rect 19420 -1060 19460 -1000
rect 19320 -1100 19460 -1060
rect 19320 -1160 19360 -1100
rect 19420 -1160 19460 -1100
rect 19320 -1200 19460 -1160
rect 19320 -1260 19360 -1200
rect 19420 -1260 19460 -1200
rect 19320 -1300 19460 -1260
rect 19320 -1360 19360 -1300
rect 19420 -1360 19460 -1300
rect 19320 -1380 19460 -1360
rect 19490 -1000 19630 -980
rect 19490 -1060 19530 -1000
rect 19590 -1060 19630 -1000
rect 19490 -1100 19630 -1060
rect 19490 -1160 19530 -1100
rect 19590 -1160 19630 -1100
rect 19490 -1200 19630 -1160
rect 19490 -1260 19530 -1200
rect 19590 -1260 19630 -1200
rect 19490 -1300 19630 -1260
rect 19490 -1360 19530 -1300
rect 19590 -1360 19630 -1300
rect 19490 -1380 19630 -1360
rect 19660 -1000 19800 -980
rect 19660 -1060 19700 -1000
rect 19760 -1060 19800 -1000
rect 19660 -1100 19800 -1060
rect 19660 -1160 19700 -1100
rect 19760 -1160 19800 -1100
rect 19660 -1200 19800 -1160
rect 19660 -1260 19700 -1200
rect 19760 -1260 19800 -1200
rect 19660 -1300 19800 -1260
rect 19660 -1360 19700 -1300
rect 19760 -1360 19800 -1300
rect 19660 -1380 19800 -1360
rect 19830 -1000 19970 -980
rect 19830 -1060 19870 -1000
rect 19930 -1060 19970 -1000
rect 19830 -1100 19970 -1060
rect 19830 -1160 19870 -1100
rect 19930 -1160 19970 -1100
rect 19830 -1200 19970 -1160
rect 19830 -1260 19870 -1200
rect 19930 -1260 19970 -1200
rect 19830 -1300 19970 -1260
rect 19830 -1360 19870 -1300
rect 19930 -1360 19970 -1300
rect 19830 -1380 19970 -1360
rect 20000 -1000 20140 -980
rect 20000 -1060 20040 -1000
rect 20100 -1060 20140 -1000
rect 20000 -1100 20140 -1060
rect 20000 -1160 20040 -1100
rect 20100 -1160 20140 -1100
rect 20000 -1200 20140 -1160
rect 20000 -1260 20040 -1200
rect 20100 -1260 20140 -1200
rect 20000 -1300 20140 -1260
rect 20000 -1360 20040 -1300
rect 20100 -1360 20140 -1300
rect 20000 -1380 20140 -1360
rect 20170 -1000 20310 -980
rect 20170 -1060 20210 -1000
rect 20270 -1060 20310 -1000
rect 20170 -1100 20310 -1060
rect 20170 -1160 20210 -1100
rect 20270 -1160 20310 -1100
rect 20170 -1200 20310 -1160
rect 20170 -1260 20210 -1200
rect 20270 -1260 20310 -1200
rect 20170 -1300 20310 -1260
rect 20170 -1360 20210 -1300
rect 20270 -1360 20310 -1300
rect 20170 -1380 20310 -1360
rect 20340 -1000 20480 -980
rect 20340 -1060 20380 -1000
rect 20440 -1060 20480 -1000
rect 20340 -1100 20480 -1060
rect 20340 -1160 20380 -1100
rect 20440 -1160 20480 -1100
rect 20340 -1200 20480 -1160
rect 20340 -1260 20380 -1200
rect 20440 -1260 20480 -1200
rect 20340 -1300 20480 -1260
rect 20340 -1360 20380 -1300
rect 20440 -1360 20480 -1300
rect 20340 -1380 20480 -1360
rect 20510 -1000 20650 -980
rect 20510 -1060 20550 -1000
rect 20610 -1060 20650 -1000
rect 20510 -1100 20650 -1060
rect 20510 -1160 20550 -1100
rect 20610 -1160 20650 -1100
rect 20510 -1200 20650 -1160
rect 20510 -1260 20550 -1200
rect 20610 -1260 20650 -1200
rect 20510 -1300 20650 -1260
rect 20510 -1360 20550 -1300
rect 20610 -1360 20650 -1300
rect 20510 -1380 20650 -1360
rect 20680 -1000 20820 -980
rect 20680 -1060 20720 -1000
rect 20780 -1060 20820 -1000
rect 20680 -1100 20820 -1060
rect 20680 -1160 20720 -1100
rect 20780 -1160 20820 -1100
rect 20680 -1200 20820 -1160
rect 20680 -1260 20720 -1200
rect 20780 -1260 20820 -1200
rect 20680 -1300 20820 -1260
rect 20680 -1360 20720 -1300
rect 20780 -1360 20820 -1300
rect 20680 -1380 20820 -1360
rect 20850 -1000 20990 -980
rect 20850 -1060 20890 -1000
rect 20950 -1060 20990 -1000
rect 20850 -1100 20990 -1060
rect 20850 -1160 20890 -1100
rect 20950 -1160 20990 -1100
rect 20850 -1200 20990 -1160
rect 20850 -1260 20890 -1200
rect 20950 -1260 20990 -1200
rect 20850 -1300 20990 -1260
rect 20850 -1360 20890 -1300
rect 20950 -1360 20990 -1300
rect 20850 -1380 20990 -1360
rect 21020 -1000 21160 -980
rect 21020 -1060 21060 -1000
rect 21120 -1060 21160 -1000
rect 21020 -1100 21160 -1060
rect 21020 -1160 21060 -1100
rect 21120 -1160 21160 -1100
rect 21020 -1200 21160 -1160
rect 21020 -1260 21060 -1200
rect 21120 -1260 21160 -1200
rect 21020 -1300 21160 -1260
rect 21020 -1360 21060 -1300
rect 21120 -1360 21160 -1300
rect 21020 -1380 21160 -1360
rect 21190 -1000 21330 -980
rect 21190 -1060 21230 -1000
rect 21290 -1060 21330 -1000
rect 21190 -1100 21330 -1060
rect 21190 -1160 21230 -1100
rect 21290 -1160 21330 -1100
rect 21190 -1200 21330 -1160
rect 21190 -1260 21230 -1200
rect 21290 -1260 21330 -1200
rect 21190 -1300 21330 -1260
rect 21190 -1360 21230 -1300
rect 21290 -1360 21330 -1300
rect 21190 -1380 21330 -1360
rect 21360 -1000 21500 -980
rect 21360 -1060 21400 -1000
rect 21460 -1060 21500 -1000
rect 21360 -1100 21500 -1060
rect 21360 -1160 21400 -1100
rect 21460 -1160 21500 -1100
rect 21360 -1200 21500 -1160
rect 21360 -1260 21400 -1200
rect 21460 -1260 21500 -1200
rect 21360 -1300 21500 -1260
rect 21360 -1360 21400 -1300
rect 21460 -1360 21500 -1300
rect 21360 -1380 21500 -1360
rect 21530 -1000 21670 -980
rect 21530 -1060 21570 -1000
rect 21630 -1060 21670 -1000
rect 21530 -1100 21670 -1060
rect 21530 -1160 21570 -1100
rect 21630 -1160 21670 -1100
rect 21530 -1200 21670 -1160
rect 21530 -1260 21570 -1200
rect 21630 -1260 21670 -1200
rect 21530 -1300 21670 -1260
rect 21530 -1360 21570 -1300
rect 21630 -1360 21670 -1300
rect 21530 -1380 21670 -1360
rect 21700 -1000 21840 -980
rect 21700 -1060 21740 -1000
rect 21800 -1060 21840 -1000
rect 21700 -1100 21840 -1060
rect 21700 -1160 21740 -1100
rect 21800 -1160 21840 -1100
rect 21700 -1200 21840 -1160
rect 21700 -1260 21740 -1200
rect 21800 -1260 21840 -1200
rect 21700 -1300 21840 -1260
rect 21700 -1360 21740 -1300
rect 21800 -1360 21840 -1300
rect 21700 -1380 21840 -1360
rect 21870 -1000 22010 -980
rect 21870 -1060 21910 -1000
rect 21970 -1060 22010 -1000
rect 21870 -1100 22010 -1060
rect 21870 -1160 21910 -1100
rect 21970 -1160 22010 -1100
rect 21870 -1200 22010 -1160
rect 21870 -1260 21910 -1200
rect 21970 -1260 22010 -1200
rect 21870 -1300 22010 -1260
rect 21870 -1360 21910 -1300
rect 21970 -1360 22010 -1300
rect 21870 -1380 22010 -1360
rect 22040 -1000 22180 -980
rect 22040 -1060 22080 -1000
rect 22140 -1060 22180 -1000
rect 22040 -1100 22180 -1060
rect 22040 -1160 22080 -1100
rect 22140 -1160 22180 -1100
rect 22040 -1200 22180 -1160
rect 22040 -1260 22080 -1200
rect 22140 -1260 22180 -1200
rect 22040 -1300 22180 -1260
rect 22040 -1360 22080 -1300
rect 22140 -1360 22180 -1300
rect 22040 -1380 22180 -1360
rect 22210 -1000 22350 -980
rect 22210 -1060 22250 -1000
rect 22310 -1060 22350 -1000
rect 22210 -1100 22350 -1060
rect 22210 -1160 22250 -1100
rect 22310 -1160 22350 -1100
rect 22210 -1200 22350 -1160
rect 22210 -1260 22250 -1200
rect 22310 -1260 22350 -1200
rect 22210 -1300 22350 -1260
rect 22210 -1360 22250 -1300
rect 22310 -1360 22350 -1300
rect 22210 -1380 22350 -1360
rect 22380 -1000 22520 -980
rect 22380 -1060 22420 -1000
rect 22480 -1060 22520 -1000
rect 22380 -1100 22520 -1060
rect 22380 -1160 22420 -1100
rect 22480 -1160 22520 -1100
rect 22380 -1200 22520 -1160
rect 22380 -1260 22420 -1200
rect 22480 -1260 22520 -1200
rect 22380 -1300 22520 -1260
rect 22380 -1360 22420 -1300
rect 22480 -1360 22520 -1300
rect 22380 -1380 22520 -1360
rect 22550 -1000 22690 -980
rect 22550 -1060 22590 -1000
rect 22650 -1060 22690 -1000
rect 22550 -1100 22690 -1060
rect 22550 -1160 22590 -1100
rect 22650 -1160 22690 -1100
rect 22550 -1200 22690 -1160
rect 22550 -1260 22590 -1200
rect 22650 -1260 22690 -1200
rect 22550 -1300 22690 -1260
rect 22550 -1360 22590 -1300
rect 22650 -1360 22690 -1300
rect 22550 -1380 22690 -1360
rect 22720 -1000 22860 -980
rect 22720 -1060 22760 -1000
rect 22820 -1060 22860 -1000
rect 22720 -1100 22860 -1060
rect 22720 -1160 22760 -1100
rect 22820 -1160 22860 -1100
rect 22720 -1200 22860 -1160
rect 22720 -1260 22760 -1200
rect 22820 -1260 22860 -1200
rect 22720 -1300 22860 -1260
rect 22720 -1360 22760 -1300
rect 22820 -1360 22860 -1300
rect 22720 -1380 22860 -1360
rect 22890 -1000 23030 -980
rect 22890 -1060 22930 -1000
rect 22990 -1060 23030 -1000
rect 22890 -1100 23030 -1060
rect 22890 -1160 22930 -1100
rect 22990 -1160 23030 -1100
rect 22890 -1200 23030 -1160
rect 22890 -1260 22930 -1200
rect 22990 -1260 23030 -1200
rect 22890 -1300 23030 -1260
rect 22890 -1360 22930 -1300
rect 22990 -1360 23030 -1300
rect 22890 -1380 23030 -1360
rect 23060 -1000 23200 -980
rect 23060 -1060 23100 -1000
rect 23160 -1060 23200 -1000
rect 23060 -1100 23200 -1060
rect 23060 -1160 23100 -1100
rect 23160 -1160 23200 -1100
rect 23060 -1200 23200 -1160
rect 23060 -1260 23100 -1200
rect 23160 -1260 23200 -1200
rect 23060 -1300 23200 -1260
rect 23060 -1360 23100 -1300
rect 23160 -1360 23200 -1300
rect 23060 -1380 23200 -1360
rect 23230 -1000 23370 -980
rect 23230 -1060 23270 -1000
rect 23330 -1060 23370 -1000
rect 23230 -1100 23370 -1060
rect 23230 -1160 23270 -1100
rect 23330 -1160 23370 -1100
rect 23230 -1200 23370 -1160
rect 23230 -1260 23270 -1200
rect 23330 -1260 23370 -1200
rect 23230 -1300 23370 -1260
rect 23230 -1360 23270 -1300
rect 23330 -1360 23370 -1300
rect 23230 -1380 23370 -1360
rect 23400 -1000 23540 -980
rect 23400 -1060 23440 -1000
rect 23500 -1060 23540 -1000
rect 23400 -1100 23540 -1060
rect 23400 -1160 23440 -1100
rect 23500 -1160 23540 -1100
rect 23400 -1200 23540 -1160
rect 23400 -1260 23440 -1200
rect 23500 -1260 23540 -1200
rect 23400 -1300 23540 -1260
rect 23400 -1360 23440 -1300
rect 23500 -1360 23540 -1300
rect 23400 -1380 23540 -1360
rect 23570 -1000 23710 -980
rect 23570 -1060 23610 -1000
rect 23670 -1060 23710 -1000
rect 23570 -1100 23710 -1060
rect 23570 -1160 23610 -1100
rect 23670 -1160 23710 -1100
rect 23570 -1200 23710 -1160
rect 23570 -1260 23610 -1200
rect 23670 -1260 23710 -1200
rect 23570 -1300 23710 -1260
rect 23570 -1360 23610 -1300
rect 23670 -1360 23710 -1300
rect 23570 -1380 23710 -1360
rect 23740 -1000 23880 -980
rect 23740 -1060 23780 -1000
rect 23840 -1060 23880 -1000
rect 23740 -1100 23880 -1060
rect 23740 -1160 23780 -1100
rect 23840 -1160 23880 -1100
rect 23740 -1200 23880 -1160
rect 23740 -1260 23780 -1200
rect 23840 -1260 23880 -1200
rect 23740 -1300 23880 -1260
rect 23740 -1360 23780 -1300
rect 23840 -1360 23880 -1300
rect 23740 -1380 23880 -1360
rect 23910 -1000 24050 -980
rect 23910 -1060 23950 -1000
rect 24010 -1060 24050 -1000
rect 23910 -1100 24050 -1060
rect 23910 -1160 23950 -1100
rect 24010 -1160 24050 -1100
rect 23910 -1200 24050 -1160
rect 23910 -1260 23950 -1200
rect 24010 -1260 24050 -1200
rect 23910 -1300 24050 -1260
rect 23910 -1360 23950 -1300
rect 24010 -1360 24050 -1300
rect 23910 -1380 24050 -1360
rect 24080 -1000 24220 -980
rect 24080 -1060 24120 -1000
rect 24180 -1060 24220 -1000
rect 24080 -1100 24220 -1060
rect 24080 -1160 24120 -1100
rect 24180 -1160 24220 -1100
rect 24080 -1200 24220 -1160
rect 24080 -1260 24120 -1200
rect 24180 -1260 24220 -1200
rect 24080 -1300 24220 -1260
rect 24080 -1360 24120 -1300
rect 24180 -1360 24220 -1300
rect 24080 -1380 24220 -1360
rect 24250 -1000 24390 -980
rect 24250 -1060 24290 -1000
rect 24350 -1060 24390 -1000
rect 24250 -1100 24390 -1060
rect 24250 -1160 24290 -1100
rect 24350 -1160 24390 -1100
rect 24250 -1200 24390 -1160
rect 24250 -1260 24290 -1200
rect 24350 -1260 24390 -1200
rect 24250 -1300 24390 -1260
rect 24250 -1360 24290 -1300
rect 24350 -1360 24390 -1300
rect 24250 -1380 24390 -1360
rect 24420 -1000 24560 -980
rect 24420 -1060 24460 -1000
rect 24520 -1060 24560 -1000
rect 24420 -1100 24560 -1060
rect 24420 -1160 24460 -1100
rect 24520 -1160 24560 -1100
rect 24420 -1200 24560 -1160
rect 24420 -1260 24460 -1200
rect 24520 -1260 24560 -1200
rect 24420 -1300 24560 -1260
rect 24420 -1360 24460 -1300
rect 24520 -1360 24560 -1300
rect 24420 -1380 24560 -1360
rect 24590 -1000 24730 -980
rect 24590 -1060 24630 -1000
rect 24690 -1060 24730 -1000
rect 24590 -1100 24730 -1060
rect 24590 -1160 24630 -1100
rect 24690 -1160 24730 -1100
rect 24590 -1200 24730 -1160
rect 24590 -1260 24630 -1200
rect 24690 -1260 24730 -1200
rect 24590 -1300 24730 -1260
rect 24590 -1360 24630 -1300
rect 24690 -1360 24730 -1300
rect 24590 -1380 24730 -1360
rect 24760 -1000 24900 -980
rect 24760 -1060 24800 -1000
rect 24860 -1060 24900 -1000
rect 24760 -1100 24900 -1060
rect 24760 -1160 24800 -1100
rect 24860 -1160 24900 -1100
rect 24760 -1200 24900 -1160
rect 24760 -1260 24800 -1200
rect 24860 -1260 24900 -1200
rect 24760 -1300 24900 -1260
rect 24760 -1360 24800 -1300
rect 24860 -1360 24900 -1300
rect 24760 -1380 24900 -1360
rect 24930 -1000 25070 -980
rect 24930 -1060 24970 -1000
rect 25030 -1060 25070 -1000
rect 24930 -1100 25070 -1060
rect 24930 -1160 24970 -1100
rect 25030 -1160 25070 -1100
rect 24930 -1200 25070 -1160
rect 24930 -1260 24970 -1200
rect 25030 -1260 25070 -1200
rect 24930 -1300 25070 -1260
rect 24930 -1360 24970 -1300
rect 25030 -1360 25070 -1300
rect 24930 -1380 25070 -1360
rect 25100 -1000 25240 -980
rect 25100 -1060 25140 -1000
rect 25200 -1060 25240 -1000
rect 25100 -1100 25240 -1060
rect 25100 -1160 25140 -1100
rect 25200 -1160 25240 -1100
rect 25100 -1200 25240 -1160
rect 25100 -1260 25140 -1200
rect 25200 -1260 25240 -1200
rect 25100 -1300 25240 -1260
rect 25100 -1360 25140 -1300
rect 25200 -1360 25240 -1300
rect 25100 -1380 25240 -1360
rect 25270 -1000 25410 -980
rect 25270 -1060 25310 -1000
rect 25370 -1060 25410 -1000
rect 25270 -1100 25410 -1060
rect 25270 -1160 25310 -1100
rect 25370 -1160 25410 -1100
rect 25270 -1200 25410 -1160
rect 25270 -1260 25310 -1200
rect 25370 -1260 25410 -1200
rect 25270 -1300 25410 -1260
rect 25270 -1360 25310 -1300
rect 25370 -1360 25410 -1300
rect 25270 -1380 25410 -1360
rect 25440 -1000 25580 -980
rect 25440 -1060 25480 -1000
rect 25540 -1060 25580 -1000
rect 25440 -1100 25580 -1060
rect 25440 -1160 25480 -1100
rect 25540 -1160 25580 -1100
rect 25440 -1200 25580 -1160
rect 25440 -1260 25480 -1200
rect 25540 -1260 25580 -1200
rect 25440 -1300 25580 -1260
rect 25440 -1360 25480 -1300
rect 25540 -1360 25580 -1300
rect 25440 -1380 25580 -1360
rect 25610 -1000 25750 -980
rect 25610 -1060 25650 -1000
rect 25710 -1060 25750 -1000
rect 25610 -1100 25750 -1060
rect 25610 -1160 25650 -1100
rect 25710 -1160 25750 -1100
rect 25610 -1200 25750 -1160
rect 25610 -1260 25650 -1200
rect 25710 -1260 25750 -1200
rect 25610 -1300 25750 -1260
rect 25610 -1360 25650 -1300
rect 25710 -1360 25750 -1300
rect 25610 -1380 25750 -1360
rect 25780 -1000 25920 -980
rect 25780 -1060 25820 -1000
rect 25880 -1060 25920 -1000
rect 25780 -1100 25920 -1060
rect 25780 -1160 25820 -1100
rect 25880 -1160 25920 -1100
rect 25780 -1200 25920 -1160
rect 25780 -1260 25820 -1200
rect 25880 -1260 25920 -1200
rect 25780 -1300 25920 -1260
rect 25780 -1360 25820 -1300
rect 25880 -1360 25920 -1300
rect 25780 -1380 25920 -1360
rect 25950 -1000 26090 -980
rect 25950 -1060 25990 -1000
rect 26050 -1060 26090 -1000
rect 25950 -1100 26090 -1060
rect 25950 -1160 25990 -1100
rect 26050 -1160 26090 -1100
rect 25950 -1200 26090 -1160
rect 25950 -1260 25990 -1200
rect 26050 -1260 26090 -1200
rect 25950 -1300 26090 -1260
rect 25950 -1360 25990 -1300
rect 26050 -1360 26090 -1300
rect 25950 -1380 26090 -1360
rect 26120 -1000 26260 -980
rect 26120 -1060 26160 -1000
rect 26220 -1060 26260 -1000
rect 26120 -1100 26260 -1060
rect 26120 -1160 26160 -1100
rect 26220 -1160 26260 -1100
rect 26120 -1200 26260 -1160
rect 26120 -1260 26160 -1200
rect 26220 -1260 26260 -1200
rect 26120 -1300 26260 -1260
rect 26120 -1360 26160 -1300
rect 26220 -1360 26260 -1300
rect 26120 -1380 26260 -1360
rect 26290 -1000 26430 -980
rect 26290 -1060 26330 -1000
rect 26390 -1060 26430 -1000
rect 26290 -1100 26430 -1060
rect 26290 -1160 26330 -1100
rect 26390 -1160 26430 -1100
rect 26290 -1200 26430 -1160
rect 26290 -1260 26330 -1200
rect 26390 -1260 26430 -1200
rect 26290 -1300 26430 -1260
rect 26290 -1360 26330 -1300
rect 26390 -1360 26430 -1300
rect 26290 -1380 26430 -1360
rect 26460 -1000 26600 -980
rect 26460 -1060 26500 -1000
rect 26560 -1060 26600 -1000
rect 26460 -1100 26600 -1060
rect 26460 -1160 26500 -1100
rect 26560 -1160 26600 -1100
rect 26460 -1200 26600 -1160
rect 26460 -1260 26500 -1200
rect 26560 -1260 26600 -1200
rect 26460 -1300 26600 -1260
rect 26460 -1360 26500 -1300
rect 26560 -1360 26600 -1300
rect 26460 -1380 26600 -1360
rect 26630 -1000 26770 -980
rect 26630 -1060 26670 -1000
rect 26730 -1060 26770 -1000
rect 26630 -1100 26770 -1060
rect 26630 -1160 26670 -1100
rect 26730 -1160 26770 -1100
rect 26630 -1200 26770 -1160
rect 26630 -1260 26670 -1200
rect 26730 -1260 26770 -1200
rect 26630 -1300 26770 -1260
rect 26630 -1360 26670 -1300
rect 26730 -1360 26770 -1300
rect 26630 -1380 26770 -1360
rect 26800 -1000 26940 -980
rect 26800 -1060 26840 -1000
rect 26900 -1060 26940 -1000
rect 26800 -1100 26940 -1060
rect 26800 -1160 26840 -1100
rect 26900 -1160 26940 -1100
rect 26800 -1200 26940 -1160
rect 26800 -1260 26840 -1200
rect 26900 -1260 26940 -1200
rect 26800 -1300 26940 -1260
rect 26800 -1360 26840 -1300
rect 26900 -1360 26940 -1300
rect 26800 -1380 26940 -1360
rect 26970 -1000 27110 -980
rect 26970 -1060 27010 -1000
rect 27070 -1060 27110 -1000
rect 26970 -1100 27110 -1060
rect 26970 -1160 27010 -1100
rect 27070 -1160 27110 -1100
rect 26970 -1200 27110 -1160
rect 26970 -1260 27010 -1200
rect 27070 -1260 27110 -1200
rect 26970 -1300 27110 -1260
rect 26970 -1360 27010 -1300
rect 27070 -1360 27110 -1300
rect 26970 -1380 27110 -1360
rect 27140 -1000 27280 -980
rect 27140 -1060 27180 -1000
rect 27240 -1060 27280 -1000
rect 27140 -1100 27280 -1060
rect 27140 -1160 27180 -1100
rect 27240 -1160 27280 -1100
rect 27140 -1200 27280 -1160
rect 27140 -1260 27180 -1200
rect 27240 -1260 27280 -1200
rect 27140 -1300 27280 -1260
rect 27140 -1360 27180 -1300
rect 27240 -1360 27280 -1300
rect 27140 -1380 27280 -1360
rect 27310 -1000 27450 -980
rect 27310 -1060 27350 -1000
rect 27410 -1060 27450 -1000
rect 27310 -1100 27450 -1060
rect 27310 -1160 27350 -1100
rect 27410 -1160 27450 -1100
rect 27310 -1200 27450 -1160
rect 27310 -1260 27350 -1200
rect 27410 -1260 27450 -1200
rect 27310 -1300 27450 -1260
rect 27310 -1360 27350 -1300
rect 27410 -1360 27450 -1300
rect 27310 -1380 27450 -1360
rect 27480 -1000 27620 -980
rect 27480 -1060 27520 -1000
rect 27580 -1060 27620 -1000
rect 27480 -1100 27620 -1060
rect 27480 -1160 27520 -1100
rect 27580 -1160 27620 -1100
rect 27480 -1200 27620 -1160
rect 27480 -1260 27520 -1200
rect 27580 -1260 27620 -1200
rect 27480 -1300 27620 -1260
rect 27480 -1360 27520 -1300
rect 27580 -1360 27620 -1300
rect 27480 -1380 27620 -1360
rect 27650 -1000 27790 -980
rect 27650 -1060 27690 -1000
rect 27750 -1060 27790 -1000
rect 27650 -1100 27790 -1060
rect 27650 -1160 27690 -1100
rect 27750 -1160 27790 -1100
rect 27650 -1200 27790 -1160
rect 27650 -1260 27690 -1200
rect 27750 -1260 27790 -1200
rect 27650 -1300 27790 -1260
rect 27650 -1360 27690 -1300
rect 27750 -1360 27790 -1300
rect 27650 -1380 27790 -1360
rect 27820 -1000 27960 -980
rect 27820 -1060 27860 -1000
rect 27920 -1060 27960 -1000
rect 27820 -1100 27960 -1060
rect 27820 -1160 27860 -1100
rect 27920 -1160 27960 -1100
rect 27820 -1200 27960 -1160
rect 27820 -1260 27860 -1200
rect 27920 -1260 27960 -1200
rect 27820 -1300 27960 -1260
rect 27820 -1360 27860 -1300
rect 27920 -1360 27960 -1300
rect 27820 -1380 27960 -1360
rect 27990 -1000 28130 -980
rect 27990 -1060 28030 -1000
rect 28090 -1060 28130 -1000
rect 27990 -1100 28130 -1060
rect 27990 -1160 28030 -1100
rect 28090 -1160 28130 -1100
rect 27990 -1200 28130 -1160
rect 27990 -1260 28030 -1200
rect 28090 -1260 28130 -1200
rect 27990 -1300 28130 -1260
rect 27990 -1360 28030 -1300
rect 28090 -1360 28130 -1300
rect 27990 -1380 28130 -1360
rect 28160 -1000 28300 -980
rect 28160 -1060 28200 -1000
rect 28260 -1060 28300 -1000
rect 28160 -1100 28300 -1060
rect 28160 -1160 28200 -1100
rect 28260 -1160 28300 -1100
rect 28160 -1200 28300 -1160
rect 28160 -1260 28200 -1200
rect 28260 -1260 28300 -1200
rect 28160 -1300 28300 -1260
rect 28160 -1360 28200 -1300
rect 28260 -1360 28300 -1300
rect 28160 -1380 28300 -1360
rect 28330 -1000 28470 -980
rect 28330 -1060 28370 -1000
rect 28430 -1060 28470 -1000
rect 28330 -1100 28470 -1060
rect 28330 -1160 28370 -1100
rect 28430 -1160 28470 -1100
rect 28330 -1200 28470 -1160
rect 28330 -1260 28370 -1200
rect 28430 -1260 28470 -1200
rect 28330 -1300 28470 -1260
rect 28330 -1360 28370 -1300
rect 28430 -1360 28470 -1300
rect 28330 -1380 28470 -1360
rect 28500 -1000 28640 -980
rect 28500 -1060 28540 -1000
rect 28600 -1060 28640 -1000
rect 28500 -1100 28640 -1060
rect 28500 -1160 28540 -1100
rect 28600 -1160 28640 -1100
rect 28500 -1200 28640 -1160
rect 28500 -1260 28540 -1200
rect 28600 -1260 28640 -1200
rect 28500 -1300 28640 -1260
rect 28500 -1360 28540 -1300
rect 28600 -1360 28640 -1300
rect 28500 -1380 28640 -1360
rect 28670 -1000 28810 -980
rect 28670 -1060 28710 -1000
rect 28770 -1060 28810 -1000
rect 28670 -1100 28810 -1060
rect 28670 -1160 28710 -1100
rect 28770 -1160 28810 -1100
rect 28670 -1200 28810 -1160
rect 28670 -1260 28710 -1200
rect 28770 -1260 28810 -1200
rect 28670 -1300 28810 -1260
rect 28670 -1360 28710 -1300
rect 28770 -1360 28810 -1300
rect 28670 -1380 28810 -1360
rect 28840 -1000 28980 -980
rect 28840 -1060 28880 -1000
rect 28940 -1060 28980 -1000
rect 28840 -1100 28980 -1060
rect 28840 -1160 28880 -1100
rect 28940 -1160 28980 -1100
rect 28840 -1200 28980 -1160
rect 28840 -1260 28880 -1200
rect 28940 -1260 28980 -1200
rect 28840 -1300 28980 -1260
rect 28840 -1360 28880 -1300
rect 28940 -1360 28980 -1300
rect 28840 -1380 28980 -1360
rect 29010 -1000 29150 -980
rect 29010 -1060 29050 -1000
rect 29110 -1060 29150 -1000
rect 29010 -1100 29150 -1060
rect 29010 -1160 29050 -1100
rect 29110 -1160 29150 -1100
rect 29010 -1200 29150 -1160
rect 29010 -1260 29050 -1200
rect 29110 -1260 29150 -1200
rect 29010 -1300 29150 -1260
rect 29010 -1360 29050 -1300
rect 29110 -1360 29150 -1300
rect 29010 -1380 29150 -1360
rect 29180 -1000 29320 -980
rect 29180 -1060 29220 -1000
rect 29280 -1060 29320 -1000
rect 29180 -1100 29320 -1060
rect 29180 -1160 29220 -1100
rect 29280 -1160 29320 -1100
rect 29180 -1200 29320 -1160
rect 29180 -1260 29220 -1200
rect 29280 -1260 29320 -1200
rect 29180 -1300 29320 -1260
rect 29180 -1360 29220 -1300
rect 29280 -1360 29320 -1300
rect 29180 -1380 29320 -1360
rect 29350 -1000 29490 -980
rect 29350 -1060 29390 -1000
rect 29450 -1060 29490 -1000
rect 29350 -1100 29490 -1060
rect 29350 -1160 29390 -1100
rect 29450 -1160 29490 -1100
rect 29350 -1200 29490 -1160
rect 29350 -1260 29390 -1200
rect 29450 -1260 29490 -1200
rect 29350 -1300 29490 -1260
rect 29350 -1360 29390 -1300
rect 29450 -1360 29490 -1300
rect 29350 -1380 29490 -1360
rect 29520 -1000 29660 -980
rect 29520 -1060 29560 -1000
rect 29620 -1060 29660 -1000
rect 29520 -1100 29660 -1060
rect 29520 -1160 29560 -1100
rect 29620 -1160 29660 -1100
rect 29520 -1200 29660 -1160
rect 29520 -1260 29560 -1200
rect 29620 -1260 29660 -1200
rect 29520 -1300 29660 -1260
rect 29520 -1360 29560 -1300
rect 29620 -1360 29660 -1300
rect 29520 -1380 29660 -1360
rect 29690 -1000 29830 -980
rect 29690 -1060 29730 -1000
rect 29790 -1060 29830 -1000
rect 29690 -1100 29830 -1060
rect 29690 -1160 29730 -1100
rect 29790 -1160 29830 -1100
rect 29690 -1200 29830 -1160
rect 29690 -1260 29730 -1200
rect 29790 -1260 29830 -1200
rect 29690 -1300 29830 -1260
rect 29690 -1360 29730 -1300
rect 29790 -1360 29830 -1300
rect 29690 -1380 29830 -1360
rect 29860 -1000 30000 -980
rect 29860 -1060 29900 -1000
rect 29960 -1060 30000 -1000
rect 29860 -1100 30000 -1060
rect 29860 -1160 29900 -1100
rect 29960 -1160 30000 -1100
rect 29860 -1200 30000 -1160
rect 29860 -1260 29900 -1200
rect 29960 -1260 30000 -1200
rect 29860 -1300 30000 -1260
rect 29860 -1360 29900 -1300
rect 29960 -1360 30000 -1300
rect 29860 -1380 30000 -1360
rect 30030 -1000 30170 -980
rect 30030 -1060 30070 -1000
rect 30130 -1060 30170 -1000
rect 30030 -1100 30170 -1060
rect 30030 -1160 30070 -1100
rect 30130 -1160 30170 -1100
rect 30030 -1200 30170 -1160
rect 30030 -1260 30070 -1200
rect 30130 -1260 30170 -1200
rect 30030 -1300 30170 -1260
rect 30030 -1360 30070 -1300
rect 30130 -1360 30170 -1300
rect 30030 -1380 30170 -1360
rect 30200 -1000 30340 -980
rect 30200 -1060 30240 -1000
rect 30300 -1060 30340 -1000
rect 30200 -1100 30340 -1060
rect 30200 -1160 30240 -1100
rect 30300 -1160 30340 -1100
rect 30200 -1200 30340 -1160
rect 30200 -1260 30240 -1200
rect 30300 -1260 30340 -1200
rect 30200 -1300 30340 -1260
rect 30200 -1360 30240 -1300
rect 30300 -1360 30340 -1300
rect 30200 -1380 30340 -1360
rect 30370 -1000 30510 -980
rect 30370 -1060 30410 -1000
rect 30470 -1060 30510 -1000
rect 30370 -1100 30510 -1060
rect 30370 -1160 30410 -1100
rect 30470 -1160 30510 -1100
rect 30370 -1200 30510 -1160
rect 30370 -1260 30410 -1200
rect 30470 -1260 30510 -1200
rect 30370 -1300 30510 -1260
rect 30370 -1360 30410 -1300
rect 30470 -1360 30510 -1300
rect 30370 -1380 30510 -1360
rect 30540 -1000 30680 -980
rect 30540 -1060 30580 -1000
rect 30640 -1060 30680 -1000
rect 30540 -1100 30680 -1060
rect 30540 -1160 30580 -1100
rect 30640 -1160 30680 -1100
rect 30540 -1200 30680 -1160
rect 30540 -1260 30580 -1200
rect 30640 -1260 30680 -1200
rect 30540 -1300 30680 -1260
rect 30540 -1360 30580 -1300
rect 30640 -1360 30680 -1300
rect 30540 -1380 30680 -1360
rect 30710 -1000 30850 -980
rect 30710 -1060 30750 -1000
rect 30810 -1060 30850 -1000
rect 30710 -1100 30850 -1060
rect 30710 -1160 30750 -1100
rect 30810 -1160 30850 -1100
rect 30710 -1200 30850 -1160
rect 30710 -1260 30750 -1200
rect 30810 -1260 30850 -1200
rect 30710 -1300 30850 -1260
rect 30710 -1360 30750 -1300
rect 30810 -1360 30850 -1300
rect 30710 -1380 30850 -1360
rect 30880 -1000 31020 -980
rect 30880 -1060 30920 -1000
rect 30980 -1060 31020 -1000
rect 30880 -1100 31020 -1060
rect 30880 -1160 30920 -1100
rect 30980 -1160 31020 -1100
rect 30880 -1200 31020 -1160
rect 30880 -1260 30920 -1200
rect 30980 -1260 31020 -1200
rect 30880 -1300 31020 -1260
rect 30880 -1360 30920 -1300
rect 30980 -1360 31020 -1300
rect 30880 -1380 31020 -1360
rect 31050 -1000 31190 -980
rect 31050 -1060 31090 -1000
rect 31150 -1060 31190 -1000
rect 31050 -1100 31190 -1060
rect 31050 -1160 31090 -1100
rect 31150 -1160 31190 -1100
rect 31050 -1200 31190 -1160
rect 31050 -1260 31090 -1200
rect 31150 -1260 31190 -1200
rect 31050 -1300 31190 -1260
rect 31050 -1360 31090 -1300
rect 31150 -1360 31190 -1300
rect 31050 -1380 31190 -1360
rect 31220 -1000 31360 -980
rect 31220 -1060 31260 -1000
rect 31320 -1060 31360 -1000
rect 31220 -1100 31360 -1060
rect 31220 -1160 31260 -1100
rect 31320 -1160 31360 -1100
rect 31220 -1200 31360 -1160
rect 31220 -1260 31260 -1200
rect 31320 -1260 31360 -1200
rect 31220 -1300 31360 -1260
rect 31220 -1360 31260 -1300
rect 31320 -1360 31360 -1300
rect 31220 -1380 31360 -1360
rect 31390 -1000 31530 -980
rect 31390 -1060 31430 -1000
rect 31490 -1060 31530 -1000
rect 31390 -1100 31530 -1060
rect 31390 -1160 31430 -1100
rect 31490 -1160 31530 -1100
rect 31390 -1200 31530 -1160
rect 31390 -1260 31430 -1200
rect 31490 -1260 31530 -1200
rect 31390 -1300 31530 -1260
rect 31390 -1360 31430 -1300
rect 31490 -1360 31530 -1300
rect 31390 -1380 31530 -1360
rect 31560 -1000 31700 -980
rect 31560 -1060 31600 -1000
rect 31660 -1060 31700 -1000
rect 31560 -1100 31700 -1060
rect 31560 -1160 31600 -1100
rect 31660 -1160 31700 -1100
rect 31560 -1200 31700 -1160
rect 31560 -1260 31600 -1200
rect 31660 -1260 31700 -1200
rect 31560 -1300 31700 -1260
rect 31560 -1360 31600 -1300
rect 31660 -1360 31700 -1300
rect 31560 -1380 31700 -1360
rect 31730 -1000 31870 -980
rect 31730 -1060 31770 -1000
rect 31830 -1060 31870 -1000
rect 31730 -1100 31870 -1060
rect 31730 -1160 31770 -1100
rect 31830 -1160 31870 -1100
rect 31730 -1200 31870 -1160
rect 31730 -1260 31770 -1200
rect 31830 -1260 31870 -1200
rect 31730 -1300 31870 -1260
rect 31730 -1360 31770 -1300
rect 31830 -1360 31870 -1300
rect 31730 -1380 31870 -1360
rect 31900 -1000 32040 -980
rect 31900 -1060 31940 -1000
rect 32000 -1060 32040 -1000
rect 31900 -1100 32040 -1060
rect 31900 -1160 31940 -1100
rect 32000 -1160 32040 -1100
rect 31900 -1200 32040 -1160
rect 31900 -1260 31940 -1200
rect 32000 -1260 32040 -1200
rect 31900 -1300 32040 -1260
rect 31900 -1360 31940 -1300
rect 32000 -1360 32040 -1300
rect 31900 -1380 32040 -1360
rect 32070 -1000 32210 -980
rect 32070 -1060 32110 -1000
rect 32170 -1060 32210 -1000
rect 32070 -1100 32210 -1060
rect 32070 -1160 32110 -1100
rect 32170 -1160 32210 -1100
rect 32070 -1200 32210 -1160
rect 32070 -1260 32110 -1200
rect 32170 -1260 32210 -1200
rect 32070 -1300 32210 -1260
rect 32070 -1360 32110 -1300
rect 32170 -1360 32210 -1300
rect 32070 -1380 32210 -1360
rect 32240 -1000 32380 -980
rect 32240 -1060 32280 -1000
rect 32340 -1060 32380 -1000
rect 32240 -1100 32380 -1060
rect 32240 -1160 32280 -1100
rect 32340 -1160 32380 -1100
rect 32240 -1200 32380 -1160
rect 32240 -1260 32280 -1200
rect 32340 -1260 32380 -1200
rect 32240 -1300 32380 -1260
rect 32240 -1360 32280 -1300
rect 32340 -1360 32380 -1300
rect 32240 -1380 32380 -1360
rect 32410 -1000 32550 -980
rect 32410 -1060 32450 -1000
rect 32510 -1060 32550 -1000
rect 32410 -1100 32550 -1060
rect 32410 -1160 32450 -1100
rect 32510 -1160 32550 -1100
rect 32410 -1200 32550 -1160
rect 32410 -1260 32450 -1200
rect 32510 -1260 32550 -1200
rect 32410 -1300 32550 -1260
rect 32410 -1360 32450 -1300
rect 32510 -1360 32550 -1300
rect 32410 -1380 32550 -1360
rect 32580 -1000 32720 -980
rect 32580 -1060 32620 -1000
rect 32680 -1060 32720 -1000
rect 32580 -1100 32720 -1060
rect 32580 -1160 32620 -1100
rect 32680 -1160 32720 -1100
rect 32580 -1200 32720 -1160
rect 32580 -1260 32620 -1200
rect 32680 -1260 32720 -1200
rect 32580 -1300 32720 -1260
rect 32580 -1360 32620 -1300
rect 32680 -1360 32720 -1300
rect 32580 -1380 32720 -1360
rect 32750 -1000 32890 -980
rect 32750 -1060 32790 -1000
rect 32850 -1060 32890 -1000
rect 32750 -1100 32890 -1060
rect 32750 -1160 32790 -1100
rect 32850 -1160 32890 -1100
rect 32750 -1200 32890 -1160
rect 32750 -1260 32790 -1200
rect 32850 -1260 32890 -1200
rect 32750 -1300 32890 -1260
rect 32750 -1360 32790 -1300
rect 32850 -1360 32890 -1300
rect 32750 -1380 32890 -1360
rect 32920 -1000 33060 -980
rect 32920 -1060 32960 -1000
rect 33020 -1060 33060 -1000
rect 32920 -1100 33060 -1060
rect 32920 -1160 32960 -1100
rect 33020 -1160 33060 -1100
rect 32920 -1200 33060 -1160
rect 32920 -1260 32960 -1200
rect 33020 -1260 33060 -1200
rect 32920 -1300 33060 -1260
rect 32920 -1360 32960 -1300
rect 33020 -1360 33060 -1300
rect 32920 -1380 33060 -1360
rect 33090 -1000 33230 -980
rect 33090 -1060 33130 -1000
rect 33190 -1060 33230 -1000
rect 33090 -1100 33230 -1060
rect 33090 -1160 33130 -1100
rect 33190 -1160 33230 -1100
rect 33090 -1200 33230 -1160
rect 33090 -1260 33130 -1200
rect 33190 -1260 33230 -1200
rect 33090 -1300 33230 -1260
rect 33090 -1360 33130 -1300
rect 33190 -1360 33230 -1300
rect 33090 -1380 33230 -1360
rect 33260 -1000 33400 -980
rect 33260 -1060 33300 -1000
rect 33360 -1060 33400 -1000
rect 33260 -1100 33400 -1060
rect 33260 -1160 33300 -1100
rect 33360 -1160 33400 -1100
rect 33260 -1200 33400 -1160
rect 33260 -1260 33300 -1200
rect 33360 -1260 33400 -1200
rect 33260 -1300 33400 -1260
rect 33260 -1360 33300 -1300
rect 33360 -1360 33400 -1300
rect 33260 -1380 33400 -1360
rect 33430 -1000 33570 -980
rect 33430 -1060 33470 -1000
rect 33530 -1060 33570 -1000
rect 33430 -1100 33570 -1060
rect 33430 -1160 33470 -1100
rect 33530 -1160 33570 -1100
rect 33430 -1200 33570 -1160
rect 33430 -1260 33470 -1200
rect 33530 -1260 33570 -1200
rect 33430 -1300 33570 -1260
rect 33430 -1360 33470 -1300
rect 33530 -1360 33570 -1300
rect 33430 -1380 33570 -1360
rect 33600 -1000 33740 -980
rect 33600 -1060 33640 -1000
rect 33700 -1060 33740 -1000
rect 33600 -1100 33740 -1060
rect 33600 -1160 33640 -1100
rect 33700 -1160 33740 -1100
rect 33600 -1200 33740 -1160
rect 33600 -1260 33640 -1200
rect 33700 -1260 33740 -1200
rect 33600 -1300 33740 -1260
rect 33600 -1360 33640 -1300
rect 33700 -1360 33740 -1300
rect 33600 -1380 33740 -1360
rect 33770 -1000 33910 -980
rect 33770 -1060 33810 -1000
rect 33870 -1060 33910 -1000
rect 33770 -1100 33910 -1060
rect 33770 -1160 33810 -1100
rect 33870 -1160 33910 -1100
rect 33770 -1200 33910 -1160
rect 33770 -1260 33810 -1200
rect 33870 -1260 33910 -1200
rect 33770 -1300 33910 -1260
rect 33770 -1360 33810 -1300
rect 33870 -1360 33910 -1300
rect 33770 -1380 33910 -1360
rect 33940 -1000 34080 -980
rect 33940 -1060 33980 -1000
rect 34040 -1060 34080 -1000
rect 33940 -1100 34080 -1060
rect 33940 -1160 33980 -1100
rect 34040 -1160 34080 -1100
rect 33940 -1200 34080 -1160
rect 33940 -1260 33980 -1200
rect 34040 -1260 34080 -1200
rect 33940 -1300 34080 -1260
rect 33940 -1360 33980 -1300
rect 34040 -1360 34080 -1300
rect 33940 -1380 34080 -1360
rect 34110 -1000 34250 -980
rect 34110 -1060 34150 -1000
rect 34210 -1060 34250 -1000
rect 34110 -1100 34250 -1060
rect 34110 -1160 34150 -1100
rect 34210 -1160 34250 -1100
rect 34110 -1200 34250 -1160
rect 34110 -1260 34150 -1200
rect 34210 -1260 34250 -1200
rect 34110 -1300 34250 -1260
rect 34110 -1360 34150 -1300
rect 34210 -1360 34250 -1300
rect 34110 -1380 34250 -1360
rect 34280 -1000 34420 -980
rect 34280 -1060 34320 -1000
rect 34380 -1060 34420 -1000
rect 34280 -1100 34420 -1060
rect 34280 -1160 34320 -1100
rect 34380 -1160 34420 -1100
rect 34280 -1200 34420 -1160
rect 34280 -1260 34320 -1200
rect 34380 -1260 34420 -1200
rect 34280 -1300 34420 -1260
rect 34280 -1360 34320 -1300
rect 34380 -1360 34420 -1300
rect 34280 -1380 34420 -1360
rect 34450 -1000 34590 -980
rect 34450 -1060 34490 -1000
rect 34550 -1060 34590 -1000
rect 34450 -1100 34590 -1060
rect 34450 -1160 34490 -1100
rect 34550 -1160 34590 -1100
rect 34450 -1200 34590 -1160
rect 34450 -1260 34490 -1200
rect 34550 -1260 34590 -1200
rect 34450 -1300 34590 -1260
rect 34450 -1360 34490 -1300
rect 34550 -1360 34590 -1300
rect 34450 -1380 34590 -1360
rect 34620 -1000 34760 -980
rect 34620 -1060 34660 -1000
rect 34720 -1060 34760 -1000
rect 34620 -1100 34760 -1060
rect 34620 -1160 34660 -1100
rect 34720 -1160 34760 -1100
rect 34620 -1200 34760 -1160
rect 34620 -1260 34660 -1200
rect 34720 -1260 34760 -1200
rect 34620 -1300 34760 -1260
rect 34620 -1360 34660 -1300
rect 34720 -1360 34760 -1300
rect 34620 -1380 34760 -1360
rect 34790 -1000 34930 -980
rect 34790 -1060 34830 -1000
rect 34890 -1060 34930 -1000
rect 34790 -1100 34930 -1060
rect 34790 -1160 34830 -1100
rect 34890 -1160 34930 -1100
rect 34790 -1200 34930 -1160
rect 34790 -1260 34830 -1200
rect 34890 -1260 34930 -1200
rect 34790 -1300 34930 -1260
rect 34790 -1360 34830 -1300
rect 34890 -1360 34930 -1300
rect 34790 -1380 34930 -1360
rect 34960 -1000 35100 -980
rect 34960 -1060 35000 -1000
rect 35060 -1060 35100 -1000
rect 34960 -1100 35100 -1060
rect 34960 -1160 35000 -1100
rect 35060 -1160 35100 -1100
rect 34960 -1200 35100 -1160
rect 34960 -1260 35000 -1200
rect 35060 -1260 35100 -1200
rect 34960 -1300 35100 -1260
rect 34960 -1360 35000 -1300
rect 35060 -1360 35100 -1300
rect 34960 -1380 35100 -1360
rect 35130 -1000 35270 -980
rect 35130 -1060 35170 -1000
rect 35230 -1060 35270 -1000
rect 35130 -1100 35270 -1060
rect 35130 -1160 35170 -1100
rect 35230 -1160 35270 -1100
rect 35130 -1200 35270 -1160
rect 35130 -1260 35170 -1200
rect 35230 -1260 35270 -1200
rect 35130 -1300 35270 -1260
rect 35130 -1360 35170 -1300
rect 35230 -1360 35270 -1300
rect 35130 -1380 35270 -1360
rect 35300 -1000 35440 -980
rect 35300 -1060 35340 -1000
rect 35400 -1060 35440 -1000
rect 35300 -1100 35440 -1060
rect 35300 -1160 35340 -1100
rect 35400 -1160 35440 -1100
rect 35300 -1200 35440 -1160
rect 35300 -1260 35340 -1200
rect 35400 -1260 35440 -1200
rect 35300 -1300 35440 -1260
rect 35300 -1360 35340 -1300
rect 35400 -1360 35440 -1300
rect 35300 -1380 35440 -1360
rect 35470 -1000 35610 -980
rect 35470 -1060 35510 -1000
rect 35570 -1060 35610 -1000
rect 35470 -1100 35610 -1060
rect 35470 -1160 35510 -1100
rect 35570 -1160 35610 -1100
rect 35470 -1200 35610 -1160
rect 35470 -1260 35510 -1200
rect 35570 -1260 35610 -1200
rect 35470 -1300 35610 -1260
rect 35470 -1360 35510 -1300
rect 35570 -1360 35610 -1300
rect 35470 -1380 35610 -1360
rect 35640 -1000 35780 -980
rect 35640 -1060 35680 -1000
rect 35740 -1060 35780 -1000
rect 35640 -1100 35780 -1060
rect 35640 -1160 35680 -1100
rect 35740 -1160 35780 -1100
rect 35640 -1200 35780 -1160
rect 35640 -1260 35680 -1200
rect 35740 -1260 35780 -1200
rect 35640 -1300 35780 -1260
rect 35640 -1360 35680 -1300
rect 35740 -1360 35780 -1300
rect 35640 -1380 35780 -1360
rect 35810 -1000 35950 -980
rect 35810 -1060 35850 -1000
rect 35910 -1060 35950 -1000
rect 35810 -1100 35950 -1060
rect 35810 -1160 35850 -1100
rect 35910 -1160 35950 -1100
rect 35810 -1200 35950 -1160
rect 35810 -1260 35850 -1200
rect 35910 -1260 35950 -1200
rect 35810 -1300 35950 -1260
rect 35810 -1360 35850 -1300
rect 35910 -1360 35950 -1300
rect 35810 -1380 35950 -1360
rect 35980 -1000 36120 -980
rect 35980 -1060 36020 -1000
rect 36080 -1060 36120 -1000
rect 35980 -1100 36120 -1060
rect 35980 -1160 36020 -1100
rect 36080 -1160 36120 -1100
rect 35980 -1200 36120 -1160
rect 35980 -1260 36020 -1200
rect 36080 -1260 36120 -1200
rect 35980 -1300 36120 -1260
rect 35980 -1360 36020 -1300
rect 36080 -1360 36120 -1300
rect 35980 -1380 36120 -1360
rect 36150 -1000 36290 -980
rect 36150 -1060 36190 -1000
rect 36250 -1060 36290 -1000
rect 36150 -1100 36290 -1060
rect 36150 -1160 36190 -1100
rect 36250 -1160 36290 -1100
rect 36150 -1200 36290 -1160
rect 36150 -1260 36190 -1200
rect 36250 -1260 36290 -1200
rect 36150 -1300 36290 -1260
rect 36150 -1360 36190 -1300
rect 36250 -1360 36290 -1300
rect 36150 -1380 36290 -1360
rect 36320 -1000 36460 -980
rect 36320 -1060 36360 -1000
rect 36420 -1060 36460 -1000
rect 36320 -1100 36460 -1060
rect 36320 -1160 36360 -1100
rect 36420 -1160 36460 -1100
rect 36320 -1200 36460 -1160
rect 36320 -1260 36360 -1200
rect 36420 -1260 36460 -1200
rect 36320 -1300 36460 -1260
rect 36320 -1360 36360 -1300
rect 36420 -1360 36460 -1300
rect 36320 -1380 36460 -1360
rect 36490 -1000 36630 -980
rect 36490 -1060 36530 -1000
rect 36590 -1060 36630 -1000
rect 36490 -1100 36630 -1060
rect 36490 -1160 36530 -1100
rect 36590 -1160 36630 -1100
rect 36490 -1200 36630 -1160
rect 36490 -1260 36530 -1200
rect 36590 -1260 36630 -1200
rect 36490 -1300 36630 -1260
rect 36490 -1360 36530 -1300
rect 36590 -1360 36630 -1300
rect 36490 -1380 36630 -1360
rect 36660 -1000 36800 -980
rect 36660 -1060 36700 -1000
rect 36760 -1060 36800 -1000
rect 36660 -1100 36800 -1060
rect 36660 -1160 36700 -1100
rect 36760 -1160 36800 -1100
rect 36660 -1200 36800 -1160
rect 36660 -1260 36700 -1200
rect 36760 -1260 36800 -1200
rect 36660 -1300 36800 -1260
rect 36660 -1360 36700 -1300
rect 36760 -1360 36800 -1300
rect 36660 -1380 36800 -1360
rect 36830 -1000 36970 -980
rect 36830 -1060 36870 -1000
rect 36930 -1060 36970 -1000
rect 36830 -1100 36970 -1060
rect 36830 -1160 36870 -1100
rect 36930 -1160 36970 -1100
rect 36830 -1200 36970 -1160
rect 36830 -1260 36870 -1200
rect 36930 -1260 36970 -1200
rect 36830 -1300 36970 -1260
rect 36830 -1360 36870 -1300
rect 36930 -1360 36970 -1300
rect 36830 -1380 36970 -1360
rect 37000 -1000 37140 -980
rect 37000 -1060 37040 -1000
rect 37100 -1060 37140 -1000
rect 37000 -1100 37140 -1060
rect 37000 -1160 37040 -1100
rect 37100 -1160 37140 -1100
rect 37000 -1200 37140 -1160
rect 37000 -1260 37040 -1200
rect 37100 -1260 37140 -1200
rect 37000 -1300 37140 -1260
rect 37000 -1360 37040 -1300
rect 37100 -1360 37140 -1300
rect 37000 -1380 37140 -1360
rect 37170 -1000 37310 -980
rect 37170 -1060 37210 -1000
rect 37270 -1060 37310 -1000
rect 37170 -1100 37310 -1060
rect 37170 -1160 37210 -1100
rect 37270 -1160 37310 -1100
rect 37170 -1200 37310 -1160
rect 37170 -1260 37210 -1200
rect 37270 -1260 37310 -1200
rect 37170 -1300 37310 -1260
rect 37170 -1360 37210 -1300
rect 37270 -1360 37310 -1300
rect 37170 -1380 37310 -1360
rect 37340 -1000 37480 -980
rect 37340 -1060 37380 -1000
rect 37440 -1060 37480 -1000
rect 37340 -1100 37480 -1060
rect 37340 -1160 37380 -1100
rect 37440 -1160 37480 -1100
rect 37340 -1200 37480 -1160
rect 37340 -1260 37380 -1200
rect 37440 -1260 37480 -1200
rect 37340 -1300 37480 -1260
rect 37340 -1360 37380 -1300
rect 37440 -1360 37480 -1300
rect 37340 -1380 37480 -1360
rect 37510 -1000 37650 -980
rect 37510 -1060 37550 -1000
rect 37610 -1060 37650 -1000
rect 37510 -1100 37650 -1060
rect 37510 -1160 37550 -1100
rect 37610 -1160 37650 -1100
rect 37510 -1200 37650 -1160
rect 37510 -1260 37550 -1200
rect 37610 -1260 37650 -1200
rect 37510 -1300 37650 -1260
rect 37510 -1360 37550 -1300
rect 37610 -1360 37650 -1300
rect 37510 -1380 37650 -1360
rect 37680 -1000 37820 -980
rect 37680 -1060 37720 -1000
rect 37780 -1060 37820 -1000
rect 37680 -1100 37820 -1060
rect 37680 -1160 37720 -1100
rect 37780 -1160 37820 -1100
rect 37680 -1200 37820 -1160
rect 37680 -1260 37720 -1200
rect 37780 -1260 37820 -1200
rect 37680 -1300 37820 -1260
rect 37680 -1360 37720 -1300
rect 37780 -1360 37820 -1300
rect 37680 -1380 37820 -1360
rect 37850 -1000 37990 -980
rect 37850 -1060 37890 -1000
rect 37950 -1060 37990 -1000
rect 37850 -1100 37990 -1060
rect 37850 -1160 37890 -1100
rect 37950 -1160 37990 -1100
rect 37850 -1200 37990 -1160
rect 37850 -1260 37890 -1200
rect 37950 -1260 37990 -1200
rect 37850 -1300 37990 -1260
rect 37850 -1360 37890 -1300
rect 37950 -1360 37990 -1300
rect 37850 -1380 37990 -1360
rect 38020 -1000 38160 -980
rect 38020 -1060 38060 -1000
rect 38120 -1060 38160 -1000
rect 38020 -1100 38160 -1060
rect 38020 -1160 38060 -1100
rect 38120 -1160 38160 -1100
rect 38020 -1200 38160 -1160
rect 38020 -1260 38060 -1200
rect 38120 -1260 38160 -1200
rect 38020 -1300 38160 -1260
rect 38020 -1360 38060 -1300
rect 38120 -1360 38160 -1300
rect 38020 -1380 38160 -1360
rect 38190 -1000 38330 -980
rect 38190 -1060 38230 -1000
rect 38290 -1060 38330 -1000
rect 38190 -1100 38330 -1060
rect 38190 -1160 38230 -1100
rect 38290 -1160 38330 -1100
rect 38190 -1200 38330 -1160
rect 38190 -1260 38230 -1200
rect 38290 -1260 38330 -1200
rect 38190 -1300 38330 -1260
rect 38190 -1360 38230 -1300
rect 38290 -1360 38330 -1300
rect 38190 -1380 38330 -1360
rect 38360 -1000 38500 -980
rect 38360 -1060 38400 -1000
rect 38460 -1060 38500 -1000
rect 38360 -1100 38500 -1060
rect 38360 -1160 38400 -1100
rect 38460 -1160 38500 -1100
rect 38360 -1200 38500 -1160
rect 38360 -1260 38400 -1200
rect 38460 -1260 38500 -1200
rect 38360 -1300 38500 -1260
rect 38360 -1360 38400 -1300
rect 38460 -1360 38500 -1300
rect 38360 -1380 38500 -1360
rect 38530 -1000 38670 -980
rect 38530 -1060 38570 -1000
rect 38630 -1060 38670 -1000
rect 38530 -1100 38670 -1060
rect 38530 -1160 38570 -1100
rect 38630 -1160 38670 -1100
rect 38530 -1200 38670 -1160
rect 38530 -1260 38570 -1200
rect 38630 -1260 38670 -1200
rect 38530 -1300 38670 -1260
rect 38530 -1360 38570 -1300
rect 38630 -1360 38670 -1300
rect 38530 -1380 38670 -1360
rect 38700 -1000 38840 -980
rect 38700 -1060 38740 -1000
rect 38800 -1060 38840 -1000
rect 38700 -1100 38840 -1060
rect 38700 -1160 38740 -1100
rect 38800 -1160 38840 -1100
rect 38700 -1200 38840 -1160
rect 38700 -1260 38740 -1200
rect 38800 -1260 38840 -1200
rect 38700 -1300 38840 -1260
rect 38700 -1360 38740 -1300
rect 38800 -1360 38840 -1300
rect 38700 -1380 38840 -1360
rect 38870 -1000 39010 -980
rect 38870 -1060 38910 -1000
rect 38970 -1060 39010 -1000
rect 38870 -1100 39010 -1060
rect 38870 -1160 38910 -1100
rect 38970 -1160 39010 -1100
rect 38870 -1200 39010 -1160
rect 38870 -1260 38910 -1200
rect 38970 -1260 39010 -1200
rect 38870 -1300 39010 -1260
rect 38870 -1360 38910 -1300
rect 38970 -1360 39010 -1300
rect 38870 -1380 39010 -1360
rect 39040 -1000 39180 -980
rect 39040 -1060 39080 -1000
rect 39140 -1060 39180 -1000
rect 39040 -1100 39180 -1060
rect 39040 -1160 39080 -1100
rect 39140 -1160 39180 -1100
rect 39040 -1200 39180 -1160
rect 39040 -1260 39080 -1200
rect 39140 -1260 39180 -1200
rect 39040 -1300 39180 -1260
rect 39040 -1360 39080 -1300
rect 39140 -1360 39180 -1300
rect 39040 -1380 39180 -1360
rect 39210 -1000 39350 -980
rect 39210 -1060 39250 -1000
rect 39310 -1060 39350 -1000
rect 39210 -1100 39350 -1060
rect 39210 -1160 39250 -1100
rect 39310 -1160 39350 -1100
rect 39210 -1200 39350 -1160
rect 39210 -1260 39250 -1200
rect 39310 -1260 39350 -1200
rect 39210 -1300 39350 -1260
rect 39210 -1360 39250 -1300
rect 39310 -1360 39350 -1300
rect 39210 -1380 39350 -1360
rect 39380 -1000 39520 -980
rect 39380 -1060 39420 -1000
rect 39480 -1060 39520 -1000
rect 39380 -1100 39520 -1060
rect 39380 -1160 39420 -1100
rect 39480 -1160 39520 -1100
rect 39380 -1200 39520 -1160
rect 39380 -1260 39420 -1200
rect 39480 -1260 39520 -1200
rect 39380 -1300 39520 -1260
rect 39380 -1360 39420 -1300
rect 39480 -1360 39520 -1300
rect 39380 -1380 39520 -1360
rect 39550 -1000 39690 -980
rect 39550 -1060 39590 -1000
rect 39650 -1060 39690 -1000
rect 39550 -1100 39690 -1060
rect 39550 -1160 39590 -1100
rect 39650 -1160 39690 -1100
rect 39550 -1200 39690 -1160
rect 39550 -1260 39590 -1200
rect 39650 -1260 39690 -1200
rect 39550 -1300 39690 -1260
rect 39550 -1360 39590 -1300
rect 39650 -1360 39690 -1300
rect 39550 -1380 39690 -1360
rect 39720 -1000 39860 -980
rect 39720 -1060 39760 -1000
rect 39820 -1060 39860 -1000
rect 39720 -1100 39860 -1060
rect 39720 -1160 39760 -1100
rect 39820 -1160 39860 -1100
rect 39720 -1200 39860 -1160
rect 39720 -1260 39760 -1200
rect 39820 -1260 39860 -1200
rect 39720 -1300 39860 -1260
rect 39720 -1360 39760 -1300
rect 39820 -1360 39860 -1300
rect 39720 -1380 39860 -1360
rect 39890 -1000 40030 -980
rect 39890 -1060 39930 -1000
rect 39990 -1060 40030 -1000
rect 39890 -1100 40030 -1060
rect 39890 -1160 39930 -1100
rect 39990 -1160 40030 -1100
rect 39890 -1200 40030 -1160
rect 39890 -1260 39930 -1200
rect 39990 -1260 40030 -1200
rect 39890 -1300 40030 -1260
rect 39890 -1360 39930 -1300
rect 39990 -1360 40030 -1300
rect 39890 -1380 40030 -1360
rect 40060 -1000 40200 -980
rect 40060 -1060 40100 -1000
rect 40160 -1060 40200 -1000
rect 40060 -1100 40200 -1060
rect 40060 -1160 40100 -1100
rect 40160 -1160 40200 -1100
rect 40060 -1200 40200 -1160
rect 40060 -1260 40100 -1200
rect 40160 -1260 40200 -1200
rect 40060 -1300 40200 -1260
rect 40060 -1360 40100 -1300
rect 40160 -1360 40200 -1300
rect 40060 -1380 40200 -1360
rect 40230 -1000 40370 -980
rect 40230 -1060 40270 -1000
rect 40330 -1060 40370 -1000
rect 40230 -1100 40370 -1060
rect 40230 -1160 40270 -1100
rect 40330 -1160 40370 -1100
rect 40230 -1200 40370 -1160
rect 40230 -1260 40270 -1200
rect 40330 -1260 40370 -1200
rect 40230 -1300 40370 -1260
rect 40230 -1360 40270 -1300
rect 40330 -1360 40370 -1300
rect 40230 -1380 40370 -1360
rect 40400 -1000 40540 -980
rect 40400 -1060 40440 -1000
rect 40500 -1060 40540 -1000
rect 40400 -1100 40540 -1060
rect 40400 -1160 40440 -1100
rect 40500 -1160 40540 -1100
rect 40400 -1200 40540 -1160
rect 40400 -1260 40440 -1200
rect 40500 -1260 40540 -1200
rect 40400 -1300 40540 -1260
rect 40400 -1360 40440 -1300
rect 40500 -1360 40540 -1300
rect 40400 -1380 40540 -1360
rect 40570 -1000 40710 -980
rect 40570 -1060 40610 -1000
rect 40670 -1060 40710 -1000
rect 40570 -1100 40710 -1060
rect 40570 -1160 40610 -1100
rect 40670 -1160 40710 -1100
rect 40570 -1200 40710 -1160
rect 40570 -1260 40610 -1200
rect 40670 -1260 40710 -1200
rect 40570 -1300 40710 -1260
rect 40570 -1360 40610 -1300
rect 40670 -1360 40710 -1300
rect 40570 -1380 40710 -1360
rect 40740 -1000 40880 -980
rect 40740 -1060 40780 -1000
rect 40840 -1060 40880 -1000
rect 40740 -1100 40880 -1060
rect 40740 -1160 40780 -1100
rect 40840 -1160 40880 -1100
rect 40740 -1200 40880 -1160
rect 40740 -1260 40780 -1200
rect 40840 -1260 40880 -1200
rect 40740 -1300 40880 -1260
rect 40740 -1360 40780 -1300
rect 40840 -1360 40880 -1300
rect 40740 -1380 40880 -1360
rect 40910 -1000 41050 -980
rect 40910 -1060 40950 -1000
rect 41010 -1060 41050 -1000
rect 40910 -1100 41050 -1060
rect 40910 -1160 40950 -1100
rect 41010 -1160 41050 -1100
rect 40910 -1200 41050 -1160
rect 40910 -1260 40950 -1200
rect 41010 -1260 41050 -1200
rect 40910 -1300 41050 -1260
rect 40910 -1360 40950 -1300
rect 41010 -1360 41050 -1300
rect 40910 -1380 41050 -1360
rect 41080 -1000 41220 -980
rect 41080 -1060 41120 -1000
rect 41180 -1060 41220 -1000
rect 41080 -1100 41220 -1060
rect 41080 -1160 41120 -1100
rect 41180 -1160 41220 -1100
rect 41080 -1200 41220 -1160
rect 41080 -1260 41120 -1200
rect 41180 -1260 41220 -1200
rect 41080 -1300 41220 -1260
rect 41080 -1360 41120 -1300
rect 41180 -1360 41220 -1300
rect 41080 -1380 41220 -1360
rect 41250 -1000 41390 -980
rect 41250 -1060 41290 -1000
rect 41350 -1060 41390 -1000
rect 41250 -1100 41390 -1060
rect 41250 -1160 41290 -1100
rect 41350 -1160 41390 -1100
rect 41250 -1200 41390 -1160
rect 41250 -1260 41290 -1200
rect 41350 -1260 41390 -1200
rect 41250 -1300 41390 -1260
rect 41250 -1360 41290 -1300
rect 41350 -1360 41390 -1300
rect 41250 -1380 41390 -1360
rect 41420 -1000 41560 -980
rect 41420 -1060 41460 -1000
rect 41520 -1060 41560 -1000
rect 41420 -1100 41560 -1060
rect 41420 -1160 41460 -1100
rect 41520 -1160 41560 -1100
rect 41420 -1200 41560 -1160
rect 41420 -1260 41460 -1200
rect 41520 -1260 41560 -1200
rect 41420 -1300 41560 -1260
rect 41420 -1360 41460 -1300
rect 41520 -1360 41560 -1300
rect 41420 -1380 41560 -1360
rect 41590 -1000 41730 -980
rect 41590 -1060 41630 -1000
rect 41690 -1060 41730 -1000
rect 41590 -1100 41730 -1060
rect 41590 -1160 41630 -1100
rect 41690 -1160 41730 -1100
rect 41590 -1200 41730 -1160
rect 41590 -1260 41630 -1200
rect 41690 -1260 41730 -1200
rect 41590 -1300 41730 -1260
rect 41590 -1360 41630 -1300
rect 41690 -1360 41730 -1300
rect 41590 -1380 41730 -1360
rect 41760 -1000 41900 -980
rect 41760 -1060 41800 -1000
rect 41860 -1060 41900 -1000
rect 41760 -1100 41900 -1060
rect 41760 -1160 41800 -1100
rect 41860 -1160 41900 -1100
rect 41760 -1200 41900 -1160
rect 41760 -1260 41800 -1200
rect 41860 -1260 41900 -1200
rect 41760 -1300 41900 -1260
rect 41760 -1360 41800 -1300
rect 41860 -1360 41900 -1300
rect 41760 -1380 41900 -1360
rect 41930 -1000 42070 -980
rect 41930 -1060 41970 -1000
rect 42030 -1060 42070 -1000
rect 41930 -1100 42070 -1060
rect 41930 -1160 41970 -1100
rect 42030 -1160 42070 -1100
rect 41930 -1200 42070 -1160
rect 41930 -1260 41970 -1200
rect 42030 -1260 42070 -1200
rect 41930 -1300 42070 -1260
rect 41930 -1360 41970 -1300
rect 42030 -1360 42070 -1300
rect 41930 -1380 42070 -1360
rect 42100 -1000 42240 -980
rect 42100 -1060 42140 -1000
rect 42200 -1060 42240 -1000
rect 42100 -1100 42240 -1060
rect 42100 -1160 42140 -1100
rect 42200 -1160 42240 -1100
rect 42100 -1200 42240 -1160
rect 42100 -1260 42140 -1200
rect 42200 -1260 42240 -1200
rect 42100 -1300 42240 -1260
rect 42100 -1360 42140 -1300
rect 42200 -1360 42240 -1300
rect 42100 -1380 42240 -1360
rect 42270 -1000 42410 -980
rect 42270 -1060 42310 -1000
rect 42370 -1060 42410 -1000
rect 42270 -1100 42410 -1060
rect 42270 -1160 42310 -1100
rect 42370 -1160 42410 -1100
rect 42270 -1200 42410 -1160
rect 42270 -1260 42310 -1200
rect 42370 -1260 42410 -1200
rect 42270 -1300 42410 -1260
rect 42270 -1360 42310 -1300
rect 42370 -1360 42410 -1300
rect 42270 -1380 42410 -1360
rect 42440 -1000 42580 -980
rect 42440 -1060 42480 -1000
rect 42540 -1060 42580 -1000
rect 42440 -1100 42580 -1060
rect 42440 -1160 42480 -1100
rect 42540 -1160 42580 -1100
rect 42440 -1200 42580 -1160
rect 42440 -1260 42480 -1200
rect 42540 -1260 42580 -1200
rect 42440 -1300 42580 -1260
rect 42440 -1360 42480 -1300
rect 42540 -1360 42580 -1300
rect 42440 -1380 42580 -1360
rect 42610 -1000 42750 -980
rect 42610 -1060 42650 -1000
rect 42710 -1060 42750 -1000
rect 42610 -1100 42750 -1060
rect 42610 -1160 42650 -1100
rect 42710 -1160 42750 -1100
rect 42610 -1200 42750 -1160
rect 42610 -1260 42650 -1200
rect 42710 -1260 42750 -1200
rect 42610 -1300 42750 -1260
rect 42610 -1360 42650 -1300
rect 42710 -1360 42750 -1300
rect 42610 -1380 42750 -1360
rect 42780 -1000 42920 -980
rect 42780 -1060 42820 -1000
rect 42880 -1060 42920 -1000
rect 42780 -1100 42920 -1060
rect 42780 -1160 42820 -1100
rect 42880 -1160 42920 -1100
rect 42780 -1200 42920 -1160
rect 42780 -1260 42820 -1200
rect 42880 -1260 42920 -1200
rect 42780 -1300 42920 -1260
rect 42780 -1360 42820 -1300
rect 42880 -1360 42920 -1300
rect 42780 -1380 42920 -1360
rect 42950 -1000 43090 -980
rect 42950 -1060 42990 -1000
rect 43050 -1060 43090 -1000
rect 42950 -1100 43090 -1060
rect 42950 -1160 42990 -1100
rect 43050 -1160 43090 -1100
rect 42950 -1200 43090 -1160
rect 42950 -1260 42990 -1200
rect 43050 -1260 43090 -1200
rect 42950 -1300 43090 -1260
rect 42950 -1360 42990 -1300
rect 43050 -1360 43090 -1300
rect 42950 -1380 43090 -1360
rect 43120 -1000 43260 -980
rect 43120 -1060 43160 -1000
rect 43220 -1060 43260 -1000
rect 43120 -1100 43260 -1060
rect 43120 -1160 43160 -1100
rect 43220 -1160 43260 -1100
rect 43120 -1200 43260 -1160
rect 43120 -1260 43160 -1200
rect 43220 -1260 43260 -1200
rect 43120 -1300 43260 -1260
rect 43120 -1360 43160 -1300
rect 43220 -1360 43260 -1300
rect 43120 -1380 43260 -1360
rect 43290 -1000 43430 -980
rect 43290 -1060 43330 -1000
rect 43390 -1060 43430 -1000
rect 43290 -1100 43430 -1060
rect 43290 -1160 43330 -1100
rect 43390 -1160 43430 -1100
rect 43290 -1200 43430 -1160
rect 43290 -1260 43330 -1200
rect 43390 -1260 43430 -1200
rect 43290 -1300 43430 -1260
rect 43290 -1360 43330 -1300
rect 43390 -1360 43430 -1300
rect 43290 -1380 43430 -1360
rect 43460 -1000 43600 -980
rect 43460 -1060 43500 -1000
rect 43560 -1060 43600 -1000
rect 43460 -1100 43600 -1060
rect 43460 -1160 43500 -1100
rect 43560 -1160 43600 -1100
rect 43460 -1200 43600 -1160
rect 43460 -1260 43500 -1200
rect 43560 -1260 43600 -1200
rect 43460 -1300 43600 -1260
rect 43460 -1360 43500 -1300
rect 43560 -1360 43600 -1300
rect 43460 -1380 43600 -1360
rect 43630 -1000 43770 -980
rect 43630 -1060 43670 -1000
rect 43730 -1060 43770 -1000
rect 43630 -1100 43770 -1060
rect 43630 -1160 43670 -1100
rect 43730 -1160 43770 -1100
rect 43630 -1200 43770 -1160
rect 43630 -1260 43670 -1200
rect 43730 -1260 43770 -1200
rect 43630 -1300 43770 -1260
rect 43630 -1360 43670 -1300
rect 43730 -1360 43770 -1300
rect 43630 -1380 43770 -1360
rect 43800 -1000 43940 -980
rect 43800 -1060 43840 -1000
rect 43900 -1060 43940 -1000
rect 43800 -1100 43940 -1060
rect 43800 -1160 43840 -1100
rect 43900 -1160 43940 -1100
rect 43800 -1200 43940 -1160
rect 43800 -1260 43840 -1200
rect 43900 -1260 43940 -1200
rect 43800 -1300 43940 -1260
rect 43800 -1360 43840 -1300
rect 43900 -1360 43940 -1300
rect 43800 -1380 43940 -1360
rect 43970 -1000 44110 -980
rect 43970 -1060 44010 -1000
rect 44070 -1060 44110 -1000
rect 43970 -1100 44110 -1060
rect 43970 -1160 44010 -1100
rect 44070 -1160 44110 -1100
rect 43970 -1200 44110 -1160
rect 43970 -1260 44010 -1200
rect 44070 -1260 44110 -1200
rect 43970 -1300 44110 -1260
rect 43970 -1360 44010 -1300
rect 44070 -1360 44110 -1300
rect 43970 -1380 44110 -1360
rect 44140 -1000 44280 -980
rect 44140 -1060 44180 -1000
rect 44240 -1060 44280 -1000
rect 44140 -1100 44280 -1060
rect 44140 -1160 44180 -1100
rect 44240 -1160 44280 -1100
rect 44140 -1200 44280 -1160
rect 44140 -1260 44180 -1200
rect 44240 -1260 44280 -1200
rect 44140 -1300 44280 -1260
rect 44140 -1360 44180 -1300
rect 44240 -1360 44280 -1300
rect 44140 -1380 44280 -1360
rect 44310 -1000 44450 -980
rect 44310 -1060 44350 -1000
rect 44410 -1060 44450 -1000
rect 44310 -1100 44450 -1060
rect 44310 -1160 44350 -1100
rect 44410 -1160 44450 -1100
rect 44310 -1200 44450 -1160
rect 44310 -1260 44350 -1200
rect 44410 -1260 44450 -1200
rect 44310 -1300 44450 -1260
rect 44310 -1360 44350 -1300
rect 44410 -1360 44450 -1300
rect 44310 -1380 44450 -1360
rect 44480 -1000 44620 -980
rect 44480 -1060 44520 -1000
rect 44580 -1060 44620 -1000
rect 44480 -1100 44620 -1060
rect 44480 -1160 44520 -1100
rect 44580 -1160 44620 -1100
rect 44480 -1200 44620 -1160
rect 44480 -1260 44520 -1200
rect 44580 -1260 44620 -1200
rect 44480 -1300 44620 -1260
rect 44480 -1360 44520 -1300
rect 44580 -1360 44620 -1300
rect 44480 -1380 44620 -1360
rect 44650 -1000 44790 -980
rect 44650 -1060 44690 -1000
rect 44750 -1060 44790 -1000
rect 44650 -1100 44790 -1060
rect 44650 -1160 44690 -1100
rect 44750 -1160 44790 -1100
rect 44650 -1200 44790 -1160
rect 44650 -1260 44690 -1200
rect 44750 -1260 44790 -1200
rect 44650 -1300 44790 -1260
rect 44650 -1360 44690 -1300
rect 44750 -1360 44790 -1300
rect 44650 -1380 44790 -1360
rect 44820 -1000 44960 -980
rect 44820 -1060 44860 -1000
rect 44920 -1060 44960 -1000
rect 44820 -1100 44960 -1060
rect 44820 -1160 44860 -1100
rect 44920 -1160 44960 -1100
rect 44820 -1200 44960 -1160
rect 44820 -1260 44860 -1200
rect 44920 -1260 44960 -1200
rect 44820 -1300 44960 -1260
rect 44820 -1360 44860 -1300
rect 44920 -1360 44960 -1300
rect 44820 -1380 44960 -1360
rect 44990 -1000 45130 -980
rect 44990 -1060 45030 -1000
rect 45090 -1060 45130 -1000
rect 44990 -1100 45130 -1060
rect 44990 -1160 45030 -1100
rect 45090 -1160 45130 -1100
rect 44990 -1200 45130 -1160
rect 44990 -1260 45030 -1200
rect 45090 -1260 45130 -1200
rect 44990 -1300 45130 -1260
rect 44990 -1360 45030 -1300
rect 45090 -1360 45130 -1300
rect 44990 -1380 45130 -1360
rect 45160 -1000 45300 -980
rect 45160 -1060 45200 -1000
rect 45260 -1060 45300 -1000
rect 45160 -1100 45300 -1060
rect 45160 -1160 45200 -1100
rect 45260 -1160 45300 -1100
rect 45160 -1200 45300 -1160
rect 45160 -1260 45200 -1200
rect 45260 -1260 45300 -1200
rect 45160 -1300 45300 -1260
rect 45160 -1360 45200 -1300
rect 45260 -1360 45300 -1300
rect 45160 -1380 45300 -1360
rect 45330 -1000 45470 -980
rect 45330 -1060 45370 -1000
rect 45430 -1060 45470 -1000
rect 45330 -1100 45470 -1060
rect 45330 -1160 45370 -1100
rect 45430 -1160 45470 -1100
rect 45330 -1200 45470 -1160
rect 45330 -1260 45370 -1200
rect 45430 -1260 45470 -1200
rect 45330 -1300 45470 -1260
rect 45330 -1360 45370 -1300
rect 45430 -1360 45470 -1300
rect 45330 -1380 45470 -1360
rect 45500 -1000 45640 -980
rect 45500 -1060 45540 -1000
rect 45600 -1060 45640 -1000
rect 45500 -1100 45640 -1060
rect 45500 -1160 45540 -1100
rect 45600 -1160 45640 -1100
rect 45500 -1200 45640 -1160
rect 45500 -1260 45540 -1200
rect 45600 -1260 45640 -1200
rect 45500 -1300 45640 -1260
rect 45500 -1360 45540 -1300
rect 45600 -1360 45640 -1300
rect 45500 -1380 45640 -1360
rect 45670 -1000 45810 -980
rect 45670 -1060 45710 -1000
rect 45770 -1060 45810 -1000
rect 45670 -1100 45810 -1060
rect 45670 -1160 45710 -1100
rect 45770 -1160 45810 -1100
rect 45670 -1200 45810 -1160
rect 45670 -1260 45710 -1200
rect 45770 -1260 45810 -1200
rect 45670 -1300 45810 -1260
rect 45670 -1360 45710 -1300
rect 45770 -1360 45810 -1300
rect 45670 -1380 45810 -1360
rect 45840 -1000 45980 -980
rect 45840 -1060 45880 -1000
rect 45940 -1060 45980 -1000
rect 45840 -1100 45980 -1060
rect 45840 -1160 45880 -1100
rect 45940 -1160 45980 -1100
rect 45840 -1200 45980 -1160
rect 45840 -1260 45880 -1200
rect 45940 -1260 45980 -1200
rect 45840 -1300 45980 -1260
rect 45840 -1360 45880 -1300
rect 45940 -1360 45980 -1300
rect 45840 -1380 45980 -1360
rect 46010 -1000 46150 -980
rect 46010 -1060 46050 -1000
rect 46110 -1060 46150 -1000
rect 46010 -1100 46150 -1060
rect 46010 -1160 46050 -1100
rect 46110 -1160 46150 -1100
rect 46010 -1200 46150 -1160
rect 46010 -1260 46050 -1200
rect 46110 -1260 46150 -1200
rect 46010 -1300 46150 -1260
rect 46010 -1360 46050 -1300
rect 46110 -1360 46150 -1300
rect 46010 -1380 46150 -1360
rect 46180 -1000 46320 -980
rect 46180 -1060 46220 -1000
rect 46280 -1060 46320 -1000
rect 46180 -1100 46320 -1060
rect 46180 -1160 46220 -1100
rect 46280 -1160 46320 -1100
rect 46180 -1200 46320 -1160
rect 46180 -1260 46220 -1200
rect 46280 -1260 46320 -1200
rect 46180 -1300 46320 -1260
rect 46180 -1360 46220 -1300
rect 46280 -1360 46320 -1300
rect 46180 -1380 46320 -1360
rect 46350 -1000 46490 -980
rect 46350 -1060 46390 -1000
rect 46450 -1060 46490 -1000
rect 46350 -1100 46490 -1060
rect 46350 -1160 46390 -1100
rect 46450 -1160 46490 -1100
rect 46350 -1200 46490 -1160
rect 46350 -1260 46390 -1200
rect 46450 -1260 46490 -1200
rect 46350 -1300 46490 -1260
rect 46350 -1360 46390 -1300
rect 46450 -1360 46490 -1300
rect 46350 -1380 46490 -1360
rect 46520 -1000 46660 -980
rect 46520 -1060 46560 -1000
rect 46620 -1060 46660 -1000
rect 46520 -1100 46660 -1060
rect 46520 -1160 46560 -1100
rect 46620 -1160 46660 -1100
rect 46520 -1200 46660 -1160
rect 46520 -1260 46560 -1200
rect 46620 -1260 46660 -1200
rect 46520 -1300 46660 -1260
rect 46520 -1360 46560 -1300
rect 46620 -1360 46660 -1300
rect 46520 -1380 46660 -1360
rect 46690 -1000 46830 -980
rect 46690 -1060 46730 -1000
rect 46790 -1060 46830 -1000
rect 46690 -1100 46830 -1060
rect 46690 -1160 46730 -1100
rect 46790 -1160 46830 -1100
rect 46690 -1200 46830 -1160
rect 46690 -1260 46730 -1200
rect 46790 -1260 46830 -1200
rect 46690 -1300 46830 -1260
rect 46690 -1360 46730 -1300
rect 46790 -1360 46830 -1300
rect 46690 -1380 46830 -1360
rect 46860 -1000 47000 -980
rect 46860 -1060 46900 -1000
rect 46960 -1060 47000 -1000
rect 46860 -1100 47000 -1060
rect 46860 -1160 46900 -1100
rect 46960 -1160 47000 -1100
rect 46860 -1200 47000 -1160
rect 46860 -1260 46900 -1200
rect 46960 -1260 47000 -1200
rect 46860 -1300 47000 -1260
rect 46860 -1360 46900 -1300
rect 46960 -1360 47000 -1300
rect 46860 -1380 47000 -1360
rect 47030 -1000 47170 -980
rect 47030 -1060 47070 -1000
rect 47130 -1060 47170 -1000
rect 47030 -1100 47170 -1060
rect 47030 -1160 47070 -1100
rect 47130 -1160 47170 -1100
rect 47030 -1200 47170 -1160
rect 47030 -1260 47070 -1200
rect 47130 -1260 47170 -1200
rect 47030 -1300 47170 -1260
rect 47030 -1360 47070 -1300
rect 47130 -1360 47170 -1300
rect 47030 -1380 47170 -1360
rect 47200 -1000 47340 -980
rect 47200 -1060 47240 -1000
rect 47300 -1060 47340 -1000
rect 47200 -1100 47340 -1060
rect 47200 -1160 47240 -1100
rect 47300 -1160 47340 -1100
rect 47200 -1200 47340 -1160
rect 47200 -1260 47240 -1200
rect 47300 -1260 47340 -1200
rect 47200 -1300 47340 -1260
rect 47200 -1360 47240 -1300
rect 47300 -1360 47340 -1300
rect 47200 -1380 47340 -1360
rect 47370 -1000 47510 -980
rect 47370 -1060 47410 -1000
rect 47470 -1060 47510 -1000
rect 47370 -1100 47510 -1060
rect 47370 -1160 47410 -1100
rect 47470 -1160 47510 -1100
rect 47370 -1200 47510 -1160
rect 47370 -1260 47410 -1200
rect 47470 -1260 47510 -1200
rect 47370 -1300 47510 -1260
rect 47370 -1360 47410 -1300
rect 47470 -1360 47510 -1300
rect 47370 -1380 47510 -1360
rect 47540 -1000 47680 -980
rect 47540 -1060 47580 -1000
rect 47640 -1060 47680 -1000
rect 47540 -1100 47680 -1060
rect 47540 -1160 47580 -1100
rect 47640 -1160 47680 -1100
rect 47540 -1200 47680 -1160
rect 47540 -1260 47580 -1200
rect 47640 -1260 47680 -1200
rect 47540 -1300 47680 -1260
rect 47540 -1360 47580 -1300
rect 47640 -1360 47680 -1300
rect 47540 -1380 47680 -1360
rect 47710 -1000 47850 -980
rect 47710 -1060 47750 -1000
rect 47810 -1060 47850 -1000
rect 47710 -1100 47850 -1060
rect 47710 -1160 47750 -1100
rect 47810 -1160 47850 -1100
rect 47710 -1200 47850 -1160
rect 47710 -1260 47750 -1200
rect 47810 -1260 47850 -1200
rect 47710 -1300 47850 -1260
rect 47710 -1360 47750 -1300
rect 47810 -1360 47850 -1300
rect 47710 -1380 47850 -1360
rect 47880 -1000 48020 -980
rect 47880 -1060 47920 -1000
rect 47980 -1060 48020 -1000
rect 47880 -1100 48020 -1060
rect 47880 -1160 47920 -1100
rect 47980 -1160 48020 -1100
rect 47880 -1200 48020 -1160
rect 47880 -1260 47920 -1200
rect 47980 -1260 48020 -1200
rect 47880 -1300 48020 -1260
rect 47880 -1360 47920 -1300
rect 47980 -1360 48020 -1300
rect 47880 -1380 48020 -1360
rect 48050 -1000 48190 -980
rect 48050 -1060 48090 -1000
rect 48150 -1060 48190 -1000
rect 48050 -1100 48190 -1060
rect 48050 -1160 48090 -1100
rect 48150 -1160 48190 -1100
rect 48050 -1200 48190 -1160
rect 48050 -1260 48090 -1200
rect 48150 -1260 48190 -1200
rect 48050 -1300 48190 -1260
rect 48050 -1360 48090 -1300
rect 48150 -1360 48190 -1300
rect 48050 -1380 48190 -1360
rect 48220 -1000 48360 -980
rect 48220 -1060 48260 -1000
rect 48320 -1060 48360 -1000
rect 48220 -1100 48360 -1060
rect 48220 -1160 48260 -1100
rect 48320 -1160 48360 -1100
rect 48220 -1200 48360 -1160
rect 48220 -1260 48260 -1200
rect 48320 -1260 48360 -1200
rect 48220 -1300 48360 -1260
rect 48220 -1360 48260 -1300
rect 48320 -1360 48360 -1300
rect 48220 -1380 48360 -1360
rect 48390 -1000 48530 -980
rect 48390 -1060 48430 -1000
rect 48490 -1060 48530 -1000
rect 48390 -1100 48530 -1060
rect 48390 -1160 48430 -1100
rect 48490 -1160 48530 -1100
rect 48390 -1200 48530 -1160
rect 48390 -1260 48430 -1200
rect 48490 -1260 48530 -1200
rect 48390 -1300 48530 -1260
rect 48390 -1360 48430 -1300
rect 48490 -1360 48530 -1300
rect 48390 -1380 48530 -1360
rect 48560 -1000 48700 -980
rect 48560 -1060 48600 -1000
rect 48660 -1060 48700 -1000
rect 48560 -1100 48700 -1060
rect 48560 -1160 48600 -1100
rect 48660 -1160 48700 -1100
rect 48560 -1200 48700 -1160
rect 48560 -1260 48600 -1200
rect 48660 -1260 48700 -1200
rect 48560 -1300 48700 -1260
rect 48560 -1360 48600 -1300
rect 48660 -1360 48700 -1300
rect 48560 -1380 48700 -1360
rect 48730 -1000 48870 -980
rect 48730 -1060 48770 -1000
rect 48830 -1060 48870 -1000
rect 48730 -1100 48870 -1060
rect 48730 -1160 48770 -1100
rect 48830 -1160 48870 -1100
rect 48730 -1200 48870 -1160
rect 48730 -1260 48770 -1200
rect 48830 -1260 48870 -1200
rect 48730 -1300 48870 -1260
rect 48730 -1360 48770 -1300
rect 48830 -1360 48870 -1300
rect 48730 -1380 48870 -1360
rect 48900 -1000 49040 -980
rect 48900 -1060 48940 -1000
rect 49000 -1060 49040 -1000
rect 48900 -1100 49040 -1060
rect 48900 -1160 48940 -1100
rect 49000 -1160 49040 -1100
rect 48900 -1200 49040 -1160
rect 48900 -1260 48940 -1200
rect 49000 -1260 49040 -1200
rect 48900 -1300 49040 -1260
rect 48900 -1360 48940 -1300
rect 49000 -1360 49040 -1300
rect 48900 -1380 49040 -1360
rect 49070 -1000 49210 -980
rect 49070 -1060 49110 -1000
rect 49170 -1060 49210 -1000
rect 49070 -1100 49210 -1060
rect 49070 -1160 49110 -1100
rect 49170 -1160 49210 -1100
rect 49070 -1200 49210 -1160
rect 49070 -1260 49110 -1200
rect 49170 -1260 49210 -1200
rect 49070 -1300 49210 -1260
rect 49070 -1360 49110 -1300
rect 49170 -1360 49210 -1300
rect 49070 -1380 49210 -1360
rect 49240 -1000 49380 -980
rect 49240 -1060 49280 -1000
rect 49340 -1060 49380 -1000
rect 49240 -1100 49380 -1060
rect 49240 -1160 49280 -1100
rect 49340 -1160 49380 -1100
rect 49240 -1200 49380 -1160
rect 49240 -1260 49280 -1200
rect 49340 -1260 49380 -1200
rect 49240 -1300 49380 -1260
rect 49240 -1360 49280 -1300
rect 49340 -1360 49380 -1300
rect 49240 -1380 49380 -1360
rect 49410 -1000 49550 -980
rect 49410 -1060 49450 -1000
rect 49510 -1060 49550 -1000
rect 49410 -1100 49550 -1060
rect 49410 -1160 49450 -1100
rect 49510 -1160 49550 -1100
rect 49410 -1200 49550 -1160
rect 49410 -1260 49450 -1200
rect 49510 -1260 49550 -1200
rect 49410 -1300 49550 -1260
rect 49410 -1360 49450 -1300
rect 49510 -1360 49550 -1300
rect 49410 -1380 49550 -1360
rect 49580 -1000 49720 -980
rect 49580 -1060 49620 -1000
rect 49680 -1060 49720 -1000
rect 49580 -1100 49720 -1060
rect 49580 -1160 49620 -1100
rect 49680 -1160 49720 -1100
rect 49580 -1200 49720 -1160
rect 49580 -1260 49620 -1200
rect 49680 -1260 49720 -1200
rect 49580 -1300 49720 -1260
rect 49580 -1360 49620 -1300
rect 49680 -1360 49720 -1300
rect 49580 -1380 49720 -1360
rect 49750 -1000 49890 -980
rect 49750 -1060 49790 -1000
rect 49850 -1060 49890 -1000
rect 49750 -1100 49890 -1060
rect 49750 -1160 49790 -1100
rect 49850 -1160 49890 -1100
rect 49750 -1200 49890 -1160
rect 49750 -1260 49790 -1200
rect 49850 -1260 49890 -1200
rect 49750 -1300 49890 -1260
rect 49750 -1360 49790 -1300
rect 49850 -1360 49890 -1300
rect 49750 -1380 49890 -1360
rect 49920 -1000 50060 -980
rect 49920 -1060 49960 -1000
rect 50020 -1060 50060 -1000
rect 49920 -1100 50060 -1060
rect 49920 -1160 49960 -1100
rect 50020 -1160 50060 -1100
rect 49920 -1200 50060 -1160
rect 49920 -1260 49960 -1200
rect 50020 -1260 50060 -1200
rect 49920 -1300 50060 -1260
rect 49920 -1360 49960 -1300
rect 50020 -1360 50060 -1300
rect 49920 -1380 50060 -1360
rect 50090 -1000 50230 -980
rect 50090 -1060 50130 -1000
rect 50190 -1060 50230 -1000
rect 50090 -1100 50230 -1060
rect 50090 -1160 50130 -1100
rect 50190 -1160 50230 -1100
rect 50090 -1200 50230 -1160
rect 50090 -1260 50130 -1200
rect 50190 -1260 50230 -1200
rect 50090 -1300 50230 -1260
rect 50090 -1360 50130 -1300
rect 50190 -1360 50230 -1300
rect 50090 -1380 50230 -1360
rect 50260 -1000 50400 -980
rect 50260 -1060 50300 -1000
rect 50360 -1060 50400 -1000
rect 50260 -1100 50400 -1060
rect 50260 -1160 50300 -1100
rect 50360 -1160 50400 -1100
rect 50260 -1200 50400 -1160
rect 50260 -1260 50300 -1200
rect 50360 -1260 50400 -1200
rect 50260 -1300 50400 -1260
rect 50260 -1360 50300 -1300
rect 50360 -1360 50400 -1300
rect 50260 -1380 50400 -1360
rect 50430 -1000 50570 -980
rect 50430 -1060 50470 -1000
rect 50530 -1060 50570 -1000
rect 50430 -1100 50570 -1060
rect 50430 -1160 50470 -1100
rect 50530 -1160 50570 -1100
rect 50430 -1200 50570 -1160
rect 50430 -1260 50470 -1200
rect 50530 -1260 50570 -1200
rect 50430 -1300 50570 -1260
rect 50430 -1360 50470 -1300
rect 50530 -1360 50570 -1300
rect 50430 -1380 50570 -1360
rect 50600 -1000 50740 -980
rect 50600 -1060 50640 -1000
rect 50700 -1060 50740 -1000
rect 50600 -1100 50740 -1060
rect 50600 -1160 50640 -1100
rect 50700 -1160 50740 -1100
rect 50600 -1200 50740 -1160
rect 50600 -1260 50640 -1200
rect 50700 -1260 50740 -1200
rect 50600 -1300 50740 -1260
rect 50600 -1360 50640 -1300
rect 50700 -1360 50740 -1300
rect 50600 -1380 50740 -1360
rect 50770 -1000 50910 -980
rect 50770 -1060 50810 -1000
rect 50870 -1060 50910 -1000
rect 50770 -1100 50910 -1060
rect 50770 -1160 50810 -1100
rect 50870 -1160 50910 -1100
rect 50770 -1200 50910 -1160
rect 50770 -1260 50810 -1200
rect 50870 -1260 50910 -1200
rect 50770 -1300 50910 -1260
rect 50770 -1360 50810 -1300
rect 50870 -1360 50910 -1300
rect 50770 -1380 50910 -1360
rect 50940 -1000 51080 -980
rect 50940 -1060 50980 -1000
rect 51040 -1060 51080 -1000
rect 50940 -1100 51080 -1060
rect 50940 -1160 50980 -1100
rect 51040 -1160 51080 -1100
rect 50940 -1200 51080 -1160
rect 50940 -1260 50980 -1200
rect 51040 -1260 51080 -1200
rect 50940 -1300 51080 -1260
rect 50940 -1360 50980 -1300
rect 51040 -1360 51080 -1300
rect 50940 -1380 51080 -1360
rect 51110 -1000 51250 -980
rect 51110 -1060 51150 -1000
rect 51210 -1060 51250 -1000
rect 51110 -1100 51250 -1060
rect 51110 -1160 51150 -1100
rect 51210 -1160 51250 -1100
rect 51110 -1200 51250 -1160
rect 51110 -1260 51150 -1200
rect 51210 -1260 51250 -1200
rect 51110 -1300 51250 -1260
rect 51110 -1360 51150 -1300
rect 51210 -1360 51250 -1300
rect 51110 -1380 51250 -1360
rect 51280 -1000 51420 -980
rect 51280 -1060 51320 -1000
rect 51380 -1060 51420 -1000
rect 51280 -1100 51420 -1060
rect 51280 -1160 51320 -1100
rect 51380 -1160 51420 -1100
rect 51280 -1200 51420 -1160
rect 51280 -1260 51320 -1200
rect 51380 -1260 51420 -1200
rect 51280 -1300 51420 -1260
rect 51280 -1360 51320 -1300
rect 51380 -1360 51420 -1300
rect 51280 -1380 51420 -1360
rect 51450 -1000 51590 -980
rect 51450 -1060 51490 -1000
rect 51550 -1060 51590 -1000
rect 51450 -1100 51590 -1060
rect 51450 -1160 51490 -1100
rect 51550 -1160 51590 -1100
rect 51450 -1200 51590 -1160
rect 51450 -1260 51490 -1200
rect 51550 -1260 51590 -1200
rect 51450 -1300 51590 -1260
rect 51450 -1360 51490 -1300
rect 51550 -1360 51590 -1300
rect 51450 -1380 51590 -1360
rect 51620 -1000 51760 -980
rect 51620 -1060 51660 -1000
rect 51720 -1060 51760 -1000
rect 51620 -1100 51760 -1060
rect 51620 -1160 51660 -1100
rect 51720 -1160 51760 -1100
rect 51620 -1200 51760 -1160
rect 51620 -1260 51660 -1200
rect 51720 -1260 51760 -1200
rect 51620 -1300 51760 -1260
rect 51620 -1360 51660 -1300
rect 51720 -1360 51760 -1300
rect 51620 -1380 51760 -1360
rect 51790 -1000 51930 -980
rect 51790 -1060 51830 -1000
rect 51890 -1060 51930 -1000
rect 51790 -1100 51930 -1060
rect 51790 -1160 51830 -1100
rect 51890 -1160 51930 -1100
rect 51790 -1200 51930 -1160
rect 51790 -1260 51830 -1200
rect 51890 -1260 51930 -1200
rect 51790 -1300 51930 -1260
rect 51790 -1360 51830 -1300
rect 51890 -1360 51930 -1300
rect 51790 -1380 51930 -1360
rect 51960 -1000 52100 -980
rect 51960 -1060 52000 -1000
rect 52060 -1060 52100 -1000
rect 51960 -1100 52100 -1060
rect 51960 -1160 52000 -1100
rect 52060 -1160 52100 -1100
rect 51960 -1200 52100 -1160
rect 51960 -1260 52000 -1200
rect 52060 -1260 52100 -1200
rect 51960 -1300 52100 -1260
rect 51960 -1360 52000 -1300
rect 52060 -1360 52100 -1300
rect 51960 -1380 52100 -1360
rect 52130 -1000 52270 -980
rect 52130 -1060 52170 -1000
rect 52230 -1060 52270 -1000
rect 52130 -1100 52270 -1060
rect 52130 -1160 52170 -1100
rect 52230 -1160 52270 -1100
rect 52130 -1200 52270 -1160
rect 52130 -1260 52170 -1200
rect 52230 -1260 52270 -1200
rect 52130 -1300 52270 -1260
rect 52130 -1360 52170 -1300
rect 52230 -1360 52270 -1300
rect 52130 -1380 52270 -1360
rect 52300 -1000 52440 -980
rect 52300 -1060 52340 -1000
rect 52400 -1060 52440 -1000
rect 52300 -1100 52440 -1060
rect 52300 -1160 52340 -1100
rect 52400 -1160 52440 -1100
rect 52300 -1200 52440 -1160
rect 52300 -1260 52340 -1200
rect 52400 -1260 52440 -1200
rect 52300 -1300 52440 -1260
rect 52300 -1360 52340 -1300
rect 52400 -1360 52440 -1300
rect 52300 -1380 52440 -1360
rect 52470 -1000 52610 -980
rect 52470 -1060 52510 -1000
rect 52570 -1060 52610 -1000
rect 52470 -1100 52610 -1060
rect 52470 -1160 52510 -1100
rect 52570 -1160 52610 -1100
rect 52470 -1200 52610 -1160
rect 52470 -1260 52510 -1200
rect 52570 -1260 52610 -1200
rect 52470 -1300 52610 -1260
rect 52470 -1360 52510 -1300
rect 52570 -1360 52610 -1300
rect 52470 -1380 52610 -1360
rect 52640 -1000 52780 -980
rect 52640 -1060 52680 -1000
rect 52740 -1060 52780 -1000
rect 52640 -1100 52780 -1060
rect 52640 -1160 52680 -1100
rect 52740 -1160 52780 -1100
rect 52640 -1200 52780 -1160
rect 52640 -1260 52680 -1200
rect 52740 -1260 52780 -1200
rect 52640 -1300 52780 -1260
rect 52640 -1360 52680 -1300
rect 52740 -1360 52780 -1300
rect 52640 -1380 52780 -1360
rect 52810 -1000 52950 -980
rect 52810 -1060 52850 -1000
rect 52910 -1060 52950 -1000
rect 52810 -1100 52950 -1060
rect 52810 -1160 52850 -1100
rect 52910 -1160 52950 -1100
rect 52810 -1200 52950 -1160
rect 52810 -1260 52850 -1200
rect 52910 -1260 52950 -1200
rect 52810 -1300 52950 -1260
rect 52810 -1360 52850 -1300
rect 52910 -1360 52950 -1300
rect 52810 -1380 52950 -1360
rect 52980 -1000 53120 -980
rect 52980 -1060 53020 -1000
rect 53080 -1060 53120 -1000
rect 52980 -1100 53120 -1060
rect 52980 -1160 53020 -1100
rect 53080 -1160 53120 -1100
rect 52980 -1200 53120 -1160
rect 52980 -1260 53020 -1200
rect 53080 -1260 53120 -1200
rect 52980 -1300 53120 -1260
rect 52980 -1360 53020 -1300
rect 53080 -1360 53120 -1300
rect 52980 -1380 53120 -1360
rect 53150 -1000 53290 -980
rect 53150 -1060 53190 -1000
rect 53250 -1060 53290 -1000
rect 53150 -1100 53290 -1060
rect 53150 -1160 53190 -1100
rect 53250 -1160 53290 -1100
rect 53150 -1200 53290 -1160
rect 53150 -1260 53190 -1200
rect 53250 -1260 53290 -1200
rect 53150 -1300 53290 -1260
rect 53150 -1360 53190 -1300
rect 53250 -1360 53290 -1300
rect 53150 -1380 53290 -1360
rect 53320 -1000 53460 -980
rect 53320 -1060 53360 -1000
rect 53420 -1060 53460 -1000
rect 53320 -1100 53460 -1060
rect 53320 -1160 53360 -1100
rect 53420 -1160 53460 -1100
rect 53320 -1200 53460 -1160
rect 53320 -1260 53360 -1200
rect 53420 -1260 53460 -1200
rect 53320 -1300 53460 -1260
rect 53320 -1360 53360 -1300
rect 53420 -1360 53460 -1300
rect 53320 -1380 53460 -1360
rect 53490 -1000 53630 -980
rect 53490 -1060 53530 -1000
rect 53590 -1060 53630 -1000
rect 53490 -1100 53630 -1060
rect 53490 -1160 53530 -1100
rect 53590 -1160 53630 -1100
rect 53490 -1200 53630 -1160
rect 53490 -1260 53530 -1200
rect 53590 -1260 53630 -1200
rect 53490 -1300 53630 -1260
rect 53490 -1360 53530 -1300
rect 53590 -1360 53630 -1300
rect 53490 -1380 53630 -1360
rect 53660 -1000 53800 -980
rect 53660 -1060 53700 -1000
rect 53760 -1060 53800 -1000
rect 53660 -1100 53800 -1060
rect 53660 -1160 53700 -1100
rect 53760 -1160 53800 -1100
rect 53660 -1200 53800 -1160
rect 53660 -1260 53700 -1200
rect 53760 -1260 53800 -1200
rect 53660 -1300 53800 -1260
rect 53660 -1360 53700 -1300
rect 53760 -1360 53800 -1300
rect 53660 -1380 53800 -1360
rect 53830 -1000 53970 -980
rect 53830 -1060 53870 -1000
rect 53930 -1060 53970 -1000
rect 53830 -1100 53970 -1060
rect 53830 -1160 53870 -1100
rect 53930 -1160 53970 -1100
rect 53830 -1200 53970 -1160
rect 53830 -1260 53870 -1200
rect 53930 -1260 53970 -1200
rect 53830 -1300 53970 -1260
rect 53830 -1360 53870 -1300
rect 53930 -1360 53970 -1300
rect 53830 -1380 53970 -1360
rect 54000 -1000 54140 -980
rect 54000 -1060 54040 -1000
rect 54100 -1060 54140 -1000
rect 54000 -1100 54140 -1060
rect 54000 -1160 54040 -1100
rect 54100 -1160 54140 -1100
rect 54000 -1200 54140 -1160
rect 54000 -1260 54040 -1200
rect 54100 -1260 54140 -1200
rect 54000 -1300 54140 -1260
rect 54000 -1360 54040 -1300
rect 54100 -1360 54140 -1300
rect 54000 -1380 54140 -1360
rect 54170 -1000 54310 -980
rect 54170 -1060 54210 -1000
rect 54270 -1060 54310 -1000
rect 54170 -1100 54310 -1060
rect 54170 -1160 54210 -1100
rect 54270 -1160 54310 -1100
rect 54170 -1200 54310 -1160
rect 54170 -1260 54210 -1200
rect 54270 -1260 54310 -1200
rect 54170 -1300 54310 -1260
rect 54170 -1360 54210 -1300
rect 54270 -1360 54310 -1300
rect 54170 -1380 54310 -1360
rect 54340 -1000 54480 -980
rect 54340 -1060 54380 -1000
rect 54440 -1060 54480 -1000
rect 54340 -1100 54480 -1060
rect 54340 -1160 54380 -1100
rect 54440 -1160 54480 -1100
rect 54340 -1200 54480 -1160
rect 54340 -1260 54380 -1200
rect 54440 -1260 54480 -1200
rect 54340 -1300 54480 -1260
rect 54340 -1360 54380 -1300
rect 54440 -1360 54480 -1300
rect 54340 -1380 54480 -1360
rect 54510 -1000 54650 -980
rect 54510 -1060 54550 -1000
rect 54610 -1060 54650 -1000
rect 54510 -1100 54650 -1060
rect 54510 -1160 54550 -1100
rect 54610 -1160 54650 -1100
rect 54510 -1200 54650 -1160
rect 54510 -1260 54550 -1200
rect 54610 -1260 54650 -1200
rect 54510 -1300 54650 -1260
rect 54510 -1360 54550 -1300
rect 54610 -1360 54650 -1300
rect 54510 -1380 54650 -1360
rect 54680 -1000 54820 -980
rect 54680 -1060 54720 -1000
rect 54780 -1060 54820 -1000
rect 54680 -1100 54820 -1060
rect 54680 -1160 54720 -1100
rect 54780 -1160 54820 -1100
rect 54680 -1200 54820 -1160
rect 54680 -1260 54720 -1200
rect 54780 -1260 54820 -1200
rect 54680 -1300 54820 -1260
rect 54680 -1360 54720 -1300
rect 54780 -1360 54820 -1300
rect 54680 -1380 54820 -1360
rect 54850 -1000 54990 -980
rect 54850 -1060 54890 -1000
rect 54950 -1060 54990 -1000
rect 54850 -1100 54990 -1060
rect 54850 -1160 54890 -1100
rect 54950 -1160 54990 -1100
rect 54850 -1200 54990 -1160
rect 54850 -1260 54890 -1200
rect 54950 -1260 54990 -1200
rect 54850 -1300 54990 -1260
rect 54850 -1360 54890 -1300
rect 54950 -1360 54990 -1300
rect 54850 -1380 54990 -1360
rect 55020 -1000 55160 -980
rect 55020 -1060 55060 -1000
rect 55120 -1060 55160 -1000
rect 55020 -1100 55160 -1060
rect 55020 -1160 55060 -1100
rect 55120 -1160 55160 -1100
rect 55020 -1200 55160 -1160
rect 55020 -1260 55060 -1200
rect 55120 -1260 55160 -1200
rect 55020 -1300 55160 -1260
rect 55020 -1360 55060 -1300
rect 55120 -1360 55160 -1300
rect 55020 -1380 55160 -1360
rect 55190 -1000 55330 -980
rect 55190 -1060 55230 -1000
rect 55290 -1060 55330 -1000
rect 55190 -1100 55330 -1060
rect 55190 -1160 55230 -1100
rect 55290 -1160 55330 -1100
rect 55190 -1200 55330 -1160
rect 55190 -1260 55230 -1200
rect 55290 -1260 55330 -1200
rect 55190 -1300 55330 -1260
rect 55190 -1360 55230 -1300
rect 55290 -1360 55330 -1300
rect 55190 -1380 55330 -1360
rect 55360 -1000 55500 -980
rect 55360 -1060 55400 -1000
rect 55460 -1060 55500 -1000
rect 55360 -1100 55500 -1060
rect 55360 -1160 55400 -1100
rect 55460 -1160 55500 -1100
rect 55360 -1200 55500 -1160
rect 55360 -1260 55400 -1200
rect 55460 -1260 55500 -1200
rect 55360 -1300 55500 -1260
rect 55360 -1360 55400 -1300
rect 55460 -1360 55500 -1300
rect 55360 -1380 55500 -1360
rect 55530 -1000 55670 -980
rect 55530 -1060 55570 -1000
rect 55630 -1060 55670 -1000
rect 55530 -1100 55670 -1060
rect 55530 -1160 55570 -1100
rect 55630 -1160 55670 -1100
rect 55530 -1200 55670 -1160
rect 55530 -1260 55570 -1200
rect 55630 -1260 55670 -1200
rect 55530 -1300 55670 -1260
rect 55530 -1360 55570 -1300
rect 55630 -1360 55670 -1300
rect 55530 -1380 55670 -1360
rect 55700 -1000 55840 -980
rect 55700 -1060 55740 -1000
rect 55800 -1060 55840 -1000
rect 55700 -1100 55840 -1060
rect 55700 -1160 55740 -1100
rect 55800 -1160 55840 -1100
rect 55700 -1200 55840 -1160
rect 55700 -1260 55740 -1200
rect 55800 -1260 55840 -1200
rect 55700 -1300 55840 -1260
rect 55700 -1360 55740 -1300
rect 55800 -1360 55840 -1300
rect 55700 -1380 55840 -1360
rect 55870 -1000 56010 -980
rect 55870 -1060 55910 -1000
rect 55970 -1060 56010 -1000
rect 55870 -1100 56010 -1060
rect 55870 -1160 55910 -1100
rect 55970 -1160 56010 -1100
rect 55870 -1200 56010 -1160
rect 55870 -1260 55910 -1200
rect 55970 -1260 56010 -1200
rect 55870 -1300 56010 -1260
rect 55870 -1360 55910 -1300
rect 55970 -1360 56010 -1300
rect 55870 -1380 56010 -1360
rect 56040 -1000 56180 -980
rect 56040 -1060 56080 -1000
rect 56140 -1060 56180 -1000
rect 56040 -1100 56180 -1060
rect 56040 -1160 56080 -1100
rect 56140 -1160 56180 -1100
rect 56040 -1200 56180 -1160
rect 56040 -1260 56080 -1200
rect 56140 -1260 56180 -1200
rect 56040 -1300 56180 -1260
rect 56040 -1360 56080 -1300
rect 56140 -1360 56180 -1300
rect 56040 -1380 56180 -1360
rect 56210 -1000 56350 -980
rect 56210 -1060 56250 -1000
rect 56310 -1060 56350 -1000
rect 56210 -1100 56350 -1060
rect 56210 -1160 56250 -1100
rect 56310 -1160 56350 -1100
rect 56210 -1200 56350 -1160
rect 56210 -1260 56250 -1200
rect 56310 -1260 56350 -1200
rect 56210 -1300 56350 -1260
rect 56210 -1360 56250 -1300
rect 56310 -1360 56350 -1300
rect 56210 -1380 56350 -1360
rect 56380 -1000 56520 -980
rect 56380 -1060 56420 -1000
rect 56480 -1060 56520 -1000
rect 56380 -1100 56520 -1060
rect 56380 -1160 56420 -1100
rect 56480 -1160 56520 -1100
rect 56380 -1200 56520 -1160
rect 56380 -1260 56420 -1200
rect 56480 -1260 56520 -1200
rect 56380 -1300 56520 -1260
rect 56380 -1360 56420 -1300
rect 56480 -1360 56520 -1300
rect 56380 -1380 56520 -1360
rect 56550 -1000 56690 -980
rect 56550 -1060 56590 -1000
rect 56650 -1060 56690 -1000
rect 56550 -1100 56690 -1060
rect 56550 -1160 56590 -1100
rect 56650 -1160 56690 -1100
rect 56550 -1200 56690 -1160
rect 56550 -1260 56590 -1200
rect 56650 -1260 56690 -1200
rect 56550 -1300 56690 -1260
rect 56550 -1360 56590 -1300
rect 56650 -1360 56690 -1300
rect 56550 -1380 56690 -1360
rect 56720 -1000 56860 -980
rect 56720 -1060 56760 -1000
rect 56820 -1060 56860 -1000
rect 56720 -1100 56860 -1060
rect 56720 -1160 56760 -1100
rect 56820 -1160 56860 -1100
rect 56720 -1200 56860 -1160
rect 56720 -1260 56760 -1200
rect 56820 -1260 56860 -1200
rect 56720 -1300 56860 -1260
rect 56720 -1360 56760 -1300
rect 56820 -1360 56860 -1300
rect 56720 -1380 56860 -1360
rect 56890 -1000 57030 -980
rect 56890 -1060 56930 -1000
rect 56990 -1060 57030 -1000
rect 56890 -1100 57030 -1060
rect 56890 -1160 56930 -1100
rect 56990 -1160 57030 -1100
rect 56890 -1200 57030 -1160
rect 56890 -1260 56930 -1200
rect 56990 -1260 57030 -1200
rect 56890 -1300 57030 -1260
rect 56890 -1360 56930 -1300
rect 56990 -1360 57030 -1300
rect 56890 -1380 57030 -1360
rect 57060 -1000 57200 -980
rect 57060 -1060 57100 -1000
rect 57160 -1060 57200 -1000
rect 57060 -1100 57200 -1060
rect 57060 -1160 57100 -1100
rect 57160 -1160 57200 -1100
rect 57060 -1200 57200 -1160
rect 57060 -1260 57100 -1200
rect 57160 -1260 57200 -1200
rect 57060 -1300 57200 -1260
rect 57060 -1360 57100 -1300
rect 57160 -1360 57200 -1300
rect 57060 -1380 57200 -1360
rect 57230 -1000 57370 -980
rect 57230 -1060 57270 -1000
rect 57330 -1060 57370 -1000
rect 57230 -1100 57370 -1060
rect 57230 -1160 57270 -1100
rect 57330 -1160 57370 -1100
rect 57230 -1200 57370 -1160
rect 57230 -1260 57270 -1200
rect 57330 -1260 57370 -1200
rect 57230 -1300 57370 -1260
rect 57230 -1360 57270 -1300
rect 57330 -1360 57370 -1300
rect 57230 -1380 57370 -1360
rect 57400 -1000 57540 -980
rect 57400 -1060 57440 -1000
rect 57500 -1060 57540 -1000
rect 57400 -1100 57540 -1060
rect 57400 -1160 57440 -1100
rect 57500 -1160 57540 -1100
rect 57400 -1200 57540 -1160
rect 57400 -1260 57440 -1200
rect 57500 -1260 57540 -1200
rect 57400 -1300 57540 -1260
rect 57400 -1360 57440 -1300
rect 57500 -1360 57540 -1300
rect 57400 -1380 57540 -1360
rect 57570 -1000 57710 -980
rect 57570 -1060 57610 -1000
rect 57670 -1060 57710 -1000
rect 57570 -1100 57710 -1060
rect 57570 -1160 57610 -1100
rect 57670 -1160 57710 -1100
rect 57570 -1200 57710 -1160
rect 57570 -1260 57610 -1200
rect 57670 -1260 57710 -1200
rect 57570 -1300 57710 -1260
rect 57570 -1360 57610 -1300
rect 57670 -1360 57710 -1300
rect 57570 -1380 57710 -1360
rect 57740 -1000 57880 -980
rect 57740 -1060 57780 -1000
rect 57840 -1060 57880 -1000
rect 57740 -1100 57880 -1060
rect 57740 -1160 57780 -1100
rect 57840 -1160 57880 -1100
rect 57740 -1200 57880 -1160
rect 57740 -1260 57780 -1200
rect 57840 -1260 57880 -1200
rect 57740 -1300 57880 -1260
rect 57740 -1360 57780 -1300
rect 57840 -1360 57880 -1300
rect 57740 -1380 57880 -1360
rect 57910 -1000 58050 -980
rect 57910 -1060 57950 -1000
rect 58010 -1060 58050 -1000
rect 57910 -1100 58050 -1060
rect 57910 -1160 57950 -1100
rect 58010 -1160 58050 -1100
rect 57910 -1200 58050 -1160
rect 57910 -1260 57950 -1200
rect 58010 -1260 58050 -1200
rect 57910 -1300 58050 -1260
rect 57910 -1360 57950 -1300
rect 58010 -1360 58050 -1300
rect 57910 -1380 58050 -1360
rect 58080 -1000 58220 -980
rect 58080 -1060 58120 -1000
rect 58180 -1060 58220 -1000
rect 58080 -1100 58220 -1060
rect 58080 -1160 58120 -1100
rect 58180 -1160 58220 -1100
rect 58080 -1200 58220 -1160
rect 58080 -1260 58120 -1200
rect 58180 -1260 58220 -1200
rect 58080 -1300 58220 -1260
rect 58080 -1360 58120 -1300
rect 58180 -1360 58220 -1300
rect 58080 -1380 58220 -1360
rect 58250 -1000 58390 -980
rect 58250 -1060 58290 -1000
rect 58350 -1060 58390 -1000
rect 58250 -1100 58390 -1060
rect 58250 -1160 58290 -1100
rect 58350 -1160 58390 -1100
rect 58250 -1200 58390 -1160
rect 58250 -1260 58290 -1200
rect 58350 -1260 58390 -1200
rect 58250 -1300 58390 -1260
rect 58250 -1360 58290 -1300
rect 58350 -1360 58390 -1300
rect 58250 -1380 58390 -1360
rect 58420 -1000 58560 -980
rect 58420 -1060 58460 -1000
rect 58520 -1060 58560 -1000
rect 58420 -1100 58560 -1060
rect 58420 -1160 58460 -1100
rect 58520 -1160 58560 -1100
rect 58420 -1200 58560 -1160
rect 58420 -1260 58460 -1200
rect 58520 -1260 58560 -1200
rect 58420 -1300 58560 -1260
rect 58420 -1360 58460 -1300
rect 58520 -1360 58560 -1300
rect 58420 -1380 58560 -1360
rect 58590 -1000 58730 -980
rect 58590 -1060 58630 -1000
rect 58690 -1060 58730 -1000
rect 58590 -1100 58730 -1060
rect 58590 -1160 58630 -1100
rect 58690 -1160 58730 -1100
rect 58590 -1200 58730 -1160
rect 58590 -1260 58630 -1200
rect 58690 -1260 58730 -1200
rect 58590 -1300 58730 -1260
rect 58590 -1360 58630 -1300
rect 58690 -1360 58730 -1300
rect 58590 -1380 58730 -1360
rect 58760 -1000 58900 -980
rect 58760 -1060 58800 -1000
rect 58860 -1060 58900 -1000
rect 58760 -1100 58900 -1060
rect 58760 -1160 58800 -1100
rect 58860 -1160 58900 -1100
rect 58760 -1200 58900 -1160
rect 58760 -1260 58800 -1200
rect 58860 -1260 58900 -1200
rect 58760 -1300 58900 -1260
rect 58760 -1360 58800 -1300
rect 58860 -1360 58900 -1300
rect 58760 -1380 58900 -1360
rect 58930 -1000 59070 -980
rect 58930 -1060 58970 -1000
rect 59030 -1060 59070 -1000
rect 58930 -1100 59070 -1060
rect 58930 -1160 58970 -1100
rect 59030 -1160 59070 -1100
rect 58930 -1200 59070 -1160
rect 58930 -1260 58970 -1200
rect 59030 -1260 59070 -1200
rect 58930 -1300 59070 -1260
rect 58930 -1360 58970 -1300
rect 59030 -1360 59070 -1300
rect 58930 -1380 59070 -1360
rect 59100 -1000 59240 -980
rect 59100 -1060 59140 -1000
rect 59200 -1060 59240 -1000
rect 59100 -1100 59240 -1060
rect 59100 -1160 59140 -1100
rect 59200 -1160 59240 -1100
rect 59100 -1200 59240 -1160
rect 59100 -1260 59140 -1200
rect 59200 -1260 59240 -1200
rect 59100 -1300 59240 -1260
rect 59100 -1360 59140 -1300
rect 59200 -1360 59240 -1300
rect 59100 -1380 59240 -1360
rect 59270 -1000 59410 -980
rect 59270 -1060 59310 -1000
rect 59370 -1060 59410 -1000
rect 59270 -1100 59410 -1060
rect 59270 -1160 59310 -1100
rect 59370 -1160 59410 -1100
rect 59270 -1200 59410 -1160
rect 59270 -1260 59310 -1200
rect 59370 -1260 59410 -1200
rect 59270 -1300 59410 -1260
rect 59270 -1360 59310 -1300
rect 59370 -1360 59410 -1300
rect 59270 -1380 59410 -1360
rect 59440 -1000 59580 -980
rect 59440 -1060 59480 -1000
rect 59540 -1060 59580 -1000
rect 59440 -1100 59580 -1060
rect 59440 -1160 59480 -1100
rect 59540 -1160 59580 -1100
rect 59440 -1200 59580 -1160
rect 59440 -1260 59480 -1200
rect 59540 -1260 59580 -1200
rect 59440 -1300 59580 -1260
rect 59440 -1360 59480 -1300
rect 59540 -1360 59580 -1300
rect 59440 -1380 59580 -1360
rect 59610 -1000 59750 -980
rect 59610 -1060 59650 -1000
rect 59710 -1060 59750 -1000
rect 59610 -1100 59750 -1060
rect 59610 -1160 59650 -1100
rect 59710 -1160 59750 -1100
rect 59610 -1200 59750 -1160
rect 59610 -1260 59650 -1200
rect 59710 -1260 59750 -1200
rect 59610 -1300 59750 -1260
rect 59610 -1360 59650 -1300
rect 59710 -1360 59750 -1300
rect 59610 -1380 59750 -1360
rect 59780 -1000 59920 -980
rect 59780 -1060 59820 -1000
rect 59880 -1060 59920 -1000
rect 59780 -1100 59920 -1060
rect 59780 -1160 59820 -1100
rect 59880 -1160 59920 -1100
rect 59780 -1200 59920 -1160
rect 59780 -1260 59820 -1200
rect 59880 -1260 59920 -1200
rect 59780 -1300 59920 -1260
rect 59780 -1360 59820 -1300
rect 59880 -1360 59920 -1300
rect 59780 -1380 59920 -1360
rect 59950 -1000 60090 -980
rect 59950 -1060 59990 -1000
rect 60050 -1060 60090 -1000
rect 59950 -1100 60090 -1060
rect 59950 -1160 59990 -1100
rect 60050 -1160 60090 -1100
rect 59950 -1200 60090 -1160
rect 59950 -1260 59990 -1200
rect 60050 -1260 60090 -1200
rect 59950 -1300 60090 -1260
rect 59950 -1360 59990 -1300
rect 60050 -1360 60090 -1300
rect 59950 -1380 60090 -1360
rect 60120 -1000 60260 -980
rect 60120 -1060 60160 -1000
rect 60220 -1060 60260 -1000
rect 60120 -1100 60260 -1060
rect 60120 -1160 60160 -1100
rect 60220 -1160 60260 -1100
rect 60120 -1200 60260 -1160
rect 60120 -1260 60160 -1200
rect 60220 -1260 60260 -1200
rect 60120 -1300 60260 -1260
rect 60120 -1360 60160 -1300
rect 60220 -1360 60260 -1300
rect 60120 -1380 60260 -1360
rect 60290 -1000 60430 -980
rect 60290 -1060 60330 -1000
rect 60390 -1060 60430 -1000
rect 60290 -1100 60430 -1060
rect 60290 -1160 60330 -1100
rect 60390 -1160 60430 -1100
rect 60290 -1200 60430 -1160
rect 60290 -1260 60330 -1200
rect 60390 -1260 60430 -1200
rect 60290 -1300 60430 -1260
rect 60290 -1360 60330 -1300
rect 60390 -1360 60430 -1300
rect 60290 -1380 60430 -1360
rect 60460 -1000 60600 -980
rect 60460 -1060 60500 -1000
rect 60560 -1060 60600 -1000
rect 60460 -1100 60600 -1060
rect 60460 -1160 60500 -1100
rect 60560 -1160 60600 -1100
rect 60460 -1200 60600 -1160
rect 60460 -1260 60500 -1200
rect 60560 -1260 60600 -1200
rect 60460 -1300 60600 -1260
rect 60460 -1360 60500 -1300
rect 60560 -1360 60600 -1300
rect 60460 -1380 60600 -1360
rect 60630 -1000 60770 -980
rect 60630 -1060 60670 -1000
rect 60730 -1060 60770 -1000
rect 60630 -1100 60770 -1060
rect 60630 -1160 60670 -1100
rect 60730 -1160 60770 -1100
rect 60630 -1200 60770 -1160
rect 60630 -1260 60670 -1200
rect 60730 -1260 60770 -1200
rect 60630 -1300 60770 -1260
rect 60630 -1360 60670 -1300
rect 60730 -1360 60770 -1300
rect 60630 -1380 60770 -1360
rect 60800 -1000 60940 -980
rect 60800 -1060 60840 -1000
rect 60900 -1060 60940 -1000
rect 60800 -1100 60940 -1060
rect 60800 -1160 60840 -1100
rect 60900 -1160 60940 -1100
rect 60800 -1200 60940 -1160
rect 60800 -1260 60840 -1200
rect 60900 -1260 60940 -1200
rect 60800 -1300 60940 -1260
rect 60800 -1360 60840 -1300
rect 60900 -1360 60940 -1300
rect 60800 -1380 60940 -1360
rect 60970 -1000 61110 -980
rect 60970 -1060 61010 -1000
rect 61070 -1060 61110 -1000
rect 60970 -1100 61110 -1060
rect 60970 -1160 61010 -1100
rect 61070 -1160 61110 -1100
rect 60970 -1200 61110 -1160
rect 60970 -1260 61010 -1200
rect 61070 -1260 61110 -1200
rect 60970 -1300 61110 -1260
rect 60970 -1360 61010 -1300
rect 61070 -1360 61110 -1300
rect 60970 -1380 61110 -1360
rect 61140 -1000 61280 -980
rect 61140 -1060 61180 -1000
rect 61240 -1060 61280 -1000
rect 61140 -1100 61280 -1060
rect 61140 -1160 61180 -1100
rect 61240 -1160 61280 -1100
rect 61140 -1200 61280 -1160
rect 61140 -1260 61180 -1200
rect 61240 -1260 61280 -1200
rect 61140 -1300 61280 -1260
rect 61140 -1360 61180 -1300
rect 61240 -1360 61280 -1300
rect 61140 -1380 61280 -1360
rect 61310 -1000 61450 -980
rect 61310 -1060 61350 -1000
rect 61410 -1060 61450 -1000
rect 61310 -1100 61450 -1060
rect 61310 -1160 61350 -1100
rect 61410 -1160 61450 -1100
rect 61310 -1200 61450 -1160
rect 61310 -1260 61350 -1200
rect 61410 -1260 61450 -1200
rect 61310 -1300 61450 -1260
rect 61310 -1360 61350 -1300
rect 61410 -1360 61450 -1300
rect 61310 -1380 61450 -1360
rect 61480 -1000 61620 -980
rect 61480 -1060 61520 -1000
rect 61580 -1060 61620 -1000
rect 61480 -1100 61620 -1060
rect 61480 -1160 61520 -1100
rect 61580 -1160 61620 -1100
rect 61480 -1200 61620 -1160
rect 61480 -1260 61520 -1200
rect 61580 -1260 61620 -1200
rect 61480 -1300 61620 -1260
rect 61480 -1360 61520 -1300
rect 61580 -1360 61620 -1300
rect 61480 -1380 61620 -1360
rect 61650 -1000 61790 -980
rect 61650 -1060 61690 -1000
rect 61750 -1060 61790 -1000
rect 61650 -1100 61790 -1060
rect 61650 -1160 61690 -1100
rect 61750 -1160 61790 -1100
rect 61650 -1200 61790 -1160
rect 61650 -1260 61690 -1200
rect 61750 -1260 61790 -1200
rect 61650 -1300 61790 -1260
rect 61650 -1360 61690 -1300
rect 61750 -1360 61790 -1300
rect 61650 -1380 61790 -1360
rect 61820 -1000 61960 -980
rect 61820 -1060 61860 -1000
rect 61920 -1060 61960 -1000
rect 61820 -1100 61960 -1060
rect 61820 -1160 61860 -1100
rect 61920 -1160 61960 -1100
rect 61820 -1200 61960 -1160
rect 61820 -1260 61860 -1200
rect 61920 -1260 61960 -1200
rect 61820 -1300 61960 -1260
rect 61820 -1360 61860 -1300
rect 61920 -1360 61960 -1300
rect 61820 -1380 61960 -1360
rect 61990 -1000 62130 -980
rect 61990 -1060 62030 -1000
rect 62090 -1060 62130 -1000
rect 61990 -1100 62130 -1060
rect 61990 -1160 62030 -1100
rect 62090 -1160 62130 -1100
rect 61990 -1200 62130 -1160
rect 61990 -1260 62030 -1200
rect 62090 -1260 62130 -1200
rect 61990 -1300 62130 -1260
rect 61990 -1360 62030 -1300
rect 62090 -1360 62130 -1300
rect 61990 -1380 62130 -1360
rect 62160 -1000 62300 -980
rect 62160 -1060 62200 -1000
rect 62260 -1060 62300 -1000
rect 62160 -1100 62300 -1060
rect 62160 -1160 62200 -1100
rect 62260 -1160 62300 -1100
rect 62160 -1200 62300 -1160
rect 62160 -1260 62200 -1200
rect 62260 -1260 62300 -1200
rect 62160 -1300 62300 -1260
rect 62160 -1360 62200 -1300
rect 62260 -1360 62300 -1300
rect 62160 -1380 62300 -1360
rect 62330 -1000 62470 -980
rect 62330 -1060 62370 -1000
rect 62430 -1060 62470 -1000
rect 62330 -1100 62470 -1060
rect 62330 -1160 62370 -1100
rect 62430 -1160 62470 -1100
rect 62330 -1200 62470 -1160
rect 62330 -1260 62370 -1200
rect 62430 -1260 62470 -1200
rect 62330 -1300 62470 -1260
rect 62330 -1360 62370 -1300
rect 62430 -1360 62470 -1300
rect 62330 -1380 62470 -1360
rect 62500 -1000 62640 -980
rect 62500 -1060 62540 -1000
rect 62600 -1060 62640 -1000
rect 62500 -1100 62640 -1060
rect 62500 -1160 62540 -1100
rect 62600 -1160 62640 -1100
rect 62500 -1200 62640 -1160
rect 62500 -1260 62540 -1200
rect 62600 -1260 62640 -1200
rect 62500 -1300 62640 -1260
rect 62500 -1360 62540 -1300
rect 62600 -1360 62640 -1300
rect 62500 -1380 62640 -1360
rect 62670 -1000 62810 -980
rect 62670 -1060 62710 -1000
rect 62770 -1060 62810 -1000
rect 62670 -1100 62810 -1060
rect 62670 -1160 62710 -1100
rect 62770 -1160 62810 -1100
rect 62670 -1200 62810 -1160
rect 62670 -1260 62710 -1200
rect 62770 -1260 62810 -1200
rect 62670 -1300 62810 -1260
rect 62670 -1360 62710 -1300
rect 62770 -1360 62810 -1300
rect 62670 -1380 62810 -1360
rect 62840 -1000 62980 -980
rect 62840 -1060 62880 -1000
rect 62940 -1060 62980 -1000
rect 62840 -1100 62980 -1060
rect 62840 -1160 62880 -1100
rect 62940 -1160 62980 -1100
rect 62840 -1200 62980 -1160
rect 62840 -1260 62880 -1200
rect 62940 -1260 62980 -1200
rect 62840 -1300 62980 -1260
rect 62840 -1360 62880 -1300
rect 62940 -1360 62980 -1300
rect 62840 -1380 62980 -1360
rect 63010 -1000 63150 -980
rect 63010 -1060 63050 -1000
rect 63110 -1060 63150 -1000
rect 63010 -1100 63150 -1060
rect 63010 -1160 63050 -1100
rect 63110 -1160 63150 -1100
rect 63010 -1200 63150 -1160
rect 63010 -1260 63050 -1200
rect 63110 -1260 63150 -1200
rect 63010 -1300 63150 -1260
rect 63010 -1360 63050 -1300
rect 63110 -1360 63150 -1300
rect 63010 -1380 63150 -1360
rect 63180 -1000 63320 -980
rect 63180 -1060 63220 -1000
rect 63280 -1060 63320 -1000
rect 63180 -1100 63320 -1060
rect 63180 -1160 63220 -1100
rect 63280 -1160 63320 -1100
rect 63180 -1200 63320 -1160
rect 63180 -1260 63220 -1200
rect 63280 -1260 63320 -1200
rect 63180 -1300 63320 -1260
rect 63180 -1360 63220 -1300
rect 63280 -1360 63320 -1300
rect 63180 -1380 63320 -1360
rect 63350 -1000 63490 -980
rect 63350 -1060 63390 -1000
rect 63450 -1060 63490 -1000
rect 63350 -1100 63490 -1060
rect 63350 -1160 63390 -1100
rect 63450 -1160 63490 -1100
rect 63350 -1200 63490 -1160
rect 63350 -1260 63390 -1200
rect 63450 -1260 63490 -1200
rect 63350 -1300 63490 -1260
rect 63350 -1360 63390 -1300
rect 63450 -1360 63490 -1300
rect 63350 -1380 63490 -1360
rect 63520 -1000 63660 -980
rect 63520 -1060 63560 -1000
rect 63620 -1060 63660 -1000
rect 63520 -1100 63660 -1060
rect 63520 -1160 63560 -1100
rect 63620 -1160 63660 -1100
rect 63520 -1200 63660 -1160
rect 63520 -1260 63560 -1200
rect 63620 -1260 63660 -1200
rect 63520 -1300 63660 -1260
rect 63520 -1360 63560 -1300
rect 63620 -1360 63660 -1300
rect 63520 -1380 63660 -1360
rect 63690 -1000 63830 -980
rect 63690 -1060 63730 -1000
rect 63790 -1060 63830 -1000
rect 63690 -1100 63830 -1060
rect 63690 -1160 63730 -1100
rect 63790 -1160 63830 -1100
rect 63690 -1200 63830 -1160
rect 63690 -1260 63730 -1200
rect 63790 -1260 63830 -1200
rect 63690 -1300 63830 -1260
rect 63690 -1360 63730 -1300
rect 63790 -1360 63830 -1300
rect 63690 -1380 63830 -1360
rect 63860 -1000 64000 -980
rect 63860 -1060 63900 -1000
rect 63960 -1060 64000 -1000
rect 63860 -1100 64000 -1060
rect 63860 -1160 63900 -1100
rect 63960 -1160 64000 -1100
rect 63860 -1200 64000 -1160
rect 63860 -1260 63900 -1200
rect 63960 -1260 64000 -1200
rect 63860 -1300 64000 -1260
rect 63860 -1360 63900 -1300
rect 63960 -1360 64000 -1300
rect 63860 -1380 64000 -1360
rect 64030 -1000 64170 -980
rect 64030 -1060 64070 -1000
rect 64130 -1060 64170 -1000
rect 64030 -1100 64170 -1060
rect 64030 -1160 64070 -1100
rect 64130 -1160 64170 -1100
rect 64030 -1200 64170 -1160
rect 64030 -1260 64070 -1200
rect 64130 -1260 64170 -1200
rect 64030 -1300 64170 -1260
rect 64030 -1360 64070 -1300
rect 64130 -1360 64170 -1300
rect 64030 -1380 64170 -1360
rect 64200 -1000 64340 -980
rect 64200 -1060 64240 -1000
rect 64300 -1060 64340 -1000
rect 64200 -1100 64340 -1060
rect 64200 -1160 64240 -1100
rect 64300 -1160 64340 -1100
rect 64200 -1200 64340 -1160
rect 64200 -1260 64240 -1200
rect 64300 -1260 64340 -1200
rect 64200 -1300 64340 -1260
rect 64200 -1360 64240 -1300
rect 64300 -1360 64340 -1300
rect 64200 -1380 64340 -1360
rect 64370 -1000 64510 -980
rect 64370 -1060 64410 -1000
rect 64470 -1060 64510 -1000
rect 64370 -1100 64510 -1060
rect 64370 -1160 64410 -1100
rect 64470 -1160 64510 -1100
rect 64370 -1200 64510 -1160
rect 64370 -1260 64410 -1200
rect 64470 -1260 64510 -1200
rect 64370 -1300 64510 -1260
rect 64370 -1360 64410 -1300
rect 64470 -1360 64510 -1300
rect 64370 -1380 64510 -1360
rect 64540 -1000 64680 -980
rect 64540 -1060 64580 -1000
rect 64640 -1060 64680 -1000
rect 64540 -1100 64680 -1060
rect 64540 -1160 64580 -1100
rect 64640 -1160 64680 -1100
rect 64540 -1200 64680 -1160
rect 64540 -1260 64580 -1200
rect 64640 -1260 64680 -1200
rect 64540 -1300 64680 -1260
rect 64540 -1360 64580 -1300
rect 64640 -1360 64680 -1300
rect 64540 -1380 64680 -1360
rect 64710 -1000 64850 -980
rect 64710 -1060 64750 -1000
rect 64810 -1060 64850 -1000
rect 64710 -1100 64850 -1060
rect 64710 -1160 64750 -1100
rect 64810 -1160 64850 -1100
rect 64710 -1200 64850 -1160
rect 64710 -1260 64750 -1200
rect 64810 -1260 64850 -1200
rect 64710 -1300 64850 -1260
rect 64710 -1360 64750 -1300
rect 64810 -1360 64850 -1300
rect 64710 -1380 64850 -1360
rect 64880 -1000 65020 -980
rect 64880 -1060 64920 -1000
rect 64980 -1060 65020 -1000
rect 64880 -1100 65020 -1060
rect 64880 -1160 64920 -1100
rect 64980 -1160 65020 -1100
rect 64880 -1200 65020 -1160
rect 64880 -1260 64920 -1200
rect 64980 -1260 65020 -1200
rect 64880 -1300 65020 -1260
rect 64880 -1360 64920 -1300
rect 64980 -1360 65020 -1300
rect 64880 -1380 65020 -1360
rect 65050 -1000 65190 -980
rect 65050 -1060 65090 -1000
rect 65150 -1060 65190 -1000
rect 65050 -1100 65190 -1060
rect 65050 -1160 65090 -1100
rect 65150 -1160 65190 -1100
rect 65050 -1200 65190 -1160
rect 65050 -1260 65090 -1200
rect 65150 -1260 65190 -1200
rect 65050 -1300 65190 -1260
rect 65050 -1360 65090 -1300
rect 65150 -1360 65190 -1300
rect 65050 -1380 65190 -1360
rect 65220 -1000 65360 -980
rect 65220 -1060 65260 -1000
rect 65320 -1060 65360 -1000
rect 65220 -1100 65360 -1060
rect 65220 -1160 65260 -1100
rect 65320 -1160 65360 -1100
rect 65220 -1200 65360 -1160
rect 65220 -1260 65260 -1200
rect 65320 -1260 65360 -1200
rect 65220 -1300 65360 -1260
rect 65220 -1360 65260 -1300
rect 65320 -1360 65360 -1300
rect 65220 -1380 65360 -1360
rect 65390 -1000 65530 -980
rect 65390 -1060 65430 -1000
rect 65490 -1060 65530 -1000
rect 65390 -1100 65530 -1060
rect 65390 -1160 65430 -1100
rect 65490 -1160 65530 -1100
rect 65390 -1200 65530 -1160
rect 65390 -1260 65430 -1200
rect 65490 -1260 65530 -1200
rect 65390 -1300 65530 -1260
rect 65390 -1360 65430 -1300
rect 65490 -1360 65530 -1300
rect 65390 -1380 65530 -1360
rect 65560 -1000 65700 -980
rect 65560 -1060 65600 -1000
rect 65660 -1060 65700 -1000
rect 65560 -1100 65700 -1060
rect 65560 -1160 65600 -1100
rect 65660 -1160 65700 -1100
rect 65560 -1200 65700 -1160
rect 65560 -1260 65600 -1200
rect 65660 -1260 65700 -1200
rect 65560 -1300 65700 -1260
rect 65560 -1360 65600 -1300
rect 65660 -1360 65700 -1300
rect 65560 -1380 65700 -1360
rect 65730 -1000 65870 -980
rect 65730 -1060 65770 -1000
rect 65830 -1060 65870 -1000
rect 65730 -1100 65870 -1060
rect 65730 -1160 65770 -1100
rect 65830 -1160 65870 -1100
rect 65730 -1200 65870 -1160
rect 65730 -1260 65770 -1200
rect 65830 -1260 65870 -1200
rect 65730 -1300 65870 -1260
rect 65730 -1360 65770 -1300
rect 65830 -1360 65870 -1300
rect 65730 -1380 65870 -1360
rect 65900 -1000 66040 -980
rect 65900 -1060 65940 -1000
rect 66000 -1060 66040 -1000
rect 65900 -1100 66040 -1060
rect 65900 -1160 65940 -1100
rect 66000 -1160 66040 -1100
rect 65900 -1200 66040 -1160
rect 65900 -1260 65940 -1200
rect 66000 -1260 66040 -1200
rect 65900 -1300 66040 -1260
rect 65900 -1360 65940 -1300
rect 66000 -1360 66040 -1300
rect 65900 -1380 66040 -1360
rect 66070 -1000 66210 -980
rect 66070 -1060 66110 -1000
rect 66170 -1060 66210 -1000
rect 66070 -1100 66210 -1060
rect 66070 -1160 66110 -1100
rect 66170 -1160 66210 -1100
rect 66070 -1200 66210 -1160
rect 66070 -1260 66110 -1200
rect 66170 -1260 66210 -1200
rect 66070 -1300 66210 -1260
rect 66070 -1360 66110 -1300
rect 66170 -1360 66210 -1300
rect 66070 -1380 66210 -1360
rect 66240 -1000 66380 -980
rect 66240 -1060 66280 -1000
rect 66340 -1060 66380 -1000
rect 66240 -1100 66380 -1060
rect 66240 -1160 66280 -1100
rect 66340 -1160 66380 -1100
rect 66240 -1200 66380 -1160
rect 66240 -1260 66280 -1200
rect 66340 -1260 66380 -1200
rect 66240 -1300 66380 -1260
rect 66240 -1360 66280 -1300
rect 66340 -1360 66380 -1300
rect 66240 -1380 66380 -1360
rect 66410 -1000 66550 -980
rect 66410 -1060 66450 -1000
rect 66510 -1060 66550 -1000
rect 66410 -1100 66550 -1060
rect 66410 -1160 66450 -1100
rect 66510 -1160 66550 -1100
rect 66410 -1200 66550 -1160
rect 66410 -1260 66450 -1200
rect 66510 -1260 66550 -1200
rect 66410 -1300 66550 -1260
rect 66410 -1360 66450 -1300
rect 66510 -1360 66550 -1300
rect 66410 -1380 66550 -1360
rect 66580 -1000 66720 -980
rect 66580 -1060 66620 -1000
rect 66680 -1060 66720 -1000
rect 66580 -1100 66720 -1060
rect 66580 -1160 66620 -1100
rect 66680 -1160 66720 -1100
rect 66580 -1200 66720 -1160
rect 66580 -1260 66620 -1200
rect 66680 -1260 66720 -1200
rect 66580 -1300 66720 -1260
rect 66580 -1360 66620 -1300
rect 66680 -1360 66720 -1300
rect 66580 -1380 66720 -1360
rect 66750 -1000 66890 -980
rect 66750 -1060 66790 -1000
rect 66850 -1060 66890 -1000
rect 66750 -1100 66890 -1060
rect 66750 -1160 66790 -1100
rect 66850 -1160 66890 -1100
rect 66750 -1200 66890 -1160
rect 66750 -1260 66790 -1200
rect 66850 -1260 66890 -1200
rect 66750 -1300 66890 -1260
rect 66750 -1360 66790 -1300
rect 66850 -1360 66890 -1300
rect 66750 -1380 66890 -1360
rect 66920 -1000 67060 -980
rect 66920 -1060 66960 -1000
rect 67020 -1060 67060 -1000
rect 66920 -1100 67060 -1060
rect 66920 -1160 66960 -1100
rect 67020 -1160 67060 -1100
rect 66920 -1200 67060 -1160
rect 66920 -1260 66960 -1200
rect 67020 -1260 67060 -1200
rect 66920 -1300 67060 -1260
rect 66920 -1360 66960 -1300
rect 67020 -1360 67060 -1300
rect 66920 -1380 67060 -1360
rect 67090 -1000 67230 -980
rect 67090 -1060 67130 -1000
rect 67190 -1060 67230 -1000
rect 67090 -1100 67230 -1060
rect 67090 -1160 67130 -1100
rect 67190 -1160 67230 -1100
rect 67090 -1200 67230 -1160
rect 67090 -1260 67130 -1200
rect 67190 -1260 67230 -1200
rect 67090 -1300 67230 -1260
rect 67090 -1360 67130 -1300
rect 67190 -1360 67230 -1300
rect 67090 -1380 67230 -1360
rect 67260 -1000 67400 -980
rect 67260 -1060 67300 -1000
rect 67360 -1060 67400 -1000
rect 67260 -1100 67400 -1060
rect 67260 -1160 67300 -1100
rect 67360 -1160 67400 -1100
rect 67260 -1200 67400 -1160
rect 67260 -1260 67300 -1200
rect 67360 -1260 67400 -1200
rect 67260 -1300 67400 -1260
rect 67260 -1360 67300 -1300
rect 67360 -1360 67400 -1300
rect 67260 -1380 67400 -1360
rect 67430 -1000 67570 -980
rect 67430 -1060 67470 -1000
rect 67530 -1060 67570 -1000
rect 67430 -1100 67570 -1060
rect 67430 -1160 67470 -1100
rect 67530 -1160 67570 -1100
rect 67430 -1200 67570 -1160
rect 67430 -1260 67470 -1200
rect 67530 -1260 67570 -1200
rect 67430 -1300 67570 -1260
rect 67430 -1360 67470 -1300
rect 67530 -1360 67570 -1300
rect 67430 -1380 67570 -1360
rect 67600 -1000 67740 -980
rect 67600 -1060 67640 -1000
rect 67700 -1060 67740 -1000
rect 67600 -1100 67740 -1060
rect 67600 -1160 67640 -1100
rect 67700 -1160 67740 -1100
rect 67600 -1200 67740 -1160
rect 67600 -1260 67640 -1200
rect 67700 -1260 67740 -1200
rect 67600 -1300 67740 -1260
rect 67600 -1360 67640 -1300
rect 67700 -1360 67740 -1300
rect 67600 -1380 67740 -1360
rect 67770 -1000 67910 -980
rect 67770 -1060 67810 -1000
rect 67870 -1060 67910 -1000
rect 67770 -1100 67910 -1060
rect 67770 -1160 67810 -1100
rect 67870 -1160 67910 -1100
rect 67770 -1200 67910 -1160
rect 67770 -1260 67810 -1200
rect 67870 -1260 67910 -1200
rect 67770 -1300 67910 -1260
rect 67770 -1360 67810 -1300
rect 67870 -1360 67910 -1300
rect 67770 -1380 67910 -1360
rect 67940 -1000 68080 -980
rect 67940 -1060 67980 -1000
rect 68040 -1060 68080 -1000
rect 67940 -1100 68080 -1060
rect 67940 -1160 67980 -1100
rect 68040 -1160 68080 -1100
rect 67940 -1200 68080 -1160
rect 67940 -1260 67980 -1200
rect 68040 -1260 68080 -1200
rect 67940 -1300 68080 -1260
rect 67940 -1360 67980 -1300
rect 68040 -1360 68080 -1300
rect 67940 -1380 68080 -1360
rect 68110 -1000 68250 -980
rect 68110 -1060 68150 -1000
rect 68210 -1060 68250 -1000
rect 68110 -1100 68250 -1060
rect 68110 -1160 68150 -1100
rect 68210 -1160 68250 -1100
rect 68110 -1200 68250 -1160
rect 68110 -1260 68150 -1200
rect 68210 -1260 68250 -1200
rect 68110 -1300 68250 -1260
rect 68110 -1360 68150 -1300
rect 68210 -1360 68250 -1300
rect 68110 -1380 68250 -1360
rect 68280 -1000 68420 -980
rect 68280 -1060 68320 -1000
rect 68380 -1060 68420 -1000
rect 68280 -1100 68420 -1060
rect 68280 -1160 68320 -1100
rect 68380 -1160 68420 -1100
rect 68280 -1200 68420 -1160
rect 68280 -1260 68320 -1200
rect 68380 -1260 68420 -1200
rect 68280 -1300 68420 -1260
rect 68280 -1360 68320 -1300
rect 68380 -1360 68420 -1300
rect 68280 -1380 68420 -1360
rect 68450 -1000 68590 -980
rect 68450 -1060 68490 -1000
rect 68550 -1060 68590 -1000
rect 68450 -1100 68590 -1060
rect 68450 -1160 68490 -1100
rect 68550 -1160 68590 -1100
rect 68450 -1200 68590 -1160
rect 68450 -1260 68490 -1200
rect 68550 -1260 68590 -1200
rect 68450 -1300 68590 -1260
rect 68450 -1360 68490 -1300
rect 68550 -1360 68590 -1300
rect 68450 -1380 68590 -1360
rect 68620 -1000 68760 -980
rect 68620 -1060 68660 -1000
rect 68720 -1060 68760 -1000
rect 68620 -1100 68760 -1060
rect 68620 -1160 68660 -1100
rect 68720 -1160 68760 -1100
rect 68620 -1200 68760 -1160
rect 68620 -1260 68660 -1200
rect 68720 -1260 68760 -1200
rect 68620 -1300 68760 -1260
rect 68620 -1360 68660 -1300
rect 68720 -1360 68760 -1300
rect 68620 -1380 68760 -1360
rect 68790 -1000 68930 -980
rect 68790 -1060 68830 -1000
rect 68890 -1060 68930 -1000
rect 68790 -1100 68930 -1060
rect 68790 -1160 68830 -1100
rect 68890 -1160 68930 -1100
rect 68790 -1200 68930 -1160
rect 68790 -1260 68830 -1200
rect 68890 -1260 68930 -1200
rect 68790 -1300 68930 -1260
rect 68790 -1360 68830 -1300
rect 68890 -1360 68930 -1300
rect 68790 -1380 68930 -1360
rect 68960 -1000 69100 -980
rect 68960 -1060 69000 -1000
rect 69060 -1060 69100 -1000
rect 68960 -1100 69100 -1060
rect 68960 -1160 69000 -1100
rect 69060 -1160 69100 -1100
rect 68960 -1200 69100 -1160
rect 68960 -1260 69000 -1200
rect 69060 -1260 69100 -1200
rect 68960 -1300 69100 -1260
rect 68960 -1360 69000 -1300
rect 69060 -1360 69100 -1300
rect 68960 -1380 69100 -1360
rect 69130 -1000 69270 -980
rect 69130 -1060 69170 -1000
rect 69230 -1060 69270 -1000
rect 69130 -1100 69270 -1060
rect 69130 -1160 69170 -1100
rect 69230 -1160 69270 -1100
rect 69130 -1200 69270 -1160
rect 69130 -1260 69170 -1200
rect 69230 -1260 69270 -1200
rect 69130 -1300 69270 -1260
rect 69130 -1360 69170 -1300
rect 69230 -1360 69270 -1300
rect 69130 -1380 69270 -1360
rect 69300 -1000 69440 -980
rect 69300 -1060 69340 -1000
rect 69400 -1060 69440 -1000
rect 69300 -1100 69440 -1060
rect 69300 -1160 69340 -1100
rect 69400 -1160 69440 -1100
rect 69300 -1200 69440 -1160
rect 69300 -1260 69340 -1200
rect 69400 -1260 69440 -1200
rect 69300 -1300 69440 -1260
rect 69300 -1360 69340 -1300
rect 69400 -1360 69440 -1300
rect 69300 -1380 69440 -1360
rect 69470 -1000 69610 -980
rect 69470 -1060 69510 -1000
rect 69570 -1060 69610 -1000
rect 69470 -1100 69610 -1060
rect 69470 -1160 69510 -1100
rect 69570 -1160 69610 -1100
rect 69470 -1200 69610 -1160
rect 69470 -1260 69510 -1200
rect 69570 -1260 69610 -1200
rect 69470 -1300 69610 -1260
rect 69470 -1360 69510 -1300
rect 69570 -1360 69610 -1300
rect 69470 -1380 69610 -1360
rect 69640 -1000 69780 -980
rect 69640 -1060 69680 -1000
rect 69740 -1060 69780 -1000
rect 69640 -1100 69780 -1060
rect 69640 -1160 69680 -1100
rect 69740 -1160 69780 -1100
rect 69640 -1200 69780 -1160
rect 69640 -1260 69680 -1200
rect 69740 -1260 69780 -1200
rect 69640 -1300 69780 -1260
rect 69640 -1360 69680 -1300
rect 69740 -1360 69780 -1300
rect 69640 -1380 69780 -1360
rect 69810 -1000 69950 -980
rect 69810 -1060 69850 -1000
rect 69910 -1060 69950 -1000
rect 69810 -1100 69950 -1060
rect 69810 -1160 69850 -1100
rect 69910 -1160 69950 -1100
rect 69810 -1200 69950 -1160
rect 69810 -1260 69850 -1200
rect 69910 -1260 69950 -1200
rect 69810 -1300 69950 -1260
rect 69810 -1360 69850 -1300
rect 69910 -1360 69950 -1300
rect 69810 -1380 69950 -1360
rect 69980 -1000 70120 -980
rect 69980 -1060 70020 -1000
rect 70080 -1060 70120 -1000
rect 69980 -1100 70120 -1060
rect 69980 -1160 70020 -1100
rect 70080 -1160 70120 -1100
rect 69980 -1200 70120 -1160
rect 69980 -1260 70020 -1200
rect 70080 -1260 70120 -1200
rect 69980 -1300 70120 -1260
rect 69980 -1360 70020 -1300
rect 70080 -1360 70120 -1300
rect 69980 -1380 70120 -1360
rect 70150 -1000 70290 -980
rect 70150 -1060 70190 -1000
rect 70250 -1060 70290 -1000
rect 70150 -1100 70290 -1060
rect 70150 -1160 70190 -1100
rect 70250 -1160 70290 -1100
rect 70150 -1200 70290 -1160
rect 70150 -1260 70190 -1200
rect 70250 -1260 70290 -1200
rect 70150 -1300 70290 -1260
rect 70150 -1360 70190 -1300
rect 70250 -1360 70290 -1300
rect 70150 -1380 70290 -1360
rect 70320 -1000 70460 -980
rect 70320 -1060 70360 -1000
rect 70420 -1060 70460 -1000
rect 70320 -1100 70460 -1060
rect 70320 -1160 70360 -1100
rect 70420 -1160 70460 -1100
rect 70320 -1200 70460 -1160
rect 70320 -1260 70360 -1200
rect 70420 -1260 70460 -1200
rect 70320 -1300 70460 -1260
rect 70320 -1360 70360 -1300
rect 70420 -1360 70460 -1300
rect 70320 -1380 70460 -1360
rect 70490 -1000 70630 -980
rect 70490 -1060 70530 -1000
rect 70590 -1060 70630 -1000
rect 70490 -1100 70630 -1060
rect 70490 -1160 70530 -1100
rect 70590 -1160 70630 -1100
rect 70490 -1200 70630 -1160
rect 70490 -1260 70530 -1200
rect 70590 -1260 70630 -1200
rect 70490 -1300 70630 -1260
rect 70490 -1360 70530 -1300
rect 70590 -1360 70630 -1300
rect 70490 -1380 70630 -1360
rect 70660 -1000 70800 -980
rect 70660 -1060 70700 -1000
rect 70760 -1060 70800 -1000
rect 70660 -1100 70800 -1060
rect 70660 -1160 70700 -1100
rect 70760 -1160 70800 -1100
rect 70660 -1200 70800 -1160
rect 70660 -1260 70700 -1200
rect 70760 -1260 70800 -1200
rect 70660 -1300 70800 -1260
rect 70660 -1360 70700 -1300
rect 70760 -1360 70800 -1300
rect 70660 -1380 70800 -1360
rect 70830 -1000 70970 -980
rect 70830 -1060 70870 -1000
rect 70930 -1060 70970 -1000
rect 70830 -1100 70970 -1060
rect 70830 -1160 70870 -1100
rect 70930 -1160 70970 -1100
rect 70830 -1200 70970 -1160
rect 70830 -1260 70870 -1200
rect 70930 -1260 70970 -1200
rect 70830 -1300 70970 -1260
rect 70830 -1360 70870 -1300
rect 70930 -1360 70970 -1300
rect 70830 -1380 70970 -1360
rect 71000 -1000 71140 -980
rect 71000 -1060 71040 -1000
rect 71100 -1060 71140 -1000
rect 71000 -1100 71140 -1060
rect 71000 -1160 71040 -1100
rect 71100 -1160 71140 -1100
rect 71000 -1200 71140 -1160
rect 71000 -1260 71040 -1200
rect 71100 -1260 71140 -1200
rect 71000 -1300 71140 -1260
rect 71000 -1360 71040 -1300
rect 71100 -1360 71140 -1300
rect 71000 -1380 71140 -1360
rect 71170 -1000 71310 -980
rect 71170 -1060 71210 -1000
rect 71270 -1060 71310 -1000
rect 71170 -1100 71310 -1060
rect 71170 -1160 71210 -1100
rect 71270 -1160 71310 -1100
rect 71170 -1200 71310 -1160
rect 71170 -1260 71210 -1200
rect 71270 -1260 71310 -1200
rect 71170 -1300 71310 -1260
rect 71170 -1360 71210 -1300
rect 71270 -1360 71310 -1300
rect 71170 -1380 71310 -1360
rect 71340 -1000 71480 -980
rect 71340 -1060 71380 -1000
rect 71440 -1060 71480 -1000
rect 71340 -1100 71480 -1060
rect 71340 -1160 71380 -1100
rect 71440 -1160 71480 -1100
rect 71340 -1200 71480 -1160
rect 71340 -1260 71380 -1200
rect 71440 -1260 71480 -1200
rect 71340 -1300 71480 -1260
rect 71340 -1360 71380 -1300
rect 71440 -1360 71480 -1300
rect 71340 -1380 71480 -1360
rect 71510 -1000 71650 -980
rect 71510 -1060 71550 -1000
rect 71610 -1060 71650 -1000
rect 71510 -1100 71650 -1060
rect 71510 -1160 71550 -1100
rect 71610 -1160 71650 -1100
rect 71510 -1200 71650 -1160
rect 71510 -1260 71550 -1200
rect 71610 -1260 71650 -1200
rect 71510 -1300 71650 -1260
rect 71510 -1360 71550 -1300
rect 71610 -1360 71650 -1300
rect 71510 -1380 71650 -1360
rect 71680 -1000 71820 -980
rect 71680 -1060 71720 -1000
rect 71780 -1060 71820 -1000
rect 71680 -1100 71820 -1060
rect 71680 -1160 71720 -1100
rect 71780 -1160 71820 -1100
rect 71680 -1200 71820 -1160
rect 71680 -1260 71720 -1200
rect 71780 -1260 71820 -1200
rect 71680 -1300 71820 -1260
rect 71680 -1360 71720 -1300
rect 71780 -1360 71820 -1300
rect 71680 -1380 71820 -1360
rect 71850 -1000 71990 -980
rect 71850 -1060 71890 -1000
rect 71950 -1060 71990 -1000
rect 71850 -1100 71990 -1060
rect 71850 -1160 71890 -1100
rect 71950 -1160 71990 -1100
rect 71850 -1200 71990 -1160
rect 71850 -1260 71890 -1200
rect 71950 -1260 71990 -1200
rect 71850 -1300 71990 -1260
rect 71850 -1360 71890 -1300
rect 71950 -1360 71990 -1300
rect 71850 -1380 71990 -1360
rect 72020 -1000 72160 -980
rect 72020 -1060 72060 -1000
rect 72120 -1060 72160 -1000
rect 72020 -1100 72160 -1060
rect 72020 -1160 72060 -1100
rect 72120 -1160 72160 -1100
rect 72020 -1200 72160 -1160
rect 72020 -1260 72060 -1200
rect 72120 -1260 72160 -1200
rect 72020 -1300 72160 -1260
rect 72020 -1360 72060 -1300
rect 72120 -1360 72160 -1300
rect 72020 -1380 72160 -1360
rect 72190 -1000 72330 -980
rect 72190 -1060 72230 -1000
rect 72290 -1060 72330 -1000
rect 72190 -1100 72330 -1060
rect 72190 -1160 72230 -1100
rect 72290 -1160 72330 -1100
rect 72190 -1200 72330 -1160
rect 72190 -1260 72230 -1200
rect 72290 -1260 72330 -1200
rect 72190 -1300 72330 -1260
rect 72190 -1360 72230 -1300
rect 72290 -1360 72330 -1300
rect 72190 -1380 72330 -1360
rect 72360 -1000 72500 -980
rect 72360 -1060 72400 -1000
rect 72460 -1060 72500 -1000
rect 72360 -1100 72500 -1060
rect 72360 -1160 72400 -1100
rect 72460 -1160 72500 -1100
rect 72360 -1200 72500 -1160
rect 72360 -1260 72400 -1200
rect 72460 -1260 72500 -1200
rect 72360 -1300 72500 -1260
rect 72360 -1360 72400 -1300
rect 72460 -1360 72500 -1300
rect 72360 -1380 72500 -1360
rect 72530 -1000 72670 -980
rect 72530 -1060 72570 -1000
rect 72630 -1060 72670 -1000
rect 72530 -1100 72670 -1060
rect 72530 -1160 72570 -1100
rect 72630 -1160 72670 -1100
rect 72530 -1200 72670 -1160
rect 72530 -1260 72570 -1200
rect 72630 -1260 72670 -1200
rect 72530 -1300 72670 -1260
rect 72530 -1360 72570 -1300
rect 72630 -1360 72670 -1300
rect 72530 -1380 72670 -1360
rect 72700 -1000 72840 -980
rect 72700 -1060 72740 -1000
rect 72800 -1060 72840 -1000
rect 72700 -1100 72840 -1060
rect 72700 -1160 72740 -1100
rect 72800 -1160 72840 -1100
rect 72700 -1200 72840 -1160
rect 72700 -1260 72740 -1200
rect 72800 -1260 72840 -1200
rect 72700 -1300 72840 -1260
rect 72700 -1360 72740 -1300
rect 72800 -1360 72840 -1300
rect 72700 -1380 72840 -1360
rect 72870 -1000 73010 -980
rect 72870 -1060 72910 -1000
rect 72970 -1060 73010 -1000
rect 72870 -1100 73010 -1060
rect 72870 -1160 72910 -1100
rect 72970 -1160 73010 -1100
rect 72870 -1200 73010 -1160
rect 72870 -1260 72910 -1200
rect 72970 -1260 73010 -1200
rect 72870 -1300 73010 -1260
rect 72870 -1360 72910 -1300
rect 72970 -1360 73010 -1300
rect 72870 -1380 73010 -1360
rect 73040 -1000 73180 -980
rect 73040 -1060 73080 -1000
rect 73140 -1060 73180 -1000
rect 73040 -1100 73180 -1060
rect 73040 -1160 73080 -1100
rect 73140 -1160 73180 -1100
rect 73040 -1200 73180 -1160
rect 73040 -1260 73080 -1200
rect 73140 -1260 73180 -1200
rect 73040 -1300 73180 -1260
rect 73040 -1360 73080 -1300
rect 73140 -1360 73180 -1300
rect 73040 -1380 73180 -1360
rect 73210 -1000 73350 -980
rect 73210 -1060 73250 -1000
rect 73310 -1060 73350 -1000
rect 73210 -1100 73350 -1060
rect 73210 -1160 73250 -1100
rect 73310 -1160 73350 -1100
rect 73210 -1200 73350 -1160
rect 73210 -1260 73250 -1200
rect 73310 -1260 73350 -1200
rect 73210 -1300 73350 -1260
rect 73210 -1360 73250 -1300
rect 73310 -1360 73350 -1300
rect 73210 -1380 73350 -1360
rect 73380 -1000 73520 -980
rect 73380 -1060 73420 -1000
rect 73480 -1060 73520 -1000
rect 73380 -1100 73520 -1060
rect 73380 -1160 73420 -1100
rect 73480 -1160 73520 -1100
rect 73380 -1200 73520 -1160
rect 73380 -1260 73420 -1200
rect 73480 -1260 73520 -1200
rect 73380 -1300 73520 -1260
rect 73380 -1360 73420 -1300
rect 73480 -1360 73520 -1300
rect 73380 -1380 73520 -1360
rect 73550 -1000 73690 -980
rect 73550 -1060 73590 -1000
rect 73650 -1060 73690 -1000
rect 73550 -1100 73690 -1060
rect 73550 -1160 73590 -1100
rect 73650 -1160 73690 -1100
rect 73550 -1200 73690 -1160
rect 73550 -1260 73590 -1200
rect 73650 -1260 73690 -1200
rect 73550 -1300 73690 -1260
rect 73550 -1360 73590 -1300
rect 73650 -1360 73690 -1300
rect 73550 -1380 73690 -1360
rect 73720 -1000 73860 -980
rect 73720 -1060 73760 -1000
rect 73820 -1060 73860 -1000
rect 73720 -1100 73860 -1060
rect 73720 -1160 73760 -1100
rect 73820 -1160 73860 -1100
rect 73720 -1200 73860 -1160
rect 73720 -1260 73760 -1200
rect 73820 -1260 73860 -1200
rect 73720 -1300 73860 -1260
rect 73720 -1360 73760 -1300
rect 73820 -1360 73860 -1300
rect 73720 -1380 73860 -1360
rect 73890 -1000 74030 -980
rect 73890 -1060 73930 -1000
rect 73990 -1060 74030 -1000
rect 73890 -1100 74030 -1060
rect 73890 -1160 73930 -1100
rect 73990 -1160 74030 -1100
rect 73890 -1200 74030 -1160
rect 73890 -1260 73930 -1200
rect 73990 -1260 74030 -1200
rect 73890 -1300 74030 -1260
rect 73890 -1360 73930 -1300
rect 73990 -1360 74030 -1300
rect 73890 -1380 74030 -1360
rect 74060 -1000 74200 -980
rect 74060 -1060 74100 -1000
rect 74160 -1060 74200 -1000
rect 74060 -1100 74200 -1060
rect 74060 -1160 74100 -1100
rect 74160 -1160 74200 -1100
rect 74060 -1200 74200 -1160
rect 74060 -1260 74100 -1200
rect 74160 -1260 74200 -1200
rect 74060 -1300 74200 -1260
rect 74060 -1360 74100 -1300
rect 74160 -1360 74200 -1300
rect 74060 -1380 74200 -1360
rect 74230 -1000 74370 -980
rect 74230 -1060 74270 -1000
rect 74330 -1060 74370 -1000
rect 74230 -1100 74370 -1060
rect 74230 -1160 74270 -1100
rect 74330 -1160 74370 -1100
rect 74230 -1200 74370 -1160
rect 74230 -1260 74270 -1200
rect 74330 -1260 74370 -1200
rect 74230 -1300 74370 -1260
rect 74230 -1360 74270 -1300
rect 74330 -1360 74370 -1300
rect 74230 -1380 74370 -1360
rect 74400 -1000 74540 -980
rect 74400 -1060 74440 -1000
rect 74500 -1060 74540 -1000
rect 74400 -1100 74540 -1060
rect 74400 -1160 74440 -1100
rect 74500 -1160 74540 -1100
rect 74400 -1200 74540 -1160
rect 74400 -1260 74440 -1200
rect 74500 -1260 74540 -1200
rect 74400 -1300 74540 -1260
rect 74400 -1360 74440 -1300
rect 74500 -1360 74540 -1300
rect 74400 -1380 74540 -1360
rect 74570 -1000 74710 -980
rect 74570 -1060 74610 -1000
rect 74670 -1060 74710 -1000
rect 74570 -1100 74710 -1060
rect 74570 -1160 74610 -1100
rect 74670 -1160 74710 -1100
rect 74570 -1200 74710 -1160
rect 74570 -1260 74610 -1200
rect 74670 -1260 74710 -1200
rect 74570 -1300 74710 -1260
rect 74570 -1360 74610 -1300
rect 74670 -1360 74710 -1300
rect 74570 -1380 74710 -1360
rect 74740 -1000 74880 -980
rect 74740 -1060 74780 -1000
rect 74840 -1060 74880 -1000
rect 74740 -1100 74880 -1060
rect 74740 -1160 74780 -1100
rect 74840 -1160 74880 -1100
rect 74740 -1200 74880 -1160
rect 74740 -1260 74780 -1200
rect 74840 -1260 74880 -1200
rect 74740 -1300 74880 -1260
rect 74740 -1360 74780 -1300
rect 74840 -1360 74880 -1300
rect 74740 -1380 74880 -1360
rect 74910 -1000 75050 -980
rect 74910 -1060 74950 -1000
rect 75010 -1060 75050 -1000
rect 74910 -1100 75050 -1060
rect 74910 -1160 74950 -1100
rect 75010 -1160 75050 -1100
rect 74910 -1200 75050 -1160
rect 74910 -1260 74950 -1200
rect 75010 -1260 75050 -1200
rect 74910 -1300 75050 -1260
rect 74910 -1360 74950 -1300
rect 75010 -1360 75050 -1300
rect 74910 -1380 75050 -1360
rect 75080 -1000 75220 -980
rect 75080 -1060 75120 -1000
rect 75180 -1060 75220 -1000
rect 75080 -1100 75220 -1060
rect 75080 -1160 75120 -1100
rect 75180 -1160 75220 -1100
rect 75080 -1200 75220 -1160
rect 75080 -1260 75120 -1200
rect 75180 -1260 75220 -1200
rect 75080 -1300 75220 -1260
rect 75080 -1360 75120 -1300
rect 75180 -1360 75220 -1300
rect 75080 -1380 75220 -1360
rect 75250 -1000 75390 -980
rect 75250 -1060 75290 -1000
rect 75350 -1060 75390 -1000
rect 75250 -1100 75390 -1060
rect 75250 -1160 75290 -1100
rect 75350 -1160 75390 -1100
rect 75250 -1200 75390 -1160
rect 75250 -1260 75290 -1200
rect 75350 -1260 75390 -1200
rect 75250 -1300 75390 -1260
rect 75250 -1360 75290 -1300
rect 75350 -1360 75390 -1300
rect 75250 -1380 75390 -1360
rect 75420 -1000 75560 -980
rect 75420 -1060 75460 -1000
rect 75520 -1060 75560 -1000
rect 75420 -1100 75560 -1060
rect 75420 -1160 75460 -1100
rect 75520 -1160 75560 -1100
rect 75420 -1200 75560 -1160
rect 75420 -1260 75460 -1200
rect 75520 -1260 75560 -1200
rect 75420 -1300 75560 -1260
rect 75420 -1360 75460 -1300
rect 75520 -1360 75560 -1300
rect 75420 -1380 75560 -1360
rect 75590 -1000 75730 -980
rect 75590 -1060 75630 -1000
rect 75690 -1060 75730 -1000
rect 75590 -1100 75730 -1060
rect 75590 -1160 75630 -1100
rect 75690 -1160 75730 -1100
rect 75590 -1200 75730 -1160
rect 75590 -1260 75630 -1200
rect 75690 -1260 75730 -1200
rect 75590 -1300 75730 -1260
rect 75590 -1360 75630 -1300
rect 75690 -1360 75730 -1300
rect 75590 -1380 75730 -1360
rect 75760 -1000 75900 -980
rect 75760 -1060 75800 -1000
rect 75860 -1060 75900 -1000
rect 75760 -1100 75900 -1060
rect 75760 -1160 75800 -1100
rect 75860 -1160 75900 -1100
rect 75760 -1200 75900 -1160
rect 75760 -1260 75800 -1200
rect 75860 -1260 75900 -1200
rect 75760 -1300 75900 -1260
rect 75760 -1360 75800 -1300
rect 75860 -1360 75900 -1300
rect 75760 -1380 75900 -1360
rect 75930 -1000 76070 -980
rect 75930 -1060 75970 -1000
rect 76030 -1060 76070 -1000
rect 75930 -1100 76070 -1060
rect 75930 -1160 75970 -1100
rect 76030 -1160 76070 -1100
rect 75930 -1200 76070 -1160
rect 75930 -1260 75970 -1200
rect 76030 -1260 76070 -1200
rect 75930 -1300 76070 -1260
rect 75930 -1360 75970 -1300
rect 76030 -1360 76070 -1300
rect 75930 -1380 76070 -1360
rect 76100 -1000 76240 -980
rect 76100 -1060 76140 -1000
rect 76200 -1060 76240 -1000
rect 76100 -1100 76240 -1060
rect 76100 -1160 76140 -1100
rect 76200 -1160 76240 -1100
rect 76100 -1200 76240 -1160
rect 76100 -1260 76140 -1200
rect 76200 -1260 76240 -1200
rect 76100 -1300 76240 -1260
rect 76100 -1360 76140 -1300
rect 76200 -1360 76240 -1300
rect 76100 -1380 76240 -1360
rect 76270 -1000 76410 -980
rect 76270 -1060 76310 -1000
rect 76370 -1060 76410 -1000
rect 76270 -1100 76410 -1060
rect 76270 -1160 76310 -1100
rect 76370 -1160 76410 -1100
rect 76270 -1200 76410 -1160
rect 76270 -1260 76310 -1200
rect 76370 -1260 76410 -1200
rect 76270 -1300 76410 -1260
rect 76270 -1360 76310 -1300
rect 76370 -1360 76410 -1300
rect 76270 -1380 76410 -1360
rect 76440 -1000 76580 -980
rect 76440 -1060 76480 -1000
rect 76540 -1060 76580 -1000
rect 76440 -1100 76580 -1060
rect 76440 -1160 76480 -1100
rect 76540 -1160 76580 -1100
rect 76440 -1200 76580 -1160
rect 76440 -1260 76480 -1200
rect 76540 -1260 76580 -1200
rect 76440 -1300 76580 -1260
rect 76440 -1360 76480 -1300
rect 76540 -1360 76580 -1300
rect 76440 -1380 76580 -1360
rect 76610 -1000 76750 -980
rect 76610 -1060 76650 -1000
rect 76710 -1060 76750 -1000
rect 76610 -1100 76750 -1060
rect 76610 -1160 76650 -1100
rect 76710 -1160 76750 -1100
rect 76610 -1200 76750 -1160
rect 76610 -1260 76650 -1200
rect 76710 -1260 76750 -1200
rect 76610 -1300 76750 -1260
rect 76610 -1360 76650 -1300
rect 76710 -1360 76750 -1300
rect 76610 -1380 76750 -1360
rect 76780 -1000 76920 -980
rect 76780 -1060 76820 -1000
rect 76880 -1060 76920 -1000
rect 76780 -1100 76920 -1060
rect 76780 -1160 76820 -1100
rect 76880 -1160 76920 -1100
rect 76780 -1200 76920 -1160
rect 76780 -1260 76820 -1200
rect 76880 -1260 76920 -1200
rect 76780 -1300 76920 -1260
rect 76780 -1360 76820 -1300
rect 76880 -1360 76920 -1300
rect 76780 -1380 76920 -1360
rect 76950 -1000 77090 -980
rect 76950 -1060 76990 -1000
rect 77050 -1060 77090 -1000
rect 76950 -1100 77090 -1060
rect 76950 -1160 76990 -1100
rect 77050 -1160 77090 -1100
rect 76950 -1200 77090 -1160
rect 76950 -1260 76990 -1200
rect 77050 -1260 77090 -1200
rect 76950 -1300 77090 -1260
rect 76950 -1360 76990 -1300
rect 77050 -1360 77090 -1300
rect 76950 -1380 77090 -1360
rect 77120 -1000 77260 -980
rect 77120 -1060 77160 -1000
rect 77220 -1060 77260 -1000
rect 77120 -1100 77260 -1060
rect 77120 -1160 77160 -1100
rect 77220 -1160 77260 -1100
rect 77120 -1200 77260 -1160
rect 77120 -1260 77160 -1200
rect 77220 -1260 77260 -1200
rect 77120 -1300 77260 -1260
rect 77120 -1360 77160 -1300
rect 77220 -1360 77260 -1300
rect 77120 -1380 77260 -1360
rect 77290 -1000 77430 -980
rect 77290 -1060 77330 -1000
rect 77390 -1060 77430 -1000
rect 77290 -1100 77430 -1060
rect 77290 -1160 77330 -1100
rect 77390 -1160 77430 -1100
rect 77290 -1200 77430 -1160
rect 77290 -1260 77330 -1200
rect 77390 -1260 77430 -1200
rect 77290 -1300 77430 -1260
rect 77290 -1360 77330 -1300
rect 77390 -1360 77430 -1300
rect 77290 -1380 77430 -1360
rect 77460 -1000 77600 -980
rect 77460 -1060 77500 -1000
rect 77560 -1060 77600 -1000
rect 77460 -1100 77600 -1060
rect 77460 -1160 77500 -1100
rect 77560 -1160 77600 -1100
rect 77460 -1200 77600 -1160
rect 77460 -1260 77500 -1200
rect 77560 -1260 77600 -1200
rect 77460 -1300 77600 -1260
rect 77460 -1360 77500 -1300
rect 77560 -1360 77600 -1300
rect 77460 -1380 77600 -1360
rect 77630 -1000 77770 -980
rect 77630 -1060 77670 -1000
rect 77730 -1060 77770 -1000
rect 77630 -1100 77770 -1060
rect 77630 -1160 77670 -1100
rect 77730 -1160 77770 -1100
rect 77630 -1200 77770 -1160
rect 77630 -1260 77670 -1200
rect 77730 -1260 77770 -1200
rect 77630 -1300 77770 -1260
rect 77630 -1360 77670 -1300
rect 77730 -1360 77770 -1300
rect 77630 -1380 77770 -1360
rect 77800 -1000 77940 -980
rect 77800 -1060 77840 -1000
rect 77900 -1060 77940 -1000
rect 77800 -1100 77940 -1060
rect 77800 -1160 77840 -1100
rect 77900 -1160 77940 -1100
rect 77800 -1200 77940 -1160
rect 77800 -1260 77840 -1200
rect 77900 -1260 77940 -1200
rect 77800 -1300 77940 -1260
rect 77800 -1360 77840 -1300
rect 77900 -1360 77940 -1300
rect 77800 -1380 77940 -1360
rect 77970 -1000 78110 -980
rect 77970 -1060 78010 -1000
rect 78070 -1060 78110 -1000
rect 77970 -1100 78110 -1060
rect 77970 -1160 78010 -1100
rect 78070 -1160 78110 -1100
rect 77970 -1200 78110 -1160
rect 77970 -1260 78010 -1200
rect 78070 -1260 78110 -1200
rect 77970 -1300 78110 -1260
rect 77970 -1360 78010 -1300
rect 78070 -1360 78110 -1300
rect 77970 -1380 78110 -1360
rect 78140 -1000 78280 -980
rect 78140 -1060 78180 -1000
rect 78240 -1060 78280 -1000
rect 78140 -1100 78280 -1060
rect 78140 -1160 78180 -1100
rect 78240 -1160 78280 -1100
rect 78140 -1200 78280 -1160
rect 78140 -1260 78180 -1200
rect 78240 -1260 78280 -1200
rect 78140 -1300 78280 -1260
rect 78140 -1360 78180 -1300
rect 78240 -1360 78280 -1300
rect 78140 -1380 78280 -1360
rect 78310 -1000 78450 -980
rect 78310 -1060 78350 -1000
rect 78410 -1060 78450 -1000
rect 78310 -1100 78450 -1060
rect 78310 -1160 78350 -1100
rect 78410 -1160 78450 -1100
rect 78310 -1200 78450 -1160
rect 78310 -1260 78350 -1200
rect 78410 -1260 78450 -1200
rect 78310 -1300 78450 -1260
rect 78310 -1360 78350 -1300
rect 78410 -1360 78450 -1300
rect 78310 -1380 78450 -1360
rect 78480 -1000 78620 -980
rect 78480 -1060 78520 -1000
rect 78580 -1060 78620 -1000
rect 78480 -1100 78620 -1060
rect 78480 -1160 78520 -1100
rect 78580 -1160 78620 -1100
rect 78480 -1200 78620 -1160
rect 78480 -1260 78520 -1200
rect 78580 -1260 78620 -1200
rect 78480 -1300 78620 -1260
rect 78480 -1360 78520 -1300
rect 78580 -1360 78620 -1300
rect 78480 -1380 78620 -1360
rect 78650 -1000 78790 -980
rect 78650 -1060 78690 -1000
rect 78750 -1060 78790 -1000
rect 78650 -1100 78790 -1060
rect 78650 -1160 78690 -1100
rect 78750 -1160 78790 -1100
rect 78650 -1200 78790 -1160
rect 78650 -1260 78690 -1200
rect 78750 -1260 78790 -1200
rect 78650 -1300 78790 -1260
rect 78650 -1360 78690 -1300
rect 78750 -1360 78790 -1300
rect 78650 -1380 78790 -1360
rect 78820 -1000 78960 -980
rect 78820 -1060 78860 -1000
rect 78920 -1060 78960 -1000
rect 78820 -1100 78960 -1060
rect 78820 -1160 78860 -1100
rect 78920 -1160 78960 -1100
rect 78820 -1200 78960 -1160
rect 78820 -1260 78860 -1200
rect 78920 -1260 78960 -1200
rect 78820 -1300 78960 -1260
rect 78820 -1360 78860 -1300
rect 78920 -1360 78960 -1300
rect 78820 -1380 78960 -1360
rect 78990 -1000 79130 -980
rect 78990 -1060 79030 -1000
rect 79090 -1060 79130 -1000
rect 78990 -1100 79130 -1060
rect 78990 -1160 79030 -1100
rect 79090 -1160 79130 -1100
rect 78990 -1200 79130 -1160
rect 78990 -1260 79030 -1200
rect 79090 -1260 79130 -1200
rect 78990 -1300 79130 -1260
rect 78990 -1360 79030 -1300
rect 79090 -1360 79130 -1300
rect 78990 -1380 79130 -1360
rect 79160 -1000 79300 -980
rect 79160 -1060 79200 -1000
rect 79260 -1060 79300 -1000
rect 79160 -1100 79300 -1060
rect 79160 -1160 79200 -1100
rect 79260 -1160 79300 -1100
rect 79160 -1200 79300 -1160
rect 79160 -1260 79200 -1200
rect 79260 -1260 79300 -1200
rect 79160 -1300 79300 -1260
rect 79160 -1360 79200 -1300
rect 79260 -1360 79300 -1300
rect 79160 -1380 79300 -1360
rect 79330 -1000 79470 -980
rect 79330 -1060 79370 -1000
rect 79430 -1060 79470 -1000
rect 79330 -1100 79470 -1060
rect 79330 -1160 79370 -1100
rect 79430 -1160 79470 -1100
rect 79330 -1200 79470 -1160
rect 79330 -1260 79370 -1200
rect 79430 -1260 79470 -1200
rect 79330 -1300 79470 -1260
rect 79330 -1360 79370 -1300
rect 79430 -1360 79470 -1300
rect 79330 -1380 79470 -1360
rect 79500 -1000 79640 -980
rect 79500 -1060 79540 -1000
rect 79600 -1060 79640 -1000
rect 79500 -1100 79640 -1060
rect 79500 -1160 79540 -1100
rect 79600 -1160 79640 -1100
rect 79500 -1200 79640 -1160
rect 79500 -1260 79540 -1200
rect 79600 -1260 79640 -1200
rect 79500 -1300 79640 -1260
rect 79500 -1360 79540 -1300
rect 79600 -1360 79640 -1300
rect 79500 -1380 79640 -1360
rect 79670 -1000 79810 -980
rect 79670 -1060 79710 -1000
rect 79770 -1060 79810 -1000
rect 79670 -1100 79810 -1060
rect 79670 -1160 79710 -1100
rect 79770 -1160 79810 -1100
rect 79670 -1200 79810 -1160
rect 79670 -1260 79710 -1200
rect 79770 -1260 79810 -1200
rect 79670 -1300 79810 -1260
rect 79670 -1360 79710 -1300
rect 79770 -1360 79810 -1300
rect 79670 -1380 79810 -1360
rect 79840 -1000 79980 -980
rect 79840 -1060 79880 -1000
rect 79940 -1060 79980 -1000
rect 79840 -1100 79980 -1060
rect 79840 -1160 79880 -1100
rect 79940 -1160 79980 -1100
rect 79840 -1200 79980 -1160
rect 79840 -1260 79880 -1200
rect 79940 -1260 79980 -1200
rect 79840 -1300 79980 -1260
rect 79840 -1360 79880 -1300
rect 79940 -1360 79980 -1300
rect 79840 -1380 79980 -1360
rect 80010 -1000 80150 -980
rect 80010 -1060 80050 -1000
rect 80110 -1060 80150 -1000
rect 80010 -1100 80150 -1060
rect 80010 -1160 80050 -1100
rect 80110 -1160 80150 -1100
rect 80010 -1200 80150 -1160
rect 80010 -1260 80050 -1200
rect 80110 -1260 80150 -1200
rect 80010 -1300 80150 -1260
rect 80010 -1360 80050 -1300
rect 80110 -1360 80150 -1300
rect 80010 -1380 80150 -1360
rect 80180 -1000 80320 -980
rect 80180 -1060 80220 -1000
rect 80280 -1060 80320 -1000
rect 80180 -1100 80320 -1060
rect 80180 -1160 80220 -1100
rect 80280 -1160 80320 -1100
rect 80180 -1200 80320 -1160
rect 80180 -1260 80220 -1200
rect 80280 -1260 80320 -1200
rect 80180 -1300 80320 -1260
rect 80180 -1360 80220 -1300
rect 80280 -1360 80320 -1300
rect 80180 -1380 80320 -1360
rect 80350 -1000 80490 -980
rect 80350 -1060 80390 -1000
rect 80450 -1060 80490 -1000
rect 80350 -1100 80490 -1060
rect 80350 -1160 80390 -1100
rect 80450 -1160 80490 -1100
rect 80350 -1200 80490 -1160
rect 80350 -1260 80390 -1200
rect 80450 -1260 80490 -1200
rect 80350 -1300 80490 -1260
rect 80350 -1360 80390 -1300
rect 80450 -1360 80490 -1300
rect 80350 -1380 80490 -1360
rect 80520 -1000 80660 -980
rect 80520 -1060 80560 -1000
rect 80620 -1060 80660 -1000
rect 80520 -1100 80660 -1060
rect 80520 -1160 80560 -1100
rect 80620 -1160 80660 -1100
rect 80520 -1200 80660 -1160
rect 80520 -1260 80560 -1200
rect 80620 -1260 80660 -1200
rect 80520 -1300 80660 -1260
rect 80520 -1360 80560 -1300
rect 80620 -1360 80660 -1300
rect 80520 -1380 80660 -1360
rect 80690 -1000 80830 -980
rect 80690 -1060 80730 -1000
rect 80790 -1060 80830 -1000
rect 80690 -1100 80830 -1060
rect 80690 -1160 80730 -1100
rect 80790 -1160 80830 -1100
rect 80690 -1200 80830 -1160
rect 80690 -1260 80730 -1200
rect 80790 -1260 80830 -1200
rect 80690 -1300 80830 -1260
rect 80690 -1360 80730 -1300
rect 80790 -1360 80830 -1300
rect 80690 -1380 80830 -1360
rect 80860 -1000 81000 -980
rect 80860 -1060 80900 -1000
rect 80960 -1060 81000 -1000
rect 80860 -1100 81000 -1060
rect 80860 -1160 80900 -1100
rect 80960 -1160 81000 -1100
rect 80860 -1200 81000 -1160
rect 80860 -1260 80900 -1200
rect 80960 -1260 81000 -1200
rect 80860 -1300 81000 -1260
rect 80860 -1360 80900 -1300
rect 80960 -1360 81000 -1300
rect 80860 -1380 81000 -1360
rect 81030 -1000 81170 -980
rect 81030 -1060 81070 -1000
rect 81130 -1060 81170 -1000
rect 81030 -1100 81170 -1060
rect 81030 -1160 81070 -1100
rect 81130 -1160 81170 -1100
rect 81030 -1200 81170 -1160
rect 81030 -1260 81070 -1200
rect 81130 -1260 81170 -1200
rect 81030 -1300 81170 -1260
rect 81030 -1360 81070 -1300
rect 81130 -1360 81170 -1300
rect 81030 -1380 81170 -1360
rect 81200 -1000 81340 -980
rect 81200 -1060 81240 -1000
rect 81300 -1060 81340 -1000
rect 81200 -1100 81340 -1060
rect 81200 -1160 81240 -1100
rect 81300 -1160 81340 -1100
rect 81200 -1200 81340 -1160
rect 81200 -1260 81240 -1200
rect 81300 -1260 81340 -1200
rect 81200 -1300 81340 -1260
rect 81200 -1360 81240 -1300
rect 81300 -1360 81340 -1300
rect 81200 -1380 81340 -1360
rect 81370 -1000 81510 -980
rect 81370 -1060 81410 -1000
rect 81470 -1060 81510 -1000
rect 81370 -1100 81510 -1060
rect 81370 -1160 81410 -1100
rect 81470 -1160 81510 -1100
rect 81370 -1200 81510 -1160
rect 81370 -1260 81410 -1200
rect 81470 -1260 81510 -1200
rect 81370 -1300 81510 -1260
rect 81370 -1360 81410 -1300
rect 81470 -1360 81510 -1300
rect 81370 -1380 81510 -1360
rect 81540 -1000 81680 -980
rect 81540 -1060 81580 -1000
rect 81640 -1060 81680 -1000
rect 81540 -1100 81680 -1060
rect 81540 -1160 81580 -1100
rect 81640 -1160 81680 -1100
rect 81540 -1200 81680 -1160
rect 81540 -1260 81580 -1200
rect 81640 -1260 81680 -1200
rect 81540 -1300 81680 -1260
rect 81540 -1360 81580 -1300
rect 81640 -1360 81680 -1300
rect 81540 -1380 81680 -1360
rect 81710 -1000 81850 -980
rect 81710 -1060 81750 -1000
rect 81810 -1060 81850 -1000
rect 81710 -1100 81850 -1060
rect 81710 -1160 81750 -1100
rect 81810 -1160 81850 -1100
rect 81710 -1200 81850 -1160
rect 81710 -1260 81750 -1200
rect 81810 -1260 81850 -1200
rect 81710 -1300 81850 -1260
rect 81710 -1360 81750 -1300
rect 81810 -1360 81850 -1300
rect 81710 -1380 81850 -1360
rect 81880 -1000 82020 -980
rect 81880 -1060 81920 -1000
rect 81980 -1060 82020 -1000
rect 81880 -1100 82020 -1060
rect 81880 -1160 81920 -1100
rect 81980 -1160 82020 -1100
rect 81880 -1200 82020 -1160
rect 81880 -1260 81920 -1200
rect 81980 -1260 82020 -1200
rect 81880 -1300 82020 -1260
rect 81880 -1360 81920 -1300
rect 81980 -1360 82020 -1300
rect 81880 -1380 82020 -1360
rect 82050 -1000 82190 -980
rect 82050 -1060 82090 -1000
rect 82150 -1060 82190 -1000
rect 82050 -1100 82190 -1060
rect 82050 -1160 82090 -1100
rect 82150 -1160 82190 -1100
rect 82050 -1200 82190 -1160
rect 82050 -1260 82090 -1200
rect 82150 -1260 82190 -1200
rect 82050 -1300 82190 -1260
rect 82050 -1360 82090 -1300
rect 82150 -1360 82190 -1300
rect 82050 -1380 82190 -1360
rect 82220 -1000 82360 -980
rect 82220 -1060 82260 -1000
rect 82320 -1060 82360 -1000
rect 82220 -1100 82360 -1060
rect 82220 -1160 82260 -1100
rect 82320 -1160 82360 -1100
rect 82220 -1200 82360 -1160
rect 82220 -1260 82260 -1200
rect 82320 -1260 82360 -1200
rect 82220 -1300 82360 -1260
rect 82220 -1360 82260 -1300
rect 82320 -1360 82360 -1300
rect 82220 -1380 82360 -1360
rect 82390 -1000 82530 -980
rect 82390 -1060 82430 -1000
rect 82490 -1060 82530 -1000
rect 82390 -1100 82530 -1060
rect 82390 -1160 82430 -1100
rect 82490 -1160 82530 -1100
rect 82390 -1200 82530 -1160
rect 82390 -1260 82430 -1200
rect 82490 -1260 82530 -1200
rect 82390 -1300 82530 -1260
rect 82390 -1360 82430 -1300
rect 82490 -1360 82530 -1300
rect 82390 -1380 82530 -1360
rect 82560 -1000 82700 -980
rect 82560 -1060 82600 -1000
rect 82660 -1060 82700 -1000
rect 82560 -1100 82700 -1060
rect 82560 -1160 82600 -1100
rect 82660 -1160 82700 -1100
rect 82560 -1200 82700 -1160
rect 82560 -1260 82600 -1200
rect 82660 -1260 82700 -1200
rect 82560 -1300 82700 -1260
rect 82560 -1360 82600 -1300
rect 82660 -1360 82700 -1300
rect 82560 -1380 82700 -1360
rect 82730 -1000 82870 -980
rect 82730 -1060 82770 -1000
rect 82830 -1060 82870 -1000
rect 82730 -1100 82870 -1060
rect 82730 -1160 82770 -1100
rect 82830 -1160 82870 -1100
rect 82730 -1200 82870 -1160
rect 82730 -1260 82770 -1200
rect 82830 -1260 82870 -1200
rect 82730 -1300 82870 -1260
rect 82730 -1360 82770 -1300
rect 82830 -1360 82870 -1300
rect 82730 -1380 82870 -1360
rect 82900 -1000 83040 -980
rect 82900 -1060 82940 -1000
rect 83000 -1060 83040 -1000
rect 82900 -1100 83040 -1060
rect 82900 -1160 82940 -1100
rect 83000 -1160 83040 -1100
rect 82900 -1200 83040 -1160
rect 82900 -1260 82940 -1200
rect 83000 -1260 83040 -1200
rect 82900 -1300 83040 -1260
rect 82900 -1360 82940 -1300
rect 83000 -1360 83040 -1300
rect 82900 -1380 83040 -1360
rect 83070 -1000 83210 -980
rect 83070 -1060 83110 -1000
rect 83170 -1060 83210 -1000
rect 83070 -1100 83210 -1060
rect 83070 -1160 83110 -1100
rect 83170 -1160 83210 -1100
rect 83070 -1200 83210 -1160
rect 83070 -1260 83110 -1200
rect 83170 -1260 83210 -1200
rect 83070 -1300 83210 -1260
rect 83070 -1360 83110 -1300
rect 83170 -1360 83210 -1300
rect 83070 -1380 83210 -1360
rect 83240 -1000 83380 -980
rect 83240 -1060 83280 -1000
rect 83340 -1060 83380 -1000
rect 83240 -1100 83380 -1060
rect 83240 -1160 83280 -1100
rect 83340 -1160 83380 -1100
rect 83240 -1200 83380 -1160
rect 83240 -1260 83280 -1200
rect 83340 -1260 83380 -1200
rect 83240 -1300 83380 -1260
rect 83240 -1360 83280 -1300
rect 83340 -1360 83380 -1300
rect 83240 -1380 83380 -1360
rect 83410 -1000 83550 -980
rect 83410 -1060 83450 -1000
rect 83510 -1060 83550 -1000
rect 83410 -1100 83550 -1060
rect 83410 -1160 83450 -1100
rect 83510 -1160 83550 -1100
rect 83410 -1200 83550 -1160
rect 83410 -1260 83450 -1200
rect 83510 -1260 83550 -1200
rect 83410 -1300 83550 -1260
rect 83410 -1360 83450 -1300
rect 83510 -1360 83550 -1300
rect 83410 -1380 83550 -1360
rect 83580 -1000 83720 -980
rect 83580 -1060 83620 -1000
rect 83680 -1060 83720 -1000
rect 83580 -1100 83720 -1060
rect 83580 -1160 83620 -1100
rect 83680 -1160 83720 -1100
rect 83580 -1200 83720 -1160
rect 83580 -1260 83620 -1200
rect 83680 -1260 83720 -1200
rect 83580 -1300 83720 -1260
rect 83580 -1360 83620 -1300
rect 83680 -1360 83720 -1300
rect 83580 -1380 83720 -1360
rect 83750 -1000 83890 -980
rect 83750 -1060 83790 -1000
rect 83850 -1060 83890 -1000
rect 83750 -1100 83890 -1060
rect 83750 -1160 83790 -1100
rect 83850 -1160 83890 -1100
rect 83750 -1200 83890 -1160
rect 83750 -1260 83790 -1200
rect 83850 -1260 83890 -1200
rect 83750 -1300 83890 -1260
rect 83750 -1360 83790 -1300
rect 83850 -1360 83890 -1300
rect 83750 -1380 83890 -1360
rect 83920 -1000 84060 -980
rect 83920 -1060 83960 -1000
rect 84020 -1060 84060 -1000
rect 83920 -1100 84060 -1060
rect 83920 -1160 83960 -1100
rect 84020 -1160 84060 -1100
rect 83920 -1200 84060 -1160
rect 83920 -1260 83960 -1200
rect 84020 -1260 84060 -1200
rect 83920 -1300 84060 -1260
rect 83920 -1360 83960 -1300
rect 84020 -1360 84060 -1300
rect 83920 -1380 84060 -1360
rect 84090 -1000 84230 -980
rect 84090 -1060 84130 -1000
rect 84190 -1060 84230 -1000
rect 84090 -1100 84230 -1060
rect 84090 -1160 84130 -1100
rect 84190 -1160 84230 -1100
rect 84090 -1200 84230 -1160
rect 84090 -1260 84130 -1200
rect 84190 -1260 84230 -1200
rect 84090 -1300 84230 -1260
rect 84090 -1360 84130 -1300
rect 84190 -1360 84230 -1300
rect 84090 -1380 84230 -1360
rect 84260 -1000 84400 -980
rect 84260 -1060 84300 -1000
rect 84360 -1060 84400 -1000
rect 84260 -1100 84400 -1060
rect 84260 -1160 84300 -1100
rect 84360 -1160 84400 -1100
rect 84260 -1200 84400 -1160
rect 84260 -1260 84300 -1200
rect 84360 -1260 84400 -1200
rect 84260 -1300 84400 -1260
rect 84260 -1360 84300 -1300
rect 84360 -1360 84400 -1300
rect 84260 -1380 84400 -1360
rect 84430 -1000 84570 -980
rect 84430 -1060 84470 -1000
rect 84530 -1060 84570 -1000
rect 84430 -1100 84570 -1060
rect 84430 -1160 84470 -1100
rect 84530 -1160 84570 -1100
rect 84430 -1200 84570 -1160
rect 84430 -1260 84470 -1200
rect 84530 -1260 84570 -1200
rect 84430 -1300 84570 -1260
rect 84430 -1360 84470 -1300
rect 84530 -1360 84570 -1300
rect 84430 -1380 84570 -1360
rect 84600 -1000 84740 -980
rect 84600 -1060 84640 -1000
rect 84700 -1060 84740 -1000
rect 84600 -1100 84740 -1060
rect 84600 -1160 84640 -1100
rect 84700 -1160 84740 -1100
rect 84600 -1200 84740 -1160
rect 84600 -1260 84640 -1200
rect 84700 -1260 84740 -1200
rect 84600 -1300 84740 -1260
rect 84600 -1360 84640 -1300
rect 84700 -1360 84740 -1300
rect 84600 -1380 84740 -1360
rect 84770 -1000 84910 -980
rect 84770 -1060 84810 -1000
rect 84870 -1060 84910 -1000
rect 84770 -1100 84910 -1060
rect 84770 -1160 84810 -1100
rect 84870 -1160 84910 -1100
rect 84770 -1200 84910 -1160
rect 84770 -1260 84810 -1200
rect 84870 -1260 84910 -1200
rect 84770 -1300 84910 -1260
rect 84770 -1360 84810 -1300
rect 84870 -1360 84910 -1300
rect 84770 -1380 84910 -1360
rect 84940 -1000 85080 -980
rect 84940 -1060 84980 -1000
rect 85040 -1060 85080 -1000
rect 84940 -1100 85080 -1060
rect 84940 -1160 84980 -1100
rect 85040 -1160 85080 -1100
rect 84940 -1200 85080 -1160
rect 84940 -1260 84980 -1200
rect 85040 -1260 85080 -1200
rect 84940 -1300 85080 -1260
rect 84940 -1360 84980 -1300
rect 85040 -1360 85080 -1300
rect 84940 -1380 85080 -1360
rect 85110 -1000 85250 -980
rect 85110 -1060 85150 -1000
rect 85210 -1060 85250 -1000
rect 85110 -1100 85250 -1060
rect 85110 -1160 85150 -1100
rect 85210 -1160 85250 -1100
rect 85110 -1200 85250 -1160
rect 85110 -1260 85150 -1200
rect 85210 -1260 85250 -1200
rect 85110 -1300 85250 -1260
rect 85110 -1360 85150 -1300
rect 85210 -1360 85250 -1300
rect 85110 -1380 85250 -1360
rect 85280 -1000 85420 -980
rect 85280 -1060 85320 -1000
rect 85380 -1060 85420 -1000
rect 85280 -1100 85420 -1060
rect 85280 -1160 85320 -1100
rect 85380 -1160 85420 -1100
rect 85280 -1200 85420 -1160
rect 85280 -1260 85320 -1200
rect 85380 -1260 85420 -1200
rect 85280 -1300 85420 -1260
rect 85280 -1360 85320 -1300
rect 85380 -1360 85420 -1300
rect 85280 -1380 85420 -1360
rect 85450 -1000 85590 -980
rect 85450 -1060 85490 -1000
rect 85550 -1060 85590 -1000
rect 85450 -1100 85590 -1060
rect 85450 -1160 85490 -1100
rect 85550 -1160 85590 -1100
rect 85450 -1200 85590 -1160
rect 85450 -1260 85490 -1200
rect 85550 -1260 85590 -1200
rect 85450 -1300 85590 -1260
rect 85450 -1360 85490 -1300
rect 85550 -1360 85590 -1300
rect 85450 -1380 85590 -1360
rect 85620 -1000 85760 -980
rect 85620 -1060 85660 -1000
rect 85720 -1060 85760 -1000
rect 85620 -1100 85760 -1060
rect 85620 -1160 85660 -1100
rect 85720 -1160 85760 -1100
rect 85620 -1200 85760 -1160
rect 85620 -1260 85660 -1200
rect 85720 -1260 85760 -1200
rect 85620 -1300 85760 -1260
rect 85620 -1360 85660 -1300
rect 85720 -1360 85760 -1300
rect 85620 -1380 85760 -1360
rect 85790 -1000 85930 -980
rect 85790 -1060 85830 -1000
rect 85890 -1060 85930 -1000
rect 85790 -1100 85930 -1060
rect 85790 -1160 85830 -1100
rect 85890 -1160 85930 -1100
rect 85790 -1200 85930 -1160
rect 85790 -1260 85830 -1200
rect 85890 -1260 85930 -1200
rect 85790 -1300 85930 -1260
rect 85790 -1360 85830 -1300
rect 85890 -1360 85930 -1300
rect 85790 -1380 85930 -1360
rect 85960 -1000 86100 -980
rect 85960 -1060 86000 -1000
rect 86060 -1060 86100 -1000
rect 85960 -1100 86100 -1060
rect 85960 -1160 86000 -1100
rect 86060 -1160 86100 -1100
rect 85960 -1200 86100 -1160
rect 85960 -1260 86000 -1200
rect 86060 -1260 86100 -1200
rect 85960 -1300 86100 -1260
rect 85960 -1360 86000 -1300
rect 86060 -1360 86100 -1300
rect 85960 -1380 86100 -1360
rect 86130 -1000 86270 -980
rect 86130 -1060 86170 -1000
rect 86230 -1060 86270 -1000
rect 86130 -1100 86270 -1060
rect 86130 -1160 86170 -1100
rect 86230 -1160 86270 -1100
rect 86130 -1200 86270 -1160
rect 86130 -1260 86170 -1200
rect 86230 -1260 86270 -1200
rect 86130 -1300 86270 -1260
rect 86130 -1360 86170 -1300
rect 86230 -1360 86270 -1300
rect 86130 -1380 86270 -1360
rect 86300 -1000 86440 -980
rect 86300 -1060 86340 -1000
rect 86400 -1060 86440 -1000
rect 86300 -1100 86440 -1060
rect 86300 -1160 86340 -1100
rect 86400 -1160 86440 -1100
rect 86300 -1200 86440 -1160
rect 86300 -1260 86340 -1200
rect 86400 -1260 86440 -1200
rect 86300 -1300 86440 -1260
rect 86300 -1360 86340 -1300
rect 86400 -1360 86440 -1300
rect 86300 -1380 86440 -1360
rect 86470 -1000 86610 -980
rect 86470 -1060 86510 -1000
rect 86570 -1060 86610 -1000
rect 86470 -1100 86610 -1060
rect 86470 -1160 86510 -1100
rect 86570 -1160 86610 -1100
rect 86470 -1200 86610 -1160
rect 86470 -1260 86510 -1200
rect 86570 -1260 86610 -1200
rect 86470 -1300 86610 -1260
rect 86470 -1360 86510 -1300
rect 86570 -1360 86610 -1300
rect 86470 -1380 86610 -1360
rect 86640 -1000 86780 -980
rect 86640 -1060 86680 -1000
rect 86740 -1060 86780 -1000
rect 86640 -1100 86780 -1060
rect 86640 -1160 86680 -1100
rect 86740 -1160 86780 -1100
rect 86640 -1200 86780 -1160
rect 86640 -1260 86680 -1200
rect 86740 -1260 86780 -1200
rect 86640 -1300 86780 -1260
rect 86640 -1360 86680 -1300
rect 86740 -1360 86780 -1300
rect 86640 -1380 86780 -1360
rect 86810 -1000 86950 -980
rect 86810 -1060 86850 -1000
rect 86910 -1060 86950 -1000
rect 86810 -1100 86950 -1060
rect 86810 -1160 86850 -1100
rect 86910 -1160 86950 -1100
rect 86810 -1200 86950 -1160
rect 86810 -1260 86850 -1200
rect 86910 -1260 86950 -1200
rect 86810 -1300 86950 -1260
rect 86810 -1360 86850 -1300
rect 86910 -1360 86950 -1300
rect 86810 -1380 86950 -1360
rect 86980 -1000 87120 -980
rect 86980 -1060 87020 -1000
rect 87080 -1060 87120 -1000
rect 86980 -1100 87120 -1060
rect 86980 -1160 87020 -1100
rect 87080 -1160 87120 -1100
rect 86980 -1200 87120 -1160
rect 86980 -1260 87020 -1200
rect 87080 -1260 87120 -1200
rect 86980 -1300 87120 -1260
rect 86980 -1360 87020 -1300
rect 87080 -1360 87120 -1300
rect 86980 -1380 87120 -1360
rect 87150 -1000 87290 -980
rect 87150 -1060 87190 -1000
rect 87250 -1060 87290 -1000
rect 87150 -1100 87290 -1060
rect 87150 -1160 87190 -1100
rect 87250 -1160 87290 -1100
rect 87150 -1200 87290 -1160
rect 87150 -1260 87190 -1200
rect 87250 -1260 87290 -1200
rect 87150 -1300 87290 -1260
rect 87150 -1360 87190 -1300
rect 87250 -1360 87290 -1300
rect 87150 -1380 87290 -1360
<< ndiffc >>
rect 543 935 577 995
rect 1311 935 1345 995
rect 5663 913 5697 973
rect 6431 913 6465 973
rect 450 20 510 80
rect 620 20 680 80
rect 790 20 850 80
rect 960 20 1020 80
rect 1130 20 1190 80
rect 1520 20 1580 80
rect 1690 20 1750 80
rect 1860 20 1920 80
rect 2030 20 2090 80
rect 2200 20 2260 80
rect 2370 20 2430 80
rect 2540 20 2600 80
rect 2710 20 2770 80
rect 2880 20 2940 80
rect 3050 20 3110 80
rect 3220 20 3280 80
rect 3390 20 3450 80
rect 3560 20 3620 80
rect 3730 20 3790 80
rect 3900 20 3960 80
rect 4070 20 4130 80
rect 4240 20 4300 80
rect 4540 20 4600 80
rect 4710 20 4770 80
rect 4880 20 4940 80
rect 5050 20 5110 80
rect 5220 20 5280 80
rect 5390 20 5450 80
rect 5560 20 5620 80
rect 5730 20 5790 80
rect 5900 20 5960 80
rect 6070 20 6130 80
rect 6240 20 6300 80
rect 6410 20 6470 80
rect 6580 20 6640 80
rect 6750 20 6810 80
rect 6920 20 6980 80
rect 7090 20 7150 80
rect 7260 20 7320 80
rect 7430 20 7490 80
rect 7600 20 7660 80
rect 7770 20 7830 80
rect 7940 20 8000 80
rect 8110 20 8170 80
rect 8280 20 8340 80
rect 8450 20 8510 80
rect 8620 20 8680 80
rect 8790 20 8850 80
rect 8960 20 9020 80
rect 9130 20 9190 80
rect 9300 20 9360 80
rect 9470 20 9530 80
rect 9640 20 9700 80
rect 9810 20 9870 80
rect 9980 20 10040 80
rect 10150 20 10210 80
rect 10320 20 10380 80
rect 10490 20 10550 80
rect 10660 20 10720 80
rect 10830 20 10890 80
rect 11000 20 11060 80
rect 11170 20 11230 80
rect 11340 20 11400 80
rect 11510 20 11570 80
rect 11680 20 11740 80
rect 11850 20 11910 80
rect 12020 20 12080 80
rect 12190 20 12250 80
rect 12360 20 12420 80
rect 12530 20 12590 80
rect 12700 20 12760 80
rect 12870 20 12930 80
rect 13040 20 13100 80
rect 13210 20 13270 80
rect 13380 20 13440 80
rect 13550 20 13610 80
rect 13720 20 13780 80
rect 13890 20 13950 80
rect 14060 20 14120 80
rect 14230 20 14290 80
rect 14400 20 14460 80
rect 14570 20 14630 80
rect 14740 20 14800 80
rect 14910 20 14970 80
rect 15080 20 15140 80
rect 15250 20 15310 80
rect 15420 20 15480 80
rect 15720 20 15780 80
rect 15890 20 15950 80
rect 16060 20 16120 80
rect 16230 20 16290 80
rect 16400 20 16460 80
rect 16570 20 16630 80
rect 16740 20 16800 80
rect 16910 20 16970 80
rect 17080 20 17140 80
rect 17250 20 17310 80
rect 17420 20 17480 80
rect 17590 20 17650 80
rect 17760 20 17820 80
rect 17930 20 17990 80
rect 18100 20 18160 80
rect 18270 20 18330 80
rect 18440 20 18500 80
rect 18610 20 18670 80
rect 18780 20 18840 80
rect 18950 20 19010 80
rect 19120 20 19180 80
rect 19290 20 19350 80
rect 19460 20 19520 80
rect 19630 20 19690 80
rect 19800 20 19860 80
rect 19970 20 20030 80
rect 20140 20 20200 80
rect 20310 20 20370 80
rect 20480 20 20540 80
rect 20650 20 20710 80
rect 20820 20 20880 80
rect 20990 20 21050 80
rect 21160 20 21220 80
rect 21330 20 21390 80
rect 21500 20 21560 80
rect 21670 20 21730 80
rect 21840 20 21900 80
rect 22010 20 22070 80
rect 22180 20 22240 80
rect 22350 20 22410 80
rect 22520 20 22580 80
rect 22690 20 22750 80
rect 22860 20 22920 80
rect 23030 20 23090 80
rect 23200 20 23260 80
rect 23370 20 23430 80
rect 23540 20 23600 80
rect 23710 20 23770 80
rect 23880 20 23940 80
rect 24050 20 24110 80
rect 24220 20 24280 80
rect 24390 20 24450 80
rect 24560 20 24620 80
rect 24730 20 24790 80
rect 24900 20 24960 80
rect 25070 20 25130 80
rect 25240 20 25300 80
rect 25410 20 25470 80
rect 25580 20 25640 80
rect 25750 20 25810 80
rect 25920 20 25980 80
rect 26090 20 26150 80
rect 26260 20 26320 80
rect 26430 20 26490 80
rect 26600 20 26660 80
rect 26770 20 26830 80
rect 26940 20 27000 80
rect 27110 20 27170 80
rect 27280 20 27340 80
rect 27450 20 27510 80
rect 27620 20 27680 80
rect 27790 20 27850 80
rect 27960 20 28020 80
rect 28130 20 28190 80
rect 28300 20 28360 80
rect 28470 20 28530 80
rect 28640 20 28700 80
rect 28810 20 28870 80
rect 28980 20 29040 80
rect 29150 20 29210 80
rect 29320 20 29380 80
rect 29490 20 29550 80
rect 29660 20 29720 80
rect 29830 20 29890 80
rect 30000 20 30060 80
rect 30170 20 30230 80
rect 30340 20 30400 80
rect 30510 20 30570 80
rect 30680 20 30740 80
rect 30850 20 30910 80
rect 31020 20 31080 80
rect 31190 20 31250 80
rect 31360 20 31420 80
rect 31530 20 31590 80
rect 31700 20 31760 80
rect 31870 20 31930 80
rect 32040 20 32100 80
rect 32210 20 32270 80
rect 32380 20 32440 80
rect 32550 20 32610 80
rect 32720 20 32780 80
rect 32890 20 32950 80
rect 33060 20 33120 80
rect 33230 20 33290 80
rect 33400 20 33460 80
rect 33570 20 33630 80
rect 33740 20 33800 80
rect 33910 20 33970 80
rect 34080 20 34140 80
rect 34250 20 34310 80
rect 34420 20 34480 80
rect 34590 20 34650 80
rect 34760 20 34820 80
rect 34930 20 34990 80
rect 35100 20 35160 80
rect 35270 20 35330 80
rect 35440 20 35500 80
rect 35610 20 35670 80
rect 35780 20 35840 80
rect 35950 20 36010 80
rect 36120 20 36180 80
rect 36290 20 36350 80
rect 36460 20 36520 80
rect 36630 20 36690 80
rect 36800 20 36860 80
rect 36970 20 37030 80
rect 37140 20 37200 80
rect 37310 20 37370 80
rect 37480 20 37540 80
rect 37650 20 37710 80
rect 37820 20 37880 80
rect 37990 20 38050 80
rect 38160 20 38220 80
rect 38330 20 38390 80
rect 38500 20 38560 80
rect 38670 20 38730 80
rect 38840 20 38900 80
rect 39010 20 39070 80
rect 39180 20 39240 80
rect 39350 20 39410 80
rect 39520 20 39580 80
rect 39690 20 39750 80
rect 39860 20 39920 80
rect 40030 20 40090 80
rect 40200 20 40260 80
rect 40370 20 40430 80
rect 40540 20 40600 80
rect 40710 20 40770 80
rect 40880 20 40940 80
rect 41050 20 41110 80
rect 41220 20 41280 80
rect 41390 20 41450 80
rect 41560 20 41620 80
rect 41730 20 41790 80
rect 41900 20 41960 80
rect 42070 20 42130 80
rect 42240 20 42300 80
rect 42410 20 42470 80
rect 42580 20 42640 80
rect 42750 20 42810 80
rect 42920 20 42980 80
rect 43090 20 43150 80
rect 43260 20 43320 80
rect 43430 20 43490 80
rect 43600 20 43660 80
rect 43770 20 43830 80
rect 43940 20 44000 80
rect 44110 20 44170 80
rect 44280 20 44340 80
rect 44450 20 44510 80
rect 44620 20 44680 80
rect 44790 20 44850 80
rect 44960 20 45020 80
rect 45130 20 45190 80
rect 45300 20 45360 80
rect 45470 20 45530 80
rect 45640 20 45700 80
rect 45810 20 45870 80
rect 45980 20 46040 80
rect 46150 20 46210 80
rect 46320 20 46380 80
rect 46490 20 46550 80
rect 46660 20 46720 80
rect 46830 20 46890 80
rect 47000 20 47060 80
rect 47170 20 47230 80
rect 47340 20 47400 80
rect 47510 20 47570 80
rect 47680 20 47740 80
rect 47850 20 47910 80
rect 48020 20 48080 80
rect 48190 20 48250 80
rect 48360 20 48420 80
rect 48530 20 48590 80
rect 48700 20 48760 80
rect 48870 20 48930 80
rect 49040 20 49100 80
rect 49210 20 49270 80
rect 49380 20 49440 80
rect 49550 20 49610 80
rect 49720 20 49780 80
rect 49890 20 49950 80
rect 50060 20 50120 80
rect 50230 20 50290 80
rect 50400 20 50460 80
rect 50570 20 50630 80
rect 50740 20 50800 80
rect 50910 20 50970 80
rect 51080 20 51140 80
rect 51250 20 51310 80
rect 51420 20 51480 80
rect 51590 20 51650 80
rect 51760 20 51820 80
rect 51930 20 51990 80
rect 52100 20 52160 80
rect 52270 20 52330 80
rect 52440 20 52500 80
rect 52610 20 52670 80
rect 52780 20 52840 80
rect 52950 20 53010 80
rect 53120 20 53180 80
rect 53290 20 53350 80
rect 53460 20 53520 80
rect 53630 20 53690 80
rect 53800 20 53860 80
rect 53970 20 54030 80
rect 54140 20 54200 80
rect 54310 20 54370 80
rect 54480 20 54540 80
rect 54650 20 54710 80
rect 54820 20 54880 80
rect 54990 20 55050 80
rect 55160 20 55220 80
rect 55330 20 55390 80
rect 55500 20 55560 80
rect 55670 20 55730 80
rect 55840 20 55900 80
rect 56010 20 56070 80
rect 56180 20 56240 80
rect 56350 20 56410 80
rect 56520 20 56580 80
rect 56690 20 56750 80
rect 56860 20 56920 80
rect 57030 20 57090 80
rect 57200 20 57260 80
rect 57370 20 57430 80
rect 57540 20 57600 80
rect 57710 20 57770 80
rect 57880 20 57940 80
rect 58050 20 58110 80
rect 58220 20 58280 80
rect 58390 20 58450 80
rect 58560 20 58620 80
rect 58730 20 58790 80
rect 58900 20 58960 80
rect 59070 20 59130 80
rect 59240 20 59300 80
rect 30 -120 90 -60
rect 200 -120 260 -60
rect 150 -730 210 -670
rect 150 -830 210 -770
rect 320 -730 380 -670
rect 320 -830 380 -770
rect 490 -730 550 -670
rect 490 -830 550 -770
rect 660 -730 720 -670
rect 660 -830 720 -770
rect 830 -730 890 -670
rect 830 -830 890 -770
rect 1000 -730 1060 -670
rect 1000 -830 1060 -770
rect 1170 -730 1230 -670
rect 1170 -830 1230 -770
rect 1340 -730 1400 -670
rect 1340 -830 1400 -770
rect 1510 -730 1570 -670
rect 1510 -830 1570 -770
rect 1680 -730 1740 -670
rect 1680 -830 1740 -770
rect 1850 -730 1910 -670
rect 1850 -830 1910 -770
rect 2020 -730 2080 -670
rect 2020 -830 2080 -770
rect 2190 -730 2250 -670
rect 2190 -830 2250 -770
rect 2360 -730 2420 -670
rect 2360 -830 2420 -770
rect 2530 -730 2590 -670
rect 2530 -830 2590 -770
rect 2700 -730 2760 -670
rect 2700 -830 2760 -770
rect 2870 -730 2930 -670
rect 2870 -830 2930 -770
rect 3040 -730 3100 -670
rect 3040 -830 3100 -770
rect 3210 -730 3270 -670
rect 3210 -830 3270 -770
rect 3380 -730 3440 -670
rect 3380 -830 3440 -770
rect 3550 -730 3610 -670
rect 3550 -830 3610 -770
rect 3720 -730 3780 -670
rect 3720 -830 3780 -770
rect 3890 -730 3950 -670
rect 3890 -830 3950 -770
rect 4060 -730 4120 -670
rect 4060 -830 4120 -770
rect 4230 -730 4290 -670
rect 4230 -830 4290 -770
rect 4400 -730 4460 -670
rect 4400 -830 4460 -770
rect 4570 -730 4630 -670
rect 4570 -830 4630 -770
rect 4740 -730 4800 -670
rect 4740 -830 4800 -770
rect 4910 -730 4970 -670
rect 4910 -830 4970 -770
rect 5080 -730 5140 -670
rect 5080 -830 5140 -770
rect 5250 -730 5310 -670
rect 5250 -830 5310 -770
rect 5420 -730 5480 -670
rect 5420 -830 5480 -770
rect 5590 -730 5650 -670
rect 5590 -830 5650 -770
rect 5760 -730 5820 -670
rect 5760 -830 5820 -770
rect 5930 -730 5990 -670
rect 5930 -830 5990 -770
rect 6100 -730 6160 -670
rect 6100 -830 6160 -770
rect 6270 -730 6330 -670
rect 6270 -830 6330 -770
rect 6440 -730 6500 -670
rect 6440 -830 6500 -770
rect 6610 -730 6670 -670
rect 6610 -830 6670 -770
rect 6780 -730 6840 -670
rect 6780 -830 6840 -770
rect 6950 -730 7010 -670
rect 6950 -830 7010 -770
rect 7120 -730 7180 -670
rect 7120 -830 7180 -770
rect 7290 -730 7350 -670
rect 7290 -830 7350 -770
rect 7460 -730 7520 -670
rect 7460 -830 7520 -770
rect 7630 -730 7690 -670
rect 7630 -830 7690 -770
rect 7800 -730 7860 -670
rect 7800 -830 7860 -770
rect 7970 -730 8030 -670
rect 7970 -830 8030 -770
rect 8140 -730 8200 -670
rect 8140 -830 8200 -770
rect 8310 -730 8370 -670
rect 8310 -830 8370 -770
rect 8480 -730 8540 -670
rect 8480 -830 8540 -770
rect 8650 -730 8710 -670
rect 8650 -830 8710 -770
rect 8820 -730 8880 -670
rect 8820 -830 8880 -770
rect 8990 -730 9050 -670
rect 8990 -830 9050 -770
rect 9160 -730 9220 -670
rect 9160 -830 9220 -770
rect 9330 -730 9390 -670
rect 9330 -830 9390 -770
rect 9500 -730 9560 -670
rect 9500 -830 9560 -770
rect 9670 -730 9730 -670
rect 9670 -830 9730 -770
rect 9840 -730 9900 -670
rect 9840 -830 9900 -770
rect 10010 -730 10070 -670
rect 10010 -830 10070 -770
rect 10180 -730 10240 -670
rect 10180 -830 10240 -770
rect 10350 -730 10410 -670
rect 10350 -830 10410 -770
rect 10520 -730 10580 -670
rect 10520 -830 10580 -770
rect 10690 -730 10750 -670
rect 10690 -830 10750 -770
rect 10860 -730 10920 -670
rect 10860 -830 10920 -770
rect 11030 -730 11090 -670
rect 11030 -830 11090 -770
rect 11200 -730 11260 -670
rect 11200 -830 11260 -770
rect 11370 -730 11430 -670
rect 11370 -830 11430 -770
rect 11540 -730 11600 -670
rect 11540 -830 11600 -770
rect 11710 -730 11770 -670
rect 11710 -830 11770 -770
rect 11880 -730 11940 -670
rect 11880 -830 11940 -770
rect 12050 -730 12110 -670
rect 12050 -830 12110 -770
rect 12220 -730 12280 -670
rect 12220 -830 12280 -770
rect 12390 -730 12450 -670
rect 12390 -830 12450 -770
rect 12560 -730 12620 -670
rect 12560 -830 12620 -770
rect 12730 -730 12790 -670
rect 12730 -830 12790 -770
rect 12900 -730 12960 -670
rect 12900 -830 12960 -770
rect 13070 -730 13130 -670
rect 13070 -830 13130 -770
rect 13240 -730 13300 -670
rect 13240 -830 13300 -770
rect 13410 -730 13470 -670
rect 13410 -830 13470 -770
rect 13580 -730 13640 -670
rect 13580 -830 13640 -770
rect 13750 -730 13810 -670
rect 13750 -830 13810 -770
rect 13920 -730 13980 -670
rect 13920 -830 13980 -770
rect 14090 -730 14150 -670
rect 14090 -830 14150 -770
rect 14260 -730 14320 -670
rect 14260 -830 14320 -770
rect 14430 -730 14490 -670
rect 14430 -830 14490 -770
rect 14600 -730 14660 -670
rect 14600 -830 14660 -770
rect 14770 -730 14830 -670
rect 14770 -830 14830 -770
rect 14940 -730 15000 -670
rect 14940 -830 15000 -770
rect 15110 -730 15170 -670
rect 15110 -830 15170 -770
rect 15280 -730 15340 -670
rect 15280 -830 15340 -770
rect 15450 -730 15510 -670
rect 15450 -830 15510 -770
rect 15620 -730 15680 -670
rect 15620 -830 15680 -770
rect 15790 -730 15850 -670
rect 15790 -830 15850 -770
rect 15960 -730 16020 -670
rect 15960 -830 16020 -770
rect 16130 -730 16190 -670
rect 16130 -830 16190 -770
rect 16300 -730 16360 -670
rect 16300 -830 16360 -770
rect 16470 -730 16530 -670
rect 16470 -830 16530 -770
rect 16640 -730 16700 -670
rect 16640 -830 16700 -770
rect 16810 -730 16870 -670
rect 16810 -830 16870 -770
rect 16980 -730 17040 -670
rect 16980 -830 17040 -770
rect 17150 -730 17210 -670
rect 17150 -830 17210 -770
rect 17320 -730 17380 -670
rect 17320 -830 17380 -770
rect 17490 -730 17550 -670
rect 17490 -830 17550 -770
rect 17660 -730 17720 -670
rect 17660 -830 17720 -770
rect 17830 -730 17890 -670
rect 17830 -830 17890 -770
rect 18000 -730 18060 -670
rect 18000 -830 18060 -770
rect 18170 -730 18230 -670
rect 18170 -830 18230 -770
rect 18340 -730 18400 -670
rect 18340 -830 18400 -770
rect 18510 -730 18570 -670
rect 18510 -830 18570 -770
rect 18680 -730 18740 -670
rect 18680 -830 18740 -770
rect 18850 -730 18910 -670
rect 18850 -830 18910 -770
rect 19020 -730 19080 -670
rect 19020 -830 19080 -770
rect 19190 -730 19250 -670
rect 19190 -830 19250 -770
rect 19360 -730 19420 -670
rect 19360 -830 19420 -770
rect 19530 -730 19590 -670
rect 19530 -830 19590 -770
rect 19700 -730 19760 -670
rect 19700 -830 19760 -770
rect 19870 -730 19930 -670
rect 19870 -830 19930 -770
rect 20040 -730 20100 -670
rect 20040 -830 20100 -770
rect 20210 -730 20270 -670
rect 20210 -830 20270 -770
rect 20380 -730 20440 -670
rect 20380 -830 20440 -770
rect 20550 -730 20610 -670
rect 20550 -830 20610 -770
rect 20720 -730 20780 -670
rect 20720 -830 20780 -770
rect 20890 -730 20950 -670
rect 20890 -830 20950 -770
rect 21060 -730 21120 -670
rect 21060 -830 21120 -770
rect 21230 -730 21290 -670
rect 21230 -830 21290 -770
rect 21400 -730 21460 -670
rect 21400 -830 21460 -770
rect 21570 -730 21630 -670
rect 21570 -830 21630 -770
rect 21740 -730 21800 -670
rect 21740 -830 21800 -770
rect 21910 -730 21970 -670
rect 21910 -830 21970 -770
rect 22080 -730 22140 -670
rect 22080 -830 22140 -770
rect 22250 -730 22310 -670
rect 22250 -830 22310 -770
rect 22420 -730 22480 -670
rect 22420 -830 22480 -770
rect 22590 -730 22650 -670
rect 22590 -830 22650 -770
rect 22760 -730 22820 -670
rect 22760 -830 22820 -770
rect 22930 -730 22990 -670
rect 22930 -830 22990 -770
rect 23100 -730 23160 -670
rect 23100 -830 23160 -770
rect 23270 -730 23330 -670
rect 23270 -830 23330 -770
rect 23440 -730 23500 -670
rect 23440 -830 23500 -770
rect 23610 -730 23670 -670
rect 23610 -830 23670 -770
rect 23780 -730 23840 -670
rect 23780 -830 23840 -770
rect 23950 -730 24010 -670
rect 23950 -830 24010 -770
rect 24120 -730 24180 -670
rect 24120 -830 24180 -770
rect 24290 -730 24350 -670
rect 24290 -830 24350 -770
rect 24460 -730 24520 -670
rect 24460 -830 24520 -770
rect 24630 -730 24690 -670
rect 24630 -830 24690 -770
rect 24800 -730 24860 -670
rect 24800 -830 24860 -770
rect 24970 -730 25030 -670
rect 24970 -830 25030 -770
rect 25140 -730 25200 -670
rect 25140 -830 25200 -770
rect 25310 -730 25370 -670
rect 25310 -830 25370 -770
rect 25480 -730 25540 -670
rect 25480 -830 25540 -770
rect 25650 -730 25710 -670
rect 25650 -830 25710 -770
rect 25820 -730 25880 -670
rect 25820 -830 25880 -770
rect 25990 -730 26050 -670
rect 25990 -830 26050 -770
rect 26160 -730 26220 -670
rect 26160 -830 26220 -770
rect 26330 -730 26390 -670
rect 26330 -830 26390 -770
rect 26500 -730 26560 -670
rect 26500 -830 26560 -770
rect 26670 -730 26730 -670
rect 26670 -830 26730 -770
rect 26840 -730 26900 -670
rect 26840 -830 26900 -770
rect 27010 -730 27070 -670
rect 27010 -830 27070 -770
rect 27180 -730 27240 -670
rect 27180 -830 27240 -770
rect 27350 -730 27410 -670
rect 27350 -830 27410 -770
rect 27520 -730 27580 -670
rect 27520 -830 27580 -770
rect 27690 -730 27750 -670
rect 27690 -830 27750 -770
rect 27860 -730 27920 -670
rect 27860 -830 27920 -770
rect 28030 -730 28090 -670
rect 28030 -830 28090 -770
rect 28200 -730 28260 -670
rect 28200 -830 28260 -770
rect 28370 -730 28430 -670
rect 28370 -830 28430 -770
rect 28540 -730 28600 -670
rect 28540 -830 28600 -770
rect 28710 -730 28770 -670
rect 28710 -830 28770 -770
rect 28880 -730 28940 -670
rect 28880 -830 28940 -770
rect 29050 -730 29110 -670
rect 29050 -830 29110 -770
rect 29220 -730 29280 -670
rect 29220 -830 29280 -770
rect 29390 -730 29450 -670
rect 29390 -830 29450 -770
rect 29560 -730 29620 -670
rect 29560 -830 29620 -770
rect 29730 -730 29790 -670
rect 29730 -830 29790 -770
rect 29900 -730 29960 -670
rect 29900 -830 29960 -770
rect 30070 -730 30130 -670
rect 30070 -830 30130 -770
rect 30240 -730 30300 -670
rect 30240 -830 30300 -770
rect 30410 -730 30470 -670
rect 30410 -830 30470 -770
rect 30580 -730 30640 -670
rect 30580 -830 30640 -770
rect 30750 -730 30810 -670
rect 30750 -830 30810 -770
rect 30920 -730 30980 -670
rect 30920 -830 30980 -770
rect 31090 -730 31150 -670
rect 31090 -830 31150 -770
rect 31260 -730 31320 -670
rect 31260 -830 31320 -770
rect 31430 -730 31490 -670
rect 31430 -830 31490 -770
rect 31600 -730 31660 -670
rect 31600 -830 31660 -770
rect 31770 -730 31830 -670
rect 31770 -830 31830 -770
rect 31940 -730 32000 -670
rect 31940 -830 32000 -770
rect 32110 -730 32170 -670
rect 32110 -830 32170 -770
rect 32280 -730 32340 -670
rect 32280 -830 32340 -770
rect 32450 -730 32510 -670
rect 32450 -830 32510 -770
rect 32620 -730 32680 -670
rect 32620 -830 32680 -770
rect 32790 -730 32850 -670
rect 32790 -830 32850 -770
rect 32960 -730 33020 -670
rect 32960 -830 33020 -770
rect 33130 -730 33190 -670
rect 33130 -830 33190 -770
rect 33300 -730 33360 -670
rect 33300 -830 33360 -770
rect 33470 -730 33530 -670
rect 33470 -830 33530 -770
rect 33640 -730 33700 -670
rect 33640 -830 33700 -770
rect 33810 -730 33870 -670
rect 33810 -830 33870 -770
rect 33980 -730 34040 -670
rect 33980 -830 34040 -770
rect 34150 -730 34210 -670
rect 34150 -830 34210 -770
rect 34320 -730 34380 -670
rect 34320 -830 34380 -770
rect 34490 -730 34550 -670
rect 34490 -830 34550 -770
rect 34660 -730 34720 -670
rect 34660 -830 34720 -770
rect 34830 -730 34890 -670
rect 34830 -830 34890 -770
rect 35000 -730 35060 -670
rect 35000 -830 35060 -770
rect 35170 -730 35230 -670
rect 35170 -830 35230 -770
rect 35340 -730 35400 -670
rect 35340 -830 35400 -770
rect 35510 -730 35570 -670
rect 35510 -830 35570 -770
rect 35680 -730 35740 -670
rect 35680 -830 35740 -770
rect 35850 -730 35910 -670
rect 35850 -830 35910 -770
rect 36020 -730 36080 -670
rect 36020 -830 36080 -770
rect 36190 -730 36250 -670
rect 36190 -830 36250 -770
rect 36360 -730 36420 -670
rect 36360 -830 36420 -770
rect 36530 -730 36590 -670
rect 36530 -830 36590 -770
rect 36700 -730 36760 -670
rect 36700 -830 36760 -770
rect 36870 -730 36930 -670
rect 36870 -830 36930 -770
rect 37040 -730 37100 -670
rect 37040 -830 37100 -770
rect 37210 -730 37270 -670
rect 37210 -830 37270 -770
rect 37380 -730 37440 -670
rect 37380 -830 37440 -770
rect 37550 -730 37610 -670
rect 37550 -830 37610 -770
rect 37720 -730 37780 -670
rect 37720 -830 37780 -770
rect 37890 -730 37950 -670
rect 37890 -830 37950 -770
rect 38060 -730 38120 -670
rect 38060 -830 38120 -770
rect 38230 -730 38290 -670
rect 38230 -830 38290 -770
rect 38400 -730 38460 -670
rect 38400 -830 38460 -770
rect 38570 -730 38630 -670
rect 38570 -830 38630 -770
rect 38740 -730 38800 -670
rect 38740 -830 38800 -770
rect 38910 -730 38970 -670
rect 38910 -830 38970 -770
rect 39080 -730 39140 -670
rect 39080 -830 39140 -770
rect 39250 -730 39310 -670
rect 39250 -830 39310 -770
rect 39420 -730 39480 -670
rect 39420 -830 39480 -770
rect 39590 -730 39650 -670
rect 39590 -830 39650 -770
rect 39760 -730 39820 -670
rect 39760 -830 39820 -770
rect 39930 -730 39990 -670
rect 39930 -830 39990 -770
rect 40100 -730 40160 -670
rect 40100 -830 40160 -770
rect 40270 -730 40330 -670
rect 40270 -830 40330 -770
rect 40440 -730 40500 -670
rect 40440 -830 40500 -770
rect 40610 -730 40670 -670
rect 40610 -830 40670 -770
rect 40780 -730 40840 -670
rect 40780 -830 40840 -770
rect 40950 -730 41010 -670
rect 40950 -830 41010 -770
rect 41120 -730 41180 -670
rect 41120 -830 41180 -770
rect 41290 -730 41350 -670
rect 41290 -830 41350 -770
rect 41460 -730 41520 -670
rect 41460 -830 41520 -770
rect 41630 -730 41690 -670
rect 41630 -830 41690 -770
rect 41800 -730 41860 -670
rect 41800 -830 41860 -770
rect 41970 -730 42030 -670
rect 41970 -830 42030 -770
rect 42140 -730 42200 -670
rect 42140 -830 42200 -770
rect 42310 -730 42370 -670
rect 42310 -830 42370 -770
rect 42480 -730 42540 -670
rect 42480 -830 42540 -770
rect 42650 -730 42710 -670
rect 42650 -830 42710 -770
rect 42820 -730 42880 -670
rect 42820 -830 42880 -770
rect 42990 -730 43050 -670
rect 42990 -830 43050 -770
rect 43160 -730 43220 -670
rect 43160 -830 43220 -770
rect 43330 -730 43390 -670
rect 43330 -830 43390 -770
rect 43500 -730 43560 -670
rect 43500 -830 43560 -770
rect 43670 -730 43730 -670
rect 43670 -830 43730 -770
rect 43840 -730 43900 -670
rect 43840 -830 43900 -770
rect 44010 -730 44070 -670
rect 44010 -830 44070 -770
rect 44180 -730 44240 -670
rect 44180 -830 44240 -770
rect 44350 -730 44410 -670
rect 44350 -830 44410 -770
rect 44520 -730 44580 -670
rect 44520 -830 44580 -770
rect 44690 -730 44750 -670
rect 44690 -830 44750 -770
rect 44860 -730 44920 -670
rect 44860 -830 44920 -770
rect 45030 -730 45090 -670
rect 45030 -830 45090 -770
rect 45200 -730 45260 -670
rect 45200 -830 45260 -770
rect 45370 -730 45430 -670
rect 45370 -830 45430 -770
rect 45540 -730 45600 -670
rect 45540 -830 45600 -770
rect 45710 -730 45770 -670
rect 45710 -830 45770 -770
rect 45880 -730 45940 -670
rect 45880 -830 45940 -770
rect 46050 -730 46110 -670
rect 46050 -830 46110 -770
rect 46220 -730 46280 -670
rect 46220 -830 46280 -770
rect 46390 -730 46450 -670
rect 46390 -830 46450 -770
rect 46560 -730 46620 -670
rect 46560 -830 46620 -770
rect 46730 -730 46790 -670
rect 46730 -830 46790 -770
rect 46900 -730 46960 -670
rect 46900 -830 46960 -770
rect 47070 -730 47130 -670
rect 47070 -830 47130 -770
rect 47240 -730 47300 -670
rect 47240 -830 47300 -770
rect 47410 -730 47470 -670
rect 47410 -830 47470 -770
rect 47580 -730 47640 -670
rect 47580 -830 47640 -770
rect 47750 -730 47810 -670
rect 47750 -830 47810 -770
rect 47920 -730 47980 -670
rect 47920 -830 47980 -770
rect 48090 -730 48150 -670
rect 48090 -830 48150 -770
rect 48260 -730 48320 -670
rect 48260 -830 48320 -770
rect 48430 -730 48490 -670
rect 48430 -830 48490 -770
rect 48600 -730 48660 -670
rect 48600 -830 48660 -770
rect 48770 -730 48830 -670
rect 48770 -830 48830 -770
rect 48940 -730 49000 -670
rect 48940 -830 49000 -770
rect 49110 -730 49170 -670
rect 49110 -830 49170 -770
rect 49280 -730 49340 -670
rect 49280 -830 49340 -770
rect 49450 -730 49510 -670
rect 49450 -830 49510 -770
rect 49620 -730 49680 -670
rect 49620 -830 49680 -770
rect 49790 -730 49850 -670
rect 49790 -830 49850 -770
rect 49960 -730 50020 -670
rect 49960 -830 50020 -770
rect 50130 -730 50190 -670
rect 50130 -830 50190 -770
rect 50300 -730 50360 -670
rect 50300 -830 50360 -770
rect 50470 -730 50530 -670
rect 50470 -830 50530 -770
rect 50640 -730 50700 -670
rect 50640 -830 50700 -770
rect 50810 -730 50870 -670
rect 50810 -830 50870 -770
rect 50980 -730 51040 -670
rect 50980 -830 51040 -770
rect 51150 -730 51210 -670
rect 51150 -830 51210 -770
rect 51320 -730 51380 -670
rect 51320 -830 51380 -770
rect 51490 -730 51550 -670
rect 51490 -830 51550 -770
rect 51660 -730 51720 -670
rect 51660 -830 51720 -770
rect 51830 -730 51890 -670
rect 51830 -830 51890 -770
rect 52000 -730 52060 -670
rect 52000 -830 52060 -770
rect 52170 -730 52230 -670
rect 52170 -830 52230 -770
rect 52340 -730 52400 -670
rect 52340 -830 52400 -770
rect 52510 -730 52570 -670
rect 52510 -830 52570 -770
rect 52680 -730 52740 -670
rect 52680 -830 52740 -770
rect 52850 -730 52910 -670
rect 52850 -830 52910 -770
rect 53020 -730 53080 -670
rect 53020 -830 53080 -770
rect 53190 -730 53250 -670
rect 53190 -830 53250 -770
rect 53360 -730 53420 -670
rect 53360 -830 53420 -770
rect 53530 -730 53590 -670
rect 53530 -830 53590 -770
rect 53700 -730 53760 -670
rect 53700 -830 53760 -770
rect 53870 -730 53930 -670
rect 53870 -830 53930 -770
rect 54040 -730 54100 -670
rect 54040 -830 54100 -770
rect 54210 -730 54270 -670
rect 54210 -830 54270 -770
rect 54380 -730 54440 -670
rect 54380 -830 54440 -770
rect 54550 -730 54610 -670
rect 54550 -830 54610 -770
rect 54720 -730 54780 -670
rect 54720 -830 54780 -770
rect 54890 -730 54950 -670
rect 54890 -830 54950 -770
rect 55060 -730 55120 -670
rect 55060 -830 55120 -770
rect 55230 -730 55290 -670
rect 55230 -830 55290 -770
rect 55400 -730 55460 -670
rect 55400 -830 55460 -770
rect 55570 -730 55630 -670
rect 55570 -830 55630 -770
rect 55740 -730 55800 -670
rect 55740 -830 55800 -770
rect 55910 -730 55970 -670
rect 55910 -830 55970 -770
rect 56080 -730 56140 -670
rect 56080 -830 56140 -770
rect 56250 -730 56310 -670
rect 56250 -830 56310 -770
rect 56420 -730 56480 -670
rect 56420 -830 56480 -770
rect 56590 -730 56650 -670
rect 56590 -830 56650 -770
rect 56760 -730 56820 -670
rect 56760 -830 56820 -770
rect 56930 -730 56990 -670
rect 56930 -830 56990 -770
rect 57100 -730 57160 -670
rect 57100 -830 57160 -770
rect 57270 -730 57330 -670
rect 57270 -830 57330 -770
rect 57440 -730 57500 -670
rect 57440 -830 57500 -770
rect 57610 -730 57670 -670
rect 57610 -830 57670 -770
rect 57780 -730 57840 -670
rect 57780 -830 57840 -770
rect 57950 -730 58010 -670
rect 57950 -830 58010 -770
rect 58120 -730 58180 -670
rect 58120 -830 58180 -770
rect 58290 -730 58350 -670
rect 58290 -830 58350 -770
rect 58460 -730 58520 -670
rect 58460 -830 58520 -770
rect 58630 -730 58690 -670
rect 58630 -830 58690 -770
rect 58800 -730 58860 -670
rect 58800 -830 58860 -770
rect 58970 -730 59030 -670
rect 58970 -830 59030 -770
rect 59140 -730 59200 -670
rect 59140 -830 59200 -770
rect 59310 -730 59370 -670
rect 59310 -830 59370 -770
rect 59480 -730 59540 -670
rect 59480 -830 59540 -770
rect 59650 -730 59710 -670
rect 59650 -830 59710 -770
rect 59820 -730 59880 -670
rect 59820 -830 59880 -770
rect 59990 -730 60050 -670
rect 59990 -830 60050 -770
rect 60160 -730 60220 -670
rect 60160 -830 60220 -770
rect 60330 -730 60390 -670
rect 60330 -830 60390 -770
rect 60500 -730 60560 -670
rect 60500 -830 60560 -770
rect 60670 -730 60730 -670
rect 60670 -830 60730 -770
rect 60840 -730 60900 -670
rect 60840 -830 60900 -770
rect 61010 -730 61070 -670
rect 61010 -830 61070 -770
rect 61180 -730 61240 -670
rect 61180 -830 61240 -770
rect 61350 -730 61410 -670
rect 61350 -830 61410 -770
rect 61520 -730 61580 -670
rect 61520 -830 61580 -770
rect 61690 -730 61750 -670
rect 61690 -830 61750 -770
rect 61860 -730 61920 -670
rect 61860 -830 61920 -770
rect 62030 -730 62090 -670
rect 62030 -830 62090 -770
rect 62200 -730 62260 -670
rect 62200 -830 62260 -770
rect 62370 -730 62430 -670
rect 62370 -830 62430 -770
rect 62540 -730 62600 -670
rect 62540 -830 62600 -770
rect 62710 -730 62770 -670
rect 62710 -830 62770 -770
rect 62880 -730 62940 -670
rect 62880 -830 62940 -770
rect 63050 -730 63110 -670
rect 63050 -830 63110 -770
rect 63220 -730 63280 -670
rect 63220 -830 63280 -770
rect 63390 -730 63450 -670
rect 63390 -830 63450 -770
rect 63560 -730 63620 -670
rect 63560 -830 63620 -770
rect 63730 -730 63790 -670
rect 63730 -830 63790 -770
rect 63900 -730 63960 -670
rect 63900 -830 63960 -770
rect 64070 -730 64130 -670
rect 64070 -830 64130 -770
rect 64240 -730 64300 -670
rect 64240 -830 64300 -770
rect 64410 -730 64470 -670
rect 64410 -830 64470 -770
rect 64580 -730 64640 -670
rect 64580 -830 64640 -770
rect 64750 -730 64810 -670
rect 64750 -830 64810 -770
rect 64920 -730 64980 -670
rect 64920 -830 64980 -770
rect 65090 -730 65150 -670
rect 65090 -830 65150 -770
rect 65260 -730 65320 -670
rect 65260 -830 65320 -770
rect 65430 -730 65490 -670
rect 65430 -830 65490 -770
rect 65600 -730 65660 -670
rect 65600 -830 65660 -770
rect 65770 -730 65830 -670
rect 65770 -830 65830 -770
rect 65940 -730 66000 -670
rect 65940 -830 66000 -770
rect 66110 -730 66170 -670
rect 66110 -830 66170 -770
rect 66280 -730 66340 -670
rect 66280 -830 66340 -770
rect 66450 -730 66510 -670
rect 66450 -830 66510 -770
rect 66620 -730 66680 -670
rect 66620 -830 66680 -770
rect 66790 -730 66850 -670
rect 66790 -830 66850 -770
rect 66960 -730 67020 -670
rect 66960 -830 67020 -770
rect 67130 -730 67190 -670
rect 67130 -830 67190 -770
rect 67300 -730 67360 -670
rect 67300 -830 67360 -770
rect 67470 -730 67530 -670
rect 67470 -830 67530 -770
rect 67640 -730 67700 -670
rect 67640 -830 67700 -770
rect 67810 -730 67870 -670
rect 67810 -830 67870 -770
rect 67980 -730 68040 -670
rect 67980 -830 68040 -770
rect 68150 -730 68210 -670
rect 68150 -830 68210 -770
rect 68320 -730 68380 -670
rect 68320 -830 68380 -770
rect 68490 -730 68550 -670
rect 68490 -830 68550 -770
rect 68660 -730 68720 -670
rect 68660 -830 68720 -770
rect 68830 -730 68890 -670
rect 68830 -830 68890 -770
rect 69000 -730 69060 -670
rect 69000 -830 69060 -770
rect 69170 -730 69230 -670
rect 69170 -830 69230 -770
rect 69340 -730 69400 -670
rect 69340 -830 69400 -770
rect 69510 -730 69570 -670
rect 69510 -830 69570 -770
rect 69680 -730 69740 -670
rect 69680 -830 69740 -770
rect 69850 -730 69910 -670
rect 69850 -830 69910 -770
rect 70020 -730 70080 -670
rect 70020 -830 70080 -770
rect 70190 -730 70250 -670
rect 70190 -830 70250 -770
rect 70360 -730 70420 -670
rect 70360 -830 70420 -770
rect 70530 -730 70590 -670
rect 70530 -830 70590 -770
rect 70700 -730 70760 -670
rect 70700 -830 70760 -770
rect 70870 -730 70930 -670
rect 70870 -830 70930 -770
rect 71040 -730 71100 -670
rect 71040 -830 71100 -770
rect 71210 -730 71270 -670
rect 71210 -830 71270 -770
rect 71380 -730 71440 -670
rect 71380 -830 71440 -770
rect 71550 -730 71610 -670
rect 71550 -830 71610 -770
rect 71720 -730 71780 -670
rect 71720 -830 71780 -770
rect 71890 -730 71950 -670
rect 71890 -830 71950 -770
rect 72060 -730 72120 -670
rect 72060 -830 72120 -770
rect 72230 -730 72290 -670
rect 72230 -830 72290 -770
rect 72400 -730 72460 -670
rect 72400 -830 72460 -770
rect 72570 -730 72630 -670
rect 72570 -830 72630 -770
rect 72740 -730 72800 -670
rect 72740 -830 72800 -770
rect 72910 -730 72970 -670
rect 72910 -830 72970 -770
rect 73080 -730 73140 -670
rect 73080 -830 73140 -770
rect 73250 -730 73310 -670
rect 73250 -830 73310 -770
rect 73420 -730 73480 -670
rect 73420 -830 73480 -770
rect 73590 -730 73650 -670
rect 73590 -830 73650 -770
rect 73760 -730 73820 -670
rect 73760 -830 73820 -770
rect 73930 -730 73990 -670
rect 73930 -830 73990 -770
rect 74100 -730 74160 -670
rect 74100 -830 74160 -770
rect 74270 -730 74330 -670
rect 74270 -830 74330 -770
rect 74440 -730 74500 -670
rect 74440 -830 74500 -770
rect 74610 -730 74670 -670
rect 74610 -830 74670 -770
rect 74780 -730 74840 -670
rect 74780 -830 74840 -770
rect 74950 -730 75010 -670
rect 74950 -830 75010 -770
rect 75120 -730 75180 -670
rect 75120 -830 75180 -770
rect 75290 -730 75350 -670
rect 75290 -830 75350 -770
rect 75460 -730 75520 -670
rect 75460 -830 75520 -770
rect 75630 -730 75690 -670
rect 75630 -830 75690 -770
rect 75800 -730 75860 -670
rect 75800 -830 75860 -770
rect 75970 -730 76030 -670
rect 75970 -830 76030 -770
rect 76140 -730 76200 -670
rect 76140 -830 76200 -770
rect 76310 -730 76370 -670
rect 76310 -830 76370 -770
rect 76480 -730 76540 -670
rect 76480 -830 76540 -770
rect 76650 -730 76710 -670
rect 76650 -830 76710 -770
rect 76820 -730 76880 -670
rect 76820 -830 76880 -770
rect 76990 -730 77050 -670
rect 76990 -830 77050 -770
rect 77160 -730 77220 -670
rect 77160 -830 77220 -770
rect 77330 -730 77390 -670
rect 77330 -830 77390 -770
rect 77500 -730 77560 -670
rect 77500 -830 77560 -770
rect 77670 -730 77730 -670
rect 77670 -830 77730 -770
rect 77840 -730 77900 -670
rect 77840 -830 77900 -770
rect 78010 -730 78070 -670
rect 78010 -830 78070 -770
rect 78180 -730 78240 -670
rect 78180 -830 78240 -770
rect 78350 -730 78410 -670
rect 78350 -830 78410 -770
rect 78520 -730 78580 -670
rect 78520 -830 78580 -770
rect 78690 -730 78750 -670
rect 78690 -830 78750 -770
rect 78860 -730 78920 -670
rect 78860 -830 78920 -770
rect 79030 -730 79090 -670
rect 79030 -830 79090 -770
rect 79200 -730 79260 -670
rect 79200 -830 79260 -770
rect 79370 -730 79430 -670
rect 79370 -830 79430 -770
rect 79540 -730 79600 -670
rect 79540 -830 79600 -770
rect 79710 -730 79770 -670
rect 79710 -830 79770 -770
rect 79880 -730 79940 -670
rect 79880 -830 79940 -770
rect 80050 -730 80110 -670
rect 80050 -830 80110 -770
rect 80220 -730 80280 -670
rect 80220 -830 80280 -770
rect 80390 -730 80450 -670
rect 80390 -830 80450 -770
rect 80560 -730 80620 -670
rect 80560 -830 80620 -770
rect 80730 -730 80790 -670
rect 80730 -830 80790 -770
rect 80900 -730 80960 -670
rect 80900 -830 80960 -770
rect 81070 -730 81130 -670
rect 81070 -830 81130 -770
rect 81240 -730 81300 -670
rect 81240 -830 81300 -770
rect 81410 -730 81470 -670
rect 81410 -830 81470 -770
rect 81580 -730 81640 -670
rect 81580 -830 81640 -770
rect 81750 -730 81810 -670
rect 81750 -830 81810 -770
rect 81920 -730 81980 -670
rect 81920 -830 81980 -770
rect 82090 -730 82150 -670
rect 82090 -830 82150 -770
rect 82260 -730 82320 -670
rect 82260 -830 82320 -770
rect 82430 -730 82490 -670
rect 82430 -830 82490 -770
rect 82600 -730 82660 -670
rect 82600 -830 82660 -770
rect 82770 -730 82830 -670
rect 82770 -830 82830 -770
rect 82940 -730 83000 -670
rect 82940 -830 83000 -770
rect 83110 -730 83170 -670
rect 83110 -830 83170 -770
rect 83280 -730 83340 -670
rect 83280 -830 83340 -770
rect 83450 -730 83510 -670
rect 83450 -830 83510 -770
rect 83620 -730 83680 -670
rect 83620 -830 83680 -770
rect 83790 -730 83850 -670
rect 83790 -830 83850 -770
rect 83960 -730 84020 -670
rect 83960 -830 84020 -770
rect 84130 -730 84190 -670
rect 84130 -830 84190 -770
rect 84300 -730 84360 -670
rect 84300 -830 84360 -770
rect 84470 -730 84530 -670
rect 84470 -830 84530 -770
rect 84640 -730 84700 -670
rect 84640 -830 84700 -770
rect 84810 -730 84870 -670
rect 84810 -830 84870 -770
rect 84980 -730 85040 -670
rect 84980 -830 85040 -770
rect 85150 -730 85210 -670
rect 85150 -830 85210 -770
rect 85320 -730 85380 -670
rect 85320 -830 85380 -770
rect 85490 -730 85550 -670
rect 85490 -830 85550 -770
rect 85660 -730 85720 -670
rect 85660 -830 85720 -770
rect 85830 -730 85890 -670
rect 85830 -830 85890 -770
rect 86000 -730 86060 -670
rect 86000 -830 86060 -770
rect 86170 -730 86230 -670
rect 86170 -830 86230 -770
rect 86340 -730 86400 -670
rect 86340 -830 86400 -770
rect 86510 -730 86570 -670
rect 86510 -830 86570 -770
rect 86680 -730 86740 -670
rect 86680 -830 86740 -770
rect 86850 -730 86910 -670
rect 86850 -830 86910 -770
rect 87020 -730 87080 -670
rect 87020 -830 87080 -770
rect 87190 -730 87250 -670
rect 87190 -830 87250 -770
<< pdiffc >>
rect 30 350 90 410
rect 30 250 90 310
rect 200 350 260 410
rect 200 250 260 310
rect 450 350 510 410
rect 450 250 510 310
rect 620 350 680 410
rect 620 250 680 310
rect 790 350 850 410
rect 790 250 850 310
rect 960 350 1020 410
rect 960 250 1020 310
rect 1130 350 1190 410
rect 1130 250 1190 310
rect 1520 350 1580 410
rect 1520 250 1580 310
rect 1690 350 1750 410
rect 1690 250 1750 310
rect 1860 350 1920 410
rect 1860 250 1920 310
rect 2030 350 2090 410
rect 2030 250 2090 310
rect 2200 350 2260 410
rect 2200 250 2260 310
rect 2370 350 2430 410
rect 2370 250 2430 310
rect 2540 350 2600 410
rect 2540 250 2600 310
rect 2710 350 2770 410
rect 2710 250 2770 310
rect 2880 350 2940 410
rect 2880 250 2940 310
rect 3050 350 3110 410
rect 3050 250 3110 310
rect 3220 350 3280 410
rect 3220 250 3280 310
rect 3390 350 3450 410
rect 3390 250 3450 310
rect 3560 350 3620 410
rect 3560 250 3620 310
rect 3730 350 3790 410
rect 3730 250 3790 310
rect 3900 350 3960 410
rect 3900 250 3960 310
rect 4070 350 4130 410
rect 4070 250 4130 310
rect 4240 350 4300 410
rect 4240 250 4300 310
rect 4540 350 4600 410
rect 4540 250 4600 310
rect 4710 350 4770 410
rect 4710 250 4770 310
rect 4880 350 4940 410
rect 4880 250 4940 310
rect 5050 350 5110 410
rect 5050 250 5110 310
rect 5220 350 5280 410
rect 5220 250 5280 310
rect 5390 350 5450 410
rect 5390 250 5450 310
rect 5560 350 5620 410
rect 5560 250 5620 310
rect 5730 350 5790 410
rect 5730 250 5790 310
rect 5900 350 5960 410
rect 5900 250 5960 310
rect 6070 350 6130 410
rect 6070 250 6130 310
rect 6240 350 6300 410
rect 6240 250 6300 310
rect 6410 350 6470 410
rect 6410 250 6470 310
rect 6580 350 6640 410
rect 6580 250 6640 310
rect 6750 350 6810 410
rect 6750 250 6810 310
rect 6920 350 6980 410
rect 6920 250 6980 310
rect 7090 350 7150 410
rect 7090 250 7150 310
rect 7260 350 7320 410
rect 7260 250 7320 310
rect 7430 350 7490 410
rect 7430 250 7490 310
rect 7600 350 7660 410
rect 7600 250 7660 310
rect 7770 350 7830 410
rect 7770 250 7830 310
rect 7940 350 8000 410
rect 7940 250 8000 310
rect 8110 350 8170 410
rect 8110 250 8170 310
rect 8280 350 8340 410
rect 8280 250 8340 310
rect 8450 350 8510 410
rect 8450 250 8510 310
rect 8620 350 8680 410
rect 8620 250 8680 310
rect 8790 350 8850 410
rect 8790 250 8850 310
rect 8960 350 9020 410
rect 8960 250 9020 310
rect 9130 350 9190 410
rect 9130 250 9190 310
rect 9300 350 9360 410
rect 9300 250 9360 310
rect 9470 350 9530 410
rect 9470 250 9530 310
rect 9640 350 9700 410
rect 9640 250 9700 310
rect 9810 350 9870 410
rect 9810 250 9870 310
rect 9980 350 10040 410
rect 9980 250 10040 310
rect 10150 350 10210 410
rect 10150 250 10210 310
rect 10320 350 10380 410
rect 10320 250 10380 310
rect 10490 350 10550 410
rect 10490 250 10550 310
rect 10660 350 10720 410
rect 10660 250 10720 310
rect 10830 350 10890 410
rect 10830 250 10890 310
rect 11000 350 11060 410
rect 11000 250 11060 310
rect 11170 350 11230 410
rect 11170 250 11230 310
rect 11340 350 11400 410
rect 11340 250 11400 310
rect 11510 350 11570 410
rect 11510 250 11570 310
rect 11680 350 11740 410
rect 11680 250 11740 310
rect 11850 350 11910 410
rect 11850 250 11910 310
rect 12020 350 12080 410
rect 12020 250 12080 310
rect 12190 350 12250 410
rect 12190 250 12250 310
rect 12360 350 12420 410
rect 12360 250 12420 310
rect 12530 350 12590 410
rect 12530 250 12590 310
rect 12700 350 12760 410
rect 12700 250 12760 310
rect 12870 350 12930 410
rect 12870 250 12930 310
rect 13040 350 13100 410
rect 13040 250 13100 310
rect 13210 350 13270 410
rect 13210 250 13270 310
rect 13380 350 13440 410
rect 13380 250 13440 310
rect 13550 350 13610 410
rect 13550 250 13610 310
rect 13720 350 13780 410
rect 13720 250 13780 310
rect 13890 350 13950 410
rect 13890 250 13950 310
rect 14060 350 14120 410
rect 14060 250 14120 310
rect 14230 350 14290 410
rect 14230 250 14290 310
rect 14400 350 14460 410
rect 14400 250 14460 310
rect 14570 350 14630 410
rect 14570 250 14630 310
rect 14740 350 14800 410
rect 14740 250 14800 310
rect 14910 350 14970 410
rect 14910 250 14970 310
rect 15080 350 15140 410
rect 15080 250 15140 310
rect 15250 350 15310 410
rect 15250 250 15310 310
rect 15420 350 15480 410
rect 15420 250 15480 310
rect 15720 350 15780 410
rect 15720 250 15780 310
rect 15890 350 15950 410
rect 15890 250 15950 310
rect 16060 350 16120 410
rect 16060 250 16120 310
rect 16230 350 16290 410
rect 16230 250 16290 310
rect 16400 350 16460 410
rect 16400 250 16460 310
rect 16570 350 16630 410
rect 16570 250 16630 310
rect 16740 350 16800 410
rect 16740 250 16800 310
rect 16910 350 16970 410
rect 16910 250 16970 310
rect 17080 350 17140 410
rect 17080 250 17140 310
rect 17250 350 17310 410
rect 17250 250 17310 310
rect 17420 350 17480 410
rect 17420 250 17480 310
rect 17590 350 17650 410
rect 17590 250 17650 310
rect 17760 350 17820 410
rect 17760 250 17820 310
rect 17930 350 17990 410
rect 17930 250 17990 310
rect 18100 350 18160 410
rect 18100 250 18160 310
rect 18270 350 18330 410
rect 18270 250 18330 310
rect 18440 350 18500 410
rect 18440 250 18500 310
rect 18610 350 18670 410
rect 18610 250 18670 310
rect 18780 350 18840 410
rect 18780 250 18840 310
rect 18950 350 19010 410
rect 18950 250 19010 310
rect 19120 350 19180 410
rect 19120 250 19180 310
rect 19290 350 19350 410
rect 19290 250 19350 310
rect 19460 350 19520 410
rect 19460 250 19520 310
rect 19630 350 19690 410
rect 19630 250 19690 310
rect 19800 350 19860 410
rect 19800 250 19860 310
rect 19970 350 20030 410
rect 19970 250 20030 310
rect 20140 350 20200 410
rect 20140 250 20200 310
rect 20310 350 20370 410
rect 20310 250 20370 310
rect 20480 350 20540 410
rect 20480 250 20540 310
rect 20650 350 20710 410
rect 20650 250 20710 310
rect 20820 350 20880 410
rect 20820 250 20880 310
rect 20990 350 21050 410
rect 20990 250 21050 310
rect 21160 350 21220 410
rect 21160 250 21220 310
rect 21330 350 21390 410
rect 21330 250 21390 310
rect 21500 350 21560 410
rect 21500 250 21560 310
rect 21670 350 21730 410
rect 21670 250 21730 310
rect 21840 350 21900 410
rect 21840 250 21900 310
rect 22010 350 22070 410
rect 22010 250 22070 310
rect 22180 350 22240 410
rect 22180 250 22240 310
rect 22350 350 22410 410
rect 22350 250 22410 310
rect 22520 350 22580 410
rect 22520 250 22580 310
rect 22690 350 22750 410
rect 22690 250 22750 310
rect 22860 350 22920 410
rect 22860 250 22920 310
rect 23030 350 23090 410
rect 23030 250 23090 310
rect 23200 350 23260 410
rect 23200 250 23260 310
rect 23370 350 23430 410
rect 23370 250 23430 310
rect 23540 350 23600 410
rect 23540 250 23600 310
rect 23710 350 23770 410
rect 23710 250 23770 310
rect 23880 350 23940 410
rect 23880 250 23940 310
rect 24050 350 24110 410
rect 24050 250 24110 310
rect 24220 350 24280 410
rect 24220 250 24280 310
rect 24390 350 24450 410
rect 24390 250 24450 310
rect 24560 350 24620 410
rect 24560 250 24620 310
rect 24730 350 24790 410
rect 24730 250 24790 310
rect 24900 350 24960 410
rect 24900 250 24960 310
rect 25070 350 25130 410
rect 25070 250 25130 310
rect 25240 350 25300 410
rect 25240 250 25300 310
rect 25410 350 25470 410
rect 25410 250 25470 310
rect 25580 350 25640 410
rect 25580 250 25640 310
rect 25750 350 25810 410
rect 25750 250 25810 310
rect 25920 350 25980 410
rect 25920 250 25980 310
rect 26090 350 26150 410
rect 26090 250 26150 310
rect 26260 350 26320 410
rect 26260 250 26320 310
rect 26430 350 26490 410
rect 26430 250 26490 310
rect 26600 350 26660 410
rect 26600 250 26660 310
rect 26770 350 26830 410
rect 26770 250 26830 310
rect 26940 350 27000 410
rect 26940 250 27000 310
rect 27110 350 27170 410
rect 27110 250 27170 310
rect 27280 350 27340 410
rect 27280 250 27340 310
rect 27450 350 27510 410
rect 27450 250 27510 310
rect 27620 350 27680 410
rect 27620 250 27680 310
rect 27790 350 27850 410
rect 27790 250 27850 310
rect 27960 350 28020 410
rect 27960 250 28020 310
rect 28130 350 28190 410
rect 28130 250 28190 310
rect 28300 350 28360 410
rect 28300 250 28360 310
rect 28470 350 28530 410
rect 28470 250 28530 310
rect 28640 350 28700 410
rect 28640 250 28700 310
rect 28810 350 28870 410
rect 28810 250 28870 310
rect 28980 350 29040 410
rect 28980 250 29040 310
rect 29150 350 29210 410
rect 29150 250 29210 310
rect 29320 350 29380 410
rect 29320 250 29380 310
rect 29490 350 29550 410
rect 29490 250 29550 310
rect 29660 350 29720 410
rect 29660 250 29720 310
rect 29830 350 29890 410
rect 29830 250 29890 310
rect 30000 350 30060 410
rect 30000 250 30060 310
rect 30170 350 30230 410
rect 30170 250 30230 310
rect 30340 350 30400 410
rect 30340 250 30400 310
rect 30510 350 30570 410
rect 30510 250 30570 310
rect 30680 350 30740 410
rect 30680 250 30740 310
rect 30850 350 30910 410
rect 30850 250 30910 310
rect 31020 350 31080 410
rect 31020 250 31080 310
rect 31190 350 31250 410
rect 31190 250 31250 310
rect 31360 350 31420 410
rect 31360 250 31420 310
rect 31530 350 31590 410
rect 31530 250 31590 310
rect 31700 350 31760 410
rect 31700 250 31760 310
rect 31870 350 31930 410
rect 31870 250 31930 310
rect 32040 350 32100 410
rect 32040 250 32100 310
rect 32210 350 32270 410
rect 32210 250 32270 310
rect 32380 350 32440 410
rect 32380 250 32440 310
rect 32550 350 32610 410
rect 32550 250 32610 310
rect 32720 350 32780 410
rect 32720 250 32780 310
rect 32890 350 32950 410
rect 32890 250 32950 310
rect 33060 350 33120 410
rect 33060 250 33120 310
rect 33230 350 33290 410
rect 33230 250 33290 310
rect 33400 350 33460 410
rect 33400 250 33460 310
rect 33570 350 33630 410
rect 33570 250 33630 310
rect 33740 350 33800 410
rect 33740 250 33800 310
rect 33910 350 33970 410
rect 33910 250 33970 310
rect 34080 350 34140 410
rect 34080 250 34140 310
rect 34250 350 34310 410
rect 34250 250 34310 310
rect 34420 350 34480 410
rect 34420 250 34480 310
rect 34590 350 34650 410
rect 34590 250 34650 310
rect 34760 350 34820 410
rect 34760 250 34820 310
rect 34930 350 34990 410
rect 34930 250 34990 310
rect 35100 350 35160 410
rect 35100 250 35160 310
rect 35270 350 35330 410
rect 35270 250 35330 310
rect 35440 350 35500 410
rect 35440 250 35500 310
rect 35610 350 35670 410
rect 35610 250 35670 310
rect 35780 350 35840 410
rect 35780 250 35840 310
rect 35950 350 36010 410
rect 35950 250 36010 310
rect 36120 350 36180 410
rect 36120 250 36180 310
rect 36290 350 36350 410
rect 36290 250 36350 310
rect 36460 350 36520 410
rect 36460 250 36520 310
rect 36630 350 36690 410
rect 36630 250 36690 310
rect 36800 350 36860 410
rect 36800 250 36860 310
rect 36970 350 37030 410
rect 36970 250 37030 310
rect 37140 350 37200 410
rect 37140 250 37200 310
rect 37310 350 37370 410
rect 37310 250 37370 310
rect 37480 350 37540 410
rect 37480 250 37540 310
rect 37650 350 37710 410
rect 37650 250 37710 310
rect 37820 350 37880 410
rect 37820 250 37880 310
rect 37990 350 38050 410
rect 37990 250 38050 310
rect 38160 350 38220 410
rect 38160 250 38220 310
rect 38330 350 38390 410
rect 38330 250 38390 310
rect 38500 350 38560 410
rect 38500 250 38560 310
rect 38670 350 38730 410
rect 38670 250 38730 310
rect 38840 350 38900 410
rect 38840 250 38900 310
rect 39010 350 39070 410
rect 39010 250 39070 310
rect 39180 350 39240 410
rect 39180 250 39240 310
rect 39350 350 39410 410
rect 39350 250 39410 310
rect 39520 350 39580 410
rect 39520 250 39580 310
rect 39690 350 39750 410
rect 39690 250 39750 310
rect 39860 350 39920 410
rect 39860 250 39920 310
rect 40030 350 40090 410
rect 40030 250 40090 310
rect 40200 350 40260 410
rect 40200 250 40260 310
rect 40370 350 40430 410
rect 40370 250 40430 310
rect 40540 350 40600 410
rect 40540 250 40600 310
rect 40710 350 40770 410
rect 40710 250 40770 310
rect 40880 350 40940 410
rect 40880 250 40940 310
rect 41050 350 41110 410
rect 41050 250 41110 310
rect 41220 350 41280 410
rect 41220 250 41280 310
rect 41390 350 41450 410
rect 41390 250 41450 310
rect 41560 350 41620 410
rect 41560 250 41620 310
rect 41730 350 41790 410
rect 41730 250 41790 310
rect 41900 350 41960 410
rect 41900 250 41960 310
rect 42070 350 42130 410
rect 42070 250 42130 310
rect 42240 350 42300 410
rect 42240 250 42300 310
rect 42410 350 42470 410
rect 42410 250 42470 310
rect 42580 350 42640 410
rect 42580 250 42640 310
rect 42750 350 42810 410
rect 42750 250 42810 310
rect 42920 350 42980 410
rect 42920 250 42980 310
rect 43090 350 43150 410
rect 43090 250 43150 310
rect 43260 350 43320 410
rect 43260 250 43320 310
rect 43430 350 43490 410
rect 43430 250 43490 310
rect 43600 350 43660 410
rect 43600 250 43660 310
rect 43770 350 43830 410
rect 43770 250 43830 310
rect 43940 350 44000 410
rect 43940 250 44000 310
rect 44110 350 44170 410
rect 44110 250 44170 310
rect 44280 350 44340 410
rect 44280 250 44340 310
rect 44450 350 44510 410
rect 44450 250 44510 310
rect 44620 350 44680 410
rect 44620 250 44680 310
rect 44790 350 44850 410
rect 44790 250 44850 310
rect 44960 350 45020 410
rect 44960 250 45020 310
rect 45130 350 45190 410
rect 45130 250 45190 310
rect 45300 350 45360 410
rect 45300 250 45360 310
rect 45470 350 45530 410
rect 45470 250 45530 310
rect 45640 350 45700 410
rect 45640 250 45700 310
rect 45810 350 45870 410
rect 45810 250 45870 310
rect 45980 350 46040 410
rect 45980 250 46040 310
rect 46150 350 46210 410
rect 46150 250 46210 310
rect 46320 350 46380 410
rect 46320 250 46380 310
rect 46490 350 46550 410
rect 46490 250 46550 310
rect 46660 350 46720 410
rect 46660 250 46720 310
rect 46830 350 46890 410
rect 46830 250 46890 310
rect 47000 350 47060 410
rect 47000 250 47060 310
rect 47170 350 47230 410
rect 47170 250 47230 310
rect 47340 350 47400 410
rect 47340 250 47400 310
rect 47510 350 47570 410
rect 47510 250 47570 310
rect 47680 350 47740 410
rect 47680 250 47740 310
rect 47850 350 47910 410
rect 47850 250 47910 310
rect 48020 350 48080 410
rect 48020 250 48080 310
rect 48190 350 48250 410
rect 48190 250 48250 310
rect 48360 350 48420 410
rect 48360 250 48420 310
rect 48530 350 48590 410
rect 48530 250 48590 310
rect 48700 350 48760 410
rect 48700 250 48760 310
rect 48870 350 48930 410
rect 48870 250 48930 310
rect 49040 350 49100 410
rect 49040 250 49100 310
rect 49210 350 49270 410
rect 49210 250 49270 310
rect 49380 350 49440 410
rect 49380 250 49440 310
rect 49550 350 49610 410
rect 49550 250 49610 310
rect 49720 350 49780 410
rect 49720 250 49780 310
rect 49890 350 49950 410
rect 49890 250 49950 310
rect 50060 350 50120 410
rect 50060 250 50120 310
rect 50230 350 50290 410
rect 50230 250 50290 310
rect 50400 350 50460 410
rect 50400 250 50460 310
rect 50570 350 50630 410
rect 50570 250 50630 310
rect 50740 350 50800 410
rect 50740 250 50800 310
rect 50910 350 50970 410
rect 50910 250 50970 310
rect 51080 350 51140 410
rect 51080 250 51140 310
rect 51250 350 51310 410
rect 51250 250 51310 310
rect 51420 350 51480 410
rect 51420 250 51480 310
rect 51590 350 51650 410
rect 51590 250 51650 310
rect 51760 350 51820 410
rect 51760 250 51820 310
rect 51930 350 51990 410
rect 51930 250 51990 310
rect 52100 350 52160 410
rect 52100 250 52160 310
rect 52270 350 52330 410
rect 52270 250 52330 310
rect 52440 350 52500 410
rect 52440 250 52500 310
rect 52610 350 52670 410
rect 52610 250 52670 310
rect 52780 350 52840 410
rect 52780 250 52840 310
rect 52950 350 53010 410
rect 52950 250 53010 310
rect 53120 350 53180 410
rect 53120 250 53180 310
rect 53290 350 53350 410
rect 53290 250 53350 310
rect 53460 350 53520 410
rect 53460 250 53520 310
rect 53630 350 53690 410
rect 53630 250 53690 310
rect 53800 350 53860 410
rect 53800 250 53860 310
rect 53970 350 54030 410
rect 53970 250 54030 310
rect 54140 350 54200 410
rect 54140 250 54200 310
rect 54310 350 54370 410
rect 54310 250 54370 310
rect 54480 350 54540 410
rect 54480 250 54540 310
rect 54650 350 54710 410
rect 54650 250 54710 310
rect 54820 350 54880 410
rect 54820 250 54880 310
rect 54990 350 55050 410
rect 54990 250 55050 310
rect 55160 350 55220 410
rect 55160 250 55220 310
rect 55330 350 55390 410
rect 55330 250 55390 310
rect 55500 350 55560 410
rect 55500 250 55560 310
rect 55670 350 55730 410
rect 55670 250 55730 310
rect 55840 350 55900 410
rect 55840 250 55900 310
rect 56010 350 56070 410
rect 56010 250 56070 310
rect 56180 350 56240 410
rect 56180 250 56240 310
rect 56350 350 56410 410
rect 56350 250 56410 310
rect 56520 350 56580 410
rect 56520 250 56580 310
rect 56690 350 56750 410
rect 56690 250 56750 310
rect 56860 350 56920 410
rect 56860 250 56920 310
rect 57030 350 57090 410
rect 57030 250 57090 310
rect 57200 350 57260 410
rect 57200 250 57260 310
rect 57370 350 57430 410
rect 57370 250 57430 310
rect 57540 350 57600 410
rect 57540 250 57600 310
rect 57710 350 57770 410
rect 57710 250 57770 310
rect 57880 350 57940 410
rect 57880 250 57940 310
rect 58050 350 58110 410
rect 58050 250 58110 310
rect 58220 350 58280 410
rect 58220 250 58280 310
rect 58390 350 58450 410
rect 58390 250 58450 310
rect 58560 350 58620 410
rect 58560 250 58620 310
rect 58730 350 58790 410
rect 58730 250 58790 310
rect 58900 350 58960 410
rect 58900 250 58960 310
rect 59070 350 59130 410
rect 59070 250 59130 310
rect 59240 350 59300 410
rect 59240 250 59300 310
rect 150 -1060 210 -1000
rect 150 -1160 210 -1100
rect 150 -1260 210 -1200
rect 150 -1360 210 -1300
rect 320 -1060 380 -1000
rect 320 -1160 380 -1100
rect 320 -1260 380 -1200
rect 320 -1360 380 -1300
rect 490 -1060 550 -1000
rect 490 -1160 550 -1100
rect 490 -1260 550 -1200
rect 490 -1360 550 -1300
rect 660 -1060 720 -1000
rect 660 -1160 720 -1100
rect 660 -1260 720 -1200
rect 660 -1360 720 -1300
rect 830 -1060 890 -1000
rect 830 -1160 890 -1100
rect 830 -1260 890 -1200
rect 830 -1360 890 -1300
rect 1000 -1060 1060 -1000
rect 1000 -1160 1060 -1100
rect 1000 -1260 1060 -1200
rect 1000 -1360 1060 -1300
rect 1170 -1060 1230 -1000
rect 1170 -1160 1230 -1100
rect 1170 -1260 1230 -1200
rect 1170 -1360 1230 -1300
rect 1340 -1060 1400 -1000
rect 1340 -1160 1400 -1100
rect 1340 -1260 1400 -1200
rect 1340 -1360 1400 -1300
rect 1510 -1060 1570 -1000
rect 1510 -1160 1570 -1100
rect 1510 -1260 1570 -1200
rect 1510 -1360 1570 -1300
rect 1680 -1060 1740 -1000
rect 1680 -1160 1740 -1100
rect 1680 -1260 1740 -1200
rect 1680 -1360 1740 -1300
rect 1850 -1060 1910 -1000
rect 1850 -1160 1910 -1100
rect 1850 -1260 1910 -1200
rect 1850 -1360 1910 -1300
rect 2020 -1060 2080 -1000
rect 2020 -1160 2080 -1100
rect 2020 -1260 2080 -1200
rect 2020 -1360 2080 -1300
rect 2190 -1060 2250 -1000
rect 2190 -1160 2250 -1100
rect 2190 -1260 2250 -1200
rect 2190 -1360 2250 -1300
rect 2360 -1060 2420 -1000
rect 2360 -1160 2420 -1100
rect 2360 -1260 2420 -1200
rect 2360 -1360 2420 -1300
rect 2530 -1060 2590 -1000
rect 2530 -1160 2590 -1100
rect 2530 -1260 2590 -1200
rect 2530 -1360 2590 -1300
rect 2700 -1060 2760 -1000
rect 2700 -1160 2760 -1100
rect 2700 -1260 2760 -1200
rect 2700 -1360 2760 -1300
rect 2870 -1060 2930 -1000
rect 2870 -1160 2930 -1100
rect 2870 -1260 2930 -1200
rect 2870 -1360 2930 -1300
rect 3040 -1060 3100 -1000
rect 3040 -1160 3100 -1100
rect 3040 -1260 3100 -1200
rect 3040 -1360 3100 -1300
rect 3210 -1060 3270 -1000
rect 3210 -1160 3270 -1100
rect 3210 -1260 3270 -1200
rect 3210 -1360 3270 -1300
rect 3380 -1060 3440 -1000
rect 3380 -1160 3440 -1100
rect 3380 -1260 3440 -1200
rect 3380 -1360 3440 -1300
rect 3550 -1060 3610 -1000
rect 3550 -1160 3610 -1100
rect 3550 -1260 3610 -1200
rect 3550 -1360 3610 -1300
rect 3720 -1060 3780 -1000
rect 3720 -1160 3780 -1100
rect 3720 -1260 3780 -1200
rect 3720 -1360 3780 -1300
rect 3890 -1060 3950 -1000
rect 3890 -1160 3950 -1100
rect 3890 -1260 3950 -1200
rect 3890 -1360 3950 -1300
rect 4060 -1060 4120 -1000
rect 4060 -1160 4120 -1100
rect 4060 -1260 4120 -1200
rect 4060 -1360 4120 -1300
rect 4230 -1060 4290 -1000
rect 4230 -1160 4290 -1100
rect 4230 -1260 4290 -1200
rect 4230 -1360 4290 -1300
rect 4400 -1060 4460 -1000
rect 4400 -1160 4460 -1100
rect 4400 -1260 4460 -1200
rect 4400 -1360 4460 -1300
rect 4570 -1060 4630 -1000
rect 4570 -1160 4630 -1100
rect 4570 -1260 4630 -1200
rect 4570 -1360 4630 -1300
rect 4740 -1060 4800 -1000
rect 4740 -1160 4800 -1100
rect 4740 -1260 4800 -1200
rect 4740 -1360 4800 -1300
rect 4910 -1060 4970 -1000
rect 4910 -1160 4970 -1100
rect 4910 -1260 4970 -1200
rect 4910 -1360 4970 -1300
rect 5080 -1060 5140 -1000
rect 5080 -1160 5140 -1100
rect 5080 -1260 5140 -1200
rect 5080 -1360 5140 -1300
rect 5250 -1060 5310 -1000
rect 5250 -1160 5310 -1100
rect 5250 -1260 5310 -1200
rect 5250 -1360 5310 -1300
rect 5420 -1060 5480 -1000
rect 5420 -1160 5480 -1100
rect 5420 -1260 5480 -1200
rect 5420 -1360 5480 -1300
rect 5590 -1060 5650 -1000
rect 5590 -1160 5650 -1100
rect 5590 -1260 5650 -1200
rect 5590 -1360 5650 -1300
rect 5760 -1060 5820 -1000
rect 5760 -1160 5820 -1100
rect 5760 -1260 5820 -1200
rect 5760 -1360 5820 -1300
rect 5930 -1060 5990 -1000
rect 5930 -1160 5990 -1100
rect 5930 -1260 5990 -1200
rect 5930 -1360 5990 -1300
rect 6100 -1060 6160 -1000
rect 6100 -1160 6160 -1100
rect 6100 -1260 6160 -1200
rect 6100 -1360 6160 -1300
rect 6270 -1060 6330 -1000
rect 6270 -1160 6330 -1100
rect 6270 -1260 6330 -1200
rect 6270 -1360 6330 -1300
rect 6440 -1060 6500 -1000
rect 6440 -1160 6500 -1100
rect 6440 -1260 6500 -1200
rect 6440 -1360 6500 -1300
rect 6610 -1060 6670 -1000
rect 6610 -1160 6670 -1100
rect 6610 -1260 6670 -1200
rect 6610 -1360 6670 -1300
rect 6780 -1060 6840 -1000
rect 6780 -1160 6840 -1100
rect 6780 -1260 6840 -1200
rect 6780 -1360 6840 -1300
rect 6950 -1060 7010 -1000
rect 6950 -1160 7010 -1100
rect 6950 -1260 7010 -1200
rect 6950 -1360 7010 -1300
rect 7120 -1060 7180 -1000
rect 7120 -1160 7180 -1100
rect 7120 -1260 7180 -1200
rect 7120 -1360 7180 -1300
rect 7290 -1060 7350 -1000
rect 7290 -1160 7350 -1100
rect 7290 -1260 7350 -1200
rect 7290 -1360 7350 -1300
rect 7460 -1060 7520 -1000
rect 7460 -1160 7520 -1100
rect 7460 -1260 7520 -1200
rect 7460 -1360 7520 -1300
rect 7630 -1060 7690 -1000
rect 7630 -1160 7690 -1100
rect 7630 -1260 7690 -1200
rect 7630 -1360 7690 -1300
rect 7800 -1060 7860 -1000
rect 7800 -1160 7860 -1100
rect 7800 -1260 7860 -1200
rect 7800 -1360 7860 -1300
rect 7970 -1060 8030 -1000
rect 7970 -1160 8030 -1100
rect 7970 -1260 8030 -1200
rect 7970 -1360 8030 -1300
rect 8140 -1060 8200 -1000
rect 8140 -1160 8200 -1100
rect 8140 -1260 8200 -1200
rect 8140 -1360 8200 -1300
rect 8310 -1060 8370 -1000
rect 8310 -1160 8370 -1100
rect 8310 -1260 8370 -1200
rect 8310 -1360 8370 -1300
rect 8480 -1060 8540 -1000
rect 8480 -1160 8540 -1100
rect 8480 -1260 8540 -1200
rect 8480 -1360 8540 -1300
rect 8650 -1060 8710 -1000
rect 8650 -1160 8710 -1100
rect 8650 -1260 8710 -1200
rect 8650 -1360 8710 -1300
rect 8820 -1060 8880 -1000
rect 8820 -1160 8880 -1100
rect 8820 -1260 8880 -1200
rect 8820 -1360 8880 -1300
rect 8990 -1060 9050 -1000
rect 8990 -1160 9050 -1100
rect 8990 -1260 9050 -1200
rect 8990 -1360 9050 -1300
rect 9160 -1060 9220 -1000
rect 9160 -1160 9220 -1100
rect 9160 -1260 9220 -1200
rect 9160 -1360 9220 -1300
rect 9330 -1060 9390 -1000
rect 9330 -1160 9390 -1100
rect 9330 -1260 9390 -1200
rect 9330 -1360 9390 -1300
rect 9500 -1060 9560 -1000
rect 9500 -1160 9560 -1100
rect 9500 -1260 9560 -1200
rect 9500 -1360 9560 -1300
rect 9670 -1060 9730 -1000
rect 9670 -1160 9730 -1100
rect 9670 -1260 9730 -1200
rect 9670 -1360 9730 -1300
rect 9840 -1060 9900 -1000
rect 9840 -1160 9900 -1100
rect 9840 -1260 9900 -1200
rect 9840 -1360 9900 -1300
rect 10010 -1060 10070 -1000
rect 10010 -1160 10070 -1100
rect 10010 -1260 10070 -1200
rect 10010 -1360 10070 -1300
rect 10180 -1060 10240 -1000
rect 10180 -1160 10240 -1100
rect 10180 -1260 10240 -1200
rect 10180 -1360 10240 -1300
rect 10350 -1060 10410 -1000
rect 10350 -1160 10410 -1100
rect 10350 -1260 10410 -1200
rect 10350 -1360 10410 -1300
rect 10520 -1060 10580 -1000
rect 10520 -1160 10580 -1100
rect 10520 -1260 10580 -1200
rect 10520 -1360 10580 -1300
rect 10690 -1060 10750 -1000
rect 10690 -1160 10750 -1100
rect 10690 -1260 10750 -1200
rect 10690 -1360 10750 -1300
rect 10860 -1060 10920 -1000
rect 10860 -1160 10920 -1100
rect 10860 -1260 10920 -1200
rect 10860 -1360 10920 -1300
rect 11030 -1060 11090 -1000
rect 11030 -1160 11090 -1100
rect 11030 -1260 11090 -1200
rect 11030 -1360 11090 -1300
rect 11200 -1060 11260 -1000
rect 11200 -1160 11260 -1100
rect 11200 -1260 11260 -1200
rect 11200 -1360 11260 -1300
rect 11370 -1060 11430 -1000
rect 11370 -1160 11430 -1100
rect 11370 -1260 11430 -1200
rect 11370 -1360 11430 -1300
rect 11540 -1060 11600 -1000
rect 11540 -1160 11600 -1100
rect 11540 -1260 11600 -1200
rect 11540 -1360 11600 -1300
rect 11710 -1060 11770 -1000
rect 11710 -1160 11770 -1100
rect 11710 -1260 11770 -1200
rect 11710 -1360 11770 -1300
rect 11880 -1060 11940 -1000
rect 11880 -1160 11940 -1100
rect 11880 -1260 11940 -1200
rect 11880 -1360 11940 -1300
rect 12050 -1060 12110 -1000
rect 12050 -1160 12110 -1100
rect 12050 -1260 12110 -1200
rect 12050 -1360 12110 -1300
rect 12220 -1060 12280 -1000
rect 12220 -1160 12280 -1100
rect 12220 -1260 12280 -1200
rect 12220 -1360 12280 -1300
rect 12390 -1060 12450 -1000
rect 12390 -1160 12450 -1100
rect 12390 -1260 12450 -1200
rect 12390 -1360 12450 -1300
rect 12560 -1060 12620 -1000
rect 12560 -1160 12620 -1100
rect 12560 -1260 12620 -1200
rect 12560 -1360 12620 -1300
rect 12730 -1060 12790 -1000
rect 12730 -1160 12790 -1100
rect 12730 -1260 12790 -1200
rect 12730 -1360 12790 -1300
rect 12900 -1060 12960 -1000
rect 12900 -1160 12960 -1100
rect 12900 -1260 12960 -1200
rect 12900 -1360 12960 -1300
rect 13070 -1060 13130 -1000
rect 13070 -1160 13130 -1100
rect 13070 -1260 13130 -1200
rect 13070 -1360 13130 -1300
rect 13240 -1060 13300 -1000
rect 13240 -1160 13300 -1100
rect 13240 -1260 13300 -1200
rect 13240 -1360 13300 -1300
rect 13410 -1060 13470 -1000
rect 13410 -1160 13470 -1100
rect 13410 -1260 13470 -1200
rect 13410 -1360 13470 -1300
rect 13580 -1060 13640 -1000
rect 13580 -1160 13640 -1100
rect 13580 -1260 13640 -1200
rect 13580 -1360 13640 -1300
rect 13750 -1060 13810 -1000
rect 13750 -1160 13810 -1100
rect 13750 -1260 13810 -1200
rect 13750 -1360 13810 -1300
rect 13920 -1060 13980 -1000
rect 13920 -1160 13980 -1100
rect 13920 -1260 13980 -1200
rect 13920 -1360 13980 -1300
rect 14090 -1060 14150 -1000
rect 14090 -1160 14150 -1100
rect 14090 -1260 14150 -1200
rect 14090 -1360 14150 -1300
rect 14260 -1060 14320 -1000
rect 14260 -1160 14320 -1100
rect 14260 -1260 14320 -1200
rect 14260 -1360 14320 -1300
rect 14430 -1060 14490 -1000
rect 14430 -1160 14490 -1100
rect 14430 -1260 14490 -1200
rect 14430 -1360 14490 -1300
rect 14600 -1060 14660 -1000
rect 14600 -1160 14660 -1100
rect 14600 -1260 14660 -1200
rect 14600 -1360 14660 -1300
rect 14770 -1060 14830 -1000
rect 14770 -1160 14830 -1100
rect 14770 -1260 14830 -1200
rect 14770 -1360 14830 -1300
rect 14940 -1060 15000 -1000
rect 14940 -1160 15000 -1100
rect 14940 -1260 15000 -1200
rect 14940 -1360 15000 -1300
rect 15110 -1060 15170 -1000
rect 15110 -1160 15170 -1100
rect 15110 -1260 15170 -1200
rect 15110 -1360 15170 -1300
rect 15280 -1060 15340 -1000
rect 15280 -1160 15340 -1100
rect 15280 -1260 15340 -1200
rect 15280 -1360 15340 -1300
rect 15450 -1060 15510 -1000
rect 15450 -1160 15510 -1100
rect 15450 -1260 15510 -1200
rect 15450 -1360 15510 -1300
rect 15620 -1060 15680 -1000
rect 15620 -1160 15680 -1100
rect 15620 -1260 15680 -1200
rect 15620 -1360 15680 -1300
rect 15790 -1060 15850 -1000
rect 15790 -1160 15850 -1100
rect 15790 -1260 15850 -1200
rect 15790 -1360 15850 -1300
rect 15960 -1060 16020 -1000
rect 15960 -1160 16020 -1100
rect 15960 -1260 16020 -1200
rect 15960 -1360 16020 -1300
rect 16130 -1060 16190 -1000
rect 16130 -1160 16190 -1100
rect 16130 -1260 16190 -1200
rect 16130 -1360 16190 -1300
rect 16300 -1060 16360 -1000
rect 16300 -1160 16360 -1100
rect 16300 -1260 16360 -1200
rect 16300 -1360 16360 -1300
rect 16470 -1060 16530 -1000
rect 16470 -1160 16530 -1100
rect 16470 -1260 16530 -1200
rect 16470 -1360 16530 -1300
rect 16640 -1060 16700 -1000
rect 16640 -1160 16700 -1100
rect 16640 -1260 16700 -1200
rect 16640 -1360 16700 -1300
rect 16810 -1060 16870 -1000
rect 16810 -1160 16870 -1100
rect 16810 -1260 16870 -1200
rect 16810 -1360 16870 -1300
rect 16980 -1060 17040 -1000
rect 16980 -1160 17040 -1100
rect 16980 -1260 17040 -1200
rect 16980 -1360 17040 -1300
rect 17150 -1060 17210 -1000
rect 17150 -1160 17210 -1100
rect 17150 -1260 17210 -1200
rect 17150 -1360 17210 -1300
rect 17320 -1060 17380 -1000
rect 17320 -1160 17380 -1100
rect 17320 -1260 17380 -1200
rect 17320 -1360 17380 -1300
rect 17490 -1060 17550 -1000
rect 17490 -1160 17550 -1100
rect 17490 -1260 17550 -1200
rect 17490 -1360 17550 -1300
rect 17660 -1060 17720 -1000
rect 17660 -1160 17720 -1100
rect 17660 -1260 17720 -1200
rect 17660 -1360 17720 -1300
rect 17830 -1060 17890 -1000
rect 17830 -1160 17890 -1100
rect 17830 -1260 17890 -1200
rect 17830 -1360 17890 -1300
rect 18000 -1060 18060 -1000
rect 18000 -1160 18060 -1100
rect 18000 -1260 18060 -1200
rect 18000 -1360 18060 -1300
rect 18170 -1060 18230 -1000
rect 18170 -1160 18230 -1100
rect 18170 -1260 18230 -1200
rect 18170 -1360 18230 -1300
rect 18340 -1060 18400 -1000
rect 18340 -1160 18400 -1100
rect 18340 -1260 18400 -1200
rect 18340 -1360 18400 -1300
rect 18510 -1060 18570 -1000
rect 18510 -1160 18570 -1100
rect 18510 -1260 18570 -1200
rect 18510 -1360 18570 -1300
rect 18680 -1060 18740 -1000
rect 18680 -1160 18740 -1100
rect 18680 -1260 18740 -1200
rect 18680 -1360 18740 -1300
rect 18850 -1060 18910 -1000
rect 18850 -1160 18910 -1100
rect 18850 -1260 18910 -1200
rect 18850 -1360 18910 -1300
rect 19020 -1060 19080 -1000
rect 19020 -1160 19080 -1100
rect 19020 -1260 19080 -1200
rect 19020 -1360 19080 -1300
rect 19190 -1060 19250 -1000
rect 19190 -1160 19250 -1100
rect 19190 -1260 19250 -1200
rect 19190 -1360 19250 -1300
rect 19360 -1060 19420 -1000
rect 19360 -1160 19420 -1100
rect 19360 -1260 19420 -1200
rect 19360 -1360 19420 -1300
rect 19530 -1060 19590 -1000
rect 19530 -1160 19590 -1100
rect 19530 -1260 19590 -1200
rect 19530 -1360 19590 -1300
rect 19700 -1060 19760 -1000
rect 19700 -1160 19760 -1100
rect 19700 -1260 19760 -1200
rect 19700 -1360 19760 -1300
rect 19870 -1060 19930 -1000
rect 19870 -1160 19930 -1100
rect 19870 -1260 19930 -1200
rect 19870 -1360 19930 -1300
rect 20040 -1060 20100 -1000
rect 20040 -1160 20100 -1100
rect 20040 -1260 20100 -1200
rect 20040 -1360 20100 -1300
rect 20210 -1060 20270 -1000
rect 20210 -1160 20270 -1100
rect 20210 -1260 20270 -1200
rect 20210 -1360 20270 -1300
rect 20380 -1060 20440 -1000
rect 20380 -1160 20440 -1100
rect 20380 -1260 20440 -1200
rect 20380 -1360 20440 -1300
rect 20550 -1060 20610 -1000
rect 20550 -1160 20610 -1100
rect 20550 -1260 20610 -1200
rect 20550 -1360 20610 -1300
rect 20720 -1060 20780 -1000
rect 20720 -1160 20780 -1100
rect 20720 -1260 20780 -1200
rect 20720 -1360 20780 -1300
rect 20890 -1060 20950 -1000
rect 20890 -1160 20950 -1100
rect 20890 -1260 20950 -1200
rect 20890 -1360 20950 -1300
rect 21060 -1060 21120 -1000
rect 21060 -1160 21120 -1100
rect 21060 -1260 21120 -1200
rect 21060 -1360 21120 -1300
rect 21230 -1060 21290 -1000
rect 21230 -1160 21290 -1100
rect 21230 -1260 21290 -1200
rect 21230 -1360 21290 -1300
rect 21400 -1060 21460 -1000
rect 21400 -1160 21460 -1100
rect 21400 -1260 21460 -1200
rect 21400 -1360 21460 -1300
rect 21570 -1060 21630 -1000
rect 21570 -1160 21630 -1100
rect 21570 -1260 21630 -1200
rect 21570 -1360 21630 -1300
rect 21740 -1060 21800 -1000
rect 21740 -1160 21800 -1100
rect 21740 -1260 21800 -1200
rect 21740 -1360 21800 -1300
rect 21910 -1060 21970 -1000
rect 21910 -1160 21970 -1100
rect 21910 -1260 21970 -1200
rect 21910 -1360 21970 -1300
rect 22080 -1060 22140 -1000
rect 22080 -1160 22140 -1100
rect 22080 -1260 22140 -1200
rect 22080 -1360 22140 -1300
rect 22250 -1060 22310 -1000
rect 22250 -1160 22310 -1100
rect 22250 -1260 22310 -1200
rect 22250 -1360 22310 -1300
rect 22420 -1060 22480 -1000
rect 22420 -1160 22480 -1100
rect 22420 -1260 22480 -1200
rect 22420 -1360 22480 -1300
rect 22590 -1060 22650 -1000
rect 22590 -1160 22650 -1100
rect 22590 -1260 22650 -1200
rect 22590 -1360 22650 -1300
rect 22760 -1060 22820 -1000
rect 22760 -1160 22820 -1100
rect 22760 -1260 22820 -1200
rect 22760 -1360 22820 -1300
rect 22930 -1060 22990 -1000
rect 22930 -1160 22990 -1100
rect 22930 -1260 22990 -1200
rect 22930 -1360 22990 -1300
rect 23100 -1060 23160 -1000
rect 23100 -1160 23160 -1100
rect 23100 -1260 23160 -1200
rect 23100 -1360 23160 -1300
rect 23270 -1060 23330 -1000
rect 23270 -1160 23330 -1100
rect 23270 -1260 23330 -1200
rect 23270 -1360 23330 -1300
rect 23440 -1060 23500 -1000
rect 23440 -1160 23500 -1100
rect 23440 -1260 23500 -1200
rect 23440 -1360 23500 -1300
rect 23610 -1060 23670 -1000
rect 23610 -1160 23670 -1100
rect 23610 -1260 23670 -1200
rect 23610 -1360 23670 -1300
rect 23780 -1060 23840 -1000
rect 23780 -1160 23840 -1100
rect 23780 -1260 23840 -1200
rect 23780 -1360 23840 -1300
rect 23950 -1060 24010 -1000
rect 23950 -1160 24010 -1100
rect 23950 -1260 24010 -1200
rect 23950 -1360 24010 -1300
rect 24120 -1060 24180 -1000
rect 24120 -1160 24180 -1100
rect 24120 -1260 24180 -1200
rect 24120 -1360 24180 -1300
rect 24290 -1060 24350 -1000
rect 24290 -1160 24350 -1100
rect 24290 -1260 24350 -1200
rect 24290 -1360 24350 -1300
rect 24460 -1060 24520 -1000
rect 24460 -1160 24520 -1100
rect 24460 -1260 24520 -1200
rect 24460 -1360 24520 -1300
rect 24630 -1060 24690 -1000
rect 24630 -1160 24690 -1100
rect 24630 -1260 24690 -1200
rect 24630 -1360 24690 -1300
rect 24800 -1060 24860 -1000
rect 24800 -1160 24860 -1100
rect 24800 -1260 24860 -1200
rect 24800 -1360 24860 -1300
rect 24970 -1060 25030 -1000
rect 24970 -1160 25030 -1100
rect 24970 -1260 25030 -1200
rect 24970 -1360 25030 -1300
rect 25140 -1060 25200 -1000
rect 25140 -1160 25200 -1100
rect 25140 -1260 25200 -1200
rect 25140 -1360 25200 -1300
rect 25310 -1060 25370 -1000
rect 25310 -1160 25370 -1100
rect 25310 -1260 25370 -1200
rect 25310 -1360 25370 -1300
rect 25480 -1060 25540 -1000
rect 25480 -1160 25540 -1100
rect 25480 -1260 25540 -1200
rect 25480 -1360 25540 -1300
rect 25650 -1060 25710 -1000
rect 25650 -1160 25710 -1100
rect 25650 -1260 25710 -1200
rect 25650 -1360 25710 -1300
rect 25820 -1060 25880 -1000
rect 25820 -1160 25880 -1100
rect 25820 -1260 25880 -1200
rect 25820 -1360 25880 -1300
rect 25990 -1060 26050 -1000
rect 25990 -1160 26050 -1100
rect 25990 -1260 26050 -1200
rect 25990 -1360 26050 -1300
rect 26160 -1060 26220 -1000
rect 26160 -1160 26220 -1100
rect 26160 -1260 26220 -1200
rect 26160 -1360 26220 -1300
rect 26330 -1060 26390 -1000
rect 26330 -1160 26390 -1100
rect 26330 -1260 26390 -1200
rect 26330 -1360 26390 -1300
rect 26500 -1060 26560 -1000
rect 26500 -1160 26560 -1100
rect 26500 -1260 26560 -1200
rect 26500 -1360 26560 -1300
rect 26670 -1060 26730 -1000
rect 26670 -1160 26730 -1100
rect 26670 -1260 26730 -1200
rect 26670 -1360 26730 -1300
rect 26840 -1060 26900 -1000
rect 26840 -1160 26900 -1100
rect 26840 -1260 26900 -1200
rect 26840 -1360 26900 -1300
rect 27010 -1060 27070 -1000
rect 27010 -1160 27070 -1100
rect 27010 -1260 27070 -1200
rect 27010 -1360 27070 -1300
rect 27180 -1060 27240 -1000
rect 27180 -1160 27240 -1100
rect 27180 -1260 27240 -1200
rect 27180 -1360 27240 -1300
rect 27350 -1060 27410 -1000
rect 27350 -1160 27410 -1100
rect 27350 -1260 27410 -1200
rect 27350 -1360 27410 -1300
rect 27520 -1060 27580 -1000
rect 27520 -1160 27580 -1100
rect 27520 -1260 27580 -1200
rect 27520 -1360 27580 -1300
rect 27690 -1060 27750 -1000
rect 27690 -1160 27750 -1100
rect 27690 -1260 27750 -1200
rect 27690 -1360 27750 -1300
rect 27860 -1060 27920 -1000
rect 27860 -1160 27920 -1100
rect 27860 -1260 27920 -1200
rect 27860 -1360 27920 -1300
rect 28030 -1060 28090 -1000
rect 28030 -1160 28090 -1100
rect 28030 -1260 28090 -1200
rect 28030 -1360 28090 -1300
rect 28200 -1060 28260 -1000
rect 28200 -1160 28260 -1100
rect 28200 -1260 28260 -1200
rect 28200 -1360 28260 -1300
rect 28370 -1060 28430 -1000
rect 28370 -1160 28430 -1100
rect 28370 -1260 28430 -1200
rect 28370 -1360 28430 -1300
rect 28540 -1060 28600 -1000
rect 28540 -1160 28600 -1100
rect 28540 -1260 28600 -1200
rect 28540 -1360 28600 -1300
rect 28710 -1060 28770 -1000
rect 28710 -1160 28770 -1100
rect 28710 -1260 28770 -1200
rect 28710 -1360 28770 -1300
rect 28880 -1060 28940 -1000
rect 28880 -1160 28940 -1100
rect 28880 -1260 28940 -1200
rect 28880 -1360 28940 -1300
rect 29050 -1060 29110 -1000
rect 29050 -1160 29110 -1100
rect 29050 -1260 29110 -1200
rect 29050 -1360 29110 -1300
rect 29220 -1060 29280 -1000
rect 29220 -1160 29280 -1100
rect 29220 -1260 29280 -1200
rect 29220 -1360 29280 -1300
rect 29390 -1060 29450 -1000
rect 29390 -1160 29450 -1100
rect 29390 -1260 29450 -1200
rect 29390 -1360 29450 -1300
rect 29560 -1060 29620 -1000
rect 29560 -1160 29620 -1100
rect 29560 -1260 29620 -1200
rect 29560 -1360 29620 -1300
rect 29730 -1060 29790 -1000
rect 29730 -1160 29790 -1100
rect 29730 -1260 29790 -1200
rect 29730 -1360 29790 -1300
rect 29900 -1060 29960 -1000
rect 29900 -1160 29960 -1100
rect 29900 -1260 29960 -1200
rect 29900 -1360 29960 -1300
rect 30070 -1060 30130 -1000
rect 30070 -1160 30130 -1100
rect 30070 -1260 30130 -1200
rect 30070 -1360 30130 -1300
rect 30240 -1060 30300 -1000
rect 30240 -1160 30300 -1100
rect 30240 -1260 30300 -1200
rect 30240 -1360 30300 -1300
rect 30410 -1060 30470 -1000
rect 30410 -1160 30470 -1100
rect 30410 -1260 30470 -1200
rect 30410 -1360 30470 -1300
rect 30580 -1060 30640 -1000
rect 30580 -1160 30640 -1100
rect 30580 -1260 30640 -1200
rect 30580 -1360 30640 -1300
rect 30750 -1060 30810 -1000
rect 30750 -1160 30810 -1100
rect 30750 -1260 30810 -1200
rect 30750 -1360 30810 -1300
rect 30920 -1060 30980 -1000
rect 30920 -1160 30980 -1100
rect 30920 -1260 30980 -1200
rect 30920 -1360 30980 -1300
rect 31090 -1060 31150 -1000
rect 31090 -1160 31150 -1100
rect 31090 -1260 31150 -1200
rect 31090 -1360 31150 -1300
rect 31260 -1060 31320 -1000
rect 31260 -1160 31320 -1100
rect 31260 -1260 31320 -1200
rect 31260 -1360 31320 -1300
rect 31430 -1060 31490 -1000
rect 31430 -1160 31490 -1100
rect 31430 -1260 31490 -1200
rect 31430 -1360 31490 -1300
rect 31600 -1060 31660 -1000
rect 31600 -1160 31660 -1100
rect 31600 -1260 31660 -1200
rect 31600 -1360 31660 -1300
rect 31770 -1060 31830 -1000
rect 31770 -1160 31830 -1100
rect 31770 -1260 31830 -1200
rect 31770 -1360 31830 -1300
rect 31940 -1060 32000 -1000
rect 31940 -1160 32000 -1100
rect 31940 -1260 32000 -1200
rect 31940 -1360 32000 -1300
rect 32110 -1060 32170 -1000
rect 32110 -1160 32170 -1100
rect 32110 -1260 32170 -1200
rect 32110 -1360 32170 -1300
rect 32280 -1060 32340 -1000
rect 32280 -1160 32340 -1100
rect 32280 -1260 32340 -1200
rect 32280 -1360 32340 -1300
rect 32450 -1060 32510 -1000
rect 32450 -1160 32510 -1100
rect 32450 -1260 32510 -1200
rect 32450 -1360 32510 -1300
rect 32620 -1060 32680 -1000
rect 32620 -1160 32680 -1100
rect 32620 -1260 32680 -1200
rect 32620 -1360 32680 -1300
rect 32790 -1060 32850 -1000
rect 32790 -1160 32850 -1100
rect 32790 -1260 32850 -1200
rect 32790 -1360 32850 -1300
rect 32960 -1060 33020 -1000
rect 32960 -1160 33020 -1100
rect 32960 -1260 33020 -1200
rect 32960 -1360 33020 -1300
rect 33130 -1060 33190 -1000
rect 33130 -1160 33190 -1100
rect 33130 -1260 33190 -1200
rect 33130 -1360 33190 -1300
rect 33300 -1060 33360 -1000
rect 33300 -1160 33360 -1100
rect 33300 -1260 33360 -1200
rect 33300 -1360 33360 -1300
rect 33470 -1060 33530 -1000
rect 33470 -1160 33530 -1100
rect 33470 -1260 33530 -1200
rect 33470 -1360 33530 -1300
rect 33640 -1060 33700 -1000
rect 33640 -1160 33700 -1100
rect 33640 -1260 33700 -1200
rect 33640 -1360 33700 -1300
rect 33810 -1060 33870 -1000
rect 33810 -1160 33870 -1100
rect 33810 -1260 33870 -1200
rect 33810 -1360 33870 -1300
rect 33980 -1060 34040 -1000
rect 33980 -1160 34040 -1100
rect 33980 -1260 34040 -1200
rect 33980 -1360 34040 -1300
rect 34150 -1060 34210 -1000
rect 34150 -1160 34210 -1100
rect 34150 -1260 34210 -1200
rect 34150 -1360 34210 -1300
rect 34320 -1060 34380 -1000
rect 34320 -1160 34380 -1100
rect 34320 -1260 34380 -1200
rect 34320 -1360 34380 -1300
rect 34490 -1060 34550 -1000
rect 34490 -1160 34550 -1100
rect 34490 -1260 34550 -1200
rect 34490 -1360 34550 -1300
rect 34660 -1060 34720 -1000
rect 34660 -1160 34720 -1100
rect 34660 -1260 34720 -1200
rect 34660 -1360 34720 -1300
rect 34830 -1060 34890 -1000
rect 34830 -1160 34890 -1100
rect 34830 -1260 34890 -1200
rect 34830 -1360 34890 -1300
rect 35000 -1060 35060 -1000
rect 35000 -1160 35060 -1100
rect 35000 -1260 35060 -1200
rect 35000 -1360 35060 -1300
rect 35170 -1060 35230 -1000
rect 35170 -1160 35230 -1100
rect 35170 -1260 35230 -1200
rect 35170 -1360 35230 -1300
rect 35340 -1060 35400 -1000
rect 35340 -1160 35400 -1100
rect 35340 -1260 35400 -1200
rect 35340 -1360 35400 -1300
rect 35510 -1060 35570 -1000
rect 35510 -1160 35570 -1100
rect 35510 -1260 35570 -1200
rect 35510 -1360 35570 -1300
rect 35680 -1060 35740 -1000
rect 35680 -1160 35740 -1100
rect 35680 -1260 35740 -1200
rect 35680 -1360 35740 -1300
rect 35850 -1060 35910 -1000
rect 35850 -1160 35910 -1100
rect 35850 -1260 35910 -1200
rect 35850 -1360 35910 -1300
rect 36020 -1060 36080 -1000
rect 36020 -1160 36080 -1100
rect 36020 -1260 36080 -1200
rect 36020 -1360 36080 -1300
rect 36190 -1060 36250 -1000
rect 36190 -1160 36250 -1100
rect 36190 -1260 36250 -1200
rect 36190 -1360 36250 -1300
rect 36360 -1060 36420 -1000
rect 36360 -1160 36420 -1100
rect 36360 -1260 36420 -1200
rect 36360 -1360 36420 -1300
rect 36530 -1060 36590 -1000
rect 36530 -1160 36590 -1100
rect 36530 -1260 36590 -1200
rect 36530 -1360 36590 -1300
rect 36700 -1060 36760 -1000
rect 36700 -1160 36760 -1100
rect 36700 -1260 36760 -1200
rect 36700 -1360 36760 -1300
rect 36870 -1060 36930 -1000
rect 36870 -1160 36930 -1100
rect 36870 -1260 36930 -1200
rect 36870 -1360 36930 -1300
rect 37040 -1060 37100 -1000
rect 37040 -1160 37100 -1100
rect 37040 -1260 37100 -1200
rect 37040 -1360 37100 -1300
rect 37210 -1060 37270 -1000
rect 37210 -1160 37270 -1100
rect 37210 -1260 37270 -1200
rect 37210 -1360 37270 -1300
rect 37380 -1060 37440 -1000
rect 37380 -1160 37440 -1100
rect 37380 -1260 37440 -1200
rect 37380 -1360 37440 -1300
rect 37550 -1060 37610 -1000
rect 37550 -1160 37610 -1100
rect 37550 -1260 37610 -1200
rect 37550 -1360 37610 -1300
rect 37720 -1060 37780 -1000
rect 37720 -1160 37780 -1100
rect 37720 -1260 37780 -1200
rect 37720 -1360 37780 -1300
rect 37890 -1060 37950 -1000
rect 37890 -1160 37950 -1100
rect 37890 -1260 37950 -1200
rect 37890 -1360 37950 -1300
rect 38060 -1060 38120 -1000
rect 38060 -1160 38120 -1100
rect 38060 -1260 38120 -1200
rect 38060 -1360 38120 -1300
rect 38230 -1060 38290 -1000
rect 38230 -1160 38290 -1100
rect 38230 -1260 38290 -1200
rect 38230 -1360 38290 -1300
rect 38400 -1060 38460 -1000
rect 38400 -1160 38460 -1100
rect 38400 -1260 38460 -1200
rect 38400 -1360 38460 -1300
rect 38570 -1060 38630 -1000
rect 38570 -1160 38630 -1100
rect 38570 -1260 38630 -1200
rect 38570 -1360 38630 -1300
rect 38740 -1060 38800 -1000
rect 38740 -1160 38800 -1100
rect 38740 -1260 38800 -1200
rect 38740 -1360 38800 -1300
rect 38910 -1060 38970 -1000
rect 38910 -1160 38970 -1100
rect 38910 -1260 38970 -1200
rect 38910 -1360 38970 -1300
rect 39080 -1060 39140 -1000
rect 39080 -1160 39140 -1100
rect 39080 -1260 39140 -1200
rect 39080 -1360 39140 -1300
rect 39250 -1060 39310 -1000
rect 39250 -1160 39310 -1100
rect 39250 -1260 39310 -1200
rect 39250 -1360 39310 -1300
rect 39420 -1060 39480 -1000
rect 39420 -1160 39480 -1100
rect 39420 -1260 39480 -1200
rect 39420 -1360 39480 -1300
rect 39590 -1060 39650 -1000
rect 39590 -1160 39650 -1100
rect 39590 -1260 39650 -1200
rect 39590 -1360 39650 -1300
rect 39760 -1060 39820 -1000
rect 39760 -1160 39820 -1100
rect 39760 -1260 39820 -1200
rect 39760 -1360 39820 -1300
rect 39930 -1060 39990 -1000
rect 39930 -1160 39990 -1100
rect 39930 -1260 39990 -1200
rect 39930 -1360 39990 -1300
rect 40100 -1060 40160 -1000
rect 40100 -1160 40160 -1100
rect 40100 -1260 40160 -1200
rect 40100 -1360 40160 -1300
rect 40270 -1060 40330 -1000
rect 40270 -1160 40330 -1100
rect 40270 -1260 40330 -1200
rect 40270 -1360 40330 -1300
rect 40440 -1060 40500 -1000
rect 40440 -1160 40500 -1100
rect 40440 -1260 40500 -1200
rect 40440 -1360 40500 -1300
rect 40610 -1060 40670 -1000
rect 40610 -1160 40670 -1100
rect 40610 -1260 40670 -1200
rect 40610 -1360 40670 -1300
rect 40780 -1060 40840 -1000
rect 40780 -1160 40840 -1100
rect 40780 -1260 40840 -1200
rect 40780 -1360 40840 -1300
rect 40950 -1060 41010 -1000
rect 40950 -1160 41010 -1100
rect 40950 -1260 41010 -1200
rect 40950 -1360 41010 -1300
rect 41120 -1060 41180 -1000
rect 41120 -1160 41180 -1100
rect 41120 -1260 41180 -1200
rect 41120 -1360 41180 -1300
rect 41290 -1060 41350 -1000
rect 41290 -1160 41350 -1100
rect 41290 -1260 41350 -1200
rect 41290 -1360 41350 -1300
rect 41460 -1060 41520 -1000
rect 41460 -1160 41520 -1100
rect 41460 -1260 41520 -1200
rect 41460 -1360 41520 -1300
rect 41630 -1060 41690 -1000
rect 41630 -1160 41690 -1100
rect 41630 -1260 41690 -1200
rect 41630 -1360 41690 -1300
rect 41800 -1060 41860 -1000
rect 41800 -1160 41860 -1100
rect 41800 -1260 41860 -1200
rect 41800 -1360 41860 -1300
rect 41970 -1060 42030 -1000
rect 41970 -1160 42030 -1100
rect 41970 -1260 42030 -1200
rect 41970 -1360 42030 -1300
rect 42140 -1060 42200 -1000
rect 42140 -1160 42200 -1100
rect 42140 -1260 42200 -1200
rect 42140 -1360 42200 -1300
rect 42310 -1060 42370 -1000
rect 42310 -1160 42370 -1100
rect 42310 -1260 42370 -1200
rect 42310 -1360 42370 -1300
rect 42480 -1060 42540 -1000
rect 42480 -1160 42540 -1100
rect 42480 -1260 42540 -1200
rect 42480 -1360 42540 -1300
rect 42650 -1060 42710 -1000
rect 42650 -1160 42710 -1100
rect 42650 -1260 42710 -1200
rect 42650 -1360 42710 -1300
rect 42820 -1060 42880 -1000
rect 42820 -1160 42880 -1100
rect 42820 -1260 42880 -1200
rect 42820 -1360 42880 -1300
rect 42990 -1060 43050 -1000
rect 42990 -1160 43050 -1100
rect 42990 -1260 43050 -1200
rect 42990 -1360 43050 -1300
rect 43160 -1060 43220 -1000
rect 43160 -1160 43220 -1100
rect 43160 -1260 43220 -1200
rect 43160 -1360 43220 -1300
rect 43330 -1060 43390 -1000
rect 43330 -1160 43390 -1100
rect 43330 -1260 43390 -1200
rect 43330 -1360 43390 -1300
rect 43500 -1060 43560 -1000
rect 43500 -1160 43560 -1100
rect 43500 -1260 43560 -1200
rect 43500 -1360 43560 -1300
rect 43670 -1060 43730 -1000
rect 43670 -1160 43730 -1100
rect 43670 -1260 43730 -1200
rect 43670 -1360 43730 -1300
rect 43840 -1060 43900 -1000
rect 43840 -1160 43900 -1100
rect 43840 -1260 43900 -1200
rect 43840 -1360 43900 -1300
rect 44010 -1060 44070 -1000
rect 44010 -1160 44070 -1100
rect 44010 -1260 44070 -1200
rect 44010 -1360 44070 -1300
rect 44180 -1060 44240 -1000
rect 44180 -1160 44240 -1100
rect 44180 -1260 44240 -1200
rect 44180 -1360 44240 -1300
rect 44350 -1060 44410 -1000
rect 44350 -1160 44410 -1100
rect 44350 -1260 44410 -1200
rect 44350 -1360 44410 -1300
rect 44520 -1060 44580 -1000
rect 44520 -1160 44580 -1100
rect 44520 -1260 44580 -1200
rect 44520 -1360 44580 -1300
rect 44690 -1060 44750 -1000
rect 44690 -1160 44750 -1100
rect 44690 -1260 44750 -1200
rect 44690 -1360 44750 -1300
rect 44860 -1060 44920 -1000
rect 44860 -1160 44920 -1100
rect 44860 -1260 44920 -1200
rect 44860 -1360 44920 -1300
rect 45030 -1060 45090 -1000
rect 45030 -1160 45090 -1100
rect 45030 -1260 45090 -1200
rect 45030 -1360 45090 -1300
rect 45200 -1060 45260 -1000
rect 45200 -1160 45260 -1100
rect 45200 -1260 45260 -1200
rect 45200 -1360 45260 -1300
rect 45370 -1060 45430 -1000
rect 45370 -1160 45430 -1100
rect 45370 -1260 45430 -1200
rect 45370 -1360 45430 -1300
rect 45540 -1060 45600 -1000
rect 45540 -1160 45600 -1100
rect 45540 -1260 45600 -1200
rect 45540 -1360 45600 -1300
rect 45710 -1060 45770 -1000
rect 45710 -1160 45770 -1100
rect 45710 -1260 45770 -1200
rect 45710 -1360 45770 -1300
rect 45880 -1060 45940 -1000
rect 45880 -1160 45940 -1100
rect 45880 -1260 45940 -1200
rect 45880 -1360 45940 -1300
rect 46050 -1060 46110 -1000
rect 46050 -1160 46110 -1100
rect 46050 -1260 46110 -1200
rect 46050 -1360 46110 -1300
rect 46220 -1060 46280 -1000
rect 46220 -1160 46280 -1100
rect 46220 -1260 46280 -1200
rect 46220 -1360 46280 -1300
rect 46390 -1060 46450 -1000
rect 46390 -1160 46450 -1100
rect 46390 -1260 46450 -1200
rect 46390 -1360 46450 -1300
rect 46560 -1060 46620 -1000
rect 46560 -1160 46620 -1100
rect 46560 -1260 46620 -1200
rect 46560 -1360 46620 -1300
rect 46730 -1060 46790 -1000
rect 46730 -1160 46790 -1100
rect 46730 -1260 46790 -1200
rect 46730 -1360 46790 -1300
rect 46900 -1060 46960 -1000
rect 46900 -1160 46960 -1100
rect 46900 -1260 46960 -1200
rect 46900 -1360 46960 -1300
rect 47070 -1060 47130 -1000
rect 47070 -1160 47130 -1100
rect 47070 -1260 47130 -1200
rect 47070 -1360 47130 -1300
rect 47240 -1060 47300 -1000
rect 47240 -1160 47300 -1100
rect 47240 -1260 47300 -1200
rect 47240 -1360 47300 -1300
rect 47410 -1060 47470 -1000
rect 47410 -1160 47470 -1100
rect 47410 -1260 47470 -1200
rect 47410 -1360 47470 -1300
rect 47580 -1060 47640 -1000
rect 47580 -1160 47640 -1100
rect 47580 -1260 47640 -1200
rect 47580 -1360 47640 -1300
rect 47750 -1060 47810 -1000
rect 47750 -1160 47810 -1100
rect 47750 -1260 47810 -1200
rect 47750 -1360 47810 -1300
rect 47920 -1060 47980 -1000
rect 47920 -1160 47980 -1100
rect 47920 -1260 47980 -1200
rect 47920 -1360 47980 -1300
rect 48090 -1060 48150 -1000
rect 48090 -1160 48150 -1100
rect 48090 -1260 48150 -1200
rect 48090 -1360 48150 -1300
rect 48260 -1060 48320 -1000
rect 48260 -1160 48320 -1100
rect 48260 -1260 48320 -1200
rect 48260 -1360 48320 -1300
rect 48430 -1060 48490 -1000
rect 48430 -1160 48490 -1100
rect 48430 -1260 48490 -1200
rect 48430 -1360 48490 -1300
rect 48600 -1060 48660 -1000
rect 48600 -1160 48660 -1100
rect 48600 -1260 48660 -1200
rect 48600 -1360 48660 -1300
rect 48770 -1060 48830 -1000
rect 48770 -1160 48830 -1100
rect 48770 -1260 48830 -1200
rect 48770 -1360 48830 -1300
rect 48940 -1060 49000 -1000
rect 48940 -1160 49000 -1100
rect 48940 -1260 49000 -1200
rect 48940 -1360 49000 -1300
rect 49110 -1060 49170 -1000
rect 49110 -1160 49170 -1100
rect 49110 -1260 49170 -1200
rect 49110 -1360 49170 -1300
rect 49280 -1060 49340 -1000
rect 49280 -1160 49340 -1100
rect 49280 -1260 49340 -1200
rect 49280 -1360 49340 -1300
rect 49450 -1060 49510 -1000
rect 49450 -1160 49510 -1100
rect 49450 -1260 49510 -1200
rect 49450 -1360 49510 -1300
rect 49620 -1060 49680 -1000
rect 49620 -1160 49680 -1100
rect 49620 -1260 49680 -1200
rect 49620 -1360 49680 -1300
rect 49790 -1060 49850 -1000
rect 49790 -1160 49850 -1100
rect 49790 -1260 49850 -1200
rect 49790 -1360 49850 -1300
rect 49960 -1060 50020 -1000
rect 49960 -1160 50020 -1100
rect 49960 -1260 50020 -1200
rect 49960 -1360 50020 -1300
rect 50130 -1060 50190 -1000
rect 50130 -1160 50190 -1100
rect 50130 -1260 50190 -1200
rect 50130 -1360 50190 -1300
rect 50300 -1060 50360 -1000
rect 50300 -1160 50360 -1100
rect 50300 -1260 50360 -1200
rect 50300 -1360 50360 -1300
rect 50470 -1060 50530 -1000
rect 50470 -1160 50530 -1100
rect 50470 -1260 50530 -1200
rect 50470 -1360 50530 -1300
rect 50640 -1060 50700 -1000
rect 50640 -1160 50700 -1100
rect 50640 -1260 50700 -1200
rect 50640 -1360 50700 -1300
rect 50810 -1060 50870 -1000
rect 50810 -1160 50870 -1100
rect 50810 -1260 50870 -1200
rect 50810 -1360 50870 -1300
rect 50980 -1060 51040 -1000
rect 50980 -1160 51040 -1100
rect 50980 -1260 51040 -1200
rect 50980 -1360 51040 -1300
rect 51150 -1060 51210 -1000
rect 51150 -1160 51210 -1100
rect 51150 -1260 51210 -1200
rect 51150 -1360 51210 -1300
rect 51320 -1060 51380 -1000
rect 51320 -1160 51380 -1100
rect 51320 -1260 51380 -1200
rect 51320 -1360 51380 -1300
rect 51490 -1060 51550 -1000
rect 51490 -1160 51550 -1100
rect 51490 -1260 51550 -1200
rect 51490 -1360 51550 -1300
rect 51660 -1060 51720 -1000
rect 51660 -1160 51720 -1100
rect 51660 -1260 51720 -1200
rect 51660 -1360 51720 -1300
rect 51830 -1060 51890 -1000
rect 51830 -1160 51890 -1100
rect 51830 -1260 51890 -1200
rect 51830 -1360 51890 -1300
rect 52000 -1060 52060 -1000
rect 52000 -1160 52060 -1100
rect 52000 -1260 52060 -1200
rect 52000 -1360 52060 -1300
rect 52170 -1060 52230 -1000
rect 52170 -1160 52230 -1100
rect 52170 -1260 52230 -1200
rect 52170 -1360 52230 -1300
rect 52340 -1060 52400 -1000
rect 52340 -1160 52400 -1100
rect 52340 -1260 52400 -1200
rect 52340 -1360 52400 -1300
rect 52510 -1060 52570 -1000
rect 52510 -1160 52570 -1100
rect 52510 -1260 52570 -1200
rect 52510 -1360 52570 -1300
rect 52680 -1060 52740 -1000
rect 52680 -1160 52740 -1100
rect 52680 -1260 52740 -1200
rect 52680 -1360 52740 -1300
rect 52850 -1060 52910 -1000
rect 52850 -1160 52910 -1100
rect 52850 -1260 52910 -1200
rect 52850 -1360 52910 -1300
rect 53020 -1060 53080 -1000
rect 53020 -1160 53080 -1100
rect 53020 -1260 53080 -1200
rect 53020 -1360 53080 -1300
rect 53190 -1060 53250 -1000
rect 53190 -1160 53250 -1100
rect 53190 -1260 53250 -1200
rect 53190 -1360 53250 -1300
rect 53360 -1060 53420 -1000
rect 53360 -1160 53420 -1100
rect 53360 -1260 53420 -1200
rect 53360 -1360 53420 -1300
rect 53530 -1060 53590 -1000
rect 53530 -1160 53590 -1100
rect 53530 -1260 53590 -1200
rect 53530 -1360 53590 -1300
rect 53700 -1060 53760 -1000
rect 53700 -1160 53760 -1100
rect 53700 -1260 53760 -1200
rect 53700 -1360 53760 -1300
rect 53870 -1060 53930 -1000
rect 53870 -1160 53930 -1100
rect 53870 -1260 53930 -1200
rect 53870 -1360 53930 -1300
rect 54040 -1060 54100 -1000
rect 54040 -1160 54100 -1100
rect 54040 -1260 54100 -1200
rect 54040 -1360 54100 -1300
rect 54210 -1060 54270 -1000
rect 54210 -1160 54270 -1100
rect 54210 -1260 54270 -1200
rect 54210 -1360 54270 -1300
rect 54380 -1060 54440 -1000
rect 54380 -1160 54440 -1100
rect 54380 -1260 54440 -1200
rect 54380 -1360 54440 -1300
rect 54550 -1060 54610 -1000
rect 54550 -1160 54610 -1100
rect 54550 -1260 54610 -1200
rect 54550 -1360 54610 -1300
rect 54720 -1060 54780 -1000
rect 54720 -1160 54780 -1100
rect 54720 -1260 54780 -1200
rect 54720 -1360 54780 -1300
rect 54890 -1060 54950 -1000
rect 54890 -1160 54950 -1100
rect 54890 -1260 54950 -1200
rect 54890 -1360 54950 -1300
rect 55060 -1060 55120 -1000
rect 55060 -1160 55120 -1100
rect 55060 -1260 55120 -1200
rect 55060 -1360 55120 -1300
rect 55230 -1060 55290 -1000
rect 55230 -1160 55290 -1100
rect 55230 -1260 55290 -1200
rect 55230 -1360 55290 -1300
rect 55400 -1060 55460 -1000
rect 55400 -1160 55460 -1100
rect 55400 -1260 55460 -1200
rect 55400 -1360 55460 -1300
rect 55570 -1060 55630 -1000
rect 55570 -1160 55630 -1100
rect 55570 -1260 55630 -1200
rect 55570 -1360 55630 -1300
rect 55740 -1060 55800 -1000
rect 55740 -1160 55800 -1100
rect 55740 -1260 55800 -1200
rect 55740 -1360 55800 -1300
rect 55910 -1060 55970 -1000
rect 55910 -1160 55970 -1100
rect 55910 -1260 55970 -1200
rect 55910 -1360 55970 -1300
rect 56080 -1060 56140 -1000
rect 56080 -1160 56140 -1100
rect 56080 -1260 56140 -1200
rect 56080 -1360 56140 -1300
rect 56250 -1060 56310 -1000
rect 56250 -1160 56310 -1100
rect 56250 -1260 56310 -1200
rect 56250 -1360 56310 -1300
rect 56420 -1060 56480 -1000
rect 56420 -1160 56480 -1100
rect 56420 -1260 56480 -1200
rect 56420 -1360 56480 -1300
rect 56590 -1060 56650 -1000
rect 56590 -1160 56650 -1100
rect 56590 -1260 56650 -1200
rect 56590 -1360 56650 -1300
rect 56760 -1060 56820 -1000
rect 56760 -1160 56820 -1100
rect 56760 -1260 56820 -1200
rect 56760 -1360 56820 -1300
rect 56930 -1060 56990 -1000
rect 56930 -1160 56990 -1100
rect 56930 -1260 56990 -1200
rect 56930 -1360 56990 -1300
rect 57100 -1060 57160 -1000
rect 57100 -1160 57160 -1100
rect 57100 -1260 57160 -1200
rect 57100 -1360 57160 -1300
rect 57270 -1060 57330 -1000
rect 57270 -1160 57330 -1100
rect 57270 -1260 57330 -1200
rect 57270 -1360 57330 -1300
rect 57440 -1060 57500 -1000
rect 57440 -1160 57500 -1100
rect 57440 -1260 57500 -1200
rect 57440 -1360 57500 -1300
rect 57610 -1060 57670 -1000
rect 57610 -1160 57670 -1100
rect 57610 -1260 57670 -1200
rect 57610 -1360 57670 -1300
rect 57780 -1060 57840 -1000
rect 57780 -1160 57840 -1100
rect 57780 -1260 57840 -1200
rect 57780 -1360 57840 -1300
rect 57950 -1060 58010 -1000
rect 57950 -1160 58010 -1100
rect 57950 -1260 58010 -1200
rect 57950 -1360 58010 -1300
rect 58120 -1060 58180 -1000
rect 58120 -1160 58180 -1100
rect 58120 -1260 58180 -1200
rect 58120 -1360 58180 -1300
rect 58290 -1060 58350 -1000
rect 58290 -1160 58350 -1100
rect 58290 -1260 58350 -1200
rect 58290 -1360 58350 -1300
rect 58460 -1060 58520 -1000
rect 58460 -1160 58520 -1100
rect 58460 -1260 58520 -1200
rect 58460 -1360 58520 -1300
rect 58630 -1060 58690 -1000
rect 58630 -1160 58690 -1100
rect 58630 -1260 58690 -1200
rect 58630 -1360 58690 -1300
rect 58800 -1060 58860 -1000
rect 58800 -1160 58860 -1100
rect 58800 -1260 58860 -1200
rect 58800 -1360 58860 -1300
rect 58970 -1060 59030 -1000
rect 58970 -1160 59030 -1100
rect 58970 -1260 59030 -1200
rect 58970 -1360 59030 -1300
rect 59140 -1060 59200 -1000
rect 59140 -1160 59200 -1100
rect 59140 -1260 59200 -1200
rect 59140 -1360 59200 -1300
rect 59310 -1060 59370 -1000
rect 59310 -1160 59370 -1100
rect 59310 -1260 59370 -1200
rect 59310 -1360 59370 -1300
rect 59480 -1060 59540 -1000
rect 59480 -1160 59540 -1100
rect 59480 -1260 59540 -1200
rect 59480 -1360 59540 -1300
rect 59650 -1060 59710 -1000
rect 59650 -1160 59710 -1100
rect 59650 -1260 59710 -1200
rect 59650 -1360 59710 -1300
rect 59820 -1060 59880 -1000
rect 59820 -1160 59880 -1100
rect 59820 -1260 59880 -1200
rect 59820 -1360 59880 -1300
rect 59990 -1060 60050 -1000
rect 59990 -1160 60050 -1100
rect 59990 -1260 60050 -1200
rect 59990 -1360 60050 -1300
rect 60160 -1060 60220 -1000
rect 60160 -1160 60220 -1100
rect 60160 -1260 60220 -1200
rect 60160 -1360 60220 -1300
rect 60330 -1060 60390 -1000
rect 60330 -1160 60390 -1100
rect 60330 -1260 60390 -1200
rect 60330 -1360 60390 -1300
rect 60500 -1060 60560 -1000
rect 60500 -1160 60560 -1100
rect 60500 -1260 60560 -1200
rect 60500 -1360 60560 -1300
rect 60670 -1060 60730 -1000
rect 60670 -1160 60730 -1100
rect 60670 -1260 60730 -1200
rect 60670 -1360 60730 -1300
rect 60840 -1060 60900 -1000
rect 60840 -1160 60900 -1100
rect 60840 -1260 60900 -1200
rect 60840 -1360 60900 -1300
rect 61010 -1060 61070 -1000
rect 61010 -1160 61070 -1100
rect 61010 -1260 61070 -1200
rect 61010 -1360 61070 -1300
rect 61180 -1060 61240 -1000
rect 61180 -1160 61240 -1100
rect 61180 -1260 61240 -1200
rect 61180 -1360 61240 -1300
rect 61350 -1060 61410 -1000
rect 61350 -1160 61410 -1100
rect 61350 -1260 61410 -1200
rect 61350 -1360 61410 -1300
rect 61520 -1060 61580 -1000
rect 61520 -1160 61580 -1100
rect 61520 -1260 61580 -1200
rect 61520 -1360 61580 -1300
rect 61690 -1060 61750 -1000
rect 61690 -1160 61750 -1100
rect 61690 -1260 61750 -1200
rect 61690 -1360 61750 -1300
rect 61860 -1060 61920 -1000
rect 61860 -1160 61920 -1100
rect 61860 -1260 61920 -1200
rect 61860 -1360 61920 -1300
rect 62030 -1060 62090 -1000
rect 62030 -1160 62090 -1100
rect 62030 -1260 62090 -1200
rect 62030 -1360 62090 -1300
rect 62200 -1060 62260 -1000
rect 62200 -1160 62260 -1100
rect 62200 -1260 62260 -1200
rect 62200 -1360 62260 -1300
rect 62370 -1060 62430 -1000
rect 62370 -1160 62430 -1100
rect 62370 -1260 62430 -1200
rect 62370 -1360 62430 -1300
rect 62540 -1060 62600 -1000
rect 62540 -1160 62600 -1100
rect 62540 -1260 62600 -1200
rect 62540 -1360 62600 -1300
rect 62710 -1060 62770 -1000
rect 62710 -1160 62770 -1100
rect 62710 -1260 62770 -1200
rect 62710 -1360 62770 -1300
rect 62880 -1060 62940 -1000
rect 62880 -1160 62940 -1100
rect 62880 -1260 62940 -1200
rect 62880 -1360 62940 -1300
rect 63050 -1060 63110 -1000
rect 63050 -1160 63110 -1100
rect 63050 -1260 63110 -1200
rect 63050 -1360 63110 -1300
rect 63220 -1060 63280 -1000
rect 63220 -1160 63280 -1100
rect 63220 -1260 63280 -1200
rect 63220 -1360 63280 -1300
rect 63390 -1060 63450 -1000
rect 63390 -1160 63450 -1100
rect 63390 -1260 63450 -1200
rect 63390 -1360 63450 -1300
rect 63560 -1060 63620 -1000
rect 63560 -1160 63620 -1100
rect 63560 -1260 63620 -1200
rect 63560 -1360 63620 -1300
rect 63730 -1060 63790 -1000
rect 63730 -1160 63790 -1100
rect 63730 -1260 63790 -1200
rect 63730 -1360 63790 -1300
rect 63900 -1060 63960 -1000
rect 63900 -1160 63960 -1100
rect 63900 -1260 63960 -1200
rect 63900 -1360 63960 -1300
rect 64070 -1060 64130 -1000
rect 64070 -1160 64130 -1100
rect 64070 -1260 64130 -1200
rect 64070 -1360 64130 -1300
rect 64240 -1060 64300 -1000
rect 64240 -1160 64300 -1100
rect 64240 -1260 64300 -1200
rect 64240 -1360 64300 -1300
rect 64410 -1060 64470 -1000
rect 64410 -1160 64470 -1100
rect 64410 -1260 64470 -1200
rect 64410 -1360 64470 -1300
rect 64580 -1060 64640 -1000
rect 64580 -1160 64640 -1100
rect 64580 -1260 64640 -1200
rect 64580 -1360 64640 -1300
rect 64750 -1060 64810 -1000
rect 64750 -1160 64810 -1100
rect 64750 -1260 64810 -1200
rect 64750 -1360 64810 -1300
rect 64920 -1060 64980 -1000
rect 64920 -1160 64980 -1100
rect 64920 -1260 64980 -1200
rect 64920 -1360 64980 -1300
rect 65090 -1060 65150 -1000
rect 65090 -1160 65150 -1100
rect 65090 -1260 65150 -1200
rect 65090 -1360 65150 -1300
rect 65260 -1060 65320 -1000
rect 65260 -1160 65320 -1100
rect 65260 -1260 65320 -1200
rect 65260 -1360 65320 -1300
rect 65430 -1060 65490 -1000
rect 65430 -1160 65490 -1100
rect 65430 -1260 65490 -1200
rect 65430 -1360 65490 -1300
rect 65600 -1060 65660 -1000
rect 65600 -1160 65660 -1100
rect 65600 -1260 65660 -1200
rect 65600 -1360 65660 -1300
rect 65770 -1060 65830 -1000
rect 65770 -1160 65830 -1100
rect 65770 -1260 65830 -1200
rect 65770 -1360 65830 -1300
rect 65940 -1060 66000 -1000
rect 65940 -1160 66000 -1100
rect 65940 -1260 66000 -1200
rect 65940 -1360 66000 -1300
rect 66110 -1060 66170 -1000
rect 66110 -1160 66170 -1100
rect 66110 -1260 66170 -1200
rect 66110 -1360 66170 -1300
rect 66280 -1060 66340 -1000
rect 66280 -1160 66340 -1100
rect 66280 -1260 66340 -1200
rect 66280 -1360 66340 -1300
rect 66450 -1060 66510 -1000
rect 66450 -1160 66510 -1100
rect 66450 -1260 66510 -1200
rect 66450 -1360 66510 -1300
rect 66620 -1060 66680 -1000
rect 66620 -1160 66680 -1100
rect 66620 -1260 66680 -1200
rect 66620 -1360 66680 -1300
rect 66790 -1060 66850 -1000
rect 66790 -1160 66850 -1100
rect 66790 -1260 66850 -1200
rect 66790 -1360 66850 -1300
rect 66960 -1060 67020 -1000
rect 66960 -1160 67020 -1100
rect 66960 -1260 67020 -1200
rect 66960 -1360 67020 -1300
rect 67130 -1060 67190 -1000
rect 67130 -1160 67190 -1100
rect 67130 -1260 67190 -1200
rect 67130 -1360 67190 -1300
rect 67300 -1060 67360 -1000
rect 67300 -1160 67360 -1100
rect 67300 -1260 67360 -1200
rect 67300 -1360 67360 -1300
rect 67470 -1060 67530 -1000
rect 67470 -1160 67530 -1100
rect 67470 -1260 67530 -1200
rect 67470 -1360 67530 -1300
rect 67640 -1060 67700 -1000
rect 67640 -1160 67700 -1100
rect 67640 -1260 67700 -1200
rect 67640 -1360 67700 -1300
rect 67810 -1060 67870 -1000
rect 67810 -1160 67870 -1100
rect 67810 -1260 67870 -1200
rect 67810 -1360 67870 -1300
rect 67980 -1060 68040 -1000
rect 67980 -1160 68040 -1100
rect 67980 -1260 68040 -1200
rect 67980 -1360 68040 -1300
rect 68150 -1060 68210 -1000
rect 68150 -1160 68210 -1100
rect 68150 -1260 68210 -1200
rect 68150 -1360 68210 -1300
rect 68320 -1060 68380 -1000
rect 68320 -1160 68380 -1100
rect 68320 -1260 68380 -1200
rect 68320 -1360 68380 -1300
rect 68490 -1060 68550 -1000
rect 68490 -1160 68550 -1100
rect 68490 -1260 68550 -1200
rect 68490 -1360 68550 -1300
rect 68660 -1060 68720 -1000
rect 68660 -1160 68720 -1100
rect 68660 -1260 68720 -1200
rect 68660 -1360 68720 -1300
rect 68830 -1060 68890 -1000
rect 68830 -1160 68890 -1100
rect 68830 -1260 68890 -1200
rect 68830 -1360 68890 -1300
rect 69000 -1060 69060 -1000
rect 69000 -1160 69060 -1100
rect 69000 -1260 69060 -1200
rect 69000 -1360 69060 -1300
rect 69170 -1060 69230 -1000
rect 69170 -1160 69230 -1100
rect 69170 -1260 69230 -1200
rect 69170 -1360 69230 -1300
rect 69340 -1060 69400 -1000
rect 69340 -1160 69400 -1100
rect 69340 -1260 69400 -1200
rect 69340 -1360 69400 -1300
rect 69510 -1060 69570 -1000
rect 69510 -1160 69570 -1100
rect 69510 -1260 69570 -1200
rect 69510 -1360 69570 -1300
rect 69680 -1060 69740 -1000
rect 69680 -1160 69740 -1100
rect 69680 -1260 69740 -1200
rect 69680 -1360 69740 -1300
rect 69850 -1060 69910 -1000
rect 69850 -1160 69910 -1100
rect 69850 -1260 69910 -1200
rect 69850 -1360 69910 -1300
rect 70020 -1060 70080 -1000
rect 70020 -1160 70080 -1100
rect 70020 -1260 70080 -1200
rect 70020 -1360 70080 -1300
rect 70190 -1060 70250 -1000
rect 70190 -1160 70250 -1100
rect 70190 -1260 70250 -1200
rect 70190 -1360 70250 -1300
rect 70360 -1060 70420 -1000
rect 70360 -1160 70420 -1100
rect 70360 -1260 70420 -1200
rect 70360 -1360 70420 -1300
rect 70530 -1060 70590 -1000
rect 70530 -1160 70590 -1100
rect 70530 -1260 70590 -1200
rect 70530 -1360 70590 -1300
rect 70700 -1060 70760 -1000
rect 70700 -1160 70760 -1100
rect 70700 -1260 70760 -1200
rect 70700 -1360 70760 -1300
rect 70870 -1060 70930 -1000
rect 70870 -1160 70930 -1100
rect 70870 -1260 70930 -1200
rect 70870 -1360 70930 -1300
rect 71040 -1060 71100 -1000
rect 71040 -1160 71100 -1100
rect 71040 -1260 71100 -1200
rect 71040 -1360 71100 -1300
rect 71210 -1060 71270 -1000
rect 71210 -1160 71270 -1100
rect 71210 -1260 71270 -1200
rect 71210 -1360 71270 -1300
rect 71380 -1060 71440 -1000
rect 71380 -1160 71440 -1100
rect 71380 -1260 71440 -1200
rect 71380 -1360 71440 -1300
rect 71550 -1060 71610 -1000
rect 71550 -1160 71610 -1100
rect 71550 -1260 71610 -1200
rect 71550 -1360 71610 -1300
rect 71720 -1060 71780 -1000
rect 71720 -1160 71780 -1100
rect 71720 -1260 71780 -1200
rect 71720 -1360 71780 -1300
rect 71890 -1060 71950 -1000
rect 71890 -1160 71950 -1100
rect 71890 -1260 71950 -1200
rect 71890 -1360 71950 -1300
rect 72060 -1060 72120 -1000
rect 72060 -1160 72120 -1100
rect 72060 -1260 72120 -1200
rect 72060 -1360 72120 -1300
rect 72230 -1060 72290 -1000
rect 72230 -1160 72290 -1100
rect 72230 -1260 72290 -1200
rect 72230 -1360 72290 -1300
rect 72400 -1060 72460 -1000
rect 72400 -1160 72460 -1100
rect 72400 -1260 72460 -1200
rect 72400 -1360 72460 -1300
rect 72570 -1060 72630 -1000
rect 72570 -1160 72630 -1100
rect 72570 -1260 72630 -1200
rect 72570 -1360 72630 -1300
rect 72740 -1060 72800 -1000
rect 72740 -1160 72800 -1100
rect 72740 -1260 72800 -1200
rect 72740 -1360 72800 -1300
rect 72910 -1060 72970 -1000
rect 72910 -1160 72970 -1100
rect 72910 -1260 72970 -1200
rect 72910 -1360 72970 -1300
rect 73080 -1060 73140 -1000
rect 73080 -1160 73140 -1100
rect 73080 -1260 73140 -1200
rect 73080 -1360 73140 -1300
rect 73250 -1060 73310 -1000
rect 73250 -1160 73310 -1100
rect 73250 -1260 73310 -1200
rect 73250 -1360 73310 -1300
rect 73420 -1060 73480 -1000
rect 73420 -1160 73480 -1100
rect 73420 -1260 73480 -1200
rect 73420 -1360 73480 -1300
rect 73590 -1060 73650 -1000
rect 73590 -1160 73650 -1100
rect 73590 -1260 73650 -1200
rect 73590 -1360 73650 -1300
rect 73760 -1060 73820 -1000
rect 73760 -1160 73820 -1100
rect 73760 -1260 73820 -1200
rect 73760 -1360 73820 -1300
rect 73930 -1060 73990 -1000
rect 73930 -1160 73990 -1100
rect 73930 -1260 73990 -1200
rect 73930 -1360 73990 -1300
rect 74100 -1060 74160 -1000
rect 74100 -1160 74160 -1100
rect 74100 -1260 74160 -1200
rect 74100 -1360 74160 -1300
rect 74270 -1060 74330 -1000
rect 74270 -1160 74330 -1100
rect 74270 -1260 74330 -1200
rect 74270 -1360 74330 -1300
rect 74440 -1060 74500 -1000
rect 74440 -1160 74500 -1100
rect 74440 -1260 74500 -1200
rect 74440 -1360 74500 -1300
rect 74610 -1060 74670 -1000
rect 74610 -1160 74670 -1100
rect 74610 -1260 74670 -1200
rect 74610 -1360 74670 -1300
rect 74780 -1060 74840 -1000
rect 74780 -1160 74840 -1100
rect 74780 -1260 74840 -1200
rect 74780 -1360 74840 -1300
rect 74950 -1060 75010 -1000
rect 74950 -1160 75010 -1100
rect 74950 -1260 75010 -1200
rect 74950 -1360 75010 -1300
rect 75120 -1060 75180 -1000
rect 75120 -1160 75180 -1100
rect 75120 -1260 75180 -1200
rect 75120 -1360 75180 -1300
rect 75290 -1060 75350 -1000
rect 75290 -1160 75350 -1100
rect 75290 -1260 75350 -1200
rect 75290 -1360 75350 -1300
rect 75460 -1060 75520 -1000
rect 75460 -1160 75520 -1100
rect 75460 -1260 75520 -1200
rect 75460 -1360 75520 -1300
rect 75630 -1060 75690 -1000
rect 75630 -1160 75690 -1100
rect 75630 -1260 75690 -1200
rect 75630 -1360 75690 -1300
rect 75800 -1060 75860 -1000
rect 75800 -1160 75860 -1100
rect 75800 -1260 75860 -1200
rect 75800 -1360 75860 -1300
rect 75970 -1060 76030 -1000
rect 75970 -1160 76030 -1100
rect 75970 -1260 76030 -1200
rect 75970 -1360 76030 -1300
rect 76140 -1060 76200 -1000
rect 76140 -1160 76200 -1100
rect 76140 -1260 76200 -1200
rect 76140 -1360 76200 -1300
rect 76310 -1060 76370 -1000
rect 76310 -1160 76370 -1100
rect 76310 -1260 76370 -1200
rect 76310 -1360 76370 -1300
rect 76480 -1060 76540 -1000
rect 76480 -1160 76540 -1100
rect 76480 -1260 76540 -1200
rect 76480 -1360 76540 -1300
rect 76650 -1060 76710 -1000
rect 76650 -1160 76710 -1100
rect 76650 -1260 76710 -1200
rect 76650 -1360 76710 -1300
rect 76820 -1060 76880 -1000
rect 76820 -1160 76880 -1100
rect 76820 -1260 76880 -1200
rect 76820 -1360 76880 -1300
rect 76990 -1060 77050 -1000
rect 76990 -1160 77050 -1100
rect 76990 -1260 77050 -1200
rect 76990 -1360 77050 -1300
rect 77160 -1060 77220 -1000
rect 77160 -1160 77220 -1100
rect 77160 -1260 77220 -1200
rect 77160 -1360 77220 -1300
rect 77330 -1060 77390 -1000
rect 77330 -1160 77390 -1100
rect 77330 -1260 77390 -1200
rect 77330 -1360 77390 -1300
rect 77500 -1060 77560 -1000
rect 77500 -1160 77560 -1100
rect 77500 -1260 77560 -1200
rect 77500 -1360 77560 -1300
rect 77670 -1060 77730 -1000
rect 77670 -1160 77730 -1100
rect 77670 -1260 77730 -1200
rect 77670 -1360 77730 -1300
rect 77840 -1060 77900 -1000
rect 77840 -1160 77900 -1100
rect 77840 -1260 77900 -1200
rect 77840 -1360 77900 -1300
rect 78010 -1060 78070 -1000
rect 78010 -1160 78070 -1100
rect 78010 -1260 78070 -1200
rect 78010 -1360 78070 -1300
rect 78180 -1060 78240 -1000
rect 78180 -1160 78240 -1100
rect 78180 -1260 78240 -1200
rect 78180 -1360 78240 -1300
rect 78350 -1060 78410 -1000
rect 78350 -1160 78410 -1100
rect 78350 -1260 78410 -1200
rect 78350 -1360 78410 -1300
rect 78520 -1060 78580 -1000
rect 78520 -1160 78580 -1100
rect 78520 -1260 78580 -1200
rect 78520 -1360 78580 -1300
rect 78690 -1060 78750 -1000
rect 78690 -1160 78750 -1100
rect 78690 -1260 78750 -1200
rect 78690 -1360 78750 -1300
rect 78860 -1060 78920 -1000
rect 78860 -1160 78920 -1100
rect 78860 -1260 78920 -1200
rect 78860 -1360 78920 -1300
rect 79030 -1060 79090 -1000
rect 79030 -1160 79090 -1100
rect 79030 -1260 79090 -1200
rect 79030 -1360 79090 -1300
rect 79200 -1060 79260 -1000
rect 79200 -1160 79260 -1100
rect 79200 -1260 79260 -1200
rect 79200 -1360 79260 -1300
rect 79370 -1060 79430 -1000
rect 79370 -1160 79430 -1100
rect 79370 -1260 79430 -1200
rect 79370 -1360 79430 -1300
rect 79540 -1060 79600 -1000
rect 79540 -1160 79600 -1100
rect 79540 -1260 79600 -1200
rect 79540 -1360 79600 -1300
rect 79710 -1060 79770 -1000
rect 79710 -1160 79770 -1100
rect 79710 -1260 79770 -1200
rect 79710 -1360 79770 -1300
rect 79880 -1060 79940 -1000
rect 79880 -1160 79940 -1100
rect 79880 -1260 79940 -1200
rect 79880 -1360 79940 -1300
rect 80050 -1060 80110 -1000
rect 80050 -1160 80110 -1100
rect 80050 -1260 80110 -1200
rect 80050 -1360 80110 -1300
rect 80220 -1060 80280 -1000
rect 80220 -1160 80280 -1100
rect 80220 -1260 80280 -1200
rect 80220 -1360 80280 -1300
rect 80390 -1060 80450 -1000
rect 80390 -1160 80450 -1100
rect 80390 -1260 80450 -1200
rect 80390 -1360 80450 -1300
rect 80560 -1060 80620 -1000
rect 80560 -1160 80620 -1100
rect 80560 -1260 80620 -1200
rect 80560 -1360 80620 -1300
rect 80730 -1060 80790 -1000
rect 80730 -1160 80790 -1100
rect 80730 -1260 80790 -1200
rect 80730 -1360 80790 -1300
rect 80900 -1060 80960 -1000
rect 80900 -1160 80960 -1100
rect 80900 -1260 80960 -1200
rect 80900 -1360 80960 -1300
rect 81070 -1060 81130 -1000
rect 81070 -1160 81130 -1100
rect 81070 -1260 81130 -1200
rect 81070 -1360 81130 -1300
rect 81240 -1060 81300 -1000
rect 81240 -1160 81300 -1100
rect 81240 -1260 81300 -1200
rect 81240 -1360 81300 -1300
rect 81410 -1060 81470 -1000
rect 81410 -1160 81470 -1100
rect 81410 -1260 81470 -1200
rect 81410 -1360 81470 -1300
rect 81580 -1060 81640 -1000
rect 81580 -1160 81640 -1100
rect 81580 -1260 81640 -1200
rect 81580 -1360 81640 -1300
rect 81750 -1060 81810 -1000
rect 81750 -1160 81810 -1100
rect 81750 -1260 81810 -1200
rect 81750 -1360 81810 -1300
rect 81920 -1060 81980 -1000
rect 81920 -1160 81980 -1100
rect 81920 -1260 81980 -1200
rect 81920 -1360 81980 -1300
rect 82090 -1060 82150 -1000
rect 82090 -1160 82150 -1100
rect 82090 -1260 82150 -1200
rect 82090 -1360 82150 -1300
rect 82260 -1060 82320 -1000
rect 82260 -1160 82320 -1100
rect 82260 -1260 82320 -1200
rect 82260 -1360 82320 -1300
rect 82430 -1060 82490 -1000
rect 82430 -1160 82490 -1100
rect 82430 -1260 82490 -1200
rect 82430 -1360 82490 -1300
rect 82600 -1060 82660 -1000
rect 82600 -1160 82660 -1100
rect 82600 -1260 82660 -1200
rect 82600 -1360 82660 -1300
rect 82770 -1060 82830 -1000
rect 82770 -1160 82830 -1100
rect 82770 -1260 82830 -1200
rect 82770 -1360 82830 -1300
rect 82940 -1060 83000 -1000
rect 82940 -1160 83000 -1100
rect 82940 -1260 83000 -1200
rect 82940 -1360 83000 -1300
rect 83110 -1060 83170 -1000
rect 83110 -1160 83170 -1100
rect 83110 -1260 83170 -1200
rect 83110 -1360 83170 -1300
rect 83280 -1060 83340 -1000
rect 83280 -1160 83340 -1100
rect 83280 -1260 83340 -1200
rect 83280 -1360 83340 -1300
rect 83450 -1060 83510 -1000
rect 83450 -1160 83510 -1100
rect 83450 -1260 83510 -1200
rect 83450 -1360 83510 -1300
rect 83620 -1060 83680 -1000
rect 83620 -1160 83680 -1100
rect 83620 -1260 83680 -1200
rect 83620 -1360 83680 -1300
rect 83790 -1060 83850 -1000
rect 83790 -1160 83850 -1100
rect 83790 -1260 83850 -1200
rect 83790 -1360 83850 -1300
rect 83960 -1060 84020 -1000
rect 83960 -1160 84020 -1100
rect 83960 -1260 84020 -1200
rect 83960 -1360 84020 -1300
rect 84130 -1060 84190 -1000
rect 84130 -1160 84190 -1100
rect 84130 -1260 84190 -1200
rect 84130 -1360 84190 -1300
rect 84300 -1060 84360 -1000
rect 84300 -1160 84360 -1100
rect 84300 -1260 84360 -1200
rect 84300 -1360 84360 -1300
rect 84470 -1060 84530 -1000
rect 84470 -1160 84530 -1100
rect 84470 -1260 84530 -1200
rect 84470 -1360 84530 -1300
rect 84640 -1060 84700 -1000
rect 84640 -1160 84700 -1100
rect 84640 -1260 84700 -1200
rect 84640 -1360 84700 -1300
rect 84810 -1060 84870 -1000
rect 84810 -1160 84870 -1100
rect 84810 -1260 84870 -1200
rect 84810 -1360 84870 -1300
rect 84980 -1060 85040 -1000
rect 84980 -1160 85040 -1100
rect 84980 -1260 85040 -1200
rect 84980 -1360 85040 -1300
rect 85150 -1060 85210 -1000
rect 85150 -1160 85210 -1100
rect 85150 -1260 85210 -1200
rect 85150 -1360 85210 -1300
rect 85320 -1060 85380 -1000
rect 85320 -1160 85380 -1100
rect 85320 -1260 85380 -1200
rect 85320 -1360 85380 -1300
rect 85490 -1060 85550 -1000
rect 85490 -1160 85550 -1100
rect 85490 -1260 85550 -1200
rect 85490 -1360 85550 -1300
rect 85660 -1060 85720 -1000
rect 85660 -1160 85720 -1100
rect 85660 -1260 85720 -1200
rect 85660 -1360 85720 -1300
rect 85830 -1060 85890 -1000
rect 85830 -1160 85890 -1100
rect 85830 -1260 85890 -1200
rect 85830 -1360 85890 -1300
rect 86000 -1060 86060 -1000
rect 86000 -1160 86060 -1100
rect 86000 -1260 86060 -1200
rect 86000 -1360 86060 -1300
rect 86170 -1060 86230 -1000
rect 86170 -1160 86230 -1100
rect 86170 -1260 86230 -1200
rect 86170 -1360 86230 -1300
rect 86340 -1060 86400 -1000
rect 86340 -1160 86400 -1100
rect 86340 -1260 86400 -1200
rect 86340 -1360 86400 -1300
rect 86510 -1060 86570 -1000
rect 86510 -1160 86570 -1100
rect 86510 -1260 86570 -1200
rect 86510 -1360 86570 -1300
rect 86680 -1060 86740 -1000
rect 86680 -1160 86740 -1100
rect 86680 -1260 86740 -1200
rect 86680 -1360 86740 -1300
rect 86850 -1060 86910 -1000
rect 86850 -1160 86910 -1100
rect 86850 -1260 86910 -1200
rect 86850 -1360 86910 -1300
rect 87020 -1060 87080 -1000
rect 87020 -1160 87080 -1100
rect 87020 -1260 87080 -1200
rect 87020 -1360 87080 -1300
rect 87190 -1060 87250 -1000
rect 87190 -1160 87250 -1100
rect 87190 -1260 87250 -1200
rect 87190 -1360 87250 -1300
<< psubdiff >>
rect 409 1095 505 1129
rect 1383 1095 1479 1129
rect 409 1033 443 1095
rect 1445 1033 1479 1095
rect 409 835 443 897
rect 1445 835 1479 897
rect 409 801 505 835
rect 1383 801 1479 835
rect 5529 1073 5625 1107
rect 6503 1073 6599 1107
rect 5529 1011 5563 1073
rect 6565 1011 6599 1073
rect 5529 813 5563 875
rect 6565 813 6599 875
rect 5529 779 5625 813
rect 6503 779 6599 813
rect 2070 -260 2400 -240
rect 2070 -390 2120 -260
rect 2350 -390 2400 -260
rect 2070 -410 2400 -390
rect 5088 -268 5418 -248
rect 5088 -398 5138 -268
rect 5368 -398 5418 -268
rect 5088 -418 5418 -398
rect 7574 -268 7904 -248
rect 7574 -398 7624 -268
rect 7854 -398 7904 -268
rect 7574 -418 7904 -398
rect 8994 -268 9324 -248
rect 8994 -398 9044 -268
rect 9274 -398 9324 -268
rect 8994 -418 9324 -398
rect 13618 -264 13948 -244
rect 13618 -394 13668 -264
rect 13898 -394 13948 -264
rect 13618 -414 13948 -394
rect 16818 -264 17148 -244
rect 16818 -394 16868 -264
rect 17098 -394 17148 -264
rect 16818 -414 17148 -394
rect 20374 -264 20704 -244
rect 20374 -394 20424 -264
rect 20654 -394 20704 -264
rect 20374 -414 20704 -394
rect 25708 -264 26038 -244
rect 25708 -394 25758 -264
rect 25988 -394 26038 -264
rect 25708 -414 26038 -394
rect 28552 -264 28882 -244
rect 28552 -394 28602 -264
rect 28832 -394 28882 -264
rect 28552 -414 28882 -394
rect 32464 -264 32794 -244
rect 32464 -394 32514 -264
rect 32744 -394 32794 -264
rect 32464 -414 32794 -394
rect 34620 -264 34950 -244
rect 34620 -394 34670 -264
rect 34900 -394 34950 -264
rect 34620 -414 34950 -394
rect 37442 -264 37772 -244
rect 37442 -394 37492 -264
rect 37722 -394 37772 -264
rect 37442 -414 37772 -394
rect 40642 -264 40972 -244
rect 40642 -394 40692 -264
rect 40922 -394 40972 -264
rect 40642 -414 40972 -394
rect 45618 -264 45948 -244
rect 45618 -394 45668 -264
rect 45898 -394 45948 -264
rect 45618 -414 45948 -394
rect 48818 -264 49148 -244
rect 48818 -394 48868 -264
rect 49098 -394 49148 -264
rect 48818 -414 49148 -394
rect 50952 -264 51282 -244
rect 50952 -394 51002 -264
rect 51232 -394 51282 -264
rect 50952 -414 51282 -394
rect 54508 -264 54838 -244
rect 54508 -394 54558 -264
rect 54788 -394 54838 -264
rect 54508 -414 54838 -394
rect 57352 -264 57682 -244
rect 57352 -394 57402 -264
rect 57632 -394 57682 -264
rect 57352 -414 57682 -394
rect 61264 -264 61594 -244
rect 61264 -394 61314 -264
rect 61544 -394 61594 -264
rect 61264 -414 61594 -394
rect 64108 -264 64438 -244
rect 64108 -394 64158 -264
rect 64388 -394 64438 -264
rect 64108 -414 64438 -394
rect 67664 -264 67994 -244
rect 67664 -394 67714 -264
rect 67944 -394 67994 -264
rect 67664 -414 67994 -394
rect 70508 -264 70838 -244
rect 70508 -394 70558 -264
rect 70788 -394 70838 -264
rect 70508 -414 70838 -394
rect 74418 -264 74748 -244
rect 74418 -394 74468 -264
rect 74698 -394 74748 -264
rect 74418 -414 74748 -394
rect 78330 -264 78660 -244
rect 78330 -394 78380 -264
rect 78610 -394 78660 -264
rect 78330 -414 78660 -394
rect 82242 -264 82572 -244
rect 82242 -394 82292 -264
rect 82522 -394 82572 -264
rect 82242 -414 82572 -394
rect 86152 -264 86482 -244
rect 86152 -394 86202 -264
rect 86432 -394 86482 -264
rect 86152 -414 86482 -394
<< nsubdiff >>
rect 730 590 930 620
rect 730 520 790 590
rect 870 520 930 590
rect 730 490 930 520
rect 2110 590 2310 620
rect 2110 520 2170 590
rect 2250 520 2310 590
rect 2110 490 2310 520
rect 3490 590 3690 620
rect 3490 520 3550 590
rect 3630 520 3690 590
rect 3490 490 3690 520
rect 5150 590 5350 620
rect 5150 520 5210 590
rect 5290 520 5350 590
rect 5150 490 5350 520
rect 7980 590 8180 620
rect 7980 520 8040 590
rect 8120 520 8180 590
rect 7980 490 8180 520
rect 10740 590 10940 620
rect 10740 520 10800 590
rect 10880 520 10940 590
rect 10740 490 10940 520
rect 13370 590 13570 620
rect 13370 520 13430 590
rect 13510 520 13570 590
rect 13370 490 13570 520
rect 16410 590 16610 620
rect 16410 520 16470 590
rect 16550 520 16610 590
rect 16410 490 16610 520
rect 20480 590 20680 620
rect 20480 520 20540 590
rect 20620 520 20680 590
rect 20480 490 20680 520
rect 24620 590 24820 620
rect 24620 520 24680 590
rect 24760 520 24820 590
rect 24620 490 24820 520
rect 28700 590 28900 620
rect 28700 520 28760 590
rect 28840 520 28900 590
rect 28700 490 28900 520
rect 32850 590 33050 620
rect 32850 520 32910 590
rect 32990 520 33050 590
rect 32850 490 33050 520
rect 36720 590 36920 620
rect 36720 520 36780 590
rect 36860 520 36920 590
rect 36720 490 36920 520
rect 40860 590 41060 620
rect 40860 520 40920 590
rect 41000 520 41060 590
rect 40860 490 41060 520
rect 44850 590 45050 620
rect 44850 520 44910 590
rect 44990 520 45050 590
rect 44850 490 45050 520
rect 48930 590 49130 620
rect 48930 520 48990 590
rect 49070 520 49130 590
rect 48930 490 49130 520
rect 53020 590 53220 620
rect 53020 520 53080 590
rect 53160 520 53220 590
rect 53020 490 53220 520
rect 57180 590 57380 620
rect 57180 520 57240 590
rect 57320 520 57380 590
rect 57180 490 57380 520
rect 770 -1470 970 -1440
rect 770 -1540 830 -1470
rect 910 -1540 970 -1470
rect 770 -1570 970 -1540
rect 4940 -1470 5140 -1440
rect 4940 -1540 5000 -1470
rect 5080 -1540 5140 -1470
rect 4940 -1570 5140 -1540
rect 8970 -1470 9170 -1440
rect 8970 -1540 9030 -1470
rect 9110 -1540 9170 -1470
rect 8970 -1570 9170 -1540
rect 13000 -1470 13200 -1440
rect 13000 -1540 13060 -1470
rect 13140 -1540 13200 -1470
rect 13000 -1570 13200 -1540
rect 17040 -1470 17240 -1440
rect 17040 -1540 17100 -1470
rect 17180 -1540 17240 -1470
rect 17040 -1570 17240 -1540
rect 21140 -1470 21340 -1440
rect 21140 -1540 21200 -1470
rect 21280 -1540 21340 -1470
rect 21140 -1570 21340 -1540
rect 25250 -1470 25450 -1440
rect 25250 -1540 25310 -1470
rect 25390 -1540 25450 -1470
rect 25250 -1570 25450 -1540
rect 29350 -1470 29550 -1440
rect 29350 -1540 29410 -1470
rect 29490 -1540 29550 -1470
rect 29350 -1570 29550 -1540
rect 33380 -1470 33580 -1440
rect 33380 -1540 33440 -1470
rect 33520 -1540 33580 -1470
rect 33380 -1570 33580 -1540
rect 37490 -1470 37690 -1440
rect 37490 -1540 37550 -1470
rect 37630 -1540 37690 -1470
rect 37490 -1570 37690 -1540
rect 41590 -1470 41790 -1440
rect 41590 -1540 41650 -1470
rect 41730 -1540 41790 -1470
rect 41590 -1570 41790 -1540
rect 47040 -1470 47240 -1440
rect 47040 -1540 47100 -1470
rect 47180 -1540 47240 -1470
rect 47040 -1570 47240 -1540
rect 51120 -1470 51320 -1440
rect 51120 -1540 51180 -1470
rect 51260 -1540 51320 -1470
rect 51120 -1570 51320 -1540
rect 55230 -1470 55430 -1440
rect 55230 -1540 55290 -1470
rect 55370 -1540 55430 -1470
rect 55230 -1570 55430 -1540
rect 59260 -1470 59460 -1440
rect 59260 -1540 59320 -1470
rect 59400 -1540 59460 -1470
rect 59260 -1570 59460 -1540
rect 63360 -1470 63560 -1440
rect 63360 -1540 63420 -1470
rect 63500 -1540 63560 -1470
rect 63360 -1570 63560 -1540
rect 67470 -1470 67670 -1440
rect 67470 -1540 67530 -1470
rect 67610 -1540 67670 -1470
rect 67470 -1570 67670 -1540
rect 71500 -1470 71700 -1440
rect 71500 -1540 71560 -1470
rect 71640 -1540 71700 -1470
rect 71500 -1570 71700 -1540
rect 75750 -1470 75950 -1440
rect 75750 -1540 75810 -1470
rect 75890 -1540 75950 -1470
rect 75750 -1570 75950 -1540
rect 79710 -1470 79910 -1440
rect 79710 -1540 79770 -1470
rect 79850 -1540 79910 -1470
rect 79710 -1570 79910 -1540
rect 83890 -1470 84090 -1440
rect 83890 -1540 83950 -1470
rect 84030 -1540 84090 -1470
rect 83890 -1570 84090 -1540
rect 86450 -1474 86648 -1444
rect 86450 -1544 86508 -1474
rect 86588 -1544 86648 -1474
rect 86450 -1572 86648 -1544
<< psubdiffcont >>
rect 505 1095 1383 1129
rect 409 897 443 1033
rect 1445 897 1479 1033
rect 505 801 1383 835
rect 5625 1073 6503 1107
rect 5529 875 5563 1011
rect 6565 875 6599 1011
rect 5625 779 6503 813
rect 2120 -390 2350 -260
rect 5138 -398 5368 -268
rect 7624 -398 7854 -268
rect 9044 -398 9274 -268
rect 13668 -394 13898 -264
rect 16868 -394 17098 -264
rect 20424 -394 20654 -264
rect 25758 -394 25988 -264
rect 28602 -394 28832 -264
rect 32514 -394 32744 -264
rect 34670 -394 34900 -264
rect 37492 -394 37722 -264
rect 40692 -394 40922 -264
rect 45668 -394 45898 -264
rect 48868 -394 49098 -264
rect 51002 -394 51232 -264
rect 54558 -394 54788 -264
rect 57402 -394 57632 -264
rect 61314 -394 61544 -264
rect 64158 -394 64388 -264
rect 67714 -394 67944 -264
rect 70558 -394 70788 -264
rect 74468 -394 74698 -264
rect 78380 -394 78610 -264
rect 82292 -394 82522 -264
rect 86202 -394 86432 -264
<< nsubdiffcont >>
rect 790 520 870 590
rect 2170 520 2250 590
rect 3550 520 3630 590
rect 5210 520 5290 590
rect 8040 520 8120 590
rect 10800 520 10880 590
rect 13430 520 13510 590
rect 16470 520 16550 590
rect 20540 520 20620 590
rect 24680 520 24760 590
rect 28760 520 28840 590
rect 32910 520 32990 590
rect 36780 520 36860 590
rect 40920 520 41000 590
rect 44910 520 44990 590
rect 48990 520 49070 590
rect 53080 520 53160 590
rect 57240 520 57320 590
rect 830 -1540 910 -1470
rect 5000 -1540 5080 -1470
rect 9030 -1540 9110 -1470
rect 13060 -1540 13140 -1470
rect 17100 -1540 17180 -1470
rect 21200 -1540 21280 -1470
rect 25310 -1540 25390 -1470
rect 29410 -1540 29490 -1470
rect 33440 -1540 33520 -1470
rect 37550 -1540 37630 -1470
rect 41650 -1540 41730 -1470
rect 47100 -1540 47180 -1470
rect 51180 -1540 51260 -1470
rect 55290 -1540 55370 -1470
rect 59320 -1540 59400 -1470
rect 63420 -1540 63500 -1470
rect 67530 -1540 67610 -1470
rect 71560 -1540 71640 -1470
rect 75810 -1540 75890 -1470
rect 79770 -1540 79850 -1470
rect 83950 -1540 84030 -1470
rect 86508 -1544 86588 -1474
<< poly >>
rect 500 690 630 710
rect 500 630 520 690
rect 610 630 630 690
rect 500 610 630 630
rect 5610 690 5740 710
rect 5610 630 5630 690
rect 5720 630 5740 690
rect 130 430 160 460
rect 550 430 580 610
rect 5610 610 5740 630
rect 720 430 750 460
rect 890 430 920 460
rect 1060 430 1090 460
rect 1620 430 1650 460
rect 1790 430 1820 460
rect 1960 430 1990 460
rect 2130 430 2160 460
rect 2300 430 2330 460
rect 2470 430 2500 460
rect 2640 430 2670 460
rect 2810 430 2840 460
rect 2980 430 3010 460
rect 3150 430 3180 460
rect 3320 430 3350 460
rect 3490 430 3520 460
rect 3660 430 3690 460
rect 3830 430 3860 460
rect 4000 430 4030 460
rect 4170 430 4200 460
rect 4640 430 4670 460
rect 4810 430 4840 460
rect 4980 430 5010 460
rect 5150 430 5180 460
rect 5320 430 5350 460
rect 5490 430 5520 460
rect 5660 430 5690 610
rect 5830 430 5860 460
rect 6000 430 6030 460
rect 6170 430 6200 460
rect 6340 430 6370 460
rect 6510 430 6540 460
rect 6680 430 6710 460
rect 6850 430 6880 460
rect 7020 430 7050 460
rect 7190 430 7220 460
rect 7360 430 7390 460
rect 7530 430 7560 460
rect 7700 430 7730 460
rect 7870 430 7900 460
rect 8040 430 8070 460
rect 8210 430 8240 460
rect 8380 430 8410 460
rect 8550 430 8580 460
rect 8720 430 8750 460
rect 8890 430 8920 460
rect 9060 430 9090 460
rect 9230 430 9260 460
rect 9400 430 9430 460
rect 9570 430 9600 460
rect 9740 430 9770 460
rect 9910 430 9940 460
rect 10080 430 10110 460
rect 10250 430 10280 460
rect 10420 430 10450 460
rect 10590 430 10620 460
rect 10760 430 10790 460
rect 10930 430 10960 460
rect 11100 430 11130 460
rect 11270 430 11300 460
rect 11440 430 11470 460
rect 11610 430 11640 460
rect 11780 430 11810 460
rect 11950 430 11980 460
rect 12120 430 12150 460
rect 12290 430 12320 460
rect 12460 430 12490 460
rect 12630 430 12660 460
rect 12800 430 12830 460
rect 12970 430 13000 460
rect 13140 430 13170 460
rect 13310 430 13340 460
rect 13480 430 13510 460
rect 13650 430 13680 460
rect 13820 430 13850 460
rect 13990 430 14020 460
rect 14160 430 14190 460
rect 14330 430 14360 460
rect 14500 430 14530 460
rect 14670 430 14700 460
rect 14840 430 14870 460
rect 15010 430 15040 460
rect 15180 430 15210 460
rect 15350 430 15380 460
rect 15820 430 15850 460
rect 15990 430 16020 460
rect 16160 430 16190 460
rect 16330 430 16360 460
rect 16500 430 16530 460
rect 16670 430 16700 460
rect 16840 430 16870 460
rect 17010 430 17040 460
rect 17180 430 17210 460
rect 17350 430 17380 460
rect 17520 430 17550 460
rect 17690 430 17720 460
rect 17860 430 17890 460
rect 18030 430 18060 460
rect 18200 430 18230 460
rect 18370 430 18400 460
rect 18540 430 18570 460
rect 18710 430 18740 460
rect 18880 430 18910 460
rect 19050 430 19080 460
rect 19220 430 19250 460
rect 19390 430 19420 460
rect 19560 430 19590 460
rect 19730 430 19760 460
rect 19900 430 19930 460
rect 20070 430 20100 460
rect 20240 430 20270 460
rect 20410 430 20440 460
rect 20580 430 20610 460
rect 20750 430 20780 460
rect 20920 430 20950 460
rect 21090 430 21120 460
rect 21260 430 21290 460
rect 21430 430 21460 460
rect 21600 430 21630 460
rect 21770 430 21800 460
rect 21940 430 21970 460
rect 22110 430 22140 460
rect 22280 430 22310 460
rect 22450 430 22480 460
rect 22620 430 22650 460
rect 22790 430 22820 460
rect 22960 430 22990 460
rect 23130 430 23160 460
rect 23300 430 23330 460
rect 23470 430 23500 460
rect 23640 430 23670 460
rect 23810 430 23840 460
rect 23980 430 24010 460
rect 24150 430 24180 460
rect 24320 430 24350 460
rect 24490 430 24520 460
rect 24660 430 24690 460
rect 24830 430 24860 460
rect 25000 430 25030 460
rect 25170 430 25200 460
rect 25340 430 25370 460
rect 25510 430 25540 460
rect 25680 430 25710 460
rect 25850 430 25880 460
rect 26020 430 26050 460
rect 26190 430 26220 460
rect 26360 430 26390 460
rect 26530 430 26560 460
rect 26700 430 26730 460
rect 26870 430 26900 460
rect 27040 430 27070 460
rect 27210 430 27240 460
rect 27380 430 27410 460
rect 27550 430 27580 460
rect 27720 430 27750 460
rect 27890 430 27920 460
rect 28060 430 28090 460
rect 28230 430 28260 460
rect 28400 430 28430 460
rect 28570 430 28600 460
rect 28740 430 28770 460
rect 28910 430 28940 460
rect 29080 430 29110 460
rect 29250 430 29280 460
rect 29420 430 29450 460
rect 29590 430 29620 460
rect 29760 430 29790 460
rect 29930 430 29960 460
rect 30100 430 30130 460
rect 30270 430 30300 460
rect 30440 430 30470 460
rect 30610 430 30640 460
rect 30780 430 30810 460
rect 30950 430 30980 460
rect 31120 430 31150 460
rect 31290 430 31320 460
rect 31460 430 31490 460
rect 31630 430 31660 460
rect 31800 430 31830 460
rect 31970 430 32000 460
rect 32140 430 32170 460
rect 32310 430 32340 460
rect 32480 430 32510 460
rect 32650 430 32680 460
rect 32820 430 32850 460
rect 32990 430 33020 460
rect 33160 430 33190 460
rect 33330 430 33360 460
rect 33500 430 33530 460
rect 33670 430 33700 460
rect 33840 430 33870 460
rect 34010 430 34040 460
rect 34180 430 34210 460
rect 34350 430 34380 460
rect 34520 430 34550 460
rect 34690 430 34720 460
rect 34860 430 34890 460
rect 35030 430 35060 460
rect 35200 430 35230 460
rect 35370 430 35400 460
rect 35540 430 35570 460
rect 35710 430 35740 460
rect 35880 430 35910 460
rect 36050 430 36080 460
rect 36220 430 36250 460
rect 36390 430 36420 460
rect 36560 430 36590 460
rect 36730 430 36760 460
rect 36900 430 36930 460
rect 37070 430 37100 460
rect 37240 430 37270 460
rect 37410 430 37440 460
rect 37580 430 37610 460
rect 37750 430 37780 460
rect 37920 430 37950 460
rect 38090 430 38120 460
rect 38260 430 38290 460
rect 38430 430 38460 460
rect 38600 430 38630 460
rect 38770 430 38800 460
rect 38940 430 38970 460
rect 39110 430 39140 460
rect 39280 430 39310 460
rect 39450 430 39480 460
rect 39620 430 39650 460
rect 39790 430 39820 460
rect 39960 430 39990 460
rect 40130 430 40160 460
rect 40300 430 40330 460
rect 40470 430 40500 460
rect 40640 430 40670 460
rect 40810 430 40840 460
rect 40980 430 41010 460
rect 41150 430 41180 460
rect 41320 430 41350 460
rect 41490 430 41520 460
rect 41660 430 41690 460
rect 41830 430 41860 460
rect 42000 430 42030 460
rect 42170 430 42200 460
rect 42340 430 42370 460
rect 42510 430 42540 460
rect 42680 430 42710 460
rect 42850 430 42880 460
rect 43020 430 43050 460
rect 43190 430 43220 460
rect 43360 430 43390 460
rect 43530 430 43560 460
rect 43700 430 43730 460
rect 43870 430 43900 460
rect 44040 430 44070 460
rect 44210 430 44240 460
rect 44380 430 44410 460
rect 44550 430 44580 460
rect 44720 430 44750 460
rect 44890 430 44920 460
rect 45060 430 45090 460
rect 45230 430 45260 460
rect 45400 430 45430 460
rect 45570 430 45600 460
rect 45740 430 45770 460
rect 45910 430 45940 460
rect 46080 430 46110 460
rect 46250 430 46280 460
rect 46420 430 46450 460
rect 46590 430 46620 460
rect 46760 430 46790 460
rect 46930 430 46960 460
rect 47100 430 47130 460
rect 47270 430 47300 460
rect 47440 430 47470 460
rect 47610 430 47640 460
rect 47780 430 47810 460
rect 47950 430 47980 460
rect 48120 430 48150 460
rect 48290 430 48320 460
rect 48460 430 48490 460
rect 48630 430 48660 460
rect 48800 430 48830 460
rect 48970 430 49000 460
rect 49140 430 49170 460
rect 49310 430 49340 460
rect 49480 430 49510 460
rect 49650 430 49680 460
rect 49820 430 49850 460
rect 49990 430 50020 460
rect 50160 430 50190 460
rect 50330 430 50360 460
rect 50500 430 50530 460
rect 50670 430 50700 460
rect 50840 430 50870 460
rect 51010 430 51040 460
rect 51180 430 51210 460
rect 51350 430 51380 460
rect 51520 430 51550 460
rect 51690 430 51720 460
rect 51860 430 51890 460
rect 52030 430 52060 460
rect 52200 430 52230 460
rect 52370 430 52400 460
rect 52540 430 52570 460
rect 52710 430 52740 460
rect 52880 430 52910 460
rect 53050 430 53080 460
rect 53220 430 53250 460
rect 53390 430 53420 460
rect 53560 430 53590 460
rect 53730 430 53760 460
rect 53900 430 53930 460
rect 54070 430 54100 460
rect 54240 430 54270 460
rect 54410 430 54440 460
rect 54580 430 54610 460
rect 54750 430 54780 460
rect 54920 430 54950 460
rect 55090 430 55120 460
rect 55260 430 55290 460
rect 55430 430 55460 460
rect 55600 430 55630 460
rect 55770 430 55800 460
rect 55940 430 55970 460
rect 56110 430 56140 460
rect 56280 430 56310 460
rect 56450 430 56480 460
rect 56620 430 56650 460
rect 56790 430 56820 460
rect 56960 430 56990 460
rect 57130 430 57160 460
rect 57300 430 57330 460
rect 57470 430 57500 460
rect 57640 430 57670 460
rect 57810 430 57840 460
rect 57980 430 58010 460
rect 58150 430 58180 460
rect 58320 430 58350 460
rect 58490 430 58520 460
rect 58660 430 58690 460
rect 58830 430 58860 460
rect 59000 430 59030 460
rect 59170 430 59200 460
rect 130 130 160 230
rect 50 110 160 130
rect 50 30 70 110
rect 130 30 160 110
rect 550 100 580 230
rect 720 100 750 230
rect 890 100 920 230
rect 1060 100 1090 230
rect 1620 100 1650 230
rect 1790 100 1820 230
rect 1960 100 1990 230
rect 2130 100 2160 230
rect 2300 100 2330 230
rect 2470 100 2500 230
rect 2640 100 2670 230
rect 2810 100 2840 230
rect 2980 100 3010 230
rect 3150 100 3180 230
rect 3320 100 3350 230
rect 3490 100 3520 230
rect 3660 100 3690 230
rect 3830 100 3860 230
rect 4000 100 4030 230
rect 4170 100 4200 230
rect 4640 100 4670 230
rect 4810 100 4840 230
rect 4980 100 5010 230
rect 5150 100 5180 230
rect 5320 100 5350 230
rect 5490 100 5520 230
rect 5660 100 5690 230
rect 5830 100 5860 230
rect 6000 100 6030 230
rect 6170 100 6200 230
rect 6340 100 6370 230
rect 6510 100 6540 230
rect 6680 100 6710 230
rect 6850 100 6880 230
rect 7020 100 7050 230
rect 7190 100 7220 230
rect 7360 100 7390 230
rect 7530 100 7560 230
rect 7700 100 7730 230
rect 7870 100 7900 230
rect 8040 100 8070 230
rect 8210 100 8240 230
rect 8380 100 8410 230
rect 8550 100 8580 230
rect 8720 100 8750 230
rect 8890 100 8920 230
rect 9060 100 9090 230
rect 9230 100 9260 230
rect 9400 100 9430 230
rect 9570 100 9600 230
rect 9740 100 9770 230
rect 9910 100 9940 230
rect 10080 100 10110 230
rect 10250 100 10280 230
rect 10420 100 10450 230
rect 10590 100 10620 230
rect 10760 100 10790 230
rect 10930 100 10960 230
rect 11100 100 11130 230
rect 11270 100 11300 230
rect 11440 100 11470 230
rect 11610 100 11640 230
rect 11780 100 11810 230
rect 11950 100 11980 230
rect 12120 100 12150 230
rect 12290 100 12320 230
rect 12460 100 12490 230
rect 12630 100 12660 230
rect 12800 100 12830 230
rect 12970 100 13000 230
rect 13140 100 13170 230
rect 13310 100 13340 230
rect 13480 100 13510 230
rect 13650 100 13680 230
rect 13820 100 13850 230
rect 13990 100 14020 230
rect 14160 100 14190 230
rect 14330 100 14360 230
rect 14500 100 14530 230
rect 14670 100 14700 230
rect 14840 100 14870 230
rect 15010 100 15040 230
rect 15180 100 15210 230
rect 15350 100 15380 230
rect 15820 100 15850 230
rect 15990 100 16020 230
rect 16160 100 16190 230
rect 16330 100 16360 230
rect 16500 100 16530 230
rect 16670 100 16700 230
rect 16840 100 16870 230
rect 17010 100 17040 230
rect 17180 100 17210 230
rect 17350 100 17380 230
rect 17520 100 17550 230
rect 17690 100 17720 230
rect 17860 100 17890 230
rect 18030 100 18060 230
rect 18200 100 18230 230
rect 18370 100 18400 230
rect 18540 100 18570 230
rect 18710 100 18740 230
rect 18880 100 18910 230
rect 19050 100 19080 230
rect 19220 100 19250 230
rect 19390 100 19420 230
rect 19560 100 19590 230
rect 19730 100 19760 230
rect 19900 100 19930 230
rect 20070 100 20100 230
rect 20240 100 20270 230
rect 20410 100 20440 230
rect 20580 100 20610 230
rect 20750 100 20780 230
rect 20920 100 20950 230
rect 21090 100 21120 230
rect 21260 100 21290 230
rect 21430 100 21460 230
rect 21600 100 21630 230
rect 21770 100 21800 230
rect 21940 100 21970 230
rect 22110 100 22140 230
rect 22280 100 22310 230
rect 22450 100 22480 230
rect 22620 100 22650 230
rect 22790 100 22820 230
rect 22960 100 22990 230
rect 23130 100 23160 230
rect 23300 100 23330 230
rect 23470 100 23500 230
rect 23640 100 23670 230
rect 23810 100 23840 230
rect 23980 100 24010 230
rect 24150 100 24180 230
rect 24320 100 24350 230
rect 24490 100 24520 230
rect 24660 100 24690 230
rect 24830 100 24860 230
rect 25000 100 25030 230
rect 25170 100 25200 230
rect 25340 100 25370 230
rect 25510 100 25540 230
rect 25680 100 25710 230
rect 25850 100 25880 230
rect 26020 100 26050 230
rect 26190 100 26220 230
rect 26360 100 26390 230
rect 26530 100 26560 230
rect 26700 100 26730 230
rect 26870 100 26900 230
rect 27040 100 27070 230
rect 27210 100 27240 230
rect 27380 100 27410 230
rect 27550 100 27580 230
rect 27720 100 27750 230
rect 27890 100 27920 230
rect 28060 100 28090 230
rect 28230 100 28260 230
rect 28400 100 28430 230
rect 28570 100 28600 230
rect 28740 100 28770 230
rect 28910 100 28940 230
rect 29080 100 29110 230
rect 29250 100 29280 230
rect 29420 100 29450 230
rect 29590 100 29620 230
rect 29760 100 29790 230
rect 29930 100 29960 230
rect 30100 100 30130 230
rect 30270 100 30300 230
rect 30440 100 30470 230
rect 30610 100 30640 230
rect 30780 100 30810 230
rect 30950 100 30980 230
rect 31120 100 31150 230
rect 31290 100 31320 230
rect 31460 100 31490 230
rect 31630 100 31660 230
rect 31800 100 31830 230
rect 31970 100 32000 230
rect 32140 100 32170 230
rect 32310 100 32340 230
rect 32480 100 32510 230
rect 32650 100 32680 230
rect 32820 100 32850 230
rect 32990 100 33020 230
rect 33160 100 33190 230
rect 33330 100 33360 230
rect 33500 100 33530 230
rect 33670 100 33700 230
rect 33840 100 33870 230
rect 34010 100 34040 230
rect 34180 100 34210 230
rect 34350 100 34380 230
rect 34520 100 34550 230
rect 34690 100 34720 230
rect 34860 100 34890 230
rect 35030 100 35060 230
rect 35200 100 35230 230
rect 35370 100 35400 230
rect 35540 100 35570 230
rect 35710 100 35740 230
rect 35880 100 35910 230
rect 36050 100 36080 230
rect 36220 100 36250 230
rect 36390 100 36420 230
rect 36560 100 36590 230
rect 36730 100 36760 230
rect 36900 100 36930 230
rect 37070 100 37100 230
rect 37240 100 37270 230
rect 37410 100 37440 230
rect 37580 100 37610 230
rect 37750 100 37780 230
rect 37920 100 37950 230
rect 38090 100 38120 230
rect 38260 100 38290 230
rect 38430 100 38460 230
rect 38600 100 38630 230
rect 38770 100 38800 230
rect 38940 100 38970 230
rect 39110 100 39140 230
rect 39280 100 39310 230
rect 39450 100 39480 230
rect 39620 100 39650 230
rect 39790 100 39820 230
rect 39960 100 39990 230
rect 40130 100 40160 230
rect 40300 100 40330 230
rect 40470 100 40500 230
rect 40640 100 40670 230
rect 40810 100 40840 230
rect 40980 100 41010 230
rect 41150 100 41180 230
rect 41320 100 41350 230
rect 41490 100 41520 230
rect 41660 100 41690 230
rect 41830 100 41860 230
rect 42000 100 42030 230
rect 42170 100 42200 230
rect 42340 100 42370 230
rect 42510 100 42540 230
rect 42680 100 42710 230
rect 42850 100 42880 230
rect 43020 100 43050 230
rect 43190 100 43220 230
rect 43360 100 43390 230
rect 43530 100 43560 230
rect 43700 100 43730 230
rect 43870 100 43900 230
rect 44040 100 44070 230
rect 44210 100 44240 230
rect 44380 100 44410 230
rect 44550 100 44580 230
rect 44720 100 44750 230
rect 44890 100 44920 230
rect 45060 100 45090 230
rect 45230 100 45260 230
rect 45400 100 45430 230
rect 45570 100 45600 230
rect 45740 100 45770 230
rect 45910 100 45940 230
rect 46080 100 46110 230
rect 46250 100 46280 230
rect 46420 100 46450 230
rect 46590 100 46620 230
rect 46760 100 46790 230
rect 46930 100 46960 230
rect 47100 100 47130 230
rect 47270 100 47300 230
rect 47440 100 47470 230
rect 47610 100 47640 230
rect 47780 100 47810 230
rect 47950 100 47980 230
rect 48120 100 48150 230
rect 48290 100 48320 230
rect 48460 100 48490 230
rect 48630 100 48660 230
rect 48800 100 48830 230
rect 48970 100 49000 230
rect 49140 100 49170 230
rect 49310 100 49340 230
rect 49480 100 49510 230
rect 49650 100 49680 230
rect 49820 100 49850 230
rect 49990 100 50020 230
rect 50160 100 50190 230
rect 50330 100 50360 230
rect 50500 100 50530 230
rect 50670 100 50700 230
rect 50840 100 50870 230
rect 51010 100 51040 230
rect 51180 100 51210 230
rect 51350 100 51380 230
rect 51520 100 51550 230
rect 51690 100 51720 230
rect 51860 100 51890 230
rect 52030 100 52060 230
rect 52200 100 52230 230
rect 52370 100 52400 230
rect 52540 100 52570 230
rect 52710 100 52740 230
rect 52880 100 52910 230
rect 53050 100 53080 230
rect 53220 100 53250 230
rect 53390 100 53420 230
rect 53560 100 53590 230
rect 53730 100 53760 230
rect 53900 100 53930 230
rect 54070 100 54100 230
rect 54240 100 54270 230
rect 54410 100 54440 230
rect 54580 100 54610 230
rect 54750 100 54780 230
rect 54920 100 54950 230
rect 55090 100 55120 230
rect 55260 100 55290 230
rect 55430 100 55460 230
rect 55600 100 55630 230
rect 55770 100 55800 230
rect 55940 100 55970 230
rect 56110 100 56140 230
rect 56280 100 56310 230
rect 56450 100 56480 230
rect 56620 100 56650 230
rect 56790 100 56820 230
rect 56960 100 56990 230
rect 57130 100 57160 230
rect 57300 100 57330 230
rect 57470 100 57500 230
rect 57640 100 57670 230
rect 57810 100 57840 230
rect 57980 100 58010 230
rect 58150 100 58180 230
rect 58320 100 58350 230
rect 58490 100 58520 230
rect 58660 100 58690 230
rect 58830 100 58860 230
rect 59000 100 59030 230
rect 59170 100 59200 230
rect 50 10 160 30
rect 130 -40 160 10
rect 550 -40 580 0
rect 720 -40 750 0
rect 890 -40 920 0
rect 1060 -40 1090 0
rect 1620 -40 1650 0
rect 1790 -40 1820 0
rect 1960 -40 1990 0
rect 2130 -40 2160 0
rect 2300 -40 2330 0
rect 2470 -40 2500 0
rect 2640 -40 2670 0
rect 2810 -40 2840 0
rect 2980 -40 3010 0
rect 3150 -40 3180 0
rect 3320 -40 3350 0
rect 3490 -40 3520 0
rect 3660 -40 3690 0
rect 3830 -40 3860 0
rect 4000 -40 4030 0
rect 4170 -40 4200 0
rect 4640 -40 4670 0
rect 4810 -40 4840 0
rect 4980 -40 5010 0
rect 5150 -40 5180 0
rect 5320 -40 5350 0
rect 5490 -40 5520 0
rect 5660 -40 5690 0
rect 5830 -40 5860 0
rect 6000 -40 6030 0
rect 6170 -40 6200 0
rect 6340 -40 6370 0
rect 6510 -40 6540 0
rect 6680 -40 6710 0
rect 6850 -40 6880 0
rect 7020 -40 7050 0
rect 7190 -40 7220 0
rect 7360 -40 7390 0
rect 7530 -40 7560 0
rect 7700 -40 7730 0
rect 7870 -40 7900 0
rect 8040 -40 8070 0
rect 8210 -40 8240 0
rect 8380 -40 8410 0
rect 8550 -40 8580 0
rect 8720 -40 8750 0
rect 8890 -40 8920 0
rect 9060 -40 9090 0
rect 9230 -40 9260 0
rect 9400 -40 9430 0
rect 9570 -40 9600 0
rect 9740 -40 9770 0
rect 9910 -40 9940 0
rect 10080 -40 10110 0
rect 10250 -40 10280 0
rect 10420 -40 10450 0
rect 10590 -40 10620 0
rect 10760 -40 10790 0
rect 10930 -40 10960 0
rect 11100 -40 11130 0
rect 11270 -40 11300 0
rect 11440 -40 11470 0
rect 11610 -40 11640 0
rect 11780 -40 11810 0
rect 11950 -40 11980 0
rect 12120 -40 12150 0
rect 12290 -40 12320 0
rect 12460 -40 12490 0
rect 12630 -40 12660 0
rect 12800 -40 12830 0
rect 12970 -40 13000 0
rect 13140 -40 13170 0
rect 13310 -40 13340 0
rect 13480 -40 13510 0
rect 13650 -40 13680 0
rect 13820 -40 13850 0
rect 13990 -40 14020 0
rect 14160 -40 14190 0
rect 14330 -40 14360 0
rect 14500 -40 14530 0
rect 14670 -40 14700 0
rect 14840 -40 14870 0
rect 15010 -40 15040 0
rect 15180 -40 15210 0
rect 15350 -40 15380 0
rect 15820 -40 15850 0
rect 15990 -40 16020 0
rect 16160 -40 16190 0
rect 16330 -40 16360 0
rect 16500 -40 16530 0
rect 16670 -40 16700 0
rect 16840 -40 16870 0
rect 17010 -40 17040 0
rect 17180 -40 17210 0
rect 17350 -40 17380 0
rect 17520 -40 17550 0
rect 17690 -40 17720 0
rect 17860 -40 17890 0
rect 18030 -40 18060 0
rect 18200 -40 18230 0
rect 18370 -40 18400 0
rect 18540 -40 18570 0
rect 18710 -40 18740 0
rect 18880 -40 18910 0
rect 19050 -40 19080 0
rect 19220 -40 19250 0
rect 19390 -40 19420 0
rect 19560 -40 19590 0
rect 19730 -40 19760 0
rect 19900 -40 19930 0
rect 20070 -40 20100 0
rect 20240 -40 20270 0
rect 20410 -40 20440 0
rect 20580 -40 20610 0
rect 20750 -40 20780 0
rect 20920 -40 20950 0
rect 21090 -40 21120 0
rect 21260 -40 21290 0
rect 21430 -40 21460 0
rect 21600 -40 21630 0
rect 21770 -40 21800 0
rect 21940 -40 21970 0
rect 22110 -40 22140 0
rect 22280 -40 22310 0
rect 22450 -40 22480 0
rect 22620 -40 22650 0
rect 22790 -40 22820 0
rect 22960 -40 22990 0
rect 23130 -40 23160 0
rect 23300 -40 23330 0
rect 23470 -40 23500 0
rect 23640 -40 23670 0
rect 23810 -40 23840 0
rect 23980 -40 24010 0
rect 24150 -40 24180 0
rect 24320 -40 24350 0
rect 24490 -40 24520 0
rect 24660 -40 24690 0
rect 24830 -40 24860 0
rect 25000 -40 25030 0
rect 25170 -40 25200 0
rect 25340 -40 25370 0
rect 25510 -40 25540 0
rect 25680 -40 25710 0
rect 25850 -40 25880 0
rect 26020 -40 26050 0
rect 26190 -40 26220 0
rect 26360 -40 26390 0
rect 26530 -40 26560 0
rect 26700 -40 26730 0
rect 26870 -40 26900 0
rect 27040 -40 27070 0
rect 27210 -40 27240 0
rect 27380 -40 27410 0
rect 27550 -40 27580 0
rect 27720 -40 27750 0
rect 27890 -40 27920 0
rect 28060 -40 28090 0
rect 28230 -40 28260 0
rect 28400 -40 28430 0
rect 28570 -40 28600 0
rect 28740 -40 28770 0
rect 28910 -40 28940 0
rect 29080 -40 29110 0
rect 29250 -40 29280 0
rect 29420 -40 29450 0
rect 29590 -40 29620 0
rect 29760 -40 29790 0
rect 29930 -40 29960 0
rect 30100 -40 30130 0
rect 30270 -40 30300 0
rect 30440 -40 30470 0
rect 30610 -40 30640 0
rect 30780 -40 30810 0
rect 30950 -40 30980 0
rect 31120 -40 31150 0
rect 31290 -40 31320 0
rect 31460 -40 31490 0
rect 31630 -40 31660 0
rect 31800 -40 31830 0
rect 31970 -40 32000 0
rect 32140 -40 32170 0
rect 32310 -40 32340 0
rect 32480 -40 32510 0
rect 32650 -40 32680 0
rect 32820 -40 32850 0
rect 32990 -40 33020 0
rect 33160 -40 33190 0
rect 33330 -40 33360 0
rect 33500 -40 33530 0
rect 33670 -40 33700 0
rect 33840 -40 33870 0
rect 34010 -40 34040 0
rect 34180 -40 34210 0
rect 34350 -40 34380 0
rect 34520 -40 34550 0
rect 34690 -40 34720 0
rect 34860 -40 34890 0
rect 35030 -40 35060 0
rect 35200 -40 35230 0
rect 35370 -40 35400 0
rect 35540 -40 35570 0
rect 35710 -40 35740 0
rect 35880 -40 35910 0
rect 36050 -40 36080 0
rect 36220 -40 36250 0
rect 36390 -40 36420 0
rect 36560 -40 36590 0
rect 36730 -40 36760 0
rect 36900 -40 36930 0
rect 37070 -40 37100 0
rect 37240 -40 37270 0
rect 37410 -40 37440 0
rect 37580 -40 37610 0
rect 37750 -40 37780 0
rect 37920 -40 37950 0
rect 38090 -40 38120 0
rect 38260 -40 38290 0
rect 38430 -40 38460 0
rect 38600 -40 38630 0
rect 38770 -40 38800 0
rect 38940 -40 38970 0
rect 39110 -40 39140 0
rect 39280 -40 39310 0
rect 39450 -40 39480 0
rect 39620 -40 39650 0
rect 39790 -40 39820 0
rect 39960 -40 39990 0
rect 40130 -40 40160 0
rect 40300 -40 40330 0
rect 40470 -40 40500 0
rect 40640 -40 40670 0
rect 40810 -40 40840 0
rect 40980 -40 41010 0
rect 41150 -40 41180 0
rect 41320 -40 41350 0
rect 41490 -40 41520 0
rect 41660 -40 41690 0
rect 41830 -40 41860 0
rect 42000 -40 42030 0
rect 42170 -40 42200 0
rect 42340 -40 42370 0
rect 42510 -40 42540 0
rect 42680 -40 42710 0
rect 42850 -40 42880 0
rect 43020 -40 43050 0
rect 43190 -40 43220 0
rect 43360 -40 43390 0
rect 43530 -40 43560 0
rect 43700 -40 43730 0
rect 43870 -40 43900 0
rect 44040 -40 44070 0
rect 44210 -40 44240 0
rect 44380 -40 44410 0
rect 44550 -40 44580 0
rect 44720 -40 44750 0
rect 44890 -40 44920 0
rect 45060 -40 45090 0
rect 45230 -40 45260 0
rect 45400 -40 45430 0
rect 45570 -40 45600 0
rect 45740 -40 45770 0
rect 45910 -40 45940 0
rect 46080 -40 46110 0
rect 46250 -40 46280 0
rect 46420 -40 46450 0
rect 46590 -40 46620 0
rect 46760 -40 46790 0
rect 46930 -40 46960 0
rect 47100 -40 47130 0
rect 47270 -40 47300 0
rect 47440 -40 47470 0
rect 47610 -40 47640 0
rect 47780 -40 47810 0
rect 47950 -40 47980 0
rect 48120 -40 48150 0
rect 48290 -40 48320 0
rect 48460 -40 48490 0
rect 48630 -40 48660 0
rect 48800 -40 48830 0
rect 48970 -40 49000 0
rect 49140 -40 49170 0
rect 49310 -40 49340 0
rect 49480 -40 49510 0
rect 49650 -40 49680 0
rect 49820 -40 49850 0
rect 49990 -40 50020 0
rect 50160 -40 50190 0
rect 50330 -40 50360 0
rect 50500 -40 50530 0
rect 50670 -40 50700 0
rect 50840 -40 50870 0
rect 51010 -40 51040 0
rect 51180 -40 51210 0
rect 51350 -40 51380 0
rect 51520 -40 51550 0
rect 51690 -40 51720 0
rect 51860 -40 51890 0
rect 52030 -40 52060 0
rect 52200 -40 52230 0
rect 52370 -40 52400 0
rect 52540 -40 52570 0
rect 52710 -40 52740 0
rect 52880 -40 52910 0
rect 53050 -40 53080 0
rect 53220 -40 53250 0
rect 53390 -40 53420 0
rect 53560 -40 53590 0
rect 53730 -40 53760 0
rect 53900 -40 53930 0
rect 54070 -40 54100 0
rect 54240 -40 54270 0
rect 54410 -40 54440 0
rect 54580 -40 54610 0
rect 54750 -40 54780 0
rect 54920 -40 54950 0
rect 55090 -40 55120 0
rect 55260 -40 55290 0
rect 55430 -40 55460 0
rect 55600 -40 55630 0
rect 55770 -40 55800 0
rect 55940 -40 55970 0
rect 56110 -40 56140 0
rect 56280 -40 56310 0
rect 56450 -40 56480 0
rect 56620 -40 56650 0
rect 56790 -40 56820 0
rect 56960 -40 56990 0
rect 57130 -40 57160 0
rect 57300 -40 57330 0
rect 57470 -40 57500 0
rect 57640 -40 57670 0
rect 57810 -40 57840 0
rect 57980 -40 58010 0
rect 58150 -40 58180 0
rect 58320 -40 58350 0
rect 58490 -40 58520 0
rect 58660 -40 58690 0
rect 58830 -40 58860 0
rect 59000 -40 59030 0
rect 59170 -40 59200 0
rect 510 -60 620 -40
rect 510 -120 530 -60
rect 600 -120 620 -60
rect 510 -140 620 -120
rect 680 -60 790 -40
rect 680 -120 700 -60
rect 770 -120 790 -60
rect 680 -140 790 -120
rect 850 -60 960 -40
rect 850 -120 870 -60
rect 940 -120 960 -60
rect 850 -140 960 -120
rect 1020 -60 1130 -40
rect 1020 -120 1040 -60
rect 1110 -120 1130 -60
rect 1020 -140 1130 -120
rect 1580 -60 1690 -40
rect 1580 -120 1600 -60
rect 1670 -120 1690 -60
rect 1580 -140 1690 -120
rect 1750 -60 1860 -40
rect 1750 -120 1770 -60
rect 1840 -120 1860 -60
rect 1750 -140 1860 -120
rect 1920 -60 2030 -40
rect 1920 -120 1940 -60
rect 2010 -120 2030 -60
rect 1920 -140 2030 -120
rect 2090 -60 2200 -40
rect 2090 -120 2110 -60
rect 2180 -120 2200 -60
rect 2090 -140 2200 -120
rect 2260 -60 2370 -40
rect 2260 -120 2280 -60
rect 2350 -120 2370 -60
rect 2260 -140 2370 -120
rect 2430 -60 2540 -40
rect 2430 -120 2450 -60
rect 2520 -120 2540 -60
rect 2430 -140 2540 -120
rect 2600 -60 2710 -40
rect 2600 -120 2620 -60
rect 2690 -120 2710 -60
rect 2600 -140 2710 -120
rect 2770 -60 2880 -40
rect 2770 -120 2790 -60
rect 2860 -120 2880 -60
rect 2770 -140 2880 -120
rect 2940 -60 3050 -40
rect 2940 -120 2960 -60
rect 3030 -120 3050 -60
rect 2940 -140 3050 -120
rect 3110 -60 3220 -40
rect 3110 -120 3130 -60
rect 3200 -120 3220 -60
rect 3110 -140 3220 -120
rect 3280 -60 3390 -40
rect 3280 -120 3300 -60
rect 3370 -120 3390 -60
rect 3280 -140 3390 -120
rect 3450 -60 3560 -40
rect 3450 -120 3470 -60
rect 3540 -120 3560 -60
rect 3450 -140 3560 -120
rect 3620 -60 3730 -40
rect 3620 -120 3640 -60
rect 3710 -120 3730 -60
rect 3620 -140 3730 -120
rect 3790 -60 3900 -40
rect 3790 -120 3810 -60
rect 3880 -120 3900 -60
rect 3790 -140 3900 -120
rect 3960 -60 4070 -40
rect 3960 -120 3980 -60
rect 4050 -120 4070 -60
rect 3960 -140 4070 -120
rect 4130 -60 4240 -40
rect 4130 -120 4150 -60
rect 4220 -120 4240 -60
rect 4130 -140 4240 -120
rect 4600 -60 4710 -40
rect 4600 -120 4620 -60
rect 4690 -120 4710 -60
rect 4600 -140 4710 -120
rect 4770 -60 4880 -40
rect 4770 -120 4790 -60
rect 4860 -120 4880 -60
rect 4770 -140 4880 -120
rect 4940 -60 5050 -40
rect 4940 -120 4960 -60
rect 5030 -120 5050 -60
rect 4940 -140 5050 -120
rect 5110 -60 5220 -40
rect 5110 -120 5130 -60
rect 5200 -120 5220 -60
rect 5110 -140 5220 -120
rect 5280 -60 5390 -40
rect 5280 -120 5300 -60
rect 5370 -120 5390 -60
rect 5280 -140 5390 -120
rect 5450 -60 5560 -40
rect 5450 -120 5470 -60
rect 5540 -120 5560 -60
rect 5450 -140 5560 -120
rect 5620 -60 5730 -40
rect 5620 -120 5640 -60
rect 5710 -120 5730 -60
rect 5620 -140 5730 -120
rect 5790 -60 5900 -40
rect 5790 -120 5810 -60
rect 5880 -120 5900 -60
rect 5790 -140 5900 -120
rect 5960 -60 6070 -40
rect 5960 -120 5980 -60
rect 6050 -120 6070 -60
rect 5960 -140 6070 -120
rect 6130 -60 6240 -40
rect 6130 -120 6150 -60
rect 6220 -120 6240 -60
rect 6130 -140 6240 -120
rect 6300 -60 6410 -40
rect 6300 -120 6320 -60
rect 6390 -120 6410 -60
rect 6300 -140 6410 -120
rect 6470 -60 6580 -40
rect 6470 -120 6490 -60
rect 6560 -120 6580 -60
rect 6470 -140 6580 -120
rect 6640 -60 6750 -40
rect 6640 -120 6660 -60
rect 6730 -120 6750 -60
rect 6640 -140 6750 -120
rect 6810 -60 6920 -40
rect 6810 -120 6830 -60
rect 6900 -120 6920 -60
rect 6810 -140 6920 -120
rect 6980 -60 7090 -40
rect 6980 -120 7000 -60
rect 7070 -120 7090 -60
rect 6980 -140 7090 -120
rect 7150 -60 7260 -40
rect 7150 -120 7170 -60
rect 7240 -120 7260 -60
rect 7150 -140 7260 -120
rect 7320 -60 7430 -40
rect 7320 -120 7340 -60
rect 7410 -120 7430 -60
rect 7320 -140 7430 -120
rect 7490 -60 7600 -40
rect 7490 -120 7510 -60
rect 7580 -120 7600 -60
rect 7490 -140 7600 -120
rect 7660 -60 7770 -40
rect 7660 -120 7680 -60
rect 7750 -120 7770 -60
rect 7660 -140 7770 -120
rect 7830 -60 7940 -40
rect 7830 -120 7850 -60
rect 7920 -120 7940 -60
rect 7830 -140 7940 -120
rect 8000 -60 8110 -40
rect 8000 -120 8020 -60
rect 8090 -120 8110 -60
rect 8000 -140 8110 -120
rect 8170 -60 8280 -40
rect 8170 -120 8190 -60
rect 8260 -120 8280 -60
rect 8170 -140 8280 -120
rect 8340 -60 8450 -40
rect 8340 -120 8360 -60
rect 8430 -120 8450 -60
rect 8340 -140 8450 -120
rect 8510 -60 8620 -40
rect 8510 -120 8530 -60
rect 8600 -120 8620 -60
rect 8510 -140 8620 -120
rect 8680 -60 8790 -40
rect 8680 -120 8700 -60
rect 8770 -120 8790 -60
rect 8680 -140 8790 -120
rect 8850 -60 8960 -40
rect 8850 -120 8870 -60
rect 8940 -120 8960 -60
rect 8850 -140 8960 -120
rect 9020 -60 9130 -40
rect 9020 -120 9040 -60
rect 9110 -120 9130 -60
rect 9020 -140 9130 -120
rect 9190 -60 9300 -40
rect 9190 -120 9210 -60
rect 9280 -120 9300 -60
rect 9190 -140 9300 -120
rect 9360 -60 9470 -40
rect 9360 -120 9380 -60
rect 9450 -120 9470 -60
rect 9360 -140 9470 -120
rect 9530 -60 9640 -40
rect 9530 -120 9550 -60
rect 9620 -120 9640 -60
rect 9530 -140 9640 -120
rect 9700 -60 9810 -40
rect 9700 -120 9720 -60
rect 9790 -120 9810 -60
rect 9700 -140 9810 -120
rect 9870 -60 9980 -40
rect 9870 -120 9890 -60
rect 9960 -120 9980 -60
rect 9870 -140 9980 -120
rect 10040 -60 10150 -40
rect 10040 -120 10060 -60
rect 10130 -120 10150 -60
rect 10040 -140 10150 -120
rect 10210 -60 10320 -40
rect 10210 -120 10230 -60
rect 10300 -120 10320 -60
rect 10210 -140 10320 -120
rect 10380 -60 10490 -40
rect 10380 -120 10400 -60
rect 10470 -120 10490 -60
rect 10380 -140 10490 -120
rect 10550 -60 10660 -40
rect 10550 -120 10570 -60
rect 10640 -120 10660 -60
rect 10550 -140 10660 -120
rect 10720 -60 10830 -40
rect 10720 -120 10740 -60
rect 10810 -120 10830 -60
rect 10720 -140 10830 -120
rect 10890 -60 11000 -40
rect 10890 -120 10910 -60
rect 10980 -120 11000 -60
rect 10890 -140 11000 -120
rect 11060 -60 11170 -40
rect 11060 -120 11080 -60
rect 11150 -120 11170 -60
rect 11060 -140 11170 -120
rect 11230 -60 11340 -40
rect 11230 -120 11250 -60
rect 11320 -120 11340 -60
rect 11230 -140 11340 -120
rect 11400 -60 11510 -40
rect 11400 -120 11420 -60
rect 11490 -120 11510 -60
rect 11400 -140 11510 -120
rect 11570 -60 11680 -40
rect 11570 -120 11590 -60
rect 11660 -120 11680 -60
rect 11570 -140 11680 -120
rect 11740 -60 11850 -40
rect 11740 -120 11760 -60
rect 11830 -120 11850 -60
rect 11740 -140 11850 -120
rect 11910 -60 12020 -40
rect 11910 -120 11930 -60
rect 12000 -120 12020 -60
rect 11910 -140 12020 -120
rect 12080 -60 12190 -40
rect 12080 -120 12100 -60
rect 12170 -120 12190 -60
rect 12080 -140 12190 -120
rect 12250 -60 12360 -40
rect 12250 -120 12270 -60
rect 12340 -120 12360 -60
rect 12250 -140 12360 -120
rect 12420 -60 12530 -40
rect 12420 -120 12440 -60
rect 12510 -120 12530 -60
rect 12420 -140 12530 -120
rect 12590 -60 12700 -40
rect 12590 -120 12610 -60
rect 12680 -120 12700 -60
rect 12590 -140 12700 -120
rect 12760 -60 12870 -40
rect 12760 -120 12780 -60
rect 12850 -120 12870 -60
rect 12760 -140 12870 -120
rect 12930 -60 13040 -40
rect 12930 -120 12950 -60
rect 13020 -120 13040 -60
rect 12930 -140 13040 -120
rect 13100 -60 13210 -40
rect 13100 -120 13120 -60
rect 13190 -120 13210 -60
rect 13100 -140 13210 -120
rect 13270 -60 13380 -40
rect 13270 -120 13290 -60
rect 13360 -120 13380 -60
rect 13270 -140 13380 -120
rect 13440 -60 13550 -40
rect 13440 -120 13460 -60
rect 13530 -120 13550 -60
rect 13440 -140 13550 -120
rect 13610 -60 13720 -40
rect 13610 -120 13630 -60
rect 13700 -120 13720 -60
rect 13610 -140 13720 -120
rect 13780 -60 13890 -40
rect 13780 -120 13800 -60
rect 13870 -120 13890 -60
rect 13780 -140 13890 -120
rect 13950 -60 14060 -40
rect 13950 -120 13970 -60
rect 14040 -120 14060 -60
rect 13950 -140 14060 -120
rect 14120 -60 14230 -40
rect 14120 -120 14140 -60
rect 14210 -120 14230 -60
rect 14120 -140 14230 -120
rect 14290 -60 14400 -40
rect 14290 -120 14310 -60
rect 14380 -120 14400 -60
rect 14290 -140 14400 -120
rect 14460 -60 14570 -40
rect 14460 -120 14480 -60
rect 14550 -120 14570 -60
rect 14460 -140 14570 -120
rect 14630 -60 14740 -40
rect 14630 -120 14650 -60
rect 14720 -120 14740 -60
rect 14630 -140 14740 -120
rect 14800 -60 14910 -40
rect 14800 -120 14820 -60
rect 14890 -120 14910 -60
rect 14800 -140 14910 -120
rect 14970 -60 15080 -40
rect 14970 -120 14990 -60
rect 15060 -120 15080 -60
rect 14970 -140 15080 -120
rect 15140 -60 15250 -40
rect 15140 -120 15160 -60
rect 15230 -120 15250 -60
rect 15140 -140 15250 -120
rect 15310 -60 15420 -40
rect 15310 -120 15330 -60
rect 15400 -120 15420 -60
rect 15310 -140 15420 -120
rect 15780 -60 15890 -40
rect 15780 -120 15800 -60
rect 15870 -120 15890 -60
rect 15780 -140 15890 -120
rect 15950 -60 16060 -40
rect 15950 -120 15970 -60
rect 16040 -120 16060 -60
rect 15950 -140 16060 -120
rect 16120 -60 16230 -40
rect 16120 -120 16140 -60
rect 16210 -120 16230 -60
rect 16120 -140 16230 -120
rect 16290 -60 16400 -40
rect 16290 -120 16310 -60
rect 16380 -120 16400 -60
rect 16290 -140 16400 -120
rect 16460 -60 16570 -40
rect 16460 -120 16480 -60
rect 16550 -120 16570 -60
rect 16460 -140 16570 -120
rect 16630 -60 16740 -40
rect 16630 -120 16650 -60
rect 16720 -120 16740 -60
rect 16630 -140 16740 -120
rect 16800 -60 16910 -40
rect 16800 -120 16820 -60
rect 16890 -120 16910 -60
rect 16800 -140 16910 -120
rect 16970 -60 17080 -40
rect 16970 -120 16990 -60
rect 17060 -120 17080 -60
rect 16970 -140 17080 -120
rect 17140 -60 17250 -40
rect 17140 -120 17160 -60
rect 17230 -120 17250 -60
rect 17140 -140 17250 -120
rect 17310 -60 17420 -40
rect 17310 -120 17330 -60
rect 17400 -120 17420 -60
rect 17310 -140 17420 -120
rect 17480 -60 17590 -40
rect 17480 -120 17500 -60
rect 17570 -120 17590 -60
rect 17480 -140 17590 -120
rect 17650 -60 17760 -40
rect 17650 -120 17670 -60
rect 17740 -120 17760 -60
rect 17650 -140 17760 -120
rect 17820 -60 17930 -40
rect 17820 -120 17840 -60
rect 17910 -120 17930 -60
rect 17820 -140 17930 -120
rect 17990 -60 18100 -40
rect 17990 -120 18010 -60
rect 18080 -120 18100 -60
rect 17990 -140 18100 -120
rect 18160 -60 18270 -40
rect 18160 -120 18180 -60
rect 18250 -120 18270 -60
rect 18160 -140 18270 -120
rect 18330 -60 18440 -40
rect 18330 -120 18350 -60
rect 18420 -120 18440 -60
rect 18330 -140 18440 -120
rect 18500 -60 18610 -40
rect 18500 -120 18520 -60
rect 18590 -120 18610 -60
rect 18500 -140 18610 -120
rect 18670 -60 18780 -40
rect 18670 -120 18690 -60
rect 18760 -120 18780 -60
rect 18670 -140 18780 -120
rect 18840 -60 18950 -40
rect 18840 -120 18860 -60
rect 18930 -120 18950 -60
rect 18840 -140 18950 -120
rect 19010 -60 19120 -40
rect 19010 -120 19030 -60
rect 19100 -120 19120 -60
rect 19010 -140 19120 -120
rect 19180 -60 19290 -40
rect 19180 -120 19200 -60
rect 19270 -120 19290 -60
rect 19180 -140 19290 -120
rect 19350 -60 19460 -40
rect 19350 -120 19370 -60
rect 19440 -120 19460 -60
rect 19350 -140 19460 -120
rect 19520 -60 19630 -40
rect 19520 -120 19540 -60
rect 19610 -120 19630 -60
rect 19520 -140 19630 -120
rect 19690 -60 19800 -40
rect 19690 -120 19710 -60
rect 19780 -120 19800 -60
rect 19690 -140 19800 -120
rect 19860 -60 19970 -40
rect 19860 -120 19880 -60
rect 19950 -120 19970 -60
rect 19860 -140 19970 -120
rect 20030 -60 20140 -40
rect 20030 -120 20050 -60
rect 20120 -120 20140 -60
rect 20030 -140 20140 -120
rect 20200 -60 20310 -40
rect 20200 -120 20220 -60
rect 20290 -120 20310 -60
rect 20200 -140 20310 -120
rect 20370 -60 20480 -40
rect 20370 -120 20390 -60
rect 20460 -120 20480 -60
rect 20370 -140 20480 -120
rect 20540 -60 20650 -40
rect 20540 -120 20560 -60
rect 20630 -120 20650 -60
rect 20540 -140 20650 -120
rect 20710 -60 20820 -40
rect 20710 -120 20730 -60
rect 20800 -120 20820 -60
rect 20710 -140 20820 -120
rect 20880 -60 20990 -40
rect 20880 -120 20900 -60
rect 20970 -120 20990 -60
rect 20880 -140 20990 -120
rect 21050 -60 21160 -40
rect 21050 -120 21070 -60
rect 21140 -120 21160 -60
rect 21050 -140 21160 -120
rect 21220 -60 21330 -40
rect 21220 -120 21240 -60
rect 21310 -120 21330 -60
rect 21220 -140 21330 -120
rect 21390 -60 21500 -40
rect 21390 -120 21410 -60
rect 21480 -120 21500 -60
rect 21390 -140 21500 -120
rect 21560 -60 21670 -40
rect 21560 -120 21580 -60
rect 21650 -120 21670 -60
rect 21560 -140 21670 -120
rect 21730 -60 21840 -40
rect 21730 -120 21750 -60
rect 21820 -120 21840 -60
rect 21730 -140 21840 -120
rect 21900 -60 22010 -40
rect 21900 -120 21920 -60
rect 21990 -120 22010 -60
rect 21900 -140 22010 -120
rect 22070 -60 22180 -40
rect 22070 -120 22090 -60
rect 22160 -120 22180 -60
rect 22070 -140 22180 -120
rect 22240 -60 22350 -40
rect 22240 -120 22260 -60
rect 22330 -120 22350 -60
rect 22240 -140 22350 -120
rect 22410 -60 22520 -40
rect 22410 -120 22430 -60
rect 22500 -120 22520 -60
rect 22410 -140 22520 -120
rect 22580 -60 22690 -40
rect 22580 -120 22600 -60
rect 22670 -120 22690 -60
rect 22580 -140 22690 -120
rect 22750 -60 22860 -40
rect 22750 -120 22770 -60
rect 22840 -120 22860 -60
rect 22750 -140 22860 -120
rect 22920 -60 23030 -40
rect 22920 -120 22940 -60
rect 23010 -120 23030 -60
rect 22920 -140 23030 -120
rect 23090 -60 23200 -40
rect 23090 -120 23110 -60
rect 23180 -120 23200 -60
rect 23090 -140 23200 -120
rect 23260 -60 23370 -40
rect 23260 -120 23280 -60
rect 23350 -120 23370 -60
rect 23260 -140 23370 -120
rect 23430 -60 23540 -40
rect 23430 -120 23450 -60
rect 23520 -120 23540 -60
rect 23430 -140 23540 -120
rect 23600 -60 23710 -40
rect 23600 -120 23620 -60
rect 23690 -120 23710 -60
rect 23600 -140 23710 -120
rect 23770 -60 23880 -40
rect 23770 -120 23790 -60
rect 23860 -120 23880 -60
rect 23770 -140 23880 -120
rect 23940 -60 24050 -40
rect 23940 -120 23960 -60
rect 24030 -120 24050 -60
rect 23940 -140 24050 -120
rect 24110 -60 24220 -40
rect 24110 -120 24130 -60
rect 24200 -120 24220 -60
rect 24110 -140 24220 -120
rect 24280 -60 24390 -40
rect 24280 -120 24300 -60
rect 24370 -120 24390 -60
rect 24280 -140 24390 -120
rect 24450 -60 24560 -40
rect 24450 -120 24470 -60
rect 24540 -120 24560 -60
rect 24450 -140 24560 -120
rect 24620 -60 24730 -40
rect 24620 -120 24640 -60
rect 24710 -120 24730 -60
rect 24620 -140 24730 -120
rect 24790 -60 24900 -40
rect 24790 -120 24810 -60
rect 24880 -120 24900 -60
rect 24790 -140 24900 -120
rect 24960 -60 25070 -40
rect 24960 -120 24980 -60
rect 25050 -120 25070 -60
rect 24960 -140 25070 -120
rect 25130 -60 25240 -40
rect 25130 -120 25150 -60
rect 25220 -120 25240 -60
rect 25130 -140 25240 -120
rect 25300 -60 25410 -40
rect 25300 -120 25320 -60
rect 25390 -120 25410 -60
rect 25300 -140 25410 -120
rect 25470 -60 25580 -40
rect 25470 -120 25490 -60
rect 25560 -120 25580 -60
rect 25470 -140 25580 -120
rect 25640 -60 25750 -40
rect 25640 -120 25660 -60
rect 25730 -120 25750 -60
rect 25640 -140 25750 -120
rect 25810 -60 25920 -40
rect 25810 -120 25830 -60
rect 25900 -120 25920 -60
rect 25810 -140 25920 -120
rect 25980 -60 26090 -40
rect 25980 -120 26000 -60
rect 26070 -120 26090 -60
rect 25980 -140 26090 -120
rect 26150 -60 26260 -40
rect 26150 -120 26170 -60
rect 26240 -120 26260 -60
rect 26150 -140 26260 -120
rect 26320 -60 26430 -40
rect 26320 -120 26340 -60
rect 26410 -120 26430 -60
rect 26320 -140 26430 -120
rect 26490 -60 26600 -40
rect 26490 -120 26510 -60
rect 26580 -120 26600 -60
rect 26490 -140 26600 -120
rect 26660 -60 26770 -40
rect 26660 -120 26680 -60
rect 26750 -120 26770 -60
rect 26660 -140 26770 -120
rect 26830 -60 26940 -40
rect 26830 -120 26850 -60
rect 26920 -120 26940 -60
rect 26830 -140 26940 -120
rect 27000 -60 27110 -40
rect 27000 -120 27020 -60
rect 27090 -120 27110 -60
rect 27000 -140 27110 -120
rect 27170 -60 27280 -40
rect 27170 -120 27190 -60
rect 27260 -120 27280 -60
rect 27170 -140 27280 -120
rect 27340 -60 27450 -40
rect 27340 -120 27360 -60
rect 27430 -120 27450 -60
rect 27340 -140 27450 -120
rect 27510 -60 27620 -40
rect 27510 -120 27530 -60
rect 27600 -120 27620 -60
rect 27510 -140 27620 -120
rect 27680 -60 27790 -40
rect 27680 -120 27700 -60
rect 27770 -120 27790 -60
rect 27680 -140 27790 -120
rect 27850 -60 27960 -40
rect 27850 -120 27870 -60
rect 27940 -120 27960 -60
rect 27850 -140 27960 -120
rect 28020 -60 28130 -40
rect 28020 -120 28040 -60
rect 28110 -120 28130 -60
rect 28020 -140 28130 -120
rect 28190 -60 28300 -40
rect 28190 -120 28210 -60
rect 28280 -120 28300 -60
rect 28190 -140 28300 -120
rect 28360 -60 28470 -40
rect 28360 -120 28380 -60
rect 28450 -120 28470 -60
rect 28360 -140 28470 -120
rect 28530 -60 28640 -40
rect 28530 -120 28550 -60
rect 28620 -120 28640 -60
rect 28530 -140 28640 -120
rect 28700 -60 28810 -40
rect 28700 -120 28720 -60
rect 28790 -120 28810 -60
rect 28700 -140 28810 -120
rect 28870 -60 28980 -40
rect 28870 -120 28890 -60
rect 28960 -120 28980 -60
rect 28870 -140 28980 -120
rect 29040 -60 29150 -40
rect 29040 -120 29060 -60
rect 29130 -120 29150 -60
rect 29040 -140 29150 -120
rect 29210 -60 29320 -40
rect 29210 -120 29230 -60
rect 29300 -120 29320 -60
rect 29210 -140 29320 -120
rect 29380 -60 29490 -40
rect 29380 -120 29400 -60
rect 29470 -120 29490 -60
rect 29380 -140 29490 -120
rect 29550 -60 29660 -40
rect 29550 -120 29570 -60
rect 29640 -120 29660 -60
rect 29550 -140 29660 -120
rect 29720 -60 29830 -40
rect 29720 -120 29740 -60
rect 29810 -120 29830 -60
rect 29720 -140 29830 -120
rect 29890 -60 30000 -40
rect 29890 -120 29910 -60
rect 29980 -120 30000 -60
rect 29890 -140 30000 -120
rect 30060 -60 30170 -40
rect 30060 -120 30080 -60
rect 30150 -120 30170 -60
rect 30060 -140 30170 -120
rect 30230 -60 30340 -40
rect 30230 -120 30250 -60
rect 30320 -120 30340 -60
rect 30230 -140 30340 -120
rect 30400 -60 30510 -40
rect 30400 -120 30420 -60
rect 30490 -120 30510 -60
rect 30400 -140 30510 -120
rect 30570 -60 30680 -40
rect 30570 -120 30590 -60
rect 30660 -120 30680 -60
rect 30570 -140 30680 -120
rect 30740 -60 30850 -40
rect 30740 -120 30760 -60
rect 30830 -120 30850 -60
rect 30740 -140 30850 -120
rect 30910 -60 31020 -40
rect 30910 -120 30930 -60
rect 31000 -120 31020 -60
rect 30910 -140 31020 -120
rect 31080 -60 31190 -40
rect 31080 -120 31100 -60
rect 31170 -120 31190 -60
rect 31080 -140 31190 -120
rect 31250 -60 31360 -40
rect 31250 -120 31270 -60
rect 31340 -120 31360 -60
rect 31250 -140 31360 -120
rect 31420 -60 31530 -40
rect 31420 -120 31440 -60
rect 31510 -120 31530 -60
rect 31420 -140 31530 -120
rect 31590 -60 31700 -40
rect 31590 -120 31610 -60
rect 31680 -120 31700 -60
rect 31590 -140 31700 -120
rect 31760 -60 31870 -40
rect 31760 -120 31780 -60
rect 31850 -120 31870 -60
rect 31760 -140 31870 -120
rect 31930 -60 32040 -40
rect 31930 -120 31950 -60
rect 32020 -120 32040 -60
rect 31930 -140 32040 -120
rect 32100 -60 32210 -40
rect 32100 -120 32120 -60
rect 32190 -120 32210 -60
rect 32100 -140 32210 -120
rect 32270 -60 32380 -40
rect 32270 -120 32290 -60
rect 32360 -120 32380 -60
rect 32270 -140 32380 -120
rect 32440 -60 32550 -40
rect 32440 -120 32460 -60
rect 32530 -120 32550 -60
rect 32440 -140 32550 -120
rect 32610 -60 32720 -40
rect 32610 -120 32630 -60
rect 32700 -120 32720 -60
rect 32610 -140 32720 -120
rect 32780 -60 32890 -40
rect 32780 -120 32800 -60
rect 32870 -120 32890 -60
rect 32780 -140 32890 -120
rect 32950 -60 33060 -40
rect 32950 -120 32970 -60
rect 33040 -120 33060 -60
rect 32950 -140 33060 -120
rect 33120 -60 33230 -40
rect 33120 -120 33140 -60
rect 33210 -120 33230 -60
rect 33120 -140 33230 -120
rect 33290 -60 33400 -40
rect 33290 -120 33310 -60
rect 33380 -120 33400 -60
rect 33290 -140 33400 -120
rect 33460 -60 33570 -40
rect 33460 -120 33480 -60
rect 33550 -120 33570 -60
rect 33460 -140 33570 -120
rect 33630 -60 33740 -40
rect 33630 -120 33650 -60
rect 33720 -120 33740 -60
rect 33630 -140 33740 -120
rect 33800 -60 33910 -40
rect 33800 -120 33820 -60
rect 33890 -120 33910 -60
rect 33800 -140 33910 -120
rect 33970 -60 34080 -40
rect 33970 -120 33990 -60
rect 34060 -120 34080 -60
rect 33970 -140 34080 -120
rect 34140 -60 34250 -40
rect 34140 -120 34160 -60
rect 34230 -120 34250 -60
rect 34140 -140 34250 -120
rect 34310 -60 34420 -40
rect 34310 -120 34330 -60
rect 34400 -120 34420 -60
rect 34310 -140 34420 -120
rect 34480 -60 34590 -40
rect 34480 -120 34500 -60
rect 34570 -120 34590 -60
rect 34480 -140 34590 -120
rect 34650 -60 34760 -40
rect 34650 -120 34670 -60
rect 34740 -120 34760 -60
rect 34650 -140 34760 -120
rect 34820 -60 34930 -40
rect 34820 -120 34840 -60
rect 34910 -120 34930 -60
rect 34820 -140 34930 -120
rect 34990 -60 35100 -40
rect 34990 -120 35010 -60
rect 35080 -120 35100 -60
rect 34990 -140 35100 -120
rect 35160 -60 35270 -40
rect 35160 -120 35180 -60
rect 35250 -120 35270 -60
rect 35160 -140 35270 -120
rect 35330 -60 35440 -40
rect 35330 -120 35350 -60
rect 35420 -120 35440 -60
rect 35330 -140 35440 -120
rect 35500 -60 35610 -40
rect 35500 -120 35520 -60
rect 35590 -120 35610 -60
rect 35500 -140 35610 -120
rect 35670 -60 35780 -40
rect 35670 -120 35690 -60
rect 35760 -120 35780 -60
rect 35670 -140 35780 -120
rect 35840 -60 35950 -40
rect 35840 -120 35860 -60
rect 35930 -120 35950 -60
rect 35840 -140 35950 -120
rect 36010 -60 36120 -40
rect 36010 -120 36030 -60
rect 36100 -120 36120 -60
rect 36010 -140 36120 -120
rect 36180 -60 36290 -40
rect 36180 -120 36200 -60
rect 36270 -120 36290 -60
rect 36180 -140 36290 -120
rect 36350 -60 36460 -40
rect 36350 -120 36370 -60
rect 36440 -120 36460 -60
rect 36350 -140 36460 -120
rect 36520 -60 36630 -40
rect 36520 -120 36540 -60
rect 36610 -120 36630 -60
rect 36520 -140 36630 -120
rect 36690 -60 36800 -40
rect 36690 -120 36710 -60
rect 36780 -120 36800 -60
rect 36690 -140 36800 -120
rect 36860 -60 36970 -40
rect 36860 -120 36880 -60
rect 36950 -120 36970 -60
rect 36860 -140 36970 -120
rect 37030 -60 37140 -40
rect 37030 -120 37050 -60
rect 37120 -120 37140 -60
rect 37030 -140 37140 -120
rect 37200 -60 37310 -40
rect 37200 -120 37220 -60
rect 37290 -120 37310 -60
rect 37200 -140 37310 -120
rect 37370 -60 37480 -40
rect 37370 -120 37390 -60
rect 37460 -120 37480 -60
rect 37370 -140 37480 -120
rect 37540 -60 37650 -40
rect 37540 -120 37560 -60
rect 37630 -120 37650 -60
rect 37540 -140 37650 -120
rect 37710 -60 37820 -40
rect 37710 -120 37730 -60
rect 37800 -120 37820 -60
rect 37710 -140 37820 -120
rect 37880 -60 37990 -40
rect 37880 -120 37900 -60
rect 37970 -120 37990 -60
rect 37880 -140 37990 -120
rect 38050 -60 38160 -40
rect 38050 -120 38070 -60
rect 38140 -120 38160 -60
rect 38050 -140 38160 -120
rect 38220 -60 38330 -40
rect 38220 -120 38240 -60
rect 38310 -120 38330 -60
rect 38220 -140 38330 -120
rect 38390 -60 38500 -40
rect 38390 -120 38410 -60
rect 38480 -120 38500 -60
rect 38390 -140 38500 -120
rect 38560 -60 38670 -40
rect 38560 -120 38580 -60
rect 38650 -120 38670 -60
rect 38560 -140 38670 -120
rect 38730 -60 38840 -40
rect 38730 -120 38750 -60
rect 38820 -120 38840 -60
rect 38730 -140 38840 -120
rect 38900 -60 39010 -40
rect 38900 -120 38920 -60
rect 38990 -120 39010 -60
rect 38900 -140 39010 -120
rect 39070 -60 39180 -40
rect 39070 -120 39090 -60
rect 39160 -120 39180 -60
rect 39070 -140 39180 -120
rect 39240 -60 39350 -40
rect 39240 -120 39260 -60
rect 39330 -120 39350 -60
rect 39240 -140 39350 -120
rect 39410 -60 39520 -40
rect 39410 -120 39430 -60
rect 39500 -120 39520 -60
rect 39410 -140 39520 -120
rect 39580 -60 39690 -40
rect 39580 -120 39600 -60
rect 39670 -120 39690 -60
rect 39580 -140 39690 -120
rect 39750 -60 39860 -40
rect 39750 -120 39770 -60
rect 39840 -120 39860 -60
rect 39750 -140 39860 -120
rect 39920 -60 40030 -40
rect 39920 -120 39940 -60
rect 40010 -120 40030 -60
rect 39920 -140 40030 -120
rect 40090 -60 40200 -40
rect 40090 -120 40110 -60
rect 40180 -120 40200 -60
rect 40090 -140 40200 -120
rect 40260 -60 40370 -40
rect 40260 -120 40280 -60
rect 40350 -120 40370 -60
rect 40260 -140 40370 -120
rect 40430 -60 40540 -40
rect 40430 -120 40450 -60
rect 40520 -120 40540 -60
rect 40430 -140 40540 -120
rect 40600 -60 40710 -40
rect 40600 -120 40620 -60
rect 40690 -120 40710 -60
rect 40600 -140 40710 -120
rect 40770 -60 40880 -40
rect 40770 -120 40790 -60
rect 40860 -120 40880 -60
rect 40770 -140 40880 -120
rect 40940 -60 41050 -40
rect 40940 -120 40960 -60
rect 41030 -120 41050 -60
rect 40940 -140 41050 -120
rect 41110 -60 41220 -40
rect 41110 -120 41130 -60
rect 41200 -120 41220 -60
rect 41110 -140 41220 -120
rect 41280 -60 41390 -40
rect 41280 -120 41300 -60
rect 41370 -120 41390 -60
rect 41280 -140 41390 -120
rect 41450 -60 41560 -40
rect 41450 -120 41470 -60
rect 41540 -120 41560 -60
rect 41450 -140 41560 -120
rect 41620 -60 41730 -40
rect 41620 -120 41640 -60
rect 41710 -120 41730 -60
rect 41620 -140 41730 -120
rect 41790 -60 41900 -40
rect 41790 -120 41810 -60
rect 41880 -120 41900 -60
rect 41790 -140 41900 -120
rect 41960 -60 42070 -40
rect 41960 -120 41980 -60
rect 42050 -120 42070 -60
rect 41960 -140 42070 -120
rect 42130 -60 42240 -40
rect 42130 -120 42150 -60
rect 42220 -120 42240 -60
rect 42130 -140 42240 -120
rect 42300 -60 42410 -40
rect 42300 -120 42320 -60
rect 42390 -120 42410 -60
rect 42300 -140 42410 -120
rect 42470 -60 42580 -40
rect 42470 -120 42490 -60
rect 42560 -120 42580 -60
rect 42470 -140 42580 -120
rect 42640 -60 42750 -40
rect 42640 -120 42660 -60
rect 42730 -120 42750 -60
rect 42640 -140 42750 -120
rect 42810 -60 42920 -40
rect 42810 -120 42830 -60
rect 42900 -120 42920 -60
rect 42810 -140 42920 -120
rect 42980 -60 43090 -40
rect 42980 -120 43000 -60
rect 43070 -120 43090 -60
rect 42980 -140 43090 -120
rect 43150 -60 43260 -40
rect 43150 -120 43170 -60
rect 43240 -120 43260 -60
rect 43150 -140 43260 -120
rect 43320 -60 43430 -40
rect 43320 -120 43340 -60
rect 43410 -120 43430 -60
rect 43320 -140 43430 -120
rect 43490 -60 43600 -40
rect 43490 -120 43510 -60
rect 43580 -120 43600 -60
rect 43490 -140 43600 -120
rect 43660 -60 43770 -40
rect 43660 -120 43680 -60
rect 43750 -120 43770 -60
rect 43660 -140 43770 -120
rect 43830 -60 43940 -40
rect 43830 -120 43850 -60
rect 43920 -120 43940 -60
rect 43830 -140 43940 -120
rect 44000 -60 44110 -40
rect 44000 -120 44020 -60
rect 44090 -120 44110 -60
rect 44000 -140 44110 -120
rect 44170 -60 44280 -40
rect 44170 -120 44190 -60
rect 44260 -120 44280 -60
rect 44170 -140 44280 -120
rect 44340 -60 44450 -40
rect 44340 -120 44360 -60
rect 44430 -120 44450 -60
rect 44340 -140 44450 -120
rect 44510 -60 44620 -40
rect 44510 -120 44530 -60
rect 44600 -120 44620 -60
rect 44510 -140 44620 -120
rect 44680 -60 44790 -40
rect 44680 -120 44700 -60
rect 44770 -120 44790 -60
rect 44680 -140 44790 -120
rect 44850 -60 44960 -40
rect 44850 -120 44870 -60
rect 44940 -120 44960 -60
rect 44850 -140 44960 -120
rect 45020 -60 45130 -40
rect 45020 -120 45040 -60
rect 45110 -120 45130 -60
rect 45020 -140 45130 -120
rect 45190 -60 45300 -40
rect 45190 -120 45210 -60
rect 45280 -120 45300 -60
rect 45190 -140 45300 -120
rect 45360 -60 45470 -40
rect 45360 -120 45380 -60
rect 45450 -120 45470 -60
rect 45360 -140 45470 -120
rect 45530 -60 45640 -40
rect 45530 -120 45550 -60
rect 45620 -120 45640 -60
rect 45530 -140 45640 -120
rect 45700 -60 45810 -40
rect 45700 -120 45720 -60
rect 45790 -120 45810 -60
rect 45700 -140 45810 -120
rect 45870 -60 45980 -40
rect 45870 -120 45890 -60
rect 45960 -120 45980 -60
rect 45870 -140 45980 -120
rect 46040 -60 46150 -40
rect 46040 -120 46060 -60
rect 46130 -120 46150 -60
rect 46040 -140 46150 -120
rect 46210 -60 46320 -40
rect 46210 -120 46230 -60
rect 46300 -120 46320 -60
rect 46210 -140 46320 -120
rect 46380 -60 46490 -40
rect 46380 -120 46400 -60
rect 46470 -120 46490 -60
rect 46380 -140 46490 -120
rect 46550 -60 46660 -40
rect 46550 -120 46570 -60
rect 46640 -120 46660 -60
rect 46550 -140 46660 -120
rect 46720 -60 46830 -40
rect 46720 -120 46740 -60
rect 46810 -120 46830 -60
rect 46720 -140 46830 -120
rect 46890 -60 47000 -40
rect 46890 -120 46910 -60
rect 46980 -120 47000 -60
rect 46890 -140 47000 -120
rect 47060 -60 47170 -40
rect 47060 -120 47080 -60
rect 47150 -120 47170 -60
rect 47060 -140 47170 -120
rect 47230 -60 47340 -40
rect 47230 -120 47250 -60
rect 47320 -120 47340 -60
rect 47230 -140 47340 -120
rect 47400 -60 47510 -40
rect 47400 -120 47420 -60
rect 47490 -120 47510 -60
rect 47400 -140 47510 -120
rect 47570 -60 47680 -40
rect 47570 -120 47590 -60
rect 47660 -120 47680 -60
rect 47570 -140 47680 -120
rect 47740 -60 47850 -40
rect 47740 -120 47760 -60
rect 47830 -120 47850 -60
rect 47740 -140 47850 -120
rect 47910 -60 48020 -40
rect 47910 -120 47930 -60
rect 48000 -120 48020 -60
rect 47910 -140 48020 -120
rect 48080 -60 48190 -40
rect 48080 -120 48100 -60
rect 48170 -120 48190 -60
rect 48080 -140 48190 -120
rect 48250 -60 48360 -40
rect 48250 -120 48270 -60
rect 48340 -120 48360 -60
rect 48250 -140 48360 -120
rect 48420 -60 48530 -40
rect 48420 -120 48440 -60
rect 48510 -120 48530 -60
rect 48420 -140 48530 -120
rect 48590 -60 48700 -40
rect 48590 -120 48610 -60
rect 48680 -120 48700 -60
rect 48590 -140 48700 -120
rect 48760 -60 48870 -40
rect 48760 -120 48780 -60
rect 48850 -120 48870 -60
rect 48760 -140 48870 -120
rect 48930 -60 49040 -40
rect 48930 -120 48950 -60
rect 49020 -120 49040 -60
rect 48930 -140 49040 -120
rect 49100 -60 49210 -40
rect 49100 -120 49120 -60
rect 49190 -120 49210 -60
rect 49100 -140 49210 -120
rect 49270 -60 49380 -40
rect 49270 -120 49290 -60
rect 49360 -120 49380 -60
rect 49270 -140 49380 -120
rect 49440 -60 49550 -40
rect 49440 -120 49460 -60
rect 49530 -120 49550 -60
rect 49440 -140 49550 -120
rect 49610 -60 49720 -40
rect 49610 -120 49630 -60
rect 49700 -120 49720 -60
rect 49610 -140 49720 -120
rect 49780 -60 49890 -40
rect 49780 -120 49800 -60
rect 49870 -120 49890 -60
rect 49780 -140 49890 -120
rect 49950 -60 50060 -40
rect 49950 -120 49970 -60
rect 50040 -120 50060 -60
rect 49950 -140 50060 -120
rect 50120 -60 50230 -40
rect 50120 -120 50140 -60
rect 50210 -120 50230 -60
rect 50120 -140 50230 -120
rect 50290 -60 50400 -40
rect 50290 -120 50310 -60
rect 50380 -120 50400 -60
rect 50290 -140 50400 -120
rect 50460 -60 50570 -40
rect 50460 -120 50480 -60
rect 50550 -120 50570 -60
rect 50460 -140 50570 -120
rect 50630 -60 50740 -40
rect 50630 -120 50650 -60
rect 50720 -120 50740 -60
rect 50630 -140 50740 -120
rect 50800 -60 50910 -40
rect 50800 -120 50820 -60
rect 50890 -120 50910 -60
rect 50800 -140 50910 -120
rect 50970 -60 51080 -40
rect 50970 -120 50990 -60
rect 51060 -120 51080 -60
rect 50970 -140 51080 -120
rect 51140 -60 51250 -40
rect 51140 -120 51160 -60
rect 51230 -120 51250 -60
rect 51140 -140 51250 -120
rect 51310 -60 51420 -40
rect 51310 -120 51330 -60
rect 51400 -120 51420 -60
rect 51310 -140 51420 -120
rect 51480 -60 51590 -40
rect 51480 -120 51500 -60
rect 51570 -120 51590 -60
rect 51480 -140 51590 -120
rect 51650 -60 51760 -40
rect 51650 -120 51670 -60
rect 51740 -120 51760 -60
rect 51650 -140 51760 -120
rect 51820 -60 51930 -40
rect 51820 -120 51840 -60
rect 51910 -120 51930 -60
rect 51820 -140 51930 -120
rect 51990 -60 52100 -40
rect 51990 -120 52010 -60
rect 52080 -120 52100 -60
rect 51990 -140 52100 -120
rect 52160 -60 52270 -40
rect 52160 -120 52180 -60
rect 52250 -120 52270 -60
rect 52160 -140 52270 -120
rect 52330 -60 52440 -40
rect 52330 -120 52350 -60
rect 52420 -120 52440 -60
rect 52330 -140 52440 -120
rect 52500 -60 52610 -40
rect 52500 -120 52520 -60
rect 52590 -120 52610 -60
rect 52500 -140 52610 -120
rect 52670 -60 52780 -40
rect 52670 -120 52690 -60
rect 52760 -120 52780 -60
rect 52670 -140 52780 -120
rect 52840 -60 52950 -40
rect 52840 -120 52860 -60
rect 52930 -120 52950 -60
rect 52840 -140 52950 -120
rect 53010 -60 53120 -40
rect 53010 -120 53030 -60
rect 53100 -120 53120 -60
rect 53010 -140 53120 -120
rect 53180 -60 53290 -40
rect 53180 -120 53200 -60
rect 53270 -120 53290 -60
rect 53180 -140 53290 -120
rect 53350 -60 53460 -40
rect 53350 -120 53370 -60
rect 53440 -120 53460 -60
rect 53350 -140 53460 -120
rect 53520 -60 53630 -40
rect 53520 -120 53540 -60
rect 53610 -120 53630 -60
rect 53520 -140 53630 -120
rect 53690 -60 53800 -40
rect 53690 -120 53710 -60
rect 53780 -120 53800 -60
rect 53690 -140 53800 -120
rect 53860 -60 53970 -40
rect 53860 -120 53880 -60
rect 53950 -120 53970 -60
rect 53860 -140 53970 -120
rect 54030 -60 54140 -40
rect 54030 -120 54050 -60
rect 54120 -120 54140 -60
rect 54030 -140 54140 -120
rect 54200 -60 54310 -40
rect 54200 -120 54220 -60
rect 54290 -120 54310 -60
rect 54200 -140 54310 -120
rect 54370 -60 54480 -40
rect 54370 -120 54390 -60
rect 54460 -120 54480 -60
rect 54370 -140 54480 -120
rect 54540 -60 54650 -40
rect 54540 -120 54560 -60
rect 54630 -120 54650 -60
rect 54540 -140 54650 -120
rect 54710 -60 54820 -40
rect 54710 -120 54730 -60
rect 54800 -120 54820 -60
rect 54710 -140 54820 -120
rect 54880 -60 54990 -40
rect 54880 -120 54900 -60
rect 54970 -120 54990 -60
rect 54880 -140 54990 -120
rect 55050 -60 55160 -40
rect 55050 -120 55070 -60
rect 55140 -120 55160 -60
rect 55050 -140 55160 -120
rect 55220 -60 55330 -40
rect 55220 -120 55240 -60
rect 55310 -120 55330 -60
rect 55220 -140 55330 -120
rect 55390 -60 55500 -40
rect 55390 -120 55410 -60
rect 55480 -120 55500 -60
rect 55390 -140 55500 -120
rect 55560 -60 55670 -40
rect 55560 -120 55580 -60
rect 55650 -120 55670 -60
rect 55560 -140 55670 -120
rect 55730 -60 55840 -40
rect 55730 -120 55750 -60
rect 55820 -120 55840 -60
rect 55730 -140 55840 -120
rect 55900 -60 56010 -40
rect 55900 -120 55920 -60
rect 55990 -120 56010 -60
rect 55900 -140 56010 -120
rect 56070 -60 56180 -40
rect 56070 -120 56090 -60
rect 56160 -120 56180 -60
rect 56070 -140 56180 -120
rect 56240 -60 56350 -40
rect 56240 -120 56260 -60
rect 56330 -120 56350 -60
rect 56240 -140 56350 -120
rect 56410 -60 56520 -40
rect 56410 -120 56430 -60
rect 56500 -120 56520 -60
rect 56410 -140 56520 -120
rect 56580 -60 56690 -40
rect 56580 -120 56600 -60
rect 56670 -120 56690 -60
rect 56580 -140 56690 -120
rect 56750 -60 56860 -40
rect 56750 -120 56770 -60
rect 56840 -120 56860 -60
rect 56750 -140 56860 -120
rect 56920 -60 57030 -40
rect 56920 -120 56940 -60
rect 57010 -120 57030 -60
rect 56920 -140 57030 -120
rect 57090 -60 57200 -40
rect 57090 -120 57110 -60
rect 57180 -120 57200 -60
rect 57090 -140 57200 -120
rect 57260 -60 57370 -40
rect 57260 -120 57280 -60
rect 57350 -120 57370 -60
rect 57260 -140 57370 -120
rect 57430 -60 57540 -40
rect 57430 -120 57450 -60
rect 57520 -120 57540 -60
rect 57430 -140 57540 -120
rect 57600 -60 57710 -40
rect 57600 -120 57620 -60
rect 57690 -120 57710 -60
rect 57600 -140 57710 -120
rect 57770 -60 57880 -40
rect 57770 -120 57790 -60
rect 57860 -120 57880 -60
rect 57770 -140 57880 -120
rect 57940 -60 58050 -40
rect 57940 -120 57960 -60
rect 58030 -120 58050 -60
rect 57940 -140 58050 -120
rect 58110 -60 58220 -40
rect 58110 -120 58130 -60
rect 58200 -120 58220 -60
rect 58110 -140 58220 -120
rect 58280 -60 58390 -40
rect 58280 -120 58300 -60
rect 58370 -120 58390 -60
rect 58280 -140 58390 -120
rect 58450 -60 58560 -40
rect 58450 -120 58470 -60
rect 58540 -120 58560 -60
rect 58450 -140 58560 -120
rect 58620 -60 58730 -40
rect 58620 -120 58640 -60
rect 58710 -120 58730 -60
rect 58620 -140 58730 -120
rect 58790 -60 58900 -40
rect 58790 -120 58810 -60
rect 58880 -120 58900 -60
rect 58790 -140 58900 -120
rect 58960 -60 59070 -40
rect 58960 -120 58980 -60
rect 59050 -120 59070 -60
rect 58960 -140 59070 -120
rect 59130 -60 59240 -40
rect 59130 -120 59150 -60
rect 59220 -120 59240 -60
rect 59130 -140 59240 -120
rect 130 -170 160 -140
rect 210 -530 320 -510
rect 210 -590 230 -530
rect 300 -590 320 -530
rect 210 -610 320 -590
rect 380 -530 490 -510
rect 380 -590 400 -530
rect 470 -590 490 -530
rect 380 -610 490 -590
rect 550 -530 660 -510
rect 550 -590 570 -530
rect 640 -590 660 -530
rect 550 -610 660 -590
rect 720 -530 830 -510
rect 720 -590 740 -530
rect 810 -590 830 -530
rect 720 -610 830 -590
rect 890 -530 1000 -510
rect 890 -590 910 -530
rect 980 -590 1000 -530
rect 890 -610 1000 -590
rect 1060 -530 1170 -510
rect 1060 -590 1080 -530
rect 1150 -590 1170 -530
rect 1060 -610 1170 -590
rect 1230 -530 1340 -510
rect 1230 -590 1250 -530
rect 1320 -590 1340 -530
rect 1230 -610 1340 -590
rect 1400 -530 1510 -510
rect 1400 -590 1420 -530
rect 1490 -590 1510 -530
rect 1400 -610 1510 -590
rect 1570 -530 1680 -510
rect 1570 -590 1590 -530
rect 1660 -590 1680 -530
rect 1570 -610 1680 -590
rect 1740 -530 1850 -510
rect 1740 -590 1760 -530
rect 1830 -590 1850 -530
rect 1740 -610 1850 -590
rect 1910 -530 2020 -510
rect 1910 -590 1930 -530
rect 2000 -590 2020 -530
rect 1910 -610 2020 -590
rect 2080 -530 2190 -510
rect 2080 -590 2100 -530
rect 2170 -590 2190 -530
rect 2080 -610 2190 -590
rect 2250 -530 2360 -510
rect 2250 -590 2270 -530
rect 2340 -590 2360 -530
rect 2250 -610 2360 -590
rect 2420 -530 2530 -510
rect 2420 -590 2440 -530
rect 2510 -590 2530 -530
rect 2420 -610 2530 -590
rect 2590 -530 2700 -510
rect 2590 -590 2610 -530
rect 2680 -590 2700 -530
rect 2590 -610 2700 -590
rect 2760 -530 2870 -510
rect 2760 -590 2780 -530
rect 2850 -590 2870 -530
rect 2760 -610 2870 -590
rect 2930 -530 3040 -510
rect 2930 -590 2950 -530
rect 3020 -590 3040 -530
rect 2930 -610 3040 -590
rect 3100 -530 3210 -510
rect 3100 -590 3120 -530
rect 3190 -590 3210 -530
rect 3100 -610 3210 -590
rect 3270 -530 3380 -510
rect 3270 -590 3290 -530
rect 3360 -590 3380 -530
rect 3270 -610 3380 -590
rect 3440 -530 3550 -510
rect 3440 -590 3460 -530
rect 3530 -590 3550 -530
rect 3440 -610 3550 -590
rect 3610 -530 3720 -510
rect 3610 -590 3630 -530
rect 3700 -590 3720 -530
rect 3610 -610 3720 -590
rect 3780 -530 3890 -510
rect 3780 -590 3800 -530
rect 3870 -590 3890 -530
rect 3780 -610 3890 -590
rect 3950 -530 4060 -510
rect 3950 -590 3970 -530
rect 4040 -590 4060 -530
rect 3950 -610 4060 -590
rect 4120 -530 4230 -510
rect 4120 -590 4140 -530
rect 4210 -590 4230 -530
rect 4120 -610 4230 -590
rect 4290 -530 4400 -510
rect 4290 -590 4310 -530
rect 4380 -590 4400 -530
rect 4290 -610 4400 -590
rect 4460 -530 4570 -510
rect 4460 -590 4480 -530
rect 4550 -590 4570 -530
rect 4460 -610 4570 -590
rect 4630 -530 4740 -510
rect 4630 -590 4650 -530
rect 4720 -590 4740 -530
rect 4630 -610 4740 -590
rect 4800 -530 4910 -510
rect 4800 -590 4820 -530
rect 4890 -590 4910 -530
rect 4800 -610 4910 -590
rect 4970 -530 5080 -510
rect 4970 -590 4990 -530
rect 5060 -590 5080 -530
rect 4970 -610 5080 -590
rect 5140 -530 5250 -510
rect 5140 -590 5160 -530
rect 5230 -590 5250 -530
rect 5140 -610 5250 -590
rect 5310 -530 5420 -510
rect 5310 -590 5330 -530
rect 5400 -590 5420 -530
rect 5310 -610 5420 -590
rect 5480 -530 5590 -510
rect 5480 -590 5500 -530
rect 5570 -590 5590 -530
rect 5480 -610 5590 -590
rect 5650 -530 5760 -510
rect 5650 -590 5670 -530
rect 5740 -590 5760 -530
rect 5650 -610 5760 -590
rect 5820 -530 5930 -510
rect 5820 -590 5840 -530
rect 5910 -590 5930 -530
rect 5820 -610 5930 -590
rect 5990 -530 6100 -510
rect 5990 -590 6010 -530
rect 6080 -590 6100 -530
rect 5990 -610 6100 -590
rect 6160 -530 6270 -510
rect 6160 -590 6180 -530
rect 6250 -590 6270 -530
rect 6160 -610 6270 -590
rect 6330 -530 6440 -510
rect 6330 -590 6350 -530
rect 6420 -590 6440 -530
rect 6330 -610 6440 -590
rect 6500 -530 6610 -510
rect 6500 -590 6520 -530
rect 6590 -590 6610 -530
rect 6500 -610 6610 -590
rect 6670 -530 6780 -510
rect 6670 -590 6690 -530
rect 6760 -590 6780 -530
rect 6670 -610 6780 -590
rect 6840 -530 6950 -510
rect 6840 -590 6860 -530
rect 6930 -590 6950 -530
rect 6840 -610 6950 -590
rect 7010 -530 7120 -510
rect 7010 -590 7030 -530
rect 7100 -590 7120 -530
rect 7010 -610 7120 -590
rect 7180 -530 7290 -510
rect 7180 -590 7200 -530
rect 7270 -590 7290 -530
rect 7180 -610 7290 -590
rect 7350 -530 7460 -510
rect 7350 -590 7370 -530
rect 7440 -590 7460 -530
rect 7350 -610 7460 -590
rect 7520 -530 7630 -510
rect 7520 -590 7540 -530
rect 7610 -590 7630 -530
rect 7520 -610 7630 -590
rect 7690 -530 7800 -510
rect 7690 -590 7710 -530
rect 7780 -590 7800 -530
rect 7690 -610 7800 -590
rect 7860 -530 7970 -510
rect 7860 -590 7880 -530
rect 7950 -590 7970 -530
rect 7860 -610 7970 -590
rect 8030 -530 8140 -510
rect 8030 -590 8050 -530
rect 8120 -590 8140 -530
rect 8030 -610 8140 -590
rect 8200 -530 8310 -510
rect 8200 -590 8220 -530
rect 8290 -590 8310 -530
rect 8200 -610 8310 -590
rect 8370 -530 8480 -510
rect 8370 -590 8390 -530
rect 8460 -590 8480 -530
rect 8370 -610 8480 -590
rect 8540 -530 8650 -510
rect 8540 -590 8560 -530
rect 8630 -590 8650 -530
rect 8540 -610 8650 -590
rect 8710 -530 8820 -510
rect 8710 -590 8730 -530
rect 8800 -590 8820 -530
rect 8710 -610 8820 -590
rect 8880 -530 8990 -510
rect 8880 -590 8900 -530
rect 8970 -590 8990 -530
rect 8880 -610 8990 -590
rect 9050 -530 9160 -510
rect 9050 -590 9070 -530
rect 9140 -590 9160 -530
rect 9050 -610 9160 -590
rect 9220 -530 9330 -510
rect 9220 -590 9240 -530
rect 9310 -590 9330 -530
rect 9220 -610 9330 -590
rect 9390 -530 9500 -510
rect 9390 -590 9410 -530
rect 9480 -590 9500 -530
rect 9390 -610 9500 -590
rect 9560 -530 9670 -510
rect 9560 -590 9580 -530
rect 9650 -590 9670 -530
rect 9560 -610 9670 -590
rect 9730 -530 9840 -510
rect 9730 -590 9750 -530
rect 9820 -590 9840 -530
rect 9730 -610 9840 -590
rect 9900 -530 10010 -510
rect 9900 -590 9920 -530
rect 9990 -590 10010 -530
rect 9900 -610 10010 -590
rect 10070 -530 10180 -510
rect 10070 -590 10090 -530
rect 10160 -590 10180 -530
rect 10070 -610 10180 -590
rect 10240 -530 10350 -510
rect 10240 -590 10260 -530
rect 10330 -590 10350 -530
rect 10240 -610 10350 -590
rect 10410 -530 10520 -510
rect 10410 -590 10430 -530
rect 10500 -590 10520 -530
rect 10410 -610 10520 -590
rect 10580 -530 10690 -510
rect 10580 -590 10600 -530
rect 10670 -590 10690 -530
rect 10580 -610 10690 -590
rect 10750 -530 10860 -510
rect 10750 -590 10770 -530
rect 10840 -590 10860 -530
rect 10750 -610 10860 -590
rect 10920 -530 11030 -510
rect 10920 -590 10940 -530
rect 11010 -590 11030 -530
rect 10920 -610 11030 -590
rect 11090 -530 11200 -510
rect 11090 -590 11110 -530
rect 11180 -590 11200 -530
rect 11090 -610 11200 -590
rect 11260 -530 11370 -510
rect 11260 -590 11280 -530
rect 11350 -590 11370 -530
rect 11260 -610 11370 -590
rect 11430 -530 11540 -510
rect 11430 -590 11450 -530
rect 11520 -590 11540 -530
rect 11430 -610 11540 -590
rect 11600 -530 11710 -510
rect 11600 -590 11620 -530
rect 11690 -590 11710 -530
rect 11600 -610 11710 -590
rect 11770 -530 11880 -510
rect 11770 -590 11790 -530
rect 11860 -590 11880 -530
rect 11770 -610 11880 -590
rect 11940 -530 12050 -510
rect 11940 -590 11960 -530
rect 12030 -590 12050 -530
rect 11940 -610 12050 -590
rect 12110 -530 12220 -510
rect 12110 -590 12130 -530
rect 12200 -590 12220 -530
rect 12110 -610 12220 -590
rect 12280 -530 12390 -510
rect 12280 -590 12300 -530
rect 12370 -590 12390 -530
rect 12280 -610 12390 -590
rect 12450 -530 12560 -510
rect 12450 -590 12470 -530
rect 12540 -590 12560 -530
rect 12450 -610 12560 -590
rect 12620 -530 12730 -510
rect 12620 -590 12640 -530
rect 12710 -590 12730 -530
rect 12620 -610 12730 -590
rect 12790 -530 12900 -510
rect 12790 -590 12810 -530
rect 12880 -590 12900 -530
rect 12790 -610 12900 -590
rect 12960 -530 13070 -510
rect 12960 -590 12980 -530
rect 13050 -590 13070 -530
rect 12960 -610 13070 -590
rect 13130 -530 13240 -510
rect 13130 -590 13150 -530
rect 13220 -590 13240 -530
rect 13130 -610 13240 -590
rect 13300 -530 13410 -510
rect 13300 -590 13320 -530
rect 13390 -590 13410 -530
rect 13300 -610 13410 -590
rect 13470 -530 13580 -510
rect 13470 -590 13490 -530
rect 13560 -590 13580 -530
rect 13470 -610 13580 -590
rect 13640 -530 13750 -510
rect 13640 -590 13660 -530
rect 13730 -590 13750 -530
rect 13640 -610 13750 -590
rect 13810 -530 13920 -510
rect 13810 -590 13830 -530
rect 13900 -590 13920 -530
rect 13810 -610 13920 -590
rect 13980 -530 14090 -510
rect 13980 -590 14000 -530
rect 14070 -590 14090 -530
rect 13980 -610 14090 -590
rect 14150 -530 14260 -510
rect 14150 -590 14170 -530
rect 14240 -590 14260 -530
rect 14150 -610 14260 -590
rect 14320 -530 14430 -510
rect 14320 -590 14340 -530
rect 14410 -590 14430 -530
rect 14320 -610 14430 -590
rect 14490 -530 14600 -510
rect 14490 -590 14510 -530
rect 14580 -590 14600 -530
rect 14490 -610 14600 -590
rect 14660 -530 14770 -510
rect 14660 -590 14680 -530
rect 14750 -590 14770 -530
rect 14660 -610 14770 -590
rect 14830 -530 14940 -510
rect 14830 -590 14850 -530
rect 14920 -590 14940 -530
rect 14830 -610 14940 -590
rect 15000 -530 15110 -510
rect 15000 -590 15020 -530
rect 15090 -590 15110 -530
rect 15000 -610 15110 -590
rect 15170 -530 15280 -510
rect 15170 -590 15190 -530
rect 15260 -590 15280 -530
rect 15170 -610 15280 -590
rect 15340 -530 15450 -510
rect 15340 -590 15360 -530
rect 15430 -590 15450 -530
rect 15340 -610 15450 -590
rect 15510 -530 15620 -510
rect 15510 -590 15530 -530
rect 15600 -590 15620 -530
rect 15510 -610 15620 -590
rect 15680 -530 15790 -510
rect 15680 -590 15700 -530
rect 15770 -590 15790 -530
rect 15680 -610 15790 -590
rect 15850 -530 15960 -510
rect 15850 -590 15870 -530
rect 15940 -590 15960 -530
rect 15850 -610 15960 -590
rect 16020 -530 16130 -510
rect 16020 -590 16040 -530
rect 16110 -590 16130 -530
rect 16020 -610 16130 -590
rect 16190 -530 16300 -510
rect 16190 -590 16210 -530
rect 16280 -590 16300 -530
rect 16190 -610 16300 -590
rect 16360 -530 16470 -510
rect 16360 -590 16380 -530
rect 16450 -590 16470 -530
rect 16360 -610 16470 -590
rect 16530 -530 16640 -510
rect 16530 -590 16550 -530
rect 16620 -590 16640 -530
rect 16530 -610 16640 -590
rect 16700 -530 16810 -510
rect 16700 -590 16720 -530
rect 16790 -590 16810 -530
rect 16700 -610 16810 -590
rect 16870 -530 16980 -510
rect 16870 -590 16890 -530
rect 16960 -590 16980 -530
rect 16870 -610 16980 -590
rect 17040 -530 17150 -510
rect 17040 -590 17060 -530
rect 17130 -590 17150 -530
rect 17040 -610 17150 -590
rect 17210 -530 17320 -510
rect 17210 -590 17230 -530
rect 17300 -590 17320 -530
rect 17210 -610 17320 -590
rect 17380 -530 17490 -510
rect 17380 -590 17400 -530
rect 17470 -590 17490 -530
rect 17380 -610 17490 -590
rect 17550 -530 17660 -510
rect 17550 -590 17570 -530
rect 17640 -590 17660 -530
rect 17550 -610 17660 -590
rect 17720 -530 17830 -510
rect 17720 -590 17740 -530
rect 17810 -590 17830 -530
rect 17720 -610 17830 -590
rect 17890 -530 18000 -510
rect 17890 -590 17910 -530
rect 17980 -590 18000 -530
rect 17890 -610 18000 -590
rect 18060 -530 18170 -510
rect 18060 -590 18080 -530
rect 18150 -590 18170 -530
rect 18060 -610 18170 -590
rect 18230 -530 18340 -510
rect 18230 -590 18250 -530
rect 18320 -590 18340 -530
rect 18230 -610 18340 -590
rect 18400 -530 18510 -510
rect 18400 -590 18420 -530
rect 18490 -590 18510 -530
rect 18400 -610 18510 -590
rect 18570 -530 18680 -510
rect 18570 -590 18590 -530
rect 18660 -590 18680 -530
rect 18570 -610 18680 -590
rect 18740 -530 18850 -510
rect 18740 -590 18760 -530
rect 18830 -590 18850 -530
rect 18740 -610 18850 -590
rect 18910 -530 19020 -510
rect 18910 -590 18930 -530
rect 19000 -590 19020 -530
rect 18910 -610 19020 -590
rect 19080 -530 19190 -510
rect 19080 -590 19100 -530
rect 19170 -590 19190 -530
rect 19080 -610 19190 -590
rect 19250 -530 19360 -510
rect 19250 -590 19270 -530
rect 19340 -590 19360 -530
rect 19250 -610 19360 -590
rect 19420 -530 19530 -510
rect 19420 -590 19440 -530
rect 19510 -590 19530 -530
rect 19420 -610 19530 -590
rect 19590 -530 19700 -510
rect 19590 -590 19610 -530
rect 19680 -590 19700 -530
rect 19590 -610 19700 -590
rect 19760 -530 19870 -510
rect 19760 -590 19780 -530
rect 19850 -590 19870 -530
rect 19760 -610 19870 -590
rect 19930 -530 20040 -510
rect 19930 -590 19950 -530
rect 20020 -590 20040 -530
rect 19930 -610 20040 -590
rect 20100 -530 20210 -510
rect 20100 -590 20120 -530
rect 20190 -590 20210 -530
rect 20100 -610 20210 -590
rect 20270 -530 20380 -510
rect 20270 -590 20290 -530
rect 20360 -590 20380 -530
rect 20270 -610 20380 -590
rect 20440 -530 20550 -510
rect 20440 -590 20460 -530
rect 20530 -590 20550 -530
rect 20440 -610 20550 -590
rect 20610 -530 20720 -510
rect 20610 -590 20630 -530
rect 20700 -590 20720 -530
rect 20610 -610 20720 -590
rect 20780 -530 20890 -510
rect 20780 -590 20800 -530
rect 20870 -590 20890 -530
rect 20780 -610 20890 -590
rect 20950 -530 21060 -510
rect 20950 -590 20970 -530
rect 21040 -590 21060 -530
rect 20950 -610 21060 -590
rect 21120 -530 21230 -510
rect 21120 -590 21140 -530
rect 21210 -590 21230 -530
rect 21120 -610 21230 -590
rect 21290 -530 21400 -510
rect 21290 -590 21310 -530
rect 21380 -590 21400 -530
rect 21290 -610 21400 -590
rect 21460 -530 21570 -510
rect 21460 -590 21480 -530
rect 21550 -590 21570 -530
rect 21460 -610 21570 -590
rect 21630 -530 21740 -510
rect 21630 -590 21650 -530
rect 21720 -590 21740 -530
rect 21630 -610 21740 -590
rect 21800 -530 21910 -510
rect 21800 -590 21820 -530
rect 21890 -590 21910 -530
rect 21800 -610 21910 -590
rect 21970 -530 22080 -510
rect 21970 -590 21990 -530
rect 22060 -590 22080 -530
rect 21970 -610 22080 -590
rect 22140 -530 22250 -510
rect 22140 -590 22160 -530
rect 22230 -590 22250 -530
rect 22140 -610 22250 -590
rect 22310 -530 22420 -510
rect 22310 -590 22330 -530
rect 22400 -590 22420 -530
rect 22310 -610 22420 -590
rect 22480 -530 22590 -510
rect 22480 -590 22500 -530
rect 22570 -590 22590 -530
rect 22480 -610 22590 -590
rect 22650 -530 22760 -510
rect 22650 -590 22670 -530
rect 22740 -590 22760 -530
rect 22650 -610 22760 -590
rect 22820 -530 22930 -510
rect 22820 -590 22840 -530
rect 22910 -590 22930 -530
rect 22820 -610 22930 -590
rect 22990 -530 23100 -510
rect 22990 -590 23010 -530
rect 23080 -590 23100 -530
rect 22990 -610 23100 -590
rect 23160 -530 23270 -510
rect 23160 -590 23180 -530
rect 23250 -590 23270 -530
rect 23160 -610 23270 -590
rect 23330 -530 23440 -510
rect 23330 -590 23350 -530
rect 23420 -590 23440 -530
rect 23330 -610 23440 -590
rect 23500 -530 23610 -510
rect 23500 -590 23520 -530
rect 23590 -590 23610 -530
rect 23500 -610 23610 -590
rect 23670 -530 23780 -510
rect 23670 -590 23690 -530
rect 23760 -590 23780 -530
rect 23670 -610 23780 -590
rect 23840 -530 23950 -510
rect 23840 -590 23860 -530
rect 23930 -590 23950 -530
rect 23840 -610 23950 -590
rect 24010 -530 24120 -510
rect 24010 -590 24030 -530
rect 24100 -590 24120 -530
rect 24010 -610 24120 -590
rect 24180 -530 24290 -510
rect 24180 -590 24200 -530
rect 24270 -590 24290 -530
rect 24180 -610 24290 -590
rect 24350 -530 24460 -510
rect 24350 -590 24370 -530
rect 24440 -590 24460 -530
rect 24350 -610 24460 -590
rect 24520 -530 24630 -510
rect 24520 -590 24540 -530
rect 24610 -590 24630 -530
rect 24520 -610 24630 -590
rect 24690 -530 24800 -510
rect 24690 -590 24710 -530
rect 24780 -590 24800 -530
rect 24690 -610 24800 -590
rect 24860 -530 24970 -510
rect 24860 -590 24880 -530
rect 24950 -590 24970 -530
rect 24860 -610 24970 -590
rect 25030 -530 25140 -510
rect 25030 -590 25050 -530
rect 25120 -590 25140 -530
rect 25030 -610 25140 -590
rect 25200 -530 25310 -510
rect 25200 -590 25220 -530
rect 25290 -590 25310 -530
rect 25200 -610 25310 -590
rect 25370 -530 25480 -510
rect 25370 -590 25390 -530
rect 25460 -590 25480 -530
rect 25370 -610 25480 -590
rect 25540 -530 25650 -510
rect 25540 -590 25560 -530
rect 25630 -590 25650 -530
rect 25540 -610 25650 -590
rect 25710 -530 25820 -510
rect 25710 -590 25730 -530
rect 25800 -590 25820 -530
rect 25710 -610 25820 -590
rect 25880 -530 25990 -510
rect 25880 -590 25900 -530
rect 25970 -590 25990 -530
rect 25880 -610 25990 -590
rect 26050 -530 26160 -510
rect 26050 -590 26070 -530
rect 26140 -590 26160 -530
rect 26050 -610 26160 -590
rect 26220 -530 26330 -510
rect 26220 -590 26240 -530
rect 26310 -590 26330 -530
rect 26220 -610 26330 -590
rect 26390 -530 26500 -510
rect 26390 -590 26410 -530
rect 26480 -590 26500 -530
rect 26390 -610 26500 -590
rect 26560 -530 26670 -510
rect 26560 -590 26580 -530
rect 26650 -590 26670 -530
rect 26560 -610 26670 -590
rect 26730 -530 26840 -510
rect 26730 -590 26750 -530
rect 26820 -590 26840 -530
rect 26730 -610 26840 -590
rect 26900 -530 27010 -510
rect 26900 -590 26920 -530
rect 26990 -590 27010 -530
rect 26900 -610 27010 -590
rect 27070 -530 27180 -510
rect 27070 -590 27090 -530
rect 27160 -590 27180 -530
rect 27070 -610 27180 -590
rect 27240 -530 27350 -510
rect 27240 -590 27260 -530
rect 27330 -590 27350 -530
rect 27240 -610 27350 -590
rect 27410 -530 27520 -510
rect 27410 -590 27430 -530
rect 27500 -590 27520 -530
rect 27410 -610 27520 -590
rect 27580 -530 27690 -510
rect 27580 -590 27600 -530
rect 27670 -590 27690 -530
rect 27580 -610 27690 -590
rect 27750 -530 27860 -510
rect 27750 -590 27770 -530
rect 27840 -590 27860 -530
rect 27750 -610 27860 -590
rect 27920 -530 28030 -510
rect 27920 -590 27940 -530
rect 28010 -590 28030 -530
rect 27920 -610 28030 -590
rect 28090 -530 28200 -510
rect 28090 -590 28110 -530
rect 28180 -590 28200 -530
rect 28090 -610 28200 -590
rect 28260 -530 28370 -510
rect 28260 -590 28280 -530
rect 28350 -590 28370 -530
rect 28260 -610 28370 -590
rect 28430 -530 28540 -510
rect 28430 -590 28450 -530
rect 28520 -590 28540 -530
rect 28430 -610 28540 -590
rect 28600 -530 28710 -510
rect 28600 -590 28620 -530
rect 28690 -590 28710 -530
rect 28600 -610 28710 -590
rect 28770 -530 28880 -510
rect 28770 -590 28790 -530
rect 28860 -590 28880 -530
rect 28770 -610 28880 -590
rect 28940 -530 29050 -510
rect 28940 -590 28960 -530
rect 29030 -590 29050 -530
rect 28940 -610 29050 -590
rect 29110 -530 29220 -510
rect 29110 -590 29130 -530
rect 29200 -590 29220 -530
rect 29110 -610 29220 -590
rect 29280 -530 29390 -510
rect 29280 -590 29300 -530
rect 29370 -590 29390 -530
rect 29280 -610 29390 -590
rect 29450 -530 29560 -510
rect 29450 -590 29470 -530
rect 29540 -590 29560 -530
rect 29450 -610 29560 -590
rect 29620 -530 29730 -510
rect 29620 -590 29640 -530
rect 29710 -590 29730 -530
rect 29620 -610 29730 -590
rect 29790 -530 29900 -510
rect 29790 -590 29810 -530
rect 29880 -590 29900 -530
rect 29790 -610 29900 -590
rect 29960 -530 30070 -510
rect 29960 -590 29980 -530
rect 30050 -590 30070 -530
rect 29960 -610 30070 -590
rect 30130 -530 30240 -510
rect 30130 -590 30150 -530
rect 30220 -590 30240 -530
rect 30130 -610 30240 -590
rect 30300 -530 30410 -510
rect 30300 -590 30320 -530
rect 30390 -590 30410 -530
rect 30300 -610 30410 -590
rect 30470 -530 30580 -510
rect 30470 -590 30490 -530
rect 30560 -590 30580 -530
rect 30470 -610 30580 -590
rect 30640 -530 30750 -510
rect 30640 -590 30660 -530
rect 30730 -590 30750 -530
rect 30640 -610 30750 -590
rect 30810 -530 30920 -510
rect 30810 -590 30830 -530
rect 30900 -590 30920 -530
rect 30810 -610 30920 -590
rect 30980 -530 31090 -510
rect 30980 -590 31000 -530
rect 31070 -590 31090 -530
rect 30980 -610 31090 -590
rect 31150 -530 31260 -510
rect 31150 -590 31170 -530
rect 31240 -590 31260 -530
rect 31150 -610 31260 -590
rect 31320 -530 31430 -510
rect 31320 -590 31340 -530
rect 31410 -590 31430 -530
rect 31320 -610 31430 -590
rect 31490 -530 31600 -510
rect 31490 -590 31510 -530
rect 31580 -590 31600 -530
rect 31490 -610 31600 -590
rect 31660 -530 31770 -510
rect 31660 -590 31680 -530
rect 31750 -590 31770 -530
rect 31660 -610 31770 -590
rect 31830 -530 31940 -510
rect 31830 -590 31850 -530
rect 31920 -590 31940 -530
rect 31830 -610 31940 -590
rect 32000 -530 32110 -510
rect 32000 -590 32020 -530
rect 32090 -590 32110 -530
rect 32000 -610 32110 -590
rect 32170 -530 32280 -510
rect 32170 -590 32190 -530
rect 32260 -590 32280 -530
rect 32170 -610 32280 -590
rect 32340 -530 32450 -510
rect 32340 -590 32360 -530
rect 32430 -590 32450 -530
rect 32340 -610 32450 -590
rect 32510 -530 32620 -510
rect 32510 -590 32530 -530
rect 32600 -590 32620 -530
rect 32510 -610 32620 -590
rect 32680 -530 32790 -510
rect 32680 -590 32700 -530
rect 32770 -590 32790 -530
rect 32680 -610 32790 -590
rect 32850 -530 32960 -510
rect 32850 -590 32870 -530
rect 32940 -590 32960 -530
rect 32850 -610 32960 -590
rect 33020 -530 33130 -510
rect 33020 -590 33040 -530
rect 33110 -590 33130 -530
rect 33020 -610 33130 -590
rect 33190 -530 33300 -510
rect 33190 -590 33210 -530
rect 33280 -590 33300 -530
rect 33190 -610 33300 -590
rect 33360 -530 33470 -510
rect 33360 -590 33380 -530
rect 33450 -590 33470 -530
rect 33360 -610 33470 -590
rect 33530 -530 33640 -510
rect 33530 -590 33550 -530
rect 33620 -590 33640 -530
rect 33530 -610 33640 -590
rect 33700 -530 33810 -510
rect 33700 -590 33720 -530
rect 33790 -590 33810 -530
rect 33700 -610 33810 -590
rect 33870 -530 33980 -510
rect 33870 -590 33890 -530
rect 33960 -590 33980 -530
rect 33870 -610 33980 -590
rect 34040 -530 34150 -510
rect 34040 -590 34060 -530
rect 34130 -590 34150 -530
rect 34040 -610 34150 -590
rect 34210 -530 34320 -510
rect 34210 -590 34230 -530
rect 34300 -590 34320 -530
rect 34210 -610 34320 -590
rect 34380 -530 34490 -510
rect 34380 -590 34400 -530
rect 34470 -590 34490 -530
rect 34380 -610 34490 -590
rect 34550 -530 34660 -510
rect 34550 -590 34570 -530
rect 34640 -590 34660 -530
rect 34550 -610 34660 -590
rect 34720 -530 34830 -510
rect 34720 -590 34740 -530
rect 34810 -590 34830 -530
rect 34720 -610 34830 -590
rect 34890 -530 35000 -510
rect 34890 -590 34910 -530
rect 34980 -590 35000 -530
rect 34890 -610 35000 -590
rect 35060 -530 35170 -510
rect 35060 -590 35080 -530
rect 35150 -590 35170 -530
rect 35060 -610 35170 -590
rect 35230 -530 35340 -510
rect 35230 -590 35250 -530
rect 35320 -590 35340 -530
rect 35230 -610 35340 -590
rect 35400 -530 35510 -510
rect 35400 -590 35420 -530
rect 35490 -590 35510 -530
rect 35400 -610 35510 -590
rect 35570 -530 35680 -510
rect 35570 -590 35590 -530
rect 35660 -590 35680 -530
rect 35570 -610 35680 -590
rect 35740 -530 35850 -510
rect 35740 -590 35760 -530
rect 35830 -590 35850 -530
rect 35740 -610 35850 -590
rect 35910 -530 36020 -510
rect 35910 -590 35930 -530
rect 36000 -590 36020 -530
rect 35910 -610 36020 -590
rect 36080 -530 36190 -510
rect 36080 -590 36100 -530
rect 36170 -590 36190 -530
rect 36080 -610 36190 -590
rect 36250 -530 36360 -510
rect 36250 -590 36270 -530
rect 36340 -590 36360 -530
rect 36250 -610 36360 -590
rect 36420 -530 36530 -510
rect 36420 -590 36440 -530
rect 36510 -590 36530 -530
rect 36420 -610 36530 -590
rect 36590 -530 36700 -510
rect 36590 -590 36610 -530
rect 36680 -590 36700 -530
rect 36590 -610 36700 -590
rect 36760 -530 36870 -510
rect 36760 -590 36780 -530
rect 36850 -590 36870 -530
rect 36760 -610 36870 -590
rect 36930 -530 37040 -510
rect 36930 -590 36950 -530
rect 37020 -590 37040 -530
rect 36930 -610 37040 -590
rect 37100 -530 37210 -510
rect 37100 -590 37120 -530
rect 37190 -590 37210 -530
rect 37100 -610 37210 -590
rect 37270 -530 37380 -510
rect 37270 -590 37290 -530
rect 37360 -590 37380 -530
rect 37270 -610 37380 -590
rect 37440 -530 37550 -510
rect 37440 -590 37460 -530
rect 37530 -590 37550 -530
rect 37440 -610 37550 -590
rect 37610 -530 37720 -510
rect 37610 -590 37630 -530
rect 37700 -590 37720 -530
rect 37610 -610 37720 -590
rect 37780 -530 37890 -510
rect 37780 -590 37800 -530
rect 37870 -590 37890 -530
rect 37780 -610 37890 -590
rect 37950 -530 38060 -510
rect 37950 -590 37970 -530
rect 38040 -590 38060 -530
rect 37950 -610 38060 -590
rect 38120 -530 38230 -510
rect 38120 -590 38140 -530
rect 38210 -590 38230 -530
rect 38120 -610 38230 -590
rect 38290 -530 38400 -510
rect 38290 -590 38310 -530
rect 38380 -590 38400 -530
rect 38290 -610 38400 -590
rect 38460 -530 38570 -510
rect 38460 -590 38480 -530
rect 38550 -590 38570 -530
rect 38460 -610 38570 -590
rect 38630 -530 38740 -510
rect 38630 -590 38650 -530
rect 38720 -590 38740 -530
rect 38630 -610 38740 -590
rect 38800 -530 38910 -510
rect 38800 -590 38820 -530
rect 38890 -590 38910 -530
rect 38800 -610 38910 -590
rect 38970 -530 39080 -510
rect 38970 -590 38990 -530
rect 39060 -590 39080 -530
rect 38970 -610 39080 -590
rect 39140 -530 39250 -510
rect 39140 -590 39160 -530
rect 39230 -590 39250 -530
rect 39140 -610 39250 -590
rect 39310 -530 39420 -510
rect 39310 -590 39330 -530
rect 39400 -590 39420 -530
rect 39310 -610 39420 -590
rect 39480 -530 39590 -510
rect 39480 -590 39500 -530
rect 39570 -590 39590 -530
rect 39480 -610 39590 -590
rect 39650 -530 39760 -510
rect 39650 -590 39670 -530
rect 39740 -590 39760 -530
rect 39650 -610 39760 -590
rect 39820 -530 39930 -510
rect 39820 -590 39840 -530
rect 39910 -590 39930 -530
rect 39820 -610 39930 -590
rect 39990 -530 40100 -510
rect 39990 -590 40010 -530
rect 40080 -590 40100 -530
rect 39990 -610 40100 -590
rect 40160 -530 40270 -510
rect 40160 -590 40180 -530
rect 40250 -590 40270 -530
rect 40160 -610 40270 -590
rect 40330 -530 40440 -510
rect 40330 -590 40350 -530
rect 40420 -590 40440 -530
rect 40330 -610 40440 -590
rect 40500 -530 40610 -510
rect 40500 -590 40520 -530
rect 40590 -590 40610 -530
rect 40500 -610 40610 -590
rect 40670 -530 40780 -510
rect 40670 -590 40690 -530
rect 40760 -590 40780 -530
rect 40670 -610 40780 -590
rect 40840 -530 40950 -510
rect 40840 -590 40860 -530
rect 40930 -590 40950 -530
rect 40840 -610 40950 -590
rect 41010 -530 41120 -510
rect 41010 -590 41030 -530
rect 41100 -590 41120 -530
rect 41010 -610 41120 -590
rect 41180 -530 41290 -510
rect 41180 -590 41200 -530
rect 41270 -590 41290 -530
rect 41180 -610 41290 -590
rect 41350 -530 41460 -510
rect 41350 -590 41370 -530
rect 41440 -590 41460 -530
rect 41350 -610 41460 -590
rect 41520 -530 41630 -510
rect 41520 -590 41540 -530
rect 41610 -590 41630 -530
rect 41520 -610 41630 -590
rect 41690 -530 41800 -510
rect 41690 -590 41710 -530
rect 41780 -590 41800 -530
rect 41690 -610 41800 -590
rect 41860 -530 41970 -510
rect 41860 -590 41880 -530
rect 41950 -590 41970 -530
rect 41860 -610 41970 -590
rect 42030 -530 42140 -510
rect 42030 -590 42050 -530
rect 42120 -590 42140 -530
rect 42030 -610 42140 -590
rect 42200 -530 42310 -510
rect 42200 -590 42220 -530
rect 42290 -590 42310 -530
rect 42200 -610 42310 -590
rect 42370 -530 42480 -510
rect 42370 -590 42390 -530
rect 42460 -590 42480 -530
rect 42370 -610 42480 -590
rect 42540 -530 42650 -510
rect 42540 -590 42560 -530
rect 42630 -590 42650 -530
rect 42540 -610 42650 -590
rect 42710 -530 42820 -510
rect 42710 -590 42730 -530
rect 42800 -590 42820 -530
rect 42710 -610 42820 -590
rect 42880 -530 42990 -510
rect 42880 -590 42900 -530
rect 42970 -590 42990 -530
rect 42880 -610 42990 -590
rect 43050 -530 43160 -510
rect 43050 -590 43070 -530
rect 43140 -590 43160 -530
rect 43050 -610 43160 -590
rect 43220 -530 43330 -510
rect 43220 -590 43240 -530
rect 43310 -590 43330 -530
rect 43220 -610 43330 -590
rect 43390 -530 43500 -510
rect 43390 -590 43410 -530
rect 43480 -590 43500 -530
rect 43390 -610 43500 -590
rect 43560 -530 43670 -510
rect 43560 -590 43580 -530
rect 43650 -590 43670 -530
rect 43560 -610 43670 -590
rect 43730 -530 43840 -510
rect 43730 -590 43750 -530
rect 43820 -590 43840 -530
rect 43730 -610 43840 -590
rect 43900 -530 44010 -510
rect 43900 -590 43920 -530
rect 43990 -590 44010 -530
rect 43900 -610 44010 -590
rect 44070 -530 44180 -510
rect 44070 -590 44090 -530
rect 44160 -590 44180 -530
rect 44070 -610 44180 -590
rect 44240 -530 44350 -510
rect 44240 -590 44260 -530
rect 44330 -590 44350 -530
rect 44240 -610 44350 -590
rect 44410 -530 44520 -510
rect 44410 -590 44430 -530
rect 44500 -590 44520 -530
rect 44410 -610 44520 -590
rect 44580 -530 44690 -510
rect 44580 -590 44600 -530
rect 44670 -590 44690 -530
rect 44580 -610 44690 -590
rect 44750 -530 44860 -510
rect 44750 -590 44770 -530
rect 44840 -590 44860 -530
rect 44750 -610 44860 -590
rect 44920 -530 45030 -510
rect 44920 -590 44940 -530
rect 45010 -590 45030 -530
rect 44920 -610 45030 -590
rect 45090 -530 45200 -510
rect 45090 -590 45110 -530
rect 45180 -590 45200 -530
rect 45090 -610 45200 -590
rect 45260 -530 45370 -510
rect 45260 -590 45280 -530
rect 45350 -590 45370 -530
rect 45260 -610 45370 -590
rect 45430 -530 45540 -510
rect 45430 -590 45450 -530
rect 45520 -590 45540 -530
rect 45430 -610 45540 -590
rect 45600 -530 45710 -510
rect 45600 -590 45620 -530
rect 45690 -590 45710 -530
rect 45600 -610 45710 -590
rect 45770 -530 45880 -510
rect 45770 -590 45790 -530
rect 45860 -590 45880 -530
rect 45770 -610 45880 -590
rect 45940 -530 46050 -510
rect 45940 -590 45960 -530
rect 46030 -590 46050 -530
rect 45940 -610 46050 -590
rect 46110 -530 46220 -510
rect 46110 -590 46130 -530
rect 46200 -590 46220 -530
rect 46110 -610 46220 -590
rect 46280 -530 46390 -510
rect 46280 -590 46300 -530
rect 46370 -590 46390 -530
rect 46280 -610 46390 -590
rect 46450 -530 46560 -510
rect 46450 -590 46470 -530
rect 46540 -590 46560 -530
rect 46450 -610 46560 -590
rect 46620 -530 46730 -510
rect 46620 -590 46640 -530
rect 46710 -590 46730 -530
rect 46620 -610 46730 -590
rect 46790 -530 46900 -510
rect 46790 -590 46810 -530
rect 46880 -590 46900 -530
rect 46790 -610 46900 -590
rect 46960 -530 47070 -510
rect 46960 -590 46980 -530
rect 47050 -590 47070 -530
rect 46960 -610 47070 -590
rect 47130 -530 47240 -510
rect 47130 -590 47150 -530
rect 47220 -590 47240 -530
rect 47130 -610 47240 -590
rect 47300 -530 47410 -510
rect 47300 -590 47320 -530
rect 47390 -590 47410 -530
rect 47300 -610 47410 -590
rect 47470 -530 47580 -510
rect 47470 -590 47490 -530
rect 47560 -590 47580 -530
rect 47470 -610 47580 -590
rect 47640 -530 47750 -510
rect 47640 -590 47660 -530
rect 47730 -590 47750 -530
rect 47640 -610 47750 -590
rect 47810 -530 47920 -510
rect 47810 -590 47830 -530
rect 47900 -590 47920 -530
rect 47810 -610 47920 -590
rect 47980 -530 48090 -510
rect 47980 -590 48000 -530
rect 48070 -590 48090 -530
rect 47980 -610 48090 -590
rect 48150 -530 48260 -510
rect 48150 -590 48170 -530
rect 48240 -590 48260 -530
rect 48150 -610 48260 -590
rect 48320 -530 48430 -510
rect 48320 -590 48340 -530
rect 48410 -590 48430 -530
rect 48320 -610 48430 -590
rect 48490 -530 48600 -510
rect 48490 -590 48510 -530
rect 48580 -590 48600 -530
rect 48490 -610 48600 -590
rect 48660 -530 48770 -510
rect 48660 -590 48680 -530
rect 48750 -590 48770 -530
rect 48660 -610 48770 -590
rect 48830 -530 48940 -510
rect 48830 -590 48850 -530
rect 48920 -590 48940 -530
rect 48830 -610 48940 -590
rect 49000 -530 49110 -510
rect 49000 -590 49020 -530
rect 49090 -590 49110 -530
rect 49000 -610 49110 -590
rect 49170 -530 49280 -510
rect 49170 -590 49190 -530
rect 49260 -590 49280 -530
rect 49170 -610 49280 -590
rect 49340 -530 49450 -510
rect 49340 -590 49360 -530
rect 49430 -590 49450 -530
rect 49340 -610 49450 -590
rect 49510 -530 49620 -510
rect 49510 -590 49530 -530
rect 49600 -590 49620 -530
rect 49510 -610 49620 -590
rect 49680 -530 49790 -510
rect 49680 -590 49700 -530
rect 49770 -590 49790 -530
rect 49680 -610 49790 -590
rect 49850 -530 49960 -510
rect 49850 -590 49870 -530
rect 49940 -590 49960 -530
rect 49850 -610 49960 -590
rect 50020 -530 50130 -510
rect 50020 -590 50040 -530
rect 50110 -590 50130 -530
rect 50020 -610 50130 -590
rect 50190 -530 50300 -510
rect 50190 -590 50210 -530
rect 50280 -590 50300 -530
rect 50190 -610 50300 -590
rect 50360 -530 50470 -510
rect 50360 -590 50380 -530
rect 50450 -590 50470 -530
rect 50360 -610 50470 -590
rect 50530 -530 50640 -510
rect 50530 -590 50550 -530
rect 50620 -590 50640 -530
rect 50530 -610 50640 -590
rect 50700 -530 50810 -510
rect 50700 -590 50720 -530
rect 50790 -590 50810 -530
rect 50700 -610 50810 -590
rect 50870 -530 50980 -510
rect 50870 -590 50890 -530
rect 50960 -590 50980 -530
rect 50870 -610 50980 -590
rect 51040 -530 51150 -510
rect 51040 -590 51060 -530
rect 51130 -590 51150 -530
rect 51040 -610 51150 -590
rect 51210 -530 51320 -510
rect 51210 -590 51230 -530
rect 51300 -590 51320 -530
rect 51210 -610 51320 -590
rect 51380 -530 51490 -510
rect 51380 -590 51400 -530
rect 51470 -590 51490 -530
rect 51380 -610 51490 -590
rect 51550 -530 51660 -510
rect 51550 -590 51570 -530
rect 51640 -590 51660 -530
rect 51550 -610 51660 -590
rect 51720 -530 51830 -510
rect 51720 -590 51740 -530
rect 51810 -590 51830 -530
rect 51720 -610 51830 -590
rect 51890 -530 52000 -510
rect 51890 -590 51910 -530
rect 51980 -590 52000 -530
rect 51890 -610 52000 -590
rect 52060 -530 52170 -510
rect 52060 -590 52080 -530
rect 52150 -590 52170 -530
rect 52060 -610 52170 -590
rect 52230 -530 52340 -510
rect 52230 -590 52250 -530
rect 52320 -590 52340 -530
rect 52230 -610 52340 -590
rect 52400 -530 52510 -510
rect 52400 -590 52420 -530
rect 52490 -590 52510 -530
rect 52400 -610 52510 -590
rect 52570 -530 52680 -510
rect 52570 -590 52590 -530
rect 52660 -590 52680 -530
rect 52570 -610 52680 -590
rect 52740 -530 52850 -510
rect 52740 -590 52760 -530
rect 52830 -590 52850 -530
rect 52740 -610 52850 -590
rect 52910 -530 53020 -510
rect 52910 -590 52930 -530
rect 53000 -590 53020 -530
rect 52910 -610 53020 -590
rect 53080 -530 53190 -510
rect 53080 -590 53100 -530
rect 53170 -590 53190 -530
rect 53080 -610 53190 -590
rect 53250 -530 53360 -510
rect 53250 -590 53270 -530
rect 53340 -590 53360 -530
rect 53250 -610 53360 -590
rect 53420 -530 53530 -510
rect 53420 -590 53440 -530
rect 53510 -590 53530 -530
rect 53420 -610 53530 -590
rect 53590 -530 53700 -510
rect 53590 -590 53610 -530
rect 53680 -590 53700 -530
rect 53590 -610 53700 -590
rect 53760 -530 53870 -510
rect 53760 -590 53780 -530
rect 53850 -590 53870 -530
rect 53760 -610 53870 -590
rect 53930 -530 54040 -510
rect 53930 -590 53950 -530
rect 54020 -590 54040 -530
rect 53930 -610 54040 -590
rect 54100 -530 54210 -510
rect 54100 -590 54120 -530
rect 54190 -590 54210 -530
rect 54100 -610 54210 -590
rect 54270 -530 54380 -510
rect 54270 -590 54290 -530
rect 54360 -590 54380 -530
rect 54270 -610 54380 -590
rect 54440 -530 54550 -510
rect 54440 -590 54460 -530
rect 54530 -590 54550 -530
rect 54440 -610 54550 -590
rect 54610 -530 54720 -510
rect 54610 -590 54630 -530
rect 54700 -590 54720 -530
rect 54610 -610 54720 -590
rect 54780 -530 54890 -510
rect 54780 -590 54800 -530
rect 54870 -590 54890 -530
rect 54780 -610 54890 -590
rect 54950 -530 55060 -510
rect 54950 -590 54970 -530
rect 55040 -590 55060 -530
rect 54950 -610 55060 -590
rect 55120 -530 55230 -510
rect 55120 -590 55140 -530
rect 55210 -590 55230 -530
rect 55120 -610 55230 -590
rect 55290 -530 55400 -510
rect 55290 -590 55310 -530
rect 55380 -590 55400 -530
rect 55290 -610 55400 -590
rect 55460 -530 55570 -510
rect 55460 -590 55480 -530
rect 55550 -590 55570 -530
rect 55460 -610 55570 -590
rect 55630 -530 55740 -510
rect 55630 -590 55650 -530
rect 55720 -590 55740 -530
rect 55630 -610 55740 -590
rect 55800 -530 55910 -510
rect 55800 -590 55820 -530
rect 55890 -590 55910 -530
rect 55800 -610 55910 -590
rect 55970 -530 56080 -510
rect 55970 -590 55990 -530
rect 56060 -590 56080 -530
rect 55970 -610 56080 -590
rect 56140 -530 56250 -510
rect 56140 -590 56160 -530
rect 56230 -590 56250 -530
rect 56140 -610 56250 -590
rect 56310 -530 56420 -510
rect 56310 -590 56330 -530
rect 56400 -590 56420 -530
rect 56310 -610 56420 -590
rect 56480 -530 56590 -510
rect 56480 -590 56500 -530
rect 56570 -590 56590 -530
rect 56480 -610 56590 -590
rect 56650 -530 56760 -510
rect 56650 -590 56670 -530
rect 56740 -590 56760 -530
rect 56650 -610 56760 -590
rect 56820 -530 56930 -510
rect 56820 -590 56840 -530
rect 56910 -590 56930 -530
rect 56820 -610 56930 -590
rect 56990 -530 57100 -510
rect 56990 -590 57010 -530
rect 57080 -590 57100 -530
rect 56990 -610 57100 -590
rect 57160 -530 57270 -510
rect 57160 -590 57180 -530
rect 57250 -590 57270 -530
rect 57160 -610 57270 -590
rect 57330 -530 57440 -510
rect 57330 -590 57350 -530
rect 57420 -590 57440 -530
rect 57330 -610 57440 -590
rect 57500 -530 57610 -510
rect 57500 -590 57520 -530
rect 57590 -590 57610 -530
rect 57500 -610 57610 -590
rect 57670 -530 57780 -510
rect 57670 -590 57690 -530
rect 57760 -590 57780 -530
rect 57670 -610 57780 -590
rect 57840 -530 57950 -510
rect 57840 -590 57860 -530
rect 57930 -590 57950 -530
rect 57840 -610 57950 -590
rect 58010 -530 58120 -510
rect 58010 -590 58030 -530
rect 58100 -590 58120 -530
rect 58010 -610 58120 -590
rect 58180 -530 58290 -510
rect 58180 -590 58200 -530
rect 58270 -590 58290 -530
rect 58180 -610 58290 -590
rect 58350 -530 58460 -510
rect 58350 -590 58370 -530
rect 58440 -590 58460 -530
rect 58350 -610 58460 -590
rect 58520 -530 58630 -510
rect 58520 -590 58540 -530
rect 58610 -590 58630 -530
rect 58520 -610 58630 -590
rect 58690 -530 58800 -510
rect 58690 -590 58710 -530
rect 58780 -590 58800 -530
rect 58690 -610 58800 -590
rect 58860 -530 58970 -510
rect 58860 -590 58880 -530
rect 58950 -590 58970 -530
rect 58860 -610 58970 -590
rect 59030 -530 59140 -510
rect 59030 -590 59050 -530
rect 59120 -590 59140 -530
rect 59030 -610 59140 -590
rect 59200 -530 59310 -510
rect 59200 -590 59220 -530
rect 59290 -590 59310 -530
rect 59200 -610 59310 -590
rect 59370 -530 59480 -510
rect 59370 -590 59390 -530
rect 59460 -590 59480 -530
rect 59370 -610 59480 -590
rect 59540 -530 59650 -510
rect 59540 -590 59560 -530
rect 59630 -590 59650 -530
rect 59540 -610 59650 -590
rect 59710 -530 59820 -510
rect 59710 -590 59730 -530
rect 59800 -590 59820 -530
rect 59710 -610 59820 -590
rect 59880 -530 59990 -510
rect 59880 -590 59900 -530
rect 59970 -590 59990 -530
rect 59880 -610 59990 -590
rect 60050 -530 60160 -510
rect 60050 -590 60070 -530
rect 60140 -590 60160 -530
rect 60050 -610 60160 -590
rect 60220 -530 60330 -510
rect 60220 -590 60240 -530
rect 60310 -590 60330 -530
rect 60220 -610 60330 -590
rect 60390 -530 60500 -510
rect 60390 -590 60410 -530
rect 60480 -590 60500 -530
rect 60390 -610 60500 -590
rect 60560 -530 60670 -510
rect 60560 -590 60580 -530
rect 60650 -590 60670 -530
rect 60560 -610 60670 -590
rect 60730 -530 60840 -510
rect 60730 -590 60750 -530
rect 60820 -590 60840 -530
rect 60730 -610 60840 -590
rect 60900 -530 61010 -510
rect 60900 -590 60920 -530
rect 60990 -590 61010 -530
rect 60900 -610 61010 -590
rect 61070 -530 61180 -510
rect 61070 -590 61090 -530
rect 61160 -590 61180 -530
rect 61070 -610 61180 -590
rect 61240 -530 61350 -510
rect 61240 -590 61260 -530
rect 61330 -590 61350 -530
rect 61240 -610 61350 -590
rect 61410 -530 61520 -510
rect 61410 -590 61430 -530
rect 61500 -590 61520 -530
rect 61410 -610 61520 -590
rect 61580 -530 61690 -510
rect 61580 -590 61600 -530
rect 61670 -590 61690 -530
rect 61580 -610 61690 -590
rect 61750 -530 61860 -510
rect 61750 -590 61770 -530
rect 61840 -590 61860 -530
rect 61750 -610 61860 -590
rect 61920 -530 62030 -510
rect 61920 -590 61940 -530
rect 62010 -590 62030 -530
rect 61920 -610 62030 -590
rect 62090 -530 62200 -510
rect 62090 -590 62110 -530
rect 62180 -590 62200 -530
rect 62090 -610 62200 -590
rect 62260 -530 62370 -510
rect 62260 -590 62280 -530
rect 62350 -590 62370 -530
rect 62260 -610 62370 -590
rect 62430 -530 62540 -510
rect 62430 -590 62450 -530
rect 62520 -590 62540 -530
rect 62430 -610 62540 -590
rect 62600 -530 62710 -510
rect 62600 -590 62620 -530
rect 62690 -590 62710 -530
rect 62600 -610 62710 -590
rect 62770 -530 62880 -510
rect 62770 -590 62790 -530
rect 62860 -590 62880 -530
rect 62770 -610 62880 -590
rect 62940 -530 63050 -510
rect 62940 -590 62960 -530
rect 63030 -590 63050 -530
rect 62940 -610 63050 -590
rect 63110 -530 63220 -510
rect 63110 -590 63130 -530
rect 63200 -590 63220 -530
rect 63110 -610 63220 -590
rect 63280 -530 63390 -510
rect 63280 -590 63300 -530
rect 63370 -590 63390 -530
rect 63280 -610 63390 -590
rect 63450 -530 63560 -510
rect 63450 -590 63470 -530
rect 63540 -590 63560 -530
rect 63450 -610 63560 -590
rect 63620 -530 63730 -510
rect 63620 -590 63640 -530
rect 63710 -590 63730 -530
rect 63620 -610 63730 -590
rect 63790 -530 63900 -510
rect 63790 -590 63810 -530
rect 63880 -590 63900 -530
rect 63790 -610 63900 -590
rect 63960 -530 64070 -510
rect 63960 -590 63980 -530
rect 64050 -590 64070 -530
rect 63960 -610 64070 -590
rect 64130 -530 64240 -510
rect 64130 -590 64150 -530
rect 64220 -590 64240 -530
rect 64130 -610 64240 -590
rect 64300 -530 64410 -510
rect 64300 -590 64320 -530
rect 64390 -590 64410 -530
rect 64300 -610 64410 -590
rect 64470 -530 64580 -510
rect 64470 -590 64490 -530
rect 64560 -590 64580 -530
rect 64470 -610 64580 -590
rect 64640 -530 64750 -510
rect 64640 -590 64660 -530
rect 64730 -590 64750 -530
rect 64640 -610 64750 -590
rect 64810 -530 64920 -510
rect 64810 -590 64830 -530
rect 64900 -590 64920 -530
rect 64810 -610 64920 -590
rect 64980 -530 65090 -510
rect 64980 -590 65000 -530
rect 65070 -590 65090 -530
rect 64980 -610 65090 -590
rect 65150 -530 65260 -510
rect 65150 -590 65170 -530
rect 65240 -590 65260 -530
rect 65150 -610 65260 -590
rect 65320 -530 65430 -510
rect 65320 -590 65340 -530
rect 65410 -590 65430 -530
rect 65320 -610 65430 -590
rect 65490 -530 65600 -510
rect 65490 -590 65510 -530
rect 65580 -590 65600 -530
rect 65490 -610 65600 -590
rect 65660 -530 65770 -510
rect 65660 -590 65680 -530
rect 65750 -590 65770 -530
rect 65660 -610 65770 -590
rect 65830 -530 65940 -510
rect 65830 -590 65850 -530
rect 65920 -590 65940 -530
rect 65830 -610 65940 -590
rect 66000 -530 66110 -510
rect 66000 -590 66020 -530
rect 66090 -590 66110 -530
rect 66000 -610 66110 -590
rect 66170 -530 66280 -510
rect 66170 -590 66190 -530
rect 66260 -590 66280 -530
rect 66170 -610 66280 -590
rect 66340 -530 66450 -510
rect 66340 -590 66360 -530
rect 66430 -590 66450 -530
rect 66340 -610 66450 -590
rect 66510 -530 66620 -510
rect 66510 -590 66530 -530
rect 66600 -590 66620 -530
rect 66510 -610 66620 -590
rect 66680 -530 66790 -510
rect 66680 -590 66700 -530
rect 66770 -590 66790 -530
rect 66680 -610 66790 -590
rect 66850 -530 66960 -510
rect 66850 -590 66870 -530
rect 66940 -590 66960 -530
rect 66850 -610 66960 -590
rect 67020 -530 67130 -510
rect 67020 -590 67040 -530
rect 67110 -590 67130 -530
rect 67020 -610 67130 -590
rect 67190 -530 67300 -510
rect 67190 -590 67210 -530
rect 67280 -590 67300 -530
rect 67190 -610 67300 -590
rect 67360 -530 67470 -510
rect 67360 -590 67380 -530
rect 67450 -590 67470 -530
rect 67360 -610 67470 -590
rect 67530 -530 67640 -510
rect 67530 -590 67550 -530
rect 67620 -590 67640 -530
rect 67530 -610 67640 -590
rect 67700 -530 67810 -510
rect 67700 -590 67720 -530
rect 67790 -590 67810 -530
rect 67700 -610 67810 -590
rect 67870 -530 67980 -510
rect 67870 -590 67890 -530
rect 67960 -590 67980 -530
rect 67870 -610 67980 -590
rect 68040 -530 68150 -510
rect 68040 -590 68060 -530
rect 68130 -590 68150 -530
rect 68040 -610 68150 -590
rect 68210 -530 68320 -510
rect 68210 -590 68230 -530
rect 68300 -590 68320 -530
rect 68210 -610 68320 -590
rect 68380 -530 68490 -510
rect 68380 -590 68400 -530
rect 68470 -590 68490 -530
rect 68380 -610 68490 -590
rect 68550 -530 68660 -510
rect 68550 -590 68570 -530
rect 68640 -590 68660 -530
rect 68550 -610 68660 -590
rect 68720 -530 68830 -510
rect 68720 -590 68740 -530
rect 68810 -590 68830 -530
rect 68720 -610 68830 -590
rect 68890 -530 69000 -510
rect 68890 -590 68910 -530
rect 68980 -590 69000 -530
rect 68890 -610 69000 -590
rect 69060 -530 69170 -510
rect 69060 -590 69080 -530
rect 69150 -590 69170 -530
rect 69060 -610 69170 -590
rect 69230 -530 69340 -510
rect 69230 -590 69250 -530
rect 69320 -590 69340 -530
rect 69230 -610 69340 -590
rect 69400 -530 69510 -510
rect 69400 -590 69420 -530
rect 69490 -590 69510 -530
rect 69400 -610 69510 -590
rect 69570 -530 69680 -510
rect 69570 -590 69590 -530
rect 69660 -590 69680 -530
rect 69570 -610 69680 -590
rect 69740 -530 69850 -510
rect 69740 -590 69760 -530
rect 69830 -590 69850 -530
rect 69740 -610 69850 -590
rect 69910 -530 70020 -510
rect 69910 -590 69930 -530
rect 70000 -590 70020 -530
rect 69910 -610 70020 -590
rect 70080 -530 70190 -510
rect 70080 -590 70100 -530
rect 70170 -590 70190 -530
rect 70080 -610 70190 -590
rect 70250 -530 70360 -510
rect 70250 -590 70270 -530
rect 70340 -590 70360 -530
rect 70250 -610 70360 -590
rect 70420 -530 70530 -510
rect 70420 -590 70440 -530
rect 70510 -590 70530 -530
rect 70420 -610 70530 -590
rect 70590 -530 70700 -510
rect 70590 -590 70610 -530
rect 70680 -590 70700 -530
rect 70590 -610 70700 -590
rect 70760 -530 70870 -510
rect 70760 -590 70780 -530
rect 70850 -590 70870 -530
rect 70760 -610 70870 -590
rect 70930 -530 71040 -510
rect 70930 -590 70950 -530
rect 71020 -590 71040 -530
rect 70930 -610 71040 -590
rect 71100 -530 71210 -510
rect 71100 -590 71120 -530
rect 71190 -590 71210 -530
rect 71100 -610 71210 -590
rect 71270 -530 71380 -510
rect 71270 -590 71290 -530
rect 71360 -590 71380 -530
rect 71270 -610 71380 -590
rect 71440 -530 71550 -510
rect 71440 -590 71460 -530
rect 71530 -590 71550 -530
rect 71440 -610 71550 -590
rect 71610 -530 71720 -510
rect 71610 -590 71630 -530
rect 71700 -590 71720 -530
rect 71610 -610 71720 -590
rect 71780 -530 71890 -510
rect 71780 -590 71800 -530
rect 71870 -590 71890 -530
rect 71780 -610 71890 -590
rect 71950 -530 72060 -510
rect 71950 -590 71970 -530
rect 72040 -590 72060 -530
rect 71950 -610 72060 -590
rect 72120 -530 72230 -510
rect 72120 -590 72140 -530
rect 72210 -590 72230 -530
rect 72120 -610 72230 -590
rect 72290 -530 72400 -510
rect 72290 -590 72310 -530
rect 72380 -590 72400 -530
rect 72290 -610 72400 -590
rect 72460 -530 72570 -510
rect 72460 -590 72480 -530
rect 72550 -590 72570 -530
rect 72460 -610 72570 -590
rect 72630 -530 72740 -510
rect 72630 -590 72650 -530
rect 72720 -590 72740 -530
rect 72630 -610 72740 -590
rect 72800 -530 72910 -510
rect 72800 -590 72820 -530
rect 72890 -590 72910 -530
rect 72800 -610 72910 -590
rect 72970 -530 73080 -510
rect 72970 -590 72990 -530
rect 73060 -590 73080 -530
rect 72970 -610 73080 -590
rect 73140 -530 73250 -510
rect 73140 -590 73160 -530
rect 73230 -590 73250 -530
rect 73140 -610 73250 -590
rect 73310 -530 73420 -510
rect 73310 -590 73330 -530
rect 73400 -590 73420 -530
rect 73310 -610 73420 -590
rect 73480 -530 73590 -510
rect 73480 -590 73500 -530
rect 73570 -590 73590 -530
rect 73480 -610 73590 -590
rect 73650 -530 73760 -510
rect 73650 -590 73670 -530
rect 73740 -590 73760 -530
rect 73650 -610 73760 -590
rect 73820 -530 73930 -510
rect 73820 -590 73840 -530
rect 73910 -590 73930 -530
rect 73820 -610 73930 -590
rect 73990 -530 74100 -510
rect 73990 -590 74010 -530
rect 74080 -590 74100 -530
rect 73990 -610 74100 -590
rect 74160 -530 74270 -510
rect 74160 -590 74180 -530
rect 74250 -590 74270 -530
rect 74160 -610 74270 -590
rect 74330 -530 74440 -510
rect 74330 -590 74350 -530
rect 74420 -590 74440 -530
rect 74330 -610 74440 -590
rect 74500 -530 74610 -510
rect 74500 -590 74520 -530
rect 74590 -590 74610 -530
rect 74500 -610 74610 -590
rect 74670 -530 74780 -510
rect 74670 -590 74690 -530
rect 74760 -590 74780 -530
rect 74670 -610 74780 -590
rect 74840 -530 74950 -510
rect 74840 -590 74860 -530
rect 74930 -590 74950 -530
rect 74840 -610 74950 -590
rect 75010 -530 75120 -510
rect 75010 -590 75030 -530
rect 75100 -590 75120 -530
rect 75010 -610 75120 -590
rect 75180 -530 75290 -510
rect 75180 -590 75200 -530
rect 75270 -590 75290 -530
rect 75180 -610 75290 -590
rect 75350 -530 75460 -510
rect 75350 -590 75370 -530
rect 75440 -590 75460 -530
rect 75350 -610 75460 -590
rect 75520 -530 75630 -510
rect 75520 -590 75540 -530
rect 75610 -590 75630 -530
rect 75520 -610 75630 -590
rect 75690 -530 75800 -510
rect 75690 -590 75710 -530
rect 75780 -590 75800 -530
rect 75690 -610 75800 -590
rect 75860 -530 75970 -510
rect 75860 -590 75880 -530
rect 75950 -590 75970 -530
rect 75860 -610 75970 -590
rect 76030 -530 76140 -510
rect 76030 -590 76050 -530
rect 76120 -590 76140 -530
rect 76030 -610 76140 -590
rect 76200 -530 76310 -510
rect 76200 -590 76220 -530
rect 76290 -590 76310 -530
rect 76200 -610 76310 -590
rect 76370 -530 76480 -510
rect 76370 -590 76390 -530
rect 76460 -590 76480 -530
rect 76370 -610 76480 -590
rect 76540 -530 76650 -510
rect 76540 -590 76560 -530
rect 76630 -590 76650 -530
rect 76540 -610 76650 -590
rect 76710 -530 76820 -510
rect 76710 -590 76730 -530
rect 76800 -590 76820 -530
rect 76710 -610 76820 -590
rect 76880 -530 76990 -510
rect 76880 -590 76900 -530
rect 76970 -590 76990 -530
rect 76880 -610 76990 -590
rect 77050 -530 77160 -510
rect 77050 -590 77070 -530
rect 77140 -590 77160 -530
rect 77050 -610 77160 -590
rect 77220 -530 77330 -510
rect 77220 -590 77240 -530
rect 77310 -590 77330 -530
rect 77220 -610 77330 -590
rect 77390 -530 77500 -510
rect 77390 -590 77410 -530
rect 77480 -590 77500 -530
rect 77390 -610 77500 -590
rect 77560 -530 77670 -510
rect 77560 -590 77580 -530
rect 77650 -590 77670 -530
rect 77560 -610 77670 -590
rect 77730 -530 77840 -510
rect 77730 -590 77750 -530
rect 77820 -590 77840 -530
rect 77730 -610 77840 -590
rect 77900 -530 78010 -510
rect 77900 -590 77920 -530
rect 77990 -590 78010 -530
rect 77900 -610 78010 -590
rect 78070 -530 78180 -510
rect 78070 -590 78090 -530
rect 78160 -590 78180 -530
rect 78070 -610 78180 -590
rect 78240 -530 78350 -510
rect 78240 -590 78260 -530
rect 78330 -590 78350 -530
rect 78240 -610 78350 -590
rect 78410 -530 78520 -510
rect 78410 -590 78430 -530
rect 78500 -590 78520 -530
rect 78410 -610 78520 -590
rect 78580 -530 78690 -510
rect 78580 -590 78600 -530
rect 78670 -590 78690 -530
rect 78580 -610 78690 -590
rect 78750 -530 78860 -510
rect 78750 -590 78770 -530
rect 78840 -590 78860 -530
rect 78750 -610 78860 -590
rect 78920 -530 79030 -510
rect 78920 -590 78940 -530
rect 79010 -590 79030 -530
rect 78920 -610 79030 -590
rect 79090 -530 79200 -510
rect 79090 -590 79110 -530
rect 79180 -590 79200 -530
rect 79090 -610 79200 -590
rect 79260 -530 79370 -510
rect 79260 -590 79280 -530
rect 79350 -590 79370 -530
rect 79260 -610 79370 -590
rect 79430 -530 79540 -510
rect 79430 -590 79450 -530
rect 79520 -590 79540 -530
rect 79430 -610 79540 -590
rect 79600 -530 79710 -510
rect 79600 -590 79620 -530
rect 79690 -590 79710 -530
rect 79600 -610 79710 -590
rect 79770 -530 79880 -510
rect 79770 -590 79790 -530
rect 79860 -590 79880 -530
rect 79770 -610 79880 -590
rect 79940 -530 80050 -510
rect 79940 -590 79960 -530
rect 80030 -590 80050 -530
rect 79940 -610 80050 -590
rect 80110 -530 80220 -510
rect 80110 -590 80130 -530
rect 80200 -590 80220 -530
rect 80110 -610 80220 -590
rect 80280 -530 80390 -510
rect 80280 -590 80300 -530
rect 80370 -590 80390 -530
rect 80280 -610 80390 -590
rect 80450 -530 80560 -510
rect 80450 -590 80470 -530
rect 80540 -590 80560 -530
rect 80450 -610 80560 -590
rect 80620 -530 80730 -510
rect 80620 -590 80640 -530
rect 80710 -590 80730 -530
rect 80620 -610 80730 -590
rect 80790 -530 80900 -510
rect 80790 -590 80810 -530
rect 80880 -590 80900 -530
rect 80790 -610 80900 -590
rect 80960 -530 81070 -510
rect 80960 -590 80980 -530
rect 81050 -590 81070 -530
rect 80960 -610 81070 -590
rect 81130 -530 81240 -510
rect 81130 -590 81150 -530
rect 81220 -590 81240 -530
rect 81130 -610 81240 -590
rect 81300 -530 81410 -510
rect 81300 -590 81320 -530
rect 81390 -590 81410 -530
rect 81300 -610 81410 -590
rect 81470 -530 81580 -510
rect 81470 -590 81490 -530
rect 81560 -590 81580 -530
rect 81470 -610 81580 -590
rect 81640 -530 81750 -510
rect 81640 -590 81660 -530
rect 81730 -590 81750 -530
rect 81640 -610 81750 -590
rect 81810 -530 81920 -510
rect 81810 -590 81830 -530
rect 81900 -590 81920 -530
rect 81810 -610 81920 -590
rect 81980 -530 82090 -510
rect 81980 -590 82000 -530
rect 82070 -590 82090 -530
rect 81980 -610 82090 -590
rect 82150 -530 82260 -510
rect 82150 -590 82170 -530
rect 82240 -590 82260 -530
rect 82150 -610 82260 -590
rect 82320 -530 82430 -510
rect 82320 -590 82340 -530
rect 82410 -590 82430 -530
rect 82320 -610 82430 -590
rect 82490 -530 82600 -510
rect 82490 -590 82510 -530
rect 82580 -590 82600 -530
rect 82490 -610 82600 -590
rect 82660 -530 82770 -510
rect 82660 -590 82680 -530
rect 82750 -590 82770 -530
rect 82660 -610 82770 -590
rect 82830 -530 82940 -510
rect 82830 -590 82850 -530
rect 82920 -590 82940 -530
rect 82830 -610 82940 -590
rect 83000 -530 83110 -510
rect 83000 -590 83020 -530
rect 83090 -590 83110 -530
rect 83000 -610 83110 -590
rect 83170 -530 83280 -510
rect 83170 -590 83190 -530
rect 83260 -590 83280 -530
rect 83170 -610 83280 -590
rect 83340 -530 83450 -510
rect 83340 -590 83360 -530
rect 83430 -590 83450 -530
rect 83340 -610 83450 -590
rect 83510 -530 83620 -510
rect 83510 -590 83530 -530
rect 83600 -590 83620 -530
rect 83510 -610 83620 -590
rect 83680 -530 83790 -510
rect 83680 -590 83700 -530
rect 83770 -590 83790 -530
rect 83680 -610 83790 -590
rect 83850 -530 83960 -510
rect 83850 -590 83870 -530
rect 83940 -590 83960 -530
rect 83850 -610 83960 -590
rect 84020 -530 84130 -510
rect 84020 -590 84040 -530
rect 84110 -590 84130 -530
rect 84020 -610 84130 -590
rect 84190 -530 84300 -510
rect 84190 -590 84210 -530
rect 84280 -590 84300 -530
rect 84190 -610 84300 -590
rect 84360 -530 84470 -510
rect 84360 -590 84380 -530
rect 84450 -590 84470 -530
rect 84360 -610 84470 -590
rect 84530 -530 84640 -510
rect 84530 -590 84550 -530
rect 84620 -590 84640 -530
rect 84530 -610 84640 -590
rect 84700 -530 84810 -510
rect 84700 -590 84720 -530
rect 84790 -590 84810 -530
rect 84700 -610 84810 -590
rect 84870 -530 84980 -510
rect 84870 -590 84890 -530
rect 84960 -590 84980 -530
rect 84870 -610 84980 -590
rect 85040 -530 85150 -510
rect 85040 -590 85060 -530
rect 85130 -590 85150 -530
rect 85040 -610 85150 -590
rect 85210 -530 85320 -510
rect 85210 -590 85230 -530
rect 85300 -590 85320 -530
rect 85210 -610 85320 -590
rect 85380 -530 85490 -510
rect 85380 -590 85400 -530
rect 85470 -590 85490 -530
rect 85380 -610 85490 -590
rect 85550 -530 85660 -510
rect 85550 -590 85570 -530
rect 85640 -590 85660 -530
rect 85550 -610 85660 -590
rect 85720 -530 85830 -510
rect 85720 -590 85740 -530
rect 85810 -590 85830 -530
rect 85720 -610 85830 -590
rect 85890 -530 86000 -510
rect 85890 -590 85910 -530
rect 85980 -590 86000 -530
rect 85890 -610 86000 -590
rect 86060 -530 86170 -510
rect 86060 -590 86080 -530
rect 86150 -590 86170 -530
rect 86060 -610 86170 -590
rect 86230 -530 86340 -510
rect 86230 -590 86250 -530
rect 86320 -590 86340 -530
rect 86230 -610 86340 -590
rect 86400 -530 86510 -510
rect 86400 -590 86420 -530
rect 86490 -590 86510 -530
rect 86400 -610 86510 -590
rect 86570 -530 86680 -510
rect 86570 -590 86590 -530
rect 86660 -590 86680 -530
rect 86570 -610 86680 -590
rect 86740 -530 86850 -510
rect 86740 -590 86760 -530
rect 86830 -590 86850 -530
rect 86740 -610 86850 -590
rect 86910 -530 87020 -510
rect 86910 -590 86930 -530
rect 87000 -590 87020 -530
rect 86910 -610 87020 -590
rect 87080 -530 87190 -510
rect 87080 -590 87100 -530
rect 87170 -590 87190 -530
rect 87080 -610 87190 -590
rect 250 -650 280 -610
rect 420 -650 450 -610
rect 590 -650 620 -610
rect 760 -650 790 -610
rect 930 -650 960 -610
rect 1100 -650 1130 -610
rect 1270 -650 1300 -610
rect 1440 -650 1470 -610
rect 1610 -650 1640 -610
rect 1780 -650 1810 -610
rect 1950 -650 1980 -610
rect 2120 -650 2150 -610
rect 2290 -650 2320 -610
rect 2460 -650 2490 -610
rect 2630 -650 2660 -610
rect 2800 -650 2830 -610
rect 2970 -650 3000 -610
rect 3140 -650 3170 -610
rect 3310 -650 3340 -610
rect 3480 -650 3510 -610
rect 3650 -650 3680 -610
rect 3820 -650 3850 -610
rect 3990 -650 4020 -610
rect 4160 -650 4190 -610
rect 4330 -650 4360 -610
rect 4500 -650 4530 -610
rect 4670 -650 4700 -610
rect 4840 -650 4870 -610
rect 5010 -650 5040 -610
rect 5180 -650 5210 -610
rect 5350 -650 5380 -610
rect 5520 -650 5550 -610
rect 5690 -650 5720 -610
rect 5860 -650 5890 -610
rect 6030 -650 6060 -610
rect 6200 -650 6230 -610
rect 6370 -650 6400 -610
rect 6540 -650 6570 -610
rect 6710 -650 6740 -610
rect 6880 -650 6910 -610
rect 7050 -650 7080 -610
rect 7220 -650 7250 -610
rect 7390 -650 7420 -610
rect 7560 -650 7590 -610
rect 7730 -650 7760 -610
rect 7900 -650 7930 -610
rect 8070 -650 8100 -610
rect 8240 -650 8270 -610
rect 8410 -650 8440 -610
rect 8580 -650 8610 -610
rect 8750 -650 8780 -610
rect 8920 -650 8950 -610
rect 9090 -650 9120 -610
rect 9260 -650 9290 -610
rect 9430 -650 9460 -610
rect 9600 -650 9630 -610
rect 9770 -650 9800 -610
rect 9940 -650 9970 -610
rect 10110 -650 10140 -610
rect 10280 -650 10310 -610
rect 10450 -650 10480 -610
rect 10620 -650 10650 -610
rect 10790 -650 10820 -610
rect 10960 -650 10990 -610
rect 11130 -650 11160 -610
rect 11300 -650 11330 -610
rect 11470 -650 11500 -610
rect 11640 -650 11670 -610
rect 11810 -650 11840 -610
rect 11980 -650 12010 -610
rect 12150 -650 12180 -610
rect 12320 -650 12350 -610
rect 12490 -650 12520 -610
rect 12660 -650 12690 -610
rect 12830 -650 12860 -610
rect 13000 -650 13030 -610
rect 13170 -650 13200 -610
rect 13340 -650 13370 -610
rect 13510 -650 13540 -610
rect 13680 -650 13710 -610
rect 13850 -650 13880 -610
rect 14020 -650 14050 -610
rect 14190 -650 14220 -610
rect 14360 -650 14390 -610
rect 14530 -650 14560 -610
rect 14700 -650 14730 -610
rect 14870 -650 14900 -610
rect 15040 -650 15070 -610
rect 15210 -650 15240 -610
rect 15380 -650 15410 -610
rect 15550 -650 15580 -610
rect 15720 -650 15750 -610
rect 15890 -650 15920 -610
rect 16060 -650 16090 -610
rect 16230 -650 16260 -610
rect 16400 -650 16430 -610
rect 16570 -650 16600 -610
rect 16740 -650 16770 -610
rect 16910 -650 16940 -610
rect 17080 -650 17110 -610
rect 17250 -650 17280 -610
rect 17420 -650 17450 -610
rect 17590 -650 17620 -610
rect 17760 -650 17790 -610
rect 17930 -650 17960 -610
rect 18100 -650 18130 -610
rect 18270 -650 18300 -610
rect 18440 -650 18470 -610
rect 18610 -650 18640 -610
rect 18780 -650 18810 -610
rect 18950 -650 18980 -610
rect 19120 -650 19150 -610
rect 19290 -650 19320 -610
rect 19460 -650 19490 -610
rect 19630 -650 19660 -610
rect 19800 -650 19830 -610
rect 19970 -650 20000 -610
rect 20140 -650 20170 -610
rect 20310 -650 20340 -610
rect 20480 -650 20510 -610
rect 20650 -650 20680 -610
rect 20820 -650 20850 -610
rect 20990 -650 21020 -610
rect 21160 -650 21190 -610
rect 21330 -650 21360 -610
rect 21500 -650 21530 -610
rect 21670 -650 21700 -610
rect 21840 -650 21870 -610
rect 22010 -650 22040 -610
rect 22180 -650 22210 -610
rect 22350 -650 22380 -610
rect 22520 -650 22550 -610
rect 22690 -650 22720 -610
rect 22860 -650 22890 -610
rect 23030 -650 23060 -610
rect 23200 -650 23230 -610
rect 23370 -650 23400 -610
rect 23540 -650 23570 -610
rect 23710 -650 23740 -610
rect 23880 -650 23910 -610
rect 24050 -650 24080 -610
rect 24220 -650 24250 -610
rect 24390 -650 24420 -610
rect 24560 -650 24590 -610
rect 24730 -650 24760 -610
rect 24900 -650 24930 -610
rect 25070 -650 25100 -610
rect 25240 -650 25270 -610
rect 25410 -650 25440 -610
rect 25580 -650 25610 -610
rect 25750 -650 25780 -610
rect 25920 -650 25950 -610
rect 26090 -650 26120 -610
rect 26260 -650 26290 -610
rect 26430 -650 26460 -610
rect 26600 -650 26630 -610
rect 26770 -650 26800 -610
rect 26940 -650 26970 -610
rect 27110 -650 27140 -610
rect 27280 -650 27310 -610
rect 27450 -650 27480 -610
rect 27620 -650 27650 -610
rect 27790 -650 27820 -610
rect 27960 -650 27990 -610
rect 28130 -650 28160 -610
rect 28300 -650 28330 -610
rect 28470 -650 28500 -610
rect 28640 -650 28670 -610
rect 28810 -650 28840 -610
rect 28980 -650 29010 -610
rect 29150 -650 29180 -610
rect 29320 -650 29350 -610
rect 29490 -650 29520 -610
rect 29660 -650 29690 -610
rect 29830 -650 29860 -610
rect 30000 -650 30030 -610
rect 30170 -650 30200 -610
rect 30340 -650 30370 -610
rect 30510 -650 30540 -610
rect 30680 -650 30710 -610
rect 30850 -650 30880 -610
rect 31020 -650 31050 -610
rect 31190 -650 31220 -610
rect 31360 -650 31390 -610
rect 31530 -650 31560 -610
rect 31700 -650 31730 -610
rect 31870 -650 31900 -610
rect 32040 -650 32070 -610
rect 32210 -650 32240 -610
rect 32380 -650 32410 -610
rect 32550 -650 32580 -610
rect 32720 -650 32750 -610
rect 32890 -650 32920 -610
rect 33060 -650 33090 -610
rect 33230 -650 33260 -610
rect 33400 -650 33430 -610
rect 33570 -650 33600 -610
rect 33740 -650 33770 -610
rect 33910 -650 33940 -610
rect 34080 -650 34110 -610
rect 34250 -650 34280 -610
rect 34420 -650 34450 -610
rect 34590 -650 34620 -610
rect 34760 -650 34790 -610
rect 34930 -650 34960 -610
rect 35100 -650 35130 -610
rect 35270 -650 35300 -610
rect 35440 -650 35470 -610
rect 35610 -650 35640 -610
rect 35780 -650 35810 -610
rect 35950 -650 35980 -610
rect 36120 -650 36150 -610
rect 36290 -650 36320 -610
rect 36460 -650 36490 -610
rect 36630 -650 36660 -610
rect 36800 -650 36830 -610
rect 36970 -650 37000 -610
rect 37140 -650 37170 -610
rect 37310 -650 37340 -610
rect 37480 -650 37510 -610
rect 37650 -650 37680 -610
rect 37820 -650 37850 -610
rect 37990 -650 38020 -610
rect 38160 -650 38190 -610
rect 38330 -650 38360 -610
rect 38500 -650 38530 -610
rect 38670 -650 38700 -610
rect 38840 -650 38870 -610
rect 39010 -650 39040 -610
rect 39180 -650 39210 -610
rect 39350 -650 39380 -610
rect 39520 -650 39550 -610
rect 39690 -650 39720 -610
rect 39860 -650 39890 -610
rect 40030 -650 40060 -610
rect 40200 -650 40230 -610
rect 40370 -650 40400 -610
rect 40540 -650 40570 -610
rect 40710 -650 40740 -610
rect 40880 -650 40910 -610
rect 41050 -650 41080 -610
rect 41220 -650 41250 -610
rect 41390 -650 41420 -610
rect 41560 -650 41590 -610
rect 41730 -650 41760 -610
rect 41900 -650 41930 -610
rect 42070 -650 42100 -610
rect 42240 -650 42270 -610
rect 42410 -650 42440 -610
rect 42580 -650 42610 -610
rect 42750 -650 42780 -610
rect 42920 -650 42950 -610
rect 43090 -650 43120 -610
rect 43260 -650 43290 -610
rect 43430 -650 43460 -610
rect 43600 -650 43630 -610
rect 43770 -650 43800 -610
rect 43940 -650 43970 -610
rect 44110 -650 44140 -610
rect 44280 -650 44310 -610
rect 44450 -650 44480 -610
rect 44620 -650 44650 -610
rect 44790 -650 44820 -610
rect 44960 -650 44990 -610
rect 45130 -650 45160 -610
rect 45300 -650 45330 -610
rect 45470 -650 45500 -610
rect 45640 -650 45670 -610
rect 45810 -650 45840 -610
rect 45980 -650 46010 -610
rect 46150 -650 46180 -610
rect 46320 -650 46350 -610
rect 46490 -650 46520 -610
rect 46660 -650 46690 -610
rect 46830 -650 46860 -610
rect 47000 -650 47030 -610
rect 47170 -650 47200 -610
rect 47340 -650 47370 -610
rect 47510 -650 47540 -610
rect 47680 -650 47710 -610
rect 47850 -650 47880 -610
rect 48020 -650 48050 -610
rect 48190 -650 48220 -610
rect 48360 -650 48390 -610
rect 48530 -650 48560 -610
rect 48700 -650 48730 -610
rect 48870 -650 48900 -610
rect 49040 -650 49070 -610
rect 49210 -650 49240 -610
rect 49380 -650 49410 -610
rect 49550 -650 49580 -610
rect 49720 -650 49750 -610
rect 49890 -650 49920 -610
rect 50060 -650 50090 -610
rect 50230 -650 50260 -610
rect 50400 -650 50430 -610
rect 50570 -650 50600 -610
rect 50740 -650 50770 -610
rect 50910 -650 50940 -610
rect 51080 -650 51110 -610
rect 51250 -650 51280 -610
rect 51420 -650 51450 -610
rect 51590 -650 51620 -610
rect 51760 -650 51790 -610
rect 51930 -650 51960 -610
rect 52100 -650 52130 -610
rect 52270 -650 52300 -610
rect 52440 -650 52470 -610
rect 52610 -650 52640 -610
rect 52780 -650 52810 -610
rect 52950 -650 52980 -610
rect 53120 -650 53150 -610
rect 53290 -650 53320 -610
rect 53460 -650 53490 -610
rect 53630 -650 53660 -610
rect 53800 -650 53830 -610
rect 53970 -650 54000 -610
rect 54140 -650 54170 -610
rect 54310 -650 54340 -610
rect 54480 -650 54510 -610
rect 54650 -650 54680 -610
rect 54820 -650 54850 -610
rect 54990 -650 55020 -610
rect 55160 -650 55190 -610
rect 55330 -650 55360 -610
rect 55500 -650 55530 -610
rect 55670 -650 55700 -610
rect 55840 -650 55870 -610
rect 56010 -650 56040 -610
rect 56180 -650 56210 -610
rect 56350 -650 56380 -610
rect 56520 -650 56550 -610
rect 56690 -650 56720 -610
rect 56860 -650 56890 -610
rect 57030 -650 57060 -610
rect 57200 -650 57230 -610
rect 57370 -650 57400 -610
rect 57540 -650 57570 -610
rect 57710 -650 57740 -610
rect 57880 -650 57910 -610
rect 58050 -650 58080 -610
rect 58220 -650 58250 -610
rect 58390 -650 58420 -610
rect 58560 -650 58590 -610
rect 58730 -650 58760 -610
rect 58900 -650 58930 -610
rect 59070 -650 59100 -610
rect 59240 -650 59270 -610
rect 59410 -650 59440 -610
rect 59580 -650 59610 -610
rect 59750 -650 59780 -610
rect 59920 -650 59950 -610
rect 60090 -650 60120 -610
rect 60260 -650 60290 -610
rect 60430 -650 60460 -610
rect 60600 -650 60630 -610
rect 60770 -650 60800 -610
rect 60940 -650 60970 -610
rect 61110 -650 61140 -610
rect 61280 -650 61310 -610
rect 61450 -650 61480 -610
rect 61620 -650 61650 -610
rect 61790 -650 61820 -610
rect 61960 -650 61990 -610
rect 62130 -650 62160 -610
rect 62300 -650 62330 -610
rect 62470 -650 62500 -610
rect 62640 -650 62670 -610
rect 62810 -650 62840 -610
rect 62980 -650 63010 -610
rect 63150 -650 63180 -610
rect 63320 -650 63350 -610
rect 63490 -650 63520 -610
rect 63660 -650 63690 -610
rect 63830 -650 63860 -610
rect 64000 -650 64030 -610
rect 64170 -650 64200 -610
rect 64340 -650 64370 -610
rect 64510 -650 64540 -610
rect 64680 -650 64710 -610
rect 64850 -650 64880 -610
rect 65020 -650 65050 -610
rect 65190 -650 65220 -610
rect 65360 -650 65390 -610
rect 65530 -650 65560 -610
rect 65700 -650 65730 -610
rect 65870 -650 65900 -610
rect 66040 -650 66070 -610
rect 66210 -650 66240 -610
rect 66380 -650 66410 -610
rect 66550 -650 66580 -610
rect 66720 -650 66750 -610
rect 66890 -650 66920 -610
rect 67060 -650 67090 -610
rect 67230 -650 67260 -610
rect 67400 -650 67430 -610
rect 67570 -650 67600 -610
rect 67740 -650 67770 -610
rect 67910 -650 67940 -610
rect 68080 -650 68110 -610
rect 68250 -650 68280 -610
rect 68420 -650 68450 -610
rect 68590 -650 68620 -610
rect 68760 -650 68790 -610
rect 68930 -650 68960 -610
rect 69100 -650 69130 -610
rect 69270 -650 69300 -610
rect 69440 -650 69470 -610
rect 69610 -650 69640 -610
rect 69780 -650 69810 -610
rect 69950 -650 69980 -610
rect 70120 -650 70150 -610
rect 70290 -650 70320 -610
rect 70460 -650 70490 -610
rect 70630 -650 70660 -610
rect 70800 -650 70830 -610
rect 70970 -650 71000 -610
rect 71140 -650 71170 -610
rect 71310 -650 71340 -610
rect 71480 -650 71510 -610
rect 71650 -650 71680 -610
rect 71820 -650 71850 -610
rect 71990 -650 72020 -610
rect 72160 -650 72190 -610
rect 72330 -650 72360 -610
rect 72500 -650 72530 -610
rect 72670 -650 72700 -610
rect 72840 -650 72870 -610
rect 73010 -650 73040 -610
rect 73180 -650 73210 -610
rect 73350 -650 73380 -610
rect 73520 -650 73550 -610
rect 73690 -650 73720 -610
rect 73860 -650 73890 -610
rect 74030 -650 74060 -610
rect 74200 -650 74230 -610
rect 74370 -650 74400 -610
rect 74540 -650 74570 -610
rect 74710 -650 74740 -610
rect 74880 -650 74910 -610
rect 75050 -650 75080 -610
rect 75220 -650 75250 -610
rect 75390 -650 75420 -610
rect 75560 -650 75590 -610
rect 75730 -650 75760 -610
rect 75900 -650 75930 -610
rect 76070 -650 76100 -610
rect 76240 -650 76270 -610
rect 76410 -650 76440 -610
rect 76580 -650 76610 -610
rect 76750 -650 76780 -610
rect 76920 -650 76950 -610
rect 77090 -650 77120 -610
rect 77260 -650 77290 -610
rect 77430 -650 77460 -610
rect 77600 -650 77630 -610
rect 77770 -650 77800 -610
rect 77940 -650 77970 -610
rect 78110 -650 78140 -610
rect 78280 -650 78310 -610
rect 78450 -650 78480 -610
rect 78620 -650 78650 -610
rect 78790 -650 78820 -610
rect 78960 -650 78990 -610
rect 79130 -650 79160 -610
rect 79300 -650 79330 -610
rect 79470 -650 79500 -610
rect 79640 -650 79670 -610
rect 79810 -650 79840 -610
rect 79980 -650 80010 -610
rect 80150 -650 80180 -610
rect 80320 -650 80350 -610
rect 80490 -650 80520 -610
rect 80660 -650 80690 -610
rect 80830 -650 80860 -610
rect 81000 -650 81030 -610
rect 81170 -650 81200 -610
rect 81340 -650 81370 -610
rect 81510 -650 81540 -610
rect 81680 -650 81710 -610
rect 81850 -650 81880 -610
rect 82020 -650 82050 -610
rect 82190 -650 82220 -610
rect 82360 -650 82390 -610
rect 82530 -650 82560 -610
rect 82700 -650 82730 -610
rect 82870 -650 82900 -610
rect 83040 -650 83070 -610
rect 83210 -650 83240 -610
rect 83380 -650 83410 -610
rect 83550 -650 83580 -610
rect 83720 -650 83750 -610
rect 83890 -650 83920 -610
rect 84060 -650 84090 -610
rect 84230 -650 84260 -610
rect 84400 -650 84430 -610
rect 84570 -650 84600 -610
rect 84740 -650 84770 -610
rect 84910 -650 84940 -610
rect 85080 -650 85110 -610
rect 85250 -650 85280 -610
rect 85420 -650 85450 -610
rect 85590 -650 85620 -610
rect 85760 -650 85790 -610
rect 85930 -650 85960 -610
rect 86100 -650 86130 -610
rect 86270 -650 86300 -610
rect 86440 -650 86470 -610
rect 86610 -650 86640 -610
rect 86780 -650 86810 -610
rect 86950 -650 86980 -610
rect 87120 -650 87150 -610
rect 250 -980 280 -850
rect 420 -980 450 -850
rect 590 -980 620 -850
rect 760 -980 790 -850
rect 930 -980 960 -850
rect 1100 -980 1130 -850
rect 1270 -980 1300 -850
rect 1440 -980 1470 -850
rect 1610 -980 1640 -850
rect 1780 -980 1810 -850
rect 1950 -980 1980 -850
rect 2120 -980 2150 -850
rect 2290 -980 2320 -850
rect 2460 -980 2490 -850
rect 2630 -980 2660 -850
rect 2800 -980 2830 -850
rect 2970 -980 3000 -850
rect 3140 -980 3170 -850
rect 3310 -980 3340 -850
rect 3480 -980 3510 -850
rect 3650 -980 3680 -850
rect 3820 -980 3850 -850
rect 3990 -980 4020 -850
rect 4160 -980 4190 -850
rect 4330 -980 4360 -850
rect 4500 -980 4530 -850
rect 4670 -980 4700 -850
rect 4840 -980 4870 -850
rect 5010 -980 5040 -850
rect 5180 -980 5210 -850
rect 5350 -980 5380 -850
rect 5520 -980 5550 -850
rect 5690 -980 5720 -850
rect 5860 -980 5890 -850
rect 6030 -980 6060 -850
rect 6200 -980 6230 -850
rect 6370 -980 6400 -850
rect 6540 -980 6570 -850
rect 6710 -980 6740 -850
rect 6880 -980 6910 -850
rect 7050 -980 7080 -850
rect 7220 -980 7250 -850
rect 7390 -980 7420 -850
rect 7560 -980 7590 -850
rect 7730 -980 7760 -850
rect 7900 -980 7930 -850
rect 8070 -980 8100 -850
rect 8240 -980 8270 -850
rect 8410 -980 8440 -850
rect 8580 -980 8610 -850
rect 8750 -980 8780 -850
rect 8920 -980 8950 -850
rect 9090 -980 9120 -850
rect 9260 -980 9290 -850
rect 9430 -980 9460 -850
rect 9600 -980 9630 -850
rect 9770 -980 9800 -850
rect 9940 -980 9970 -850
rect 10110 -980 10140 -850
rect 10280 -980 10310 -850
rect 10450 -980 10480 -850
rect 10620 -980 10650 -850
rect 10790 -980 10820 -850
rect 10960 -980 10990 -850
rect 11130 -980 11160 -850
rect 11300 -980 11330 -850
rect 11470 -980 11500 -850
rect 11640 -980 11670 -850
rect 11810 -980 11840 -850
rect 11980 -980 12010 -850
rect 12150 -980 12180 -850
rect 12320 -980 12350 -850
rect 12490 -980 12520 -850
rect 12660 -980 12690 -850
rect 12830 -980 12860 -850
rect 13000 -980 13030 -850
rect 13170 -980 13200 -850
rect 13340 -980 13370 -850
rect 13510 -980 13540 -850
rect 13680 -980 13710 -850
rect 13850 -980 13880 -850
rect 14020 -980 14050 -850
rect 14190 -980 14220 -850
rect 14360 -980 14390 -850
rect 14530 -980 14560 -850
rect 14700 -980 14730 -850
rect 14870 -980 14900 -850
rect 15040 -980 15070 -850
rect 15210 -980 15240 -850
rect 15380 -980 15410 -850
rect 15550 -980 15580 -850
rect 15720 -980 15750 -850
rect 15890 -980 15920 -850
rect 16060 -980 16090 -850
rect 16230 -980 16260 -850
rect 16400 -980 16430 -850
rect 16570 -980 16600 -850
rect 16740 -980 16770 -850
rect 16910 -980 16940 -850
rect 17080 -980 17110 -850
rect 17250 -980 17280 -850
rect 17420 -980 17450 -850
rect 17590 -980 17620 -850
rect 17760 -980 17790 -850
rect 17930 -980 17960 -850
rect 18100 -980 18130 -850
rect 18270 -980 18300 -850
rect 18440 -980 18470 -850
rect 18610 -980 18640 -850
rect 18780 -980 18810 -850
rect 18950 -980 18980 -850
rect 19120 -980 19150 -850
rect 19290 -980 19320 -850
rect 19460 -980 19490 -850
rect 19630 -980 19660 -850
rect 19800 -980 19830 -850
rect 19970 -980 20000 -850
rect 20140 -980 20170 -850
rect 20310 -980 20340 -850
rect 20480 -980 20510 -850
rect 20650 -980 20680 -850
rect 20820 -980 20850 -850
rect 20990 -980 21020 -850
rect 21160 -980 21190 -850
rect 21330 -980 21360 -850
rect 21500 -980 21530 -850
rect 21670 -980 21700 -850
rect 21840 -980 21870 -850
rect 22010 -980 22040 -850
rect 22180 -980 22210 -850
rect 22350 -980 22380 -850
rect 22520 -980 22550 -850
rect 22690 -980 22720 -850
rect 22860 -980 22890 -850
rect 23030 -980 23060 -850
rect 23200 -980 23230 -850
rect 23370 -980 23400 -850
rect 23540 -980 23570 -850
rect 23710 -980 23740 -850
rect 23880 -980 23910 -850
rect 24050 -980 24080 -850
rect 24220 -980 24250 -850
rect 24390 -980 24420 -850
rect 24560 -980 24590 -850
rect 24730 -980 24760 -850
rect 24900 -980 24930 -850
rect 25070 -980 25100 -850
rect 25240 -980 25270 -850
rect 25410 -980 25440 -850
rect 25580 -980 25610 -850
rect 25750 -980 25780 -850
rect 25920 -980 25950 -850
rect 26090 -980 26120 -850
rect 26260 -980 26290 -850
rect 26430 -980 26460 -850
rect 26600 -980 26630 -850
rect 26770 -980 26800 -850
rect 26940 -980 26970 -850
rect 27110 -980 27140 -850
rect 27280 -980 27310 -850
rect 27450 -980 27480 -850
rect 27620 -980 27650 -850
rect 27790 -980 27820 -850
rect 27960 -980 27990 -850
rect 28130 -980 28160 -850
rect 28300 -980 28330 -850
rect 28470 -980 28500 -850
rect 28640 -980 28670 -850
rect 28810 -980 28840 -850
rect 28980 -980 29010 -850
rect 29150 -980 29180 -850
rect 29320 -980 29350 -850
rect 29490 -980 29520 -850
rect 29660 -980 29690 -850
rect 29830 -980 29860 -850
rect 30000 -980 30030 -850
rect 30170 -980 30200 -850
rect 30340 -980 30370 -850
rect 30510 -980 30540 -850
rect 30680 -980 30710 -850
rect 30850 -980 30880 -850
rect 31020 -980 31050 -850
rect 31190 -980 31220 -850
rect 31360 -980 31390 -850
rect 31530 -980 31560 -850
rect 31700 -980 31730 -850
rect 31870 -980 31900 -850
rect 32040 -980 32070 -850
rect 32210 -980 32240 -850
rect 32380 -980 32410 -850
rect 32550 -980 32580 -850
rect 32720 -980 32750 -850
rect 32890 -980 32920 -850
rect 33060 -980 33090 -850
rect 33230 -980 33260 -850
rect 33400 -980 33430 -850
rect 33570 -980 33600 -850
rect 33740 -980 33770 -850
rect 33910 -980 33940 -850
rect 34080 -980 34110 -850
rect 34250 -980 34280 -850
rect 34420 -980 34450 -850
rect 34590 -980 34620 -850
rect 34760 -980 34790 -850
rect 34930 -980 34960 -850
rect 35100 -980 35130 -850
rect 35270 -980 35300 -850
rect 35440 -980 35470 -850
rect 35610 -980 35640 -850
rect 35780 -980 35810 -850
rect 35950 -980 35980 -850
rect 36120 -980 36150 -850
rect 36290 -980 36320 -850
rect 36460 -980 36490 -850
rect 36630 -980 36660 -850
rect 36800 -980 36830 -850
rect 36970 -980 37000 -850
rect 37140 -980 37170 -850
rect 37310 -980 37340 -850
rect 37480 -980 37510 -850
rect 37650 -980 37680 -850
rect 37820 -980 37850 -850
rect 37990 -980 38020 -850
rect 38160 -980 38190 -850
rect 38330 -980 38360 -850
rect 38500 -980 38530 -850
rect 38670 -980 38700 -850
rect 38840 -980 38870 -850
rect 39010 -980 39040 -850
rect 39180 -980 39210 -850
rect 39350 -980 39380 -850
rect 39520 -980 39550 -850
rect 39690 -980 39720 -850
rect 39860 -980 39890 -850
rect 40030 -980 40060 -850
rect 40200 -980 40230 -850
rect 40370 -980 40400 -850
rect 40540 -980 40570 -850
rect 40710 -980 40740 -850
rect 40880 -980 40910 -850
rect 41050 -980 41080 -850
rect 41220 -980 41250 -850
rect 41390 -980 41420 -850
rect 41560 -980 41590 -850
rect 41730 -980 41760 -850
rect 41900 -980 41930 -850
rect 42070 -980 42100 -850
rect 42240 -980 42270 -850
rect 42410 -980 42440 -850
rect 42580 -980 42610 -850
rect 42750 -980 42780 -850
rect 42920 -980 42950 -850
rect 43090 -980 43120 -850
rect 43260 -980 43290 -850
rect 43430 -980 43460 -850
rect 43600 -980 43630 -850
rect 43770 -980 43800 -850
rect 43940 -980 43970 -850
rect 44110 -980 44140 -850
rect 44280 -980 44310 -850
rect 44450 -980 44480 -850
rect 44620 -980 44650 -850
rect 44790 -980 44820 -850
rect 44960 -980 44990 -850
rect 45130 -980 45160 -850
rect 45300 -980 45330 -850
rect 45470 -980 45500 -850
rect 45640 -980 45670 -850
rect 45810 -980 45840 -850
rect 45980 -980 46010 -850
rect 46150 -980 46180 -850
rect 46320 -980 46350 -850
rect 46490 -980 46520 -850
rect 46660 -980 46690 -850
rect 46830 -980 46860 -850
rect 47000 -980 47030 -850
rect 47170 -980 47200 -850
rect 47340 -980 47370 -850
rect 47510 -980 47540 -850
rect 47680 -980 47710 -850
rect 47850 -980 47880 -850
rect 48020 -980 48050 -850
rect 48190 -980 48220 -850
rect 48360 -980 48390 -850
rect 48530 -980 48560 -850
rect 48700 -980 48730 -850
rect 48870 -980 48900 -850
rect 49040 -980 49070 -850
rect 49210 -980 49240 -850
rect 49380 -980 49410 -850
rect 49550 -980 49580 -850
rect 49720 -980 49750 -850
rect 49890 -980 49920 -850
rect 50060 -980 50090 -850
rect 50230 -980 50260 -850
rect 50400 -980 50430 -850
rect 50570 -980 50600 -850
rect 50740 -980 50770 -850
rect 50910 -980 50940 -850
rect 51080 -980 51110 -850
rect 51250 -980 51280 -850
rect 51420 -980 51450 -850
rect 51590 -980 51620 -850
rect 51760 -980 51790 -850
rect 51930 -980 51960 -850
rect 52100 -980 52130 -850
rect 52270 -980 52300 -850
rect 52440 -980 52470 -850
rect 52610 -980 52640 -850
rect 52780 -980 52810 -850
rect 52950 -980 52980 -850
rect 53120 -980 53150 -850
rect 53290 -980 53320 -850
rect 53460 -980 53490 -850
rect 53630 -980 53660 -850
rect 53800 -980 53830 -850
rect 53970 -980 54000 -850
rect 54140 -980 54170 -850
rect 54310 -980 54340 -850
rect 54480 -980 54510 -850
rect 54650 -980 54680 -850
rect 54820 -980 54850 -850
rect 54990 -980 55020 -850
rect 55160 -980 55190 -850
rect 55330 -980 55360 -850
rect 55500 -980 55530 -850
rect 55670 -980 55700 -850
rect 55840 -980 55870 -850
rect 56010 -980 56040 -850
rect 56180 -980 56210 -850
rect 56350 -980 56380 -850
rect 56520 -980 56550 -850
rect 56690 -980 56720 -850
rect 56860 -980 56890 -850
rect 57030 -980 57060 -850
rect 57200 -980 57230 -850
rect 57370 -980 57400 -850
rect 57540 -980 57570 -850
rect 57710 -980 57740 -850
rect 57880 -980 57910 -850
rect 58050 -980 58080 -850
rect 58220 -980 58250 -850
rect 58390 -980 58420 -850
rect 58560 -980 58590 -850
rect 58730 -980 58760 -850
rect 58900 -980 58930 -850
rect 59070 -980 59100 -850
rect 59240 -980 59270 -850
rect 59410 -980 59440 -850
rect 59580 -980 59610 -850
rect 59750 -980 59780 -850
rect 59920 -980 59950 -850
rect 60090 -980 60120 -850
rect 60260 -980 60290 -850
rect 60430 -980 60460 -850
rect 60600 -980 60630 -850
rect 60770 -980 60800 -850
rect 60940 -980 60970 -850
rect 61110 -980 61140 -850
rect 61280 -980 61310 -850
rect 61450 -980 61480 -850
rect 61620 -980 61650 -850
rect 61790 -980 61820 -850
rect 61960 -980 61990 -850
rect 62130 -980 62160 -850
rect 62300 -980 62330 -850
rect 62470 -980 62500 -850
rect 62640 -980 62670 -850
rect 62810 -980 62840 -850
rect 62980 -980 63010 -850
rect 63150 -980 63180 -850
rect 63320 -980 63350 -850
rect 63490 -980 63520 -850
rect 63660 -980 63690 -850
rect 63830 -980 63860 -850
rect 64000 -980 64030 -850
rect 64170 -980 64200 -850
rect 64340 -980 64370 -850
rect 64510 -980 64540 -850
rect 64680 -980 64710 -850
rect 64850 -980 64880 -850
rect 65020 -980 65050 -850
rect 65190 -980 65220 -850
rect 65360 -980 65390 -850
rect 65530 -980 65560 -850
rect 65700 -980 65730 -850
rect 65870 -980 65900 -850
rect 66040 -980 66070 -850
rect 66210 -980 66240 -850
rect 66380 -980 66410 -850
rect 66550 -980 66580 -850
rect 66720 -980 66750 -850
rect 66890 -980 66920 -850
rect 67060 -980 67090 -850
rect 67230 -980 67260 -850
rect 67400 -980 67430 -850
rect 67570 -980 67600 -850
rect 67740 -980 67770 -850
rect 67910 -980 67940 -850
rect 68080 -980 68110 -850
rect 68250 -980 68280 -850
rect 68420 -980 68450 -850
rect 68590 -980 68620 -850
rect 68760 -980 68790 -850
rect 68930 -980 68960 -850
rect 69100 -980 69130 -850
rect 69270 -980 69300 -850
rect 69440 -980 69470 -850
rect 69610 -980 69640 -850
rect 69780 -980 69810 -850
rect 69950 -980 69980 -850
rect 70120 -980 70150 -850
rect 70290 -980 70320 -850
rect 70460 -980 70490 -850
rect 70630 -980 70660 -850
rect 70800 -980 70830 -850
rect 70970 -980 71000 -850
rect 71140 -980 71170 -850
rect 71310 -980 71340 -850
rect 71480 -980 71510 -850
rect 71650 -980 71680 -850
rect 71820 -980 71850 -850
rect 71990 -980 72020 -850
rect 72160 -980 72190 -850
rect 72330 -980 72360 -850
rect 72500 -980 72530 -850
rect 72670 -980 72700 -850
rect 72840 -980 72870 -850
rect 73010 -980 73040 -850
rect 73180 -980 73210 -850
rect 73350 -980 73380 -850
rect 73520 -980 73550 -850
rect 73690 -980 73720 -850
rect 73860 -980 73890 -850
rect 74030 -980 74060 -850
rect 74200 -980 74230 -850
rect 74370 -980 74400 -850
rect 74540 -980 74570 -850
rect 74710 -980 74740 -850
rect 74880 -980 74910 -850
rect 75050 -980 75080 -850
rect 75220 -980 75250 -850
rect 75390 -980 75420 -850
rect 75560 -980 75590 -850
rect 75730 -980 75760 -850
rect 75900 -980 75930 -850
rect 76070 -980 76100 -850
rect 76240 -980 76270 -850
rect 76410 -980 76440 -850
rect 76580 -980 76610 -850
rect 76750 -980 76780 -850
rect 76920 -980 76950 -850
rect 77090 -980 77120 -850
rect 77260 -980 77290 -850
rect 77430 -980 77460 -850
rect 77600 -980 77630 -850
rect 77770 -980 77800 -850
rect 77940 -980 77970 -850
rect 78110 -980 78140 -850
rect 78280 -980 78310 -850
rect 78450 -980 78480 -850
rect 78620 -980 78650 -850
rect 78790 -980 78820 -850
rect 78960 -980 78990 -850
rect 79130 -980 79160 -850
rect 79300 -980 79330 -850
rect 79470 -980 79500 -850
rect 79640 -980 79670 -850
rect 79810 -980 79840 -850
rect 79980 -980 80010 -850
rect 80150 -980 80180 -850
rect 80320 -980 80350 -850
rect 80490 -980 80520 -850
rect 80660 -980 80690 -850
rect 80830 -980 80860 -850
rect 81000 -980 81030 -850
rect 81170 -980 81200 -850
rect 81340 -980 81370 -850
rect 81510 -980 81540 -850
rect 81680 -980 81710 -850
rect 81850 -980 81880 -850
rect 82020 -980 82050 -850
rect 82190 -980 82220 -850
rect 82360 -980 82390 -850
rect 82530 -980 82560 -850
rect 82700 -980 82730 -850
rect 82870 -980 82900 -850
rect 83040 -980 83070 -850
rect 83210 -980 83240 -850
rect 83380 -980 83410 -850
rect 83550 -980 83580 -850
rect 83720 -980 83750 -850
rect 83890 -980 83920 -850
rect 84060 -980 84090 -850
rect 84230 -980 84260 -850
rect 84400 -980 84430 -850
rect 84570 -980 84600 -850
rect 84740 -980 84770 -850
rect 84910 -980 84940 -850
rect 85080 -980 85110 -850
rect 85250 -980 85280 -850
rect 85420 -980 85450 -850
rect 85590 -980 85620 -850
rect 85760 -980 85790 -850
rect 85930 -980 85960 -850
rect 86100 -980 86130 -850
rect 86270 -980 86300 -850
rect 86440 -980 86470 -850
rect 86610 -980 86640 -850
rect 86780 -980 86810 -850
rect 86950 -980 86980 -850
rect 87120 -980 87150 -850
rect 250 -1410 280 -1380
rect 420 -1410 450 -1380
rect 590 -1410 620 -1380
rect 760 -1410 790 -1380
rect 930 -1410 960 -1380
rect 1100 -1410 1130 -1380
rect 1270 -1410 1300 -1380
rect 1440 -1410 1470 -1380
rect 1610 -1410 1640 -1380
rect 1780 -1410 1810 -1380
rect 1950 -1410 1980 -1380
rect 2120 -1410 2150 -1380
rect 2290 -1410 2320 -1380
rect 2460 -1410 2490 -1380
rect 2630 -1410 2660 -1380
rect 2800 -1410 2830 -1380
rect 2970 -1410 3000 -1380
rect 3140 -1410 3170 -1380
rect 3310 -1410 3340 -1380
rect 3480 -1410 3510 -1380
rect 3650 -1410 3680 -1380
rect 3820 -1410 3850 -1380
rect 3990 -1410 4020 -1380
rect 4160 -1410 4190 -1380
rect 4330 -1410 4360 -1380
rect 4500 -1410 4530 -1380
rect 4670 -1410 4700 -1380
rect 4840 -1410 4870 -1380
rect 5010 -1410 5040 -1380
rect 5180 -1410 5210 -1380
rect 5350 -1410 5380 -1380
rect 5520 -1410 5550 -1380
rect 5690 -1410 5720 -1380
rect 5860 -1410 5890 -1380
rect 6030 -1410 6060 -1380
rect 6200 -1410 6230 -1380
rect 6370 -1410 6400 -1380
rect 6540 -1410 6570 -1380
rect 6710 -1410 6740 -1380
rect 6880 -1410 6910 -1380
rect 7050 -1410 7080 -1380
rect 7220 -1410 7250 -1380
rect 7390 -1410 7420 -1380
rect 7560 -1410 7590 -1380
rect 7730 -1410 7760 -1380
rect 7900 -1410 7930 -1380
rect 8070 -1410 8100 -1380
rect 8240 -1410 8270 -1380
rect 8410 -1410 8440 -1380
rect 8580 -1410 8610 -1380
rect 8750 -1410 8780 -1380
rect 8920 -1410 8950 -1380
rect 9090 -1410 9120 -1380
rect 9260 -1410 9290 -1380
rect 9430 -1410 9460 -1380
rect 9600 -1410 9630 -1380
rect 9770 -1410 9800 -1380
rect 9940 -1410 9970 -1380
rect 10110 -1410 10140 -1380
rect 10280 -1410 10310 -1380
rect 10450 -1410 10480 -1380
rect 10620 -1410 10650 -1380
rect 10790 -1410 10820 -1380
rect 10960 -1410 10990 -1380
rect 11130 -1410 11160 -1380
rect 11300 -1410 11330 -1380
rect 11470 -1410 11500 -1380
rect 11640 -1410 11670 -1380
rect 11810 -1410 11840 -1380
rect 11980 -1410 12010 -1380
rect 12150 -1410 12180 -1380
rect 12320 -1410 12350 -1380
rect 12490 -1410 12520 -1380
rect 12660 -1410 12690 -1380
rect 12830 -1410 12860 -1380
rect 13000 -1410 13030 -1380
rect 13170 -1410 13200 -1380
rect 13340 -1410 13370 -1380
rect 13510 -1410 13540 -1380
rect 13680 -1410 13710 -1380
rect 13850 -1410 13880 -1380
rect 14020 -1410 14050 -1380
rect 14190 -1410 14220 -1380
rect 14360 -1410 14390 -1380
rect 14530 -1410 14560 -1380
rect 14700 -1410 14730 -1380
rect 14870 -1410 14900 -1380
rect 15040 -1410 15070 -1380
rect 15210 -1410 15240 -1380
rect 15380 -1410 15410 -1380
rect 15550 -1410 15580 -1380
rect 15720 -1410 15750 -1380
rect 15890 -1410 15920 -1380
rect 16060 -1410 16090 -1380
rect 16230 -1410 16260 -1380
rect 16400 -1410 16430 -1380
rect 16570 -1410 16600 -1380
rect 16740 -1410 16770 -1380
rect 16910 -1410 16940 -1380
rect 17080 -1410 17110 -1380
rect 17250 -1410 17280 -1380
rect 17420 -1410 17450 -1380
rect 17590 -1410 17620 -1380
rect 17760 -1410 17790 -1380
rect 17930 -1410 17960 -1380
rect 18100 -1410 18130 -1380
rect 18270 -1410 18300 -1380
rect 18440 -1410 18470 -1380
rect 18610 -1410 18640 -1380
rect 18780 -1410 18810 -1380
rect 18950 -1410 18980 -1380
rect 19120 -1410 19150 -1380
rect 19290 -1410 19320 -1380
rect 19460 -1410 19490 -1380
rect 19630 -1410 19660 -1380
rect 19800 -1410 19830 -1380
rect 19970 -1410 20000 -1380
rect 20140 -1410 20170 -1380
rect 20310 -1410 20340 -1380
rect 20480 -1410 20510 -1380
rect 20650 -1410 20680 -1380
rect 20820 -1410 20850 -1380
rect 20990 -1410 21020 -1380
rect 21160 -1410 21190 -1380
rect 21330 -1410 21360 -1380
rect 21500 -1410 21530 -1380
rect 21670 -1410 21700 -1380
rect 21840 -1410 21870 -1380
rect 22010 -1410 22040 -1380
rect 22180 -1410 22210 -1380
rect 22350 -1410 22380 -1380
rect 22520 -1410 22550 -1380
rect 22690 -1410 22720 -1380
rect 22860 -1410 22890 -1380
rect 23030 -1410 23060 -1380
rect 23200 -1410 23230 -1380
rect 23370 -1410 23400 -1380
rect 23540 -1410 23570 -1380
rect 23710 -1410 23740 -1380
rect 23880 -1410 23910 -1380
rect 24050 -1410 24080 -1380
rect 24220 -1410 24250 -1380
rect 24390 -1410 24420 -1380
rect 24560 -1410 24590 -1380
rect 24730 -1410 24760 -1380
rect 24900 -1410 24930 -1380
rect 25070 -1410 25100 -1380
rect 25240 -1410 25270 -1380
rect 25410 -1410 25440 -1380
rect 25580 -1410 25610 -1380
rect 25750 -1410 25780 -1380
rect 25920 -1410 25950 -1380
rect 26090 -1410 26120 -1380
rect 26260 -1410 26290 -1380
rect 26430 -1410 26460 -1380
rect 26600 -1410 26630 -1380
rect 26770 -1410 26800 -1380
rect 26940 -1410 26970 -1380
rect 27110 -1410 27140 -1380
rect 27280 -1410 27310 -1380
rect 27450 -1410 27480 -1380
rect 27620 -1410 27650 -1380
rect 27790 -1410 27820 -1380
rect 27960 -1410 27990 -1380
rect 28130 -1410 28160 -1380
rect 28300 -1410 28330 -1380
rect 28470 -1410 28500 -1380
rect 28640 -1410 28670 -1380
rect 28810 -1410 28840 -1380
rect 28980 -1410 29010 -1380
rect 29150 -1410 29180 -1380
rect 29320 -1410 29350 -1380
rect 29490 -1410 29520 -1380
rect 29660 -1410 29690 -1380
rect 29830 -1410 29860 -1380
rect 30000 -1410 30030 -1380
rect 30170 -1410 30200 -1380
rect 30340 -1410 30370 -1380
rect 30510 -1410 30540 -1380
rect 30680 -1410 30710 -1380
rect 30850 -1410 30880 -1380
rect 31020 -1410 31050 -1380
rect 31190 -1410 31220 -1380
rect 31360 -1410 31390 -1380
rect 31530 -1410 31560 -1380
rect 31700 -1410 31730 -1380
rect 31870 -1410 31900 -1380
rect 32040 -1410 32070 -1380
rect 32210 -1410 32240 -1380
rect 32380 -1410 32410 -1380
rect 32550 -1410 32580 -1380
rect 32720 -1410 32750 -1380
rect 32890 -1410 32920 -1380
rect 33060 -1410 33090 -1380
rect 33230 -1410 33260 -1380
rect 33400 -1410 33430 -1380
rect 33570 -1410 33600 -1380
rect 33740 -1410 33770 -1380
rect 33910 -1410 33940 -1380
rect 34080 -1410 34110 -1380
rect 34250 -1410 34280 -1380
rect 34420 -1410 34450 -1380
rect 34590 -1410 34620 -1380
rect 34760 -1410 34790 -1380
rect 34930 -1410 34960 -1380
rect 35100 -1410 35130 -1380
rect 35270 -1410 35300 -1380
rect 35440 -1410 35470 -1380
rect 35610 -1410 35640 -1380
rect 35780 -1410 35810 -1380
rect 35950 -1410 35980 -1380
rect 36120 -1410 36150 -1380
rect 36290 -1410 36320 -1380
rect 36460 -1410 36490 -1380
rect 36630 -1410 36660 -1380
rect 36800 -1410 36830 -1380
rect 36970 -1410 37000 -1380
rect 37140 -1410 37170 -1380
rect 37310 -1410 37340 -1380
rect 37480 -1410 37510 -1380
rect 37650 -1410 37680 -1380
rect 37820 -1410 37850 -1380
rect 37990 -1410 38020 -1380
rect 38160 -1410 38190 -1380
rect 38330 -1410 38360 -1380
rect 38500 -1410 38530 -1380
rect 38670 -1410 38700 -1380
rect 38840 -1410 38870 -1380
rect 39010 -1410 39040 -1380
rect 39180 -1410 39210 -1380
rect 39350 -1410 39380 -1380
rect 39520 -1410 39550 -1380
rect 39690 -1410 39720 -1380
rect 39860 -1410 39890 -1380
rect 40030 -1410 40060 -1380
rect 40200 -1410 40230 -1380
rect 40370 -1410 40400 -1380
rect 40540 -1410 40570 -1380
rect 40710 -1410 40740 -1380
rect 40880 -1410 40910 -1380
rect 41050 -1410 41080 -1380
rect 41220 -1410 41250 -1380
rect 41390 -1410 41420 -1380
rect 41560 -1410 41590 -1380
rect 41730 -1410 41760 -1380
rect 41900 -1410 41930 -1380
rect 42070 -1410 42100 -1380
rect 42240 -1410 42270 -1380
rect 42410 -1410 42440 -1380
rect 42580 -1410 42610 -1380
rect 42750 -1410 42780 -1380
rect 42920 -1410 42950 -1380
rect 43090 -1410 43120 -1380
rect 43260 -1410 43290 -1380
rect 43430 -1410 43460 -1380
rect 43600 -1410 43630 -1380
rect 43770 -1410 43800 -1380
rect 43940 -1410 43970 -1380
rect 44110 -1410 44140 -1380
rect 44280 -1410 44310 -1380
rect 44450 -1410 44480 -1380
rect 44620 -1410 44650 -1380
rect 44790 -1410 44820 -1380
rect 44960 -1410 44990 -1380
rect 45130 -1410 45160 -1380
rect 45300 -1410 45330 -1380
rect 45470 -1410 45500 -1380
rect 45640 -1410 45670 -1380
rect 45810 -1410 45840 -1380
rect 45980 -1410 46010 -1380
rect 46150 -1410 46180 -1380
rect 46320 -1410 46350 -1380
rect 46490 -1410 46520 -1380
rect 46660 -1410 46690 -1380
rect 46830 -1410 46860 -1380
rect 47000 -1410 47030 -1380
rect 47170 -1410 47200 -1380
rect 47340 -1410 47370 -1380
rect 47510 -1410 47540 -1380
rect 47680 -1410 47710 -1380
rect 47850 -1410 47880 -1380
rect 48020 -1410 48050 -1380
rect 48190 -1410 48220 -1380
rect 48360 -1410 48390 -1380
rect 48530 -1410 48560 -1380
rect 48700 -1410 48730 -1380
rect 48870 -1410 48900 -1380
rect 49040 -1410 49070 -1380
rect 49210 -1410 49240 -1380
rect 49380 -1410 49410 -1380
rect 49550 -1410 49580 -1380
rect 49720 -1410 49750 -1380
rect 49890 -1410 49920 -1380
rect 50060 -1410 50090 -1380
rect 50230 -1410 50260 -1380
rect 50400 -1410 50430 -1380
rect 50570 -1410 50600 -1380
rect 50740 -1410 50770 -1380
rect 50910 -1410 50940 -1380
rect 51080 -1410 51110 -1380
rect 51250 -1410 51280 -1380
rect 51420 -1410 51450 -1380
rect 51590 -1410 51620 -1380
rect 51760 -1410 51790 -1380
rect 51930 -1410 51960 -1380
rect 52100 -1410 52130 -1380
rect 52270 -1410 52300 -1380
rect 52440 -1410 52470 -1380
rect 52610 -1410 52640 -1380
rect 52780 -1410 52810 -1380
rect 52950 -1410 52980 -1380
rect 53120 -1410 53150 -1380
rect 53290 -1410 53320 -1380
rect 53460 -1410 53490 -1380
rect 53630 -1410 53660 -1380
rect 53800 -1410 53830 -1380
rect 53970 -1410 54000 -1380
rect 54140 -1410 54170 -1380
rect 54310 -1410 54340 -1380
rect 54480 -1410 54510 -1380
rect 54650 -1410 54680 -1380
rect 54820 -1410 54850 -1380
rect 54990 -1410 55020 -1380
rect 55160 -1410 55190 -1380
rect 55330 -1410 55360 -1380
rect 55500 -1410 55530 -1380
rect 55670 -1410 55700 -1380
rect 55840 -1410 55870 -1380
rect 56010 -1410 56040 -1380
rect 56180 -1410 56210 -1380
rect 56350 -1410 56380 -1380
rect 56520 -1410 56550 -1380
rect 56690 -1410 56720 -1380
rect 56860 -1410 56890 -1380
rect 57030 -1410 57060 -1380
rect 57200 -1410 57230 -1380
rect 57370 -1410 57400 -1380
rect 57540 -1410 57570 -1380
rect 57710 -1410 57740 -1380
rect 57880 -1410 57910 -1380
rect 58050 -1410 58080 -1380
rect 58220 -1410 58250 -1380
rect 58390 -1410 58420 -1380
rect 58560 -1410 58590 -1380
rect 58730 -1410 58760 -1380
rect 58900 -1410 58930 -1380
rect 59070 -1410 59100 -1380
rect 59240 -1410 59270 -1380
rect 59410 -1410 59440 -1380
rect 59580 -1410 59610 -1380
rect 59750 -1410 59780 -1380
rect 59920 -1410 59950 -1380
rect 60090 -1410 60120 -1380
rect 60260 -1410 60290 -1380
rect 60430 -1410 60460 -1380
rect 60600 -1410 60630 -1380
rect 60770 -1410 60800 -1380
rect 60940 -1410 60970 -1380
rect 61110 -1410 61140 -1380
rect 61280 -1410 61310 -1380
rect 61450 -1410 61480 -1380
rect 61620 -1410 61650 -1380
rect 61790 -1410 61820 -1380
rect 61960 -1410 61990 -1380
rect 62130 -1410 62160 -1380
rect 62300 -1410 62330 -1380
rect 62470 -1410 62500 -1380
rect 62640 -1410 62670 -1380
rect 62810 -1410 62840 -1380
rect 62980 -1410 63010 -1380
rect 63150 -1410 63180 -1380
rect 63320 -1410 63350 -1380
rect 63490 -1410 63520 -1380
rect 63660 -1410 63690 -1380
rect 63830 -1410 63860 -1380
rect 64000 -1410 64030 -1380
rect 64170 -1410 64200 -1380
rect 64340 -1410 64370 -1380
rect 64510 -1410 64540 -1380
rect 64680 -1410 64710 -1380
rect 64850 -1410 64880 -1380
rect 65020 -1410 65050 -1380
rect 65190 -1410 65220 -1380
rect 65360 -1410 65390 -1380
rect 65530 -1410 65560 -1380
rect 65700 -1410 65730 -1380
rect 65870 -1410 65900 -1380
rect 66040 -1410 66070 -1380
rect 66210 -1410 66240 -1380
rect 66380 -1410 66410 -1380
rect 66550 -1410 66580 -1380
rect 66720 -1410 66750 -1380
rect 66890 -1410 66920 -1380
rect 67060 -1410 67090 -1380
rect 67230 -1410 67260 -1380
rect 67400 -1410 67430 -1380
rect 67570 -1410 67600 -1380
rect 67740 -1410 67770 -1380
rect 67910 -1410 67940 -1380
rect 68080 -1410 68110 -1380
rect 68250 -1410 68280 -1380
rect 68420 -1410 68450 -1380
rect 68590 -1410 68620 -1380
rect 68760 -1410 68790 -1380
rect 68930 -1410 68960 -1380
rect 69100 -1410 69130 -1380
rect 69270 -1410 69300 -1380
rect 69440 -1410 69470 -1380
rect 69610 -1410 69640 -1380
rect 69780 -1410 69810 -1380
rect 69950 -1410 69980 -1380
rect 70120 -1410 70150 -1380
rect 70290 -1410 70320 -1380
rect 70460 -1410 70490 -1380
rect 70630 -1410 70660 -1380
rect 70800 -1410 70830 -1380
rect 70970 -1410 71000 -1380
rect 71140 -1410 71170 -1380
rect 71310 -1410 71340 -1380
rect 71480 -1410 71510 -1380
rect 71650 -1410 71680 -1380
rect 71820 -1410 71850 -1380
rect 71990 -1410 72020 -1380
rect 72160 -1410 72190 -1380
rect 72330 -1410 72360 -1380
rect 72500 -1410 72530 -1380
rect 72670 -1410 72700 -1380
rect 72840 -1410 72870 -1380
rect 73010 -1410 73040 -1380
rect 73180 -1410 73210 -1380
rect 73350 -1410 73380 -1380
rect 73520 -1410 73550 -1380
rect 73690 -1410 73720 -1380
rect 73860 -1410 73890 -1380
rect 74030 -1410 74060 -1380
rect 74200 -1410 74230 -1380
rect 74370 -1410 74400 -1380
rect 74540 -1410 74570 -1380
rect 74710 -1410 74740 -1380
rect 74880 -1410 74910 -1380
rect 75050 -1410 75080 -1380
rect 75220 -1410 75250 -1380
rect 75390 -1410 75420 -1380
rect 75560 -1410 75590 -1380
rect 75730 -1410 75760 -1380
rect 75900 -1410 75930 -1380
rect 76070 -1410 76100 -1380
rect 76240 -1410 76270 -1380
rect 76410 -1410 76440 -1380
rect 76580 -1410 76610 -1380
rect 76750 -1410 76780 -1380
rect 76920 -1410 76950 -1380
rect 77090 -1410 77120 -1380
rect 77260 -1410 77290 -1380
rect 77430 -1410 77460 -1380
rect 77600 -1410 77630 -1380
rect 77770 -1410 77800 -1380
rect 77940 -1410 77970 -1380
rect 78110 -1410 78140 -1380
rect 78280 -1410 78310 -1380
rect 78450 -1410 78480 -1380
rect 78620 -1410 78650 -1380
rect 78790 -1410 78820 -1380
rect 78960 -1410 78990 -1380
rect 79130 -1410 79160 -1380
rect 79300 -1410 79330 -1380
rect 79470 -1410 79500 -1380
rect 79640 -1410 79670 -1380
rect 79810 -1410 79840 -1380
rect 79980 -1410 80010 -1380
rect 80150 -1410 80180 -1380
rect 80320 -1410 80350 -1380
rect 80490 -1410 80520 -1380
rect 80660 -1410 80690 -1380
rect 80830 -1410 80860 -1380
rect 81000 -1410 81030 -1380
rect 81170 -1410 81200 -1380
rect 81340 -1410 81370 -1380
rect 81510 -1410 81540 -1380
rect 81680 -1410 81710 -1380
rect 81850 -1410 81880 -1380
rect 82020 -1410 82050 -1380
rect 82190 -1410 82220 -1380
rect 82360 -1410 82390 -1380
rect 82530 -1410 82560 -1380
rect 82700 -1410 82730 -1380
rect 82870 -1410 82900 -1380
rect 83040 -1410 83070 -1380
rect 83210 -1410 83240 -1380
rect 83380 -1410 83410 -1380
rect 83550 -1410 83580 -1380
rect 83720 -1410 83750 -1380
rect 83890 -1410 83920 -1380
rect 84060 -1410 84090 -1380
rect 84230 -1410 84260 -1380
rect 84400 -1410 84430 -1380
rect 84570 -1410 84600 -1380
rect 84740 -1410 84770 -1380
rect 84910 -1410 84940 -1380
rect 85080 -1410 85110 -1380
rect 85250 -1410 85280 -1380
rect 85420 -1410 85450 -1380
rect 85590 -1410 85620 -1380
rect 85760 -1410 85790 -1380
rect 85930 -1410 85960 -1380
rect 86100 -1410 86130 -1380
rect 86270 -1410 86300 -1380
rect 86440 -1410 86470 -1380
rect 86610 -1410 86640 -1380
rect 86780 -1410 86810 -1380
rect 86950 -1410 86980 -1380
rect 87120 -1410 87150 -1380
<< polycont >>
rect 520 630 610 690
rect 5630 630 5720 690
rect 70 30 130 110
rect 530 -120 600 -60
rect 700 -120 770 -60
rect 870 -120 940 -60
rect 1040 -120 1110 -60
rect 1600 -120 1670 -60
rect 1770 -120 1840 -60
rect 1940 -120 2010 -60
rect 2110 -120 2180 -60
rect 2280 -120 2350 -60
rect 2450 -120 2520 -60
rect 2620 -120 2690 -60
rect 2790 -120 2860 -60
rect 2960 -120 3030 -60
rect 3130 -120 3200 -60
rect 3300 -120 3370 -60
rect 3470 -120 3540 -60
rect 3640 -120 3710 -60
rect 3810 -120 3880 -60
rect 3980 -120 4050 -60
rect 4150 -120 4220 -60
rect 4620 -120 4690 -60
rect 4790 -120 4860 -60
rect 4960 -120 5030 -60
rect 5130 -120 5200 -60
rect 5300 -120 5370 -60
rect 5470 -120 5540 -60
rect 5640 -120 5710 -60
rect 5810 -120 5880 -60
rect 5980 -120 6050 -60
rect 6150 -120 6220 -60
rect 6320 -120 6390 -60
rect 6490 -120 6560 -60
rect 6660 -120 6730 -60
rect 6830 -120 6900 -60
rect 7000 -120 7070 -60
rect 7170 -120 7240 -60
rect 7340 -120 7410 -60
rect 7510 -120 7580 -60
rect 7680 -120 7750 -60
rect 7850 -120 7920 -60
rect 8020 -120 8090 -60
rect 8190 -120 8260 -60
rect 8360 -120 8430 -60
rect 8530 -120 8600 -60
rect 8700 -120 8770 -60
rect 8870 -120 8940 -60
rect 9040 -120 9110 -60
rect 9210 -120 9280 -60
rect 9380 -120 9450 -60
rect 9550 -120 9620 -60
rect 9720 -120 9790 -60
rect 9890 -120 9960 -60
rect 10060 -120 10130 -60
rect 10230 -120 10300 -60
rect 10400 -120 10470 -60
rect 10570 -120 10640 -60
rect 10740 -120 10810 -60
rect 10910 -120 10980 -60
rect 11080 -120 11150 -60
rect 11250 -120 11320 -60
rect 11420 -120 11490 -60
rect 11590 -120 11660 -60
rect 11760 -120 11830 -60
rect 11930 -120 12000 -60
rect 12100 -120 12170 -60
rect 12270 -120 12340 -60
rect 12440 -120 12510 -60
rect 12610 -120 12680 -60
rect 12780 -120 12850 -60
rect 12950 -120 13020 -60
rect 13120 -120 13190 -60
rect 13290 -120 13360 -60
rect 13460 -120 13530 -60
rect 13630 -120 13700 -60
rect 13800 -120 13870 -60
rect 13970 -120 14040 -60
rect 14140 -120 14210 -60
rect 14310 -120 14380 -60
rect 14480 -120 14550 -60
rect 14650 -120 14720 -60
rect 14820 -120 14890 -60
rect 14990 -120 15060 -60
rect 15160 -120 15230 -60
rect 15330 -120 15400 -60
rect 15800 -120 15870 -60
rect 15970 -120 16040 -60
rect 16140 -120 16210 -60
rect 16310 -120 16380 -60
rect 16480 -120 16550 -60
rect 16650 -120 16720 -60
rect 16820 -120 16890 -60
rect 16990 -120 17060 -60
rect 17160 -120 17230 -60
rect 17330 -120 17400 -60
rect 17500 -120 17570 -60
rect 17670 -120 17740 -60
rect 17840 -120 17910 -60
rect 18010 -120 18080 -60
rect 18180 -120 18250 -60
rect 18350 -120 18420 -60
rect 18520 -120 18590 -60
rect 18690 -120 18760 -60
rect 18860 -120 18930 -60
rect 19030 -120 19100 -60
rect 19200 -120 19270 -60
rect 19370 -120 19440 -60
rect 19540 -120 19610 -60
rect 19710 -120 19780 -60
rect 19880 -120 19950 -60
rect 20050 -120 20120 -60
rect 20220 -120 20290 -60
rect 20390 -120 20460 -60
rect 20560 -120 20630 -60
rect 20730 -120 20800 -60
rect 20900 -120 20970 -60
rect 21070 -120 21140 -60
rect 21240 -120 21310 -60
rect 21410 -120 21480 -60
rect 21580 -120 21650 -60
rect 21750 -120 21820 -60
rect 21920 -120 21990 -60
rect 22090 -120 22160 -60
rect 22260 -120 22330 -60
rect 22430 -120 22500 -60
rect 22600 -120 22670 -60
rect 22770 -120 22840 -60
rect 22940 -120 23010 -60
rect 23110 -120 23180 -60
rect 23280 -120 23350 -60
rect 23450 -120 23520 -60
rect 23620 -120 23690 -60
rect 23790 -120 23860 -60
rect 23960 -120 24030 -60
rect 24130 -120 24200 -60
rect 24300 -120 24370 -60
rect 24470 -120 24540 -60
rect 24640 -120 24710 -60
rect 24810 -120 24880 -60
rect 24980 -120 25050 -60
rect 25150 -120 25220 -60
rect 25320 -120 25390 -60
rect 25490 -120 25560 -60
rect 25660 -120 25730 -60
rect 25830 -120 25900 -60
rect 26000 -120 26070 -60
rect 26170 -120 26240 -60
rect 26340 -120 26410 -60
rect 26510 -120 26580 -60
rect 26680 -120 26750 -60
rect 26850 -120 26920 -60
rect 27020 -120 27090 -60
rect 27190 -120 27260 -60
rect 27360 -120 27430 -60
rect 27530 -120 27600 -60
rect 27700 -120 27770 -60
rect 27870 -120 27940 -60
rect 28040 -120 28110 -60
rect 28210 -120 28280 -60
rect 28380 -120 28450 -60
rect 28550 -120 28620 -60
rect 28720 -120 28790 -60
rect 28890 -120 28960 -60
rect 29060 -120 29130 -60
rect 29230 -120 29300 -60
rect 29400 -120 29470 -60
rect 29570 -120 29640 -60
rect 29740 -120 29810 -60
rect 29910 -120 29980 -60
rect 30080 -120 30150 -60
rect 30250 -120 30320 -60
rect 30420 -120 30490 -60
rect 30590 -120 30660 -60
rect 30760 -120 30830 -60
rect 30930 -120 31000 -60
rect 31100 -120 31170 -60
rect 31270 -120 31340 -60
rect 31440 -120 31510 -60
rect 31610 -120 31680 -60
rect 31780 -120 31850 -60
rect 31950 -120 32020 -60
rect 32120 -120 32190 -60
rect 32290 -120 32360 -60
rect 32460 -120 32530 -60
rect 32630 -120 32700 -60
rect 32800 -120 32870 -60
rect 32970 -120 33040 -60
rect 33140 -120 33210 -60
rect 33310 -120 33380 -60
rect 33480 -120 33550 -60
rect 33650 -120 33720 -60
rect 33820 -120 33890 -60
rect 33990 -120 34060 -60
rect 34160 -120 34230 -60
rect 34330 -120 34400 -60
rect 34500 -120 34570 -60
rect 34670 -120 34740 -60
rect 34840 -120 34910 -60
rect 35010 -120 35080 -60
rect 35180 -120 35250 -60
rect 35350 -120 35420 -60
rect 35520 -120 35590 -60
rect 35690 -120 35760 -60
rect 35860 -120 35930 -60
rect 36030 -120 36100 -60
rect 36200 -120 36270 -60
rect 36370 -120 36440 -60
rect 36540 -120 36610 -60
rect 36710 -120 36780 -60
rect 36880 -120 36950 -60
rect 37050 -120 37120 -60
rect 37220 -120 37290 -60
rect 37390 -120 37460 -60
rect 37560 -120 37630 -60
rect 37730 -120 37800 -60
rect 37900 -120 37970 -60
rect 38070 -120 38140 -60
rect 38240 -120 38310 -60
rect 38410 -120 38480 -60
rect 38580 -120 38650 -60
rect 38750 -120 38820 -60
rect 38920 -120 38990 -60
rect 39090 -120 39160 -60
rect 39260 -120 39330 -60
rect 39430 -120 39500 -60
rect 39600 -120 39670 -60
rect 39770 -120 39840 -60
rect 39940 -120 40010 -60
rect 40110 -120 40180 -60
rect 40280 -120 40350 -60
rect 40450 -120 40520 -60
rect 40620 -120 40690 -60
rect 40790 -120 40860 -60
rect 40960 -120 41030 -60
rect 41130 -120 41200 -60
rect 41300 -120 41370 -60
rect 41470 -120 41540 -60
rect 41640 -120 41710 -60
rect 41810 -120 41880 -60
rect 41980 -120 42050 -60
rect 42150 -120 42220 -60
rect 42320 -120 42390 -60
rect 42490 -120 42560 -60
rect 42660 -120 42730 -60
rect 42830 -120 42900 -60
rect 43000 -120 43070 -60
rect 43170 -120 43240 -60
rect 43340 -120 43410 -60
rect 43510 -120 43580 -60
rect 43680 -120 43750 -60
rect 43850 -120 43920 -60
rect 44020 -120 44090 -60
rect 44190 -120 44260 -60
rect 44360 -120 44430 -60
rect 44530 -120 44600 -60
rect 44700 -120 44770 -60
rect 44870 -120 44940 -60
rect 45040 -120 45110 -60
rect 45210 -120 45280 -60
rect 45380 -120 45450 -60
rect 45550 -120 45620 -60
rect 45720 -120 45790 -60
rect 45890 -120 45960 -60
rect 46060 -120 46130 -60
rect 46230 -120 46300 -60
rect 46400 -120 46470 -60
rect 46570 -120 46640 -60
rect 46740 -120 46810 -60
rect 46910 -120 46980 -60
rect 47080 -120 47150 -60
rect 47250 -120 47320 -60
rect 47420 -120 47490 -60
rect 47590 -120 47660 -60
rect 47760 -120 47830 -60
rect 47930 -120 48000 -60
rect 48100 -120 48170 -60
rect 48270 -120 48340 -60
rect 48440 -120 48510 -60
rect 48610 -120 48680 -60
rect 48780 -120 48850 -60
rect 48950 -120 49020 -60
rect 49120 -120 49190 -60
rect 49290 -120 49360 -60
rect 49460 -120 49530 -60
rect 49630 -120 49700 -60
rect 49800 -120 49870 -60
rect 49970 -120 50040 -60
rect 50140 -120 50210 -60
rect 50310 -120 50380 -60
rect 50480 -120 50550 -60
rect 50650 -120 50720 -60
rect 50820 -120 50890 -60
rect 50990 -120 51060 -60
rect 51160 -120 51230 -60
rect 51330 -120 51400 -60
rect 51500 -120 51570 -60
rect 51670 -120 51740 -60
rect 51840 -120 51910 -60
rect 52010 -120 52080 -60
rect 52180 -120 52250 -60
rect 52350 -120 52420 -60
rect 52520 -120 52590 -60
rect 52690 -120 52760 -60
rect 52860 -120 52930 -60
rect 53030 -120 53100 -60
rect 53200 -120 53270 -60
rect 53370 -120 53440 -60
rect 53540 -120 53610 -60
rect 53710 -120 53780 -60
rect 53880 -120 53950 -60
rect 54050 -120 54120 -60
rect 54220 -120 54290 -60
rect 54390 -120 54460 -60
rect 54560 -120 54630 -60
rect 54730 -120 54800 -60
rect 54900 -120 54970 -60
rect 55070 -120 55140 -60
rect 55240 -120 55310 -60
rect 55410 -120 55480 -60
rect 55580 -120 55650 -60
rect 55750 -120 55820 -60
rect 55920 -120 55990 -60
rect 56090 -120 56160 -60
rect 56260 -120 56330 -60
rect 56430 -120 56500 -60
rect 56600 -120 56670 -60
rect 56770 -120 56840 -60
rect 56940 -120 57010 -60
rect 57110 -120 57180 -60
rect 57280 -120 57350 -60
rect 57450 -120 57520 -60
rect 57620 -120 57690 -60
rect 57790 -120 57860 -60
rect 57960 -120 58030 -60
rect 58130 -120 58200 -60
rect 58300 -120 58370 -60
rect 58470 -120 58540 -60
rect 58640 -120 58710 -60
rect 58810 -120 58880 -60
rect 58980 -120 59050 -60
rect 59150 -120 59220 -60
rect 230 -590 300 -530
rect 400 -590 470 -530
rect 570 -590 640 -530
rect 740 -590 810 -530
rect 910 -590 980 -530
rect 1080 -590 1150 -530
rect 1250 -590 1320 -530
rect 1420 -590 1490 -530
rect 1590 -590 1660 -530
rect 1760 -590 1830 -530
rect 1930 -590 2000 -530
rect 2100 -590 2170 -530
rect 2270 -590 2340 -530
rect 2440 -590 2510 -530
rect 2610 -590 2680 -530
rect 2780 -590 2850 -530
rect 2950 -590 3020 -530
rect 3120 -590 3190 -530
rect 3290 -590 3360 -530
rect 3460 -590 3530 -530
rect 3630 -590 3700 -530
rect 3800 -590 3870 -530
rect 3970 -590 4040 -530
rect 4140 -590 4210 -530
rect 4310 -590 4380 -530
rect 4480 -590 4550 -530
rect 4650 -590 4720 -530
rect 4820 -590 4890 -530
rect 4990 -590 5060 -530
rect 5160 -590 5230 -530
rect 5330 -590 5400 -530
rect 5500 -590 5570 -530
rect 5670 -590 5740 -530
rect 5840 -590 5910 -530
rect 6010 -590 6080 -530
rect 6180 -590 6250 -530
rect 6350 -590 6420 -530
rect 6520 -590 6590 -530
rect 6690 -590 6760 -530
rect 6860 -590 6930 -530
rect 7030 -590 7100 -530
rect 7200 -590 7270 -530
rect 7370 -590 7440 -530
rect 7540 -590 7610 -530
rect 7710 -590 7780 -530
rect 7880 -590 7950 -530
rect 8050 -590 8120 -530
rect 8220 -590 8290 -530
rect 8390 -590 8460 -530
rect 8560 -590 8630 -530
rect 8730 -590 8800 -530
rect 8900 -590 8970 -530
rect 9070 -590 9140 -530
rect 9240 -590 9310 -530
rect 9410 -590 9480 -530
rect 9580 -590 9650 -530
rect 9750 -590 9820 -530
rect 9920 -590 9990 -530
rect 10090 -590 10160 -530
rect 10260 -590 10330 -530
rect 10430 -590 10500 -530
rect 10600 -590 10670 -530
rect 10770 -590 10840 -530
rect 10940 -590 11010 -530
rect 11110 -590 11180 -530
rect 11280 -590 11350 -530
rect 11450 -590 11520 -530
rect 11620 -590 11690 -530
rect 11790 -590 11860 -530
rect 11960 -590 12030 -530
rect 12130 -590 12200 -530
rect 12300 -590 12370 -530
rect 12470 -590 12540 -530
rect 12640 -590 12710 -530
rect 12810 -590 12880 -530
rect 12980 -590 13050 -530
rect 13150 -590 13220 -530
rect 13320 -590 13390 -530
rect 13490 -590 13560 -530
rect 13660 -590 13730 -530
rect 13830 -590 13900 -530
rect 14000 -590 14070 -530
rect 14170 -590 14240 -530
rect 14340 -590 14410 -530
rect 14510 -590 14580 -530
rect 14680 -590 14750 -530
rect 14850 -590 14920 -530
rect 15020 -590 15090 -530
rect 15190 -590 15260 -530
rect 15360 -590 15430 -530
rect 15530 -590 15600 -530
rect 15700 -590 15770 -530
rect 15870 -590 15940 -530
rect 16040 -590 16110 -530
rect 16210 -590 16280 -530
rect 16380 -590 16450 -530
rect 16550 -590 16620 -530
rect 16720 -590 16790 -530
rect 16890 -590 16960 -530
rect 17060 -590 17130 -530
rect 17230 -590 17300 -530
rect 17400 -590 17470 -530
rect 17570 -590 17640 -530
rect 17740 -590 17810 -530
rect 17910 -590 17980 -530
rect 18080 -590 18150 -530
rect 18250 -590 18320 -530
rect 18420 -590 18490 -530
rect 18590 -590 18660 -530
rect 18760 -590 18830 -530
rect 18930 -590 19000 -530
rect 19100 -590 19170 -530
rect 19270 -590 19340 -530
rect 19440 -590 19510 -530
rect 19610 -590 19680 -530
rect 19780 -590 19850 -530
rect 19950 -590 20020 -530
rect 20120 -590 20190 -530
rect 20290 -590 20360 -530
rect 20460 -590 20530 -530
rect 20630 -590 20700 -530
rect 20800 -590 20870 -530
rect 20970 -590 21040 -530
rect 21140 -590 21210 -530
rect 21310 -590 21380 -530
rect 21480 -590 21550 -530
rect 21650 -590 21720 -530
rect 21820 -590 21890 -530
rect 21990 -590 22060 -530
rect 22160 -590 22230 -530
rect 22330 -590 22400 -530
rect 22500 -590 22570 -530
rect 22670 -590 22740 -530
rect 22840 -590 22910 -530
rect 23010 -590 23080 -530
rect 23180 -590 23250 -530
rect 23350 -590 23420 -530
rect 23520 -590 23590 -530
rect 23690 -590 23760 -530
rect 23860 -590 23930 -530
rect 24030 -590 24100 -530
rect 24200 -590 24270 -530
rect 24370 -590 24440 -530
rect 24540 -590 24610 -530
rect 24710 -590 24780 -530
rect 24880 -590 24950 -530
rect 25050 -590 25120 -530
rect 25220 -590 25290 -530
rect 25390 -590 25460 -530
rect 25560 -590 25630 -530
rect 25730 -590 25800 -530
rect 25900 -590 25970 -530
rect 26070 -590 26140 -530
rect 26240 -590 26310 -530
rect 26410 -590 26480 -530
rect 26580 -590 26650 -530
rect 26750 -590 26820 -530
rect 26920 -590 26990 -530
rect 27090 -590 27160 -530
rect 27260 -590 27330 -530
rect 27430 -590 27500 -530
rect 27600 -590 27670 -530
rect 27770 -590 27840 -530
rect 27940 -590 28010 -530
rect 28110 -590 28180 -530
rect 28280 -590 28350 -530
rect 28450 -590 28520 -530
rect 28620 -590 28690 -530
rect 28790 -590 28860 -530
rect 28960 -590 29030 -530
rect 29130 -590 29200 -530
rect 29300 -590 29370 -530
rect 29470 -590 29540 -530
rect 29640 -590 29710 -530
rect 29810 -590 29880 -530
rect 29980 -590 30050 -530
rect 30150 -590 30220 -530
rect 30320 -590 30390 -530
rect 30490 -590 30560 -530
rect 30660 -590 30730 -530
rect 30830 -590 30900 -530
rect 31000 -590 31070 -530
rect 31170 -590 31240 -530
rect 31340 -590 31410 -530
rect 31510 -590 31580 -530
rect 31680 -590 31750 -530
rect 31850 -590 31920 -530
rect 32020 -590 32090 -530
rect 32190 -590 32260 -530
rect 32360 -590 32430 -530
rect 32530 -590 32600 -530
rect 32700 -590 32770 -530
rect 32870 -590 32940 -530
rect 33040 -590 33110 -530
rect 33210 -590 33280 -530
rect 33380 -590 33450 -530
rect 33550 -590 33620 -530
rect 33720 -590 33790 -530
rect 33890 -590 33960 -530
rect 34060 -590 34130 -530
rect 34230 -590 34300 -530
rect 34400 -590 34470 -530
rect 34570 -590 34640 -530
rect 34740 -590 34810 -530
rect 34910 -590 34980 -530
rect 35080 -590 35150 -530
rect 35250 -590 35320 -530
rect 35420 -590 35490 -530
rect 35590 -590 35660 -530
rect 35760 -590 35830 -530
rect 35930 -590 36000 -530
rect 36100 -590 36170 -530
rect 36270 -590 36340 -530
rect 36440 -590 36510 -530
rect 36610 -590 36680 -530
rect 36780 -590 36850 -530
rect 36950 -590 37020 -530
rect 37120 -590 37190 -530
rect 37290 -590 37360 -530
rect 37460 -590 37530 -530
rect 37630 -590 37700 -530
rect 37800 -590 37870 -530
rect 37970 -590 38040 -530
rect 38140 -590 38210 -530
rect 38310 -590 38380 -530
rect 38480 -590 38550 -530
rect 38650 -590 38720 -530
rect 38820 -590 38890 -530
rect 38990 -590 39060 -530
rect 39160 -590 39230 -530
rect 39330 -590 39400 -530
rect 39500 -590 39570 -530
rect 39670 -590 39740 -530
rect 39840 -590 39910 -530
rect 40010 -590 40080 -530
rect 40180 -590 40250 -530
rect 40350 -590 40420 -530
rect 40520 -590 40590 -530
rect 40690 -590 40760 -530
rect 40860 -590 40930 -530
rect 41030 -590 41100 -530
rect 41200 -590 41270 -530
rect 41370 -590 41440 -530
rect 41540 -590 41610 -530
rect 41710 -590 41780 -530
rect 41880 -590 41950 -530
rect 42050 -590 42120 -530
rect 42220 -590 42290 -530
rect 42390 -590 42460 -530
rect 42560 -590 42630 -530
rect 42730 -590 42800 -530
rect 42900 -590 42970 -530
rect 43070 -590 43140 -530
rect 43240 -590 43310 -530
rect 43410 -590 43480 -530
rect 43580 -590 43650 -530
rect 43750 -590 43820 -530
rect 43920 -590 43990 -530
rect 44090 -590 44160 -530
rect 44260 -590 44330 -530
rect 44430 -590 44500 -530
rect 44600 -590 44670 -530
rect 44770 -590 44840 -530
rect 44940 -590 45010 -530
rect 45110 -590 45180 -530
rect 45280 -590 45350 -530
rect 45450 -590 45520 -530
rect 45620 -590 45690 -530
rect 45790 -590 45860 -530
rect 45960 -590 46030 -530
rect 46130 -590 46200 -530
rect 46300 -590 46370 -530
rect 46470 -590 46540 -530
rect 46640 -590 46710 -530
rect 46810 -590 46880 -530
rect 46980 -590 47050 -530
rect 47150 -590 47220 -530
rect 47320 -590 47390 -530
rect 47490 -590 47560 -530
rect 47660 -590 47730 -530
rect 47830 -590 47900 -530
rect 48000 -590 48070 -530
rect 48170 -590 48240 -530
rect 48340 -590 48410 -530
rect 48510 -590 48580 -530
rect 48680 -590 48750 -530
rect 48850 -590 48920 -530
rect 49020 -590 49090 -530
rect 49190 -590 49260 -530
rect 49360 -590 49430 -530
rect 49530 -590 49600 -530
rect 49700 -590 49770 -530
rect 49870 -590 49940 -530
rect 50040 -590 50110 -530
rect 50210 -590 50280 -530
rect 50380 -590 50450 -530
rect 50550 -590 50620 -530
rect 50720 -590 50790 -530
rect 50890 -590 50960 -530
rect 51060 -590 51130 -530
rect 51230 -590 51300 -530
rect 51400 -590 51470 -530
rect 51570 -590 51640 -530
rect 51740 -590 51810 -530
rect 51910 -590 51980 -530
rect 52080 -590 52150 -530
rect 52250 -590 52320 -530
rect 52420 -590 52490 -530
rect 52590 -590 52660 -530
rect 52760 -590 52830 -530
rect 52930 -590 53000 -530
rect 53100 -590 53170 -530
rect 53270 -590 53340 -530
rect 53440 -590 53510 -530
rect 53610 -590 53680 -530
rect 53780 -590 53850 -530
rect 53950 -590 54020 -530
rect 54120 -590 54190 -530
rect 54290 -590 54360 -530
rect 54460 -590 54530 -530
rect 54630 -590 54700 -530
rect 54800 -590 54870 -530
rect 54970 -590 55040 -530
rect 55140 -590 55210 -530
rect 55310 -590 55380 -530
rect 55480 -590 55550 -530
rect 55650 -590 55720 -530
rect 55820 -590 55890 -530
rect 55990 -590 56060 -530
rect 56160 -590 56230 -530
rect 56330 -590 56400 -530
rect 56500 -590 56570 -530
rect 56670 -590 56740 -530
rect 56840 -590 56910 -530
rect 57010 -590 57080 -530
rect 57180 -590 57250 -530
rect 57350 -590 57420 -530
rect 57520 -590 57590 -530
rect 57690 -590 57760 -530
rect 57860 -590 57930 -530
rect 58030 -590 58100 -530
rect 58200 -590 58270 -530
rect 58370 -590 58440 -530
rect 58540 -590 58610 -530
rect 58710 -590 58780 -530
rect 58880 -590 58950 -530
rect 59050 -590 59120 -530
rect 59220 -590 59290 -530
rect 59390 -590 59460 -530
rect 59560 -590 59630 -530
rect 59730 -590 59800 -530
rect 59900 -590 59970 -530
rect 60070 -590 60140 -530
rect 60240 -590 60310 -530
rect 60410 -590 60480 -530
rect 60580 -590 60650 -530
rect 60750 -590 60820 -530
rect 60920 -590 60990 -530
rect 61090 -590 61160 -530
rect 61260 -590 61330 -530
rect 61430 -590 61500 -530
rect 61600 -590 61670 -530
rect 61770 -590 61840 -530
rect 61940 -590 62010 -530
rect 62110 -590 62180 -530
rect 62280 -590 62350 -530
rect 62450 -590 62520 -530
rect 62620 -590 62690 -530
rect 62790 -590 62860 -530
rect 62960 -590 63030 -530
rect 63130 -590 63200 -530
rect 63300 -590 63370 -530
rect 63470 -590 63540 -530
rect 63640 -590 63710 -530
rect 63810 -590 63880 -530
rect 63980 -590 64050 -530
rect 64150 -590 64220 -530
rect 64320 -590 64390 -530
rect 64490 -590 64560 -530
rect 64660 -590 64730 -530
rect 64830 -590 64900 -530
rect 65000 -590 65070 -530
rect 65170 -590 65240 -530
rect 65340 -590 65410 -530
rect 65510 -590 65580 -530
rect 65680 -590 65750 -530
rect 65850 -590 65920 -530
rect 66020 -590 66090 -530
rect 66190 -590 66260 -530
rect 66360 -590 66430 -530
rect 66530 -590 66600 -530
rect 66700 -590 66770 -530
rect 66870 -590 66940 -530
rect 67040 -590 67110 -530
rect 67210 -590 67280 -530
rect 67380 -590 67450 -530
rect 67550 -590 67620 -530
rect 67720 -590 67790 -530
rect 67890 -590 67960 -530
rect 68060 -590 68130 -530
rect 68230 -590 68300 -530
rect 68400 -590 68470 -530
rect 68570 -590 68640 -530
rect 68740 -590 68810 -530
rect 68910 -590 68980 -530
rect 69080 -590 69150 -530
rect 69250 -590 69320 -530
rect 69420 -590 69490 -530
rect 69590 -590 69660 -530
rect 69760 -590 69830 -530
rect 69930 -590 70000 -530
rect 70100 -590 70170 -530
rect 70270 -590 70340 -530
rect 70440 -590 70510 -530
rect 70610 -590 70680 -530
rect 70780 -590 70850 -530
rect 70950 -590 71020 -530
rect 71120 -590 71190 -530
rect 71290 -590 71360 -530
rect 71460 -590 71530 -530
rect 71630 -590 71700 -530
rect 71800 -590 71870 -530
rect 71970 -590 72040 -530
rect 72140 -590 72210 -530
rect 72310 -590 72380 -530
rect 72480 -590 72550 -530
rect 72650 -590 72720 -530
rect 72820 -590 72890 -530
rect 72990 -590 73060 -530
rect 73160 -590 73230 -530
rect 73330 -590 73400 -530
rect 73500 -590 73570 -530
rect 73670 -590 73740 -530
rect 73840 -590 73910 -530
rect 74010 -590 74080 -530
rect 74180 -590 74250 -530
rect 74350 -590 74420 -530
rect 74520 -590 74590 -530
rect 74690 -590 74760 -530
rect 74860 -590 74930 -530
rect 75030 -590 75100 -530
rect 75200 -590 75270 -530
rect 75370 -590 75440 -530
rect 75540 -590 75610 -530
rect 75710 -590 75780 -530
rect 75880 -590 75950 -530
rect 76050 -590 76120 -530
rect 76220 -590 76290 -530
rect 76390 -590 76460 -530
rect 76560 -590 76630 -530
rect 76730 -590 76800 -530
rect 76900 -590 76970 -530
rect 77070 -590 77140 -530
rect 77240 -590 77310 -530
rect 77410 -590 77480 -530
rect 77580 -590 77650 -530
rect 77750 -590 77820 -530
rect 77920 -590 77990 -530
rect 78090 -590 78160 -530
rect 78260 -590 78330 -530
rect 78430 -590 78500 -530
rect 78600 -590 78670 -530
rect 78770 -590 78840 -530
rect 78940 -590 79010 -530
rect 79110 -590 79180 -530
rect 79280 -590 79350 -530
rect 79450 -590 79520 -530
rect 79620 -590 79690 -530
rect 79790 -590 79860 -530
rect 79960 -590 80030 -530
rect 80130 -590 80200 -530
rect 80300 -590 80370 -530
rect 80470 -590 80540 -530
rect 80640 -590 80710 -530
rect 80810 -590 80880 -530
rect 80980 -590 81050 -530
rect 81150 -590 81220 -530
rect 81320 -590 81390 -530
rect 81490 -590 81560 -530
rect 81660 -590 81730 -530
rect 81830 -590 81900 -530
rect 82000 -590 82070 -530
rect 82170 -590 82240 -530
rect 82340 -590 82410 -530
rect 82510 -590 82580 -530
rect 82680 -590 82750 -530
rect 82850 -590 82920 -530
rect 83020 -590 83090 -530
rect 83190 -590 83260 -530
rect 83360 -590 83430 -530
rect 83530 -590 83600 -530
rect 83700 -590 83770 -530
rect 83870 -590 83940 -530
rect 84040 -590 84110 -530
rect 84210 -590 84280 -530
rect 84380 -590 84450 -530
rect 84550 -590 84620 -530
rect 84720 -590 84790 -530
rect 84890 -590 84960 -530
rect 85060 -590 85130 -530
rect 85230 -590 85300 -530
rect 85400 -590 85470 -530
rect 85570 -590 85640 -530
rect 85740 -590 85810 -530
rect 85910 -590 85980 -530
rect 86080 -590 86150 -530
rect 86250 -590 86320 -530
rect 86420 -590 86490 -530
rect 86590 -590 86660 -530
rect 86760 -590 86830 -530
rect 86930 -590 87000 -530
rect 87100 -590 87170 -530
<< ndiffres >>
rect 634 923 1254 1007
rect 5754 901 6374 985
<< locali >>
rect 409 1095 505 1129
rect 1383 1095 1479 1129
rect 409 1033 443 1095
rect 1445 1033 1479 1095
rect 543 1010 577 1011
rect 540 995 580 1010
rect 1311 995 1345 1011
rect 540 935 543 995
rect 540 910 580 935
rect 1311 919 1345 935
rect 409 835 443 897
rect 1445 835 1479 897
rect 409 801 505 835
rect 1383 801 1479 835
rect 5529 1073 5625 1107
rect 6503 1073 6599 1107
rect 5529 1011 5563 1073
rect 6565 1011 6599 1073
rect 5663 973 5697 989
rect 6431 973 6465 989
rect 5663 897 5697 913
rect 6431 897 6465 913
rect 5529 813 5563 875
rect 6565 813 6599 875
rect 5529 779 5625 813
rect 6503 779 6599 813
rect 500 690 630 710
rect 500 630 520 690
rect 610 630 630 690
rect 500 610 630 630
rect 5610 690 5740 710
rect 5610 630 5630 690
rect 5720 630 5740 690
rect 730 590 930 620
rect 730 520 790 590
rect 870 520 930 590
rect 730 490 930 520
rect 2110 590 2310 620
rect 2110 520 2170 590
rect 2250 520 2310 590
rect 2110 490 2310 520
rect 3490 590 3690 620
rect 3490 520 3550 590
rect 3630 520 3690 590
rect 3490 490 3690 520
rect 5150 590 5350 620
rect 5610 610 5740 630
rect 5150 520 5210 590
rect 5290 520 5350 590
rect 5150 490 5350 520
rect 7980 590 8180 620
rect 7980 520 8040 590
rect 8120 520 8180 590
rect 7980 490 8180 520
rect 10740 590 10940 620
rect 10740 520 10800 590
rect 10880 520 10940 590
rect 10740 490 10940 520
rect 13370 590 13570 620
rect 13370 520 13430 590
rect 13510 520 13570 590
rect 13370 490 13570 520
rect 16410 590 16610 620
rect 16410 520 16470 590
rect 16550 520 16610 590
rect 16410 490 16610 520
rect 20480 590 20680 620
rect 20480 520 20540 590
rect 20620 520 20680 590
rect 20480 490 20680 520
rect 24620 590 24820 620
rect 24620 520 24680 590
rect 24760 520 24820 590
rect 24620 490 24820 520
rect 28700 590 28900 620
rect 28700 520 28760 590
rect 28840 520 28900 590
rect 28700 490 28900 520
rect 32850 590 33050 620
rect 32850 520 32910 590
rect 32990 520 33050 590
rect 32850 490 33050 520
rect 36720 590 36920 620
rect 36720 520 36780 590
rect 36860 520 36920 590
rect 36720 490 36920 520
rect 40860 590 41060 620
rect 40860 520 40920 590
rect 41000 520 41060 590
rect 40860 490 41060 520
rect 44850 590 45050 620
rect 44850 520 44910 590
rect 44990 520 45050 590
rect 44850 490 45050 520
rect 48930 590 49130 620
rect 48930 520 48990 590
rect 49070 520 49130 590
rect 48930 490 49130 520
rect 53020 590 53220 620
rect 53020 520 53080 590
rect 53160 520 53220 590
rect 53020 490 53220 520
rect 57180 590 57380 620
rect 57180 520 57240 590
rect 57320 520 57380 590
rect 57180 490 57380 520
rect 10 410 110 430
rect 10 350 30 410
rect 90 350 110 410
rect 10 310 110 350
rect 10 250 30 310
rect 90 250 110 310
rect 10 230 110 250
rect 180 410 280 430
rect 180 350 200 410
rect 260 350 280 410
rect 180 310 280 350
rect 180 250 200 310
rect 260 250 280 310
rect 180 230 280 250
rect 430 410 530 430
rect 430 350 450 410
rect 510 350 530 410
rect 430 310 530 350
rect 430 250 450 310
rect 510 250 530 310
rect 430 230 530 250
rect 600 410 700 430
rect 600 350 620 410
rect 680 350 700 410
rect 600 310 700 350
rect 600 250 620 310
rect 680 250 700 310
rect 600 230 700 250
rect 770 410 870 430
rect 770 350 790 410
rect 850 350 870 410
rect 770 310 870 350
rect 770 250 790 310
rect 850 250 870 310
rect 770 230 870 250
rect 940 410 1040 430
rect 940 350 960 410
rect 1020 350 1040 410
rect 940 310 1040 350
rect 940 250 960 310
rect 1020 250 1040 310
rect 940 230 1040 250
rect 1110 410 1210 430
rect 1110 350 1130 410
rect 1190 350 1210 410
rect 1110 310 1210 350
rect 1110 250 1130 310
rect 1190 250 1210 310
rect 1110 230 1210 250
rect 1500 410 1600 430
rect 1500 350 1520 410
rect 1580 350 1600 410
rect 1500 310 1600 350
rect 1500 250 1520 310
rect 1580 250 1600 310
rect 1500 230 1600 250
rect 1670 410 1770 430
rect 1670 350 1690 410
rect 1750 350 1770 410
rect 1670 310 1770 350
rect 1670 250 1690 310
rect 1750 250 1770 310
rect 1670 230 1770 250
rect 1840 410 1940 430
rect 1840 350 1860 410
rect 1920 350 1940 410
rect 1840 310 1940 350
rect 1840 250 1860 310
rect 1920 250 1940 310
rect 1840 230 1940 250
rect 2010 410 2110 430
rect 2010 350 2030 410
rect 2090 350 2110 410
rect 2010 310 2110 350
rect 2010 250 2030 310
rect 2090 250 2110 310
rect 2010 230 2110 250
rect 2180 410 2280 430
rect 2180 350 2200 410
rect 2260 350 2280 410
rect 2180 310 2280 350
rect 2180 250 2200 310
rect 2260 250 2280 310
rect 2180 230 2280 250
rect 2350 410 2450 430
rect 2350 350 2370 410
rect 2430 350 2450 410
rect 2350 310 2450 350
rect 2350 250 2370 310
rect 2430 250 2450 310
rect 2350 230 2450 250
rect 2520 410 2620 430
rect 2520 350 2540 410
rect 2600 350 2620 410
rect 2520 310 2620 350
rect 2520 250 2540 310
rect 2600 250 2620 310
rect 2520 230 2620 250
rect 2690 410 2790 430
rect 2690 350 2710 410
rect 2770 350 2790 410
rect 2690 310 2790 350
rect 2690 250 2710 310
rect 2770 250 2790 310
rect 2690 230 2790 250
rect 2860 410 2960 430
rect 2860 350 2880 410
rect 2940 350 2960 410
rect 2860 310 2960 350
rect 2860 250 2880 310
rect 2940 250 2960 310
rect 2860 230 2960 250
rect 3030 410 3130 430
rect 3030 350 3050 410
rect 3110 350 3130 410
rect 3030 310 3130 350
rect 3030 250 3050 310
rect 3110 250 3130 310
rect 3030 230 3130 250
rect 3200 410 3300 430
rect 3200 350 3220 410
rect 3280 350 3300 410
rect 3200 310 3300 350
rect 3200 250 3220 310
rect 3280 250 3300 310
rect 3200 230 3300 250
rect 3370 410 3470 430
rect 3370 350 3390 410
rect 3450 350 3470 410
rect 3370 310 3470 350
rect 3370 250 3390 310
rect 3450 250 3470 310
rect 3370 230 3470 250
rect 3540 410 3640 430
rect 3540 350 3560 410
rect 3620 350 3640 410
rect 3540 310 3640 350
rect 3540 250 3560 310
rect 3620 250 3640 310
rect 3540 230 3640 250
rect 3710 410 3810 430
rect 3710 350 3730 410
rect 3790 350 3810 410
rect 3710 310 3810 350
rect 3710 250 3730 310
rect 3790 250 3810 310
rect 3710 230 3810 250
rect 3880 410 3980 430
rect 3880 350 3900 410
rect 3960 350 3980 410
rect 3880 310 3980 350
rect 3880 250 3900 310
rect 3960 250 3980 310
rect 3880 230 3980 250
rect 4050 410 4150 430
rect 4050 350 4070 410
rect 4130 350 4150 410
rect 4050 310 4150 350
rect 4050 250 4070 310
rect 4130 250 4150 310
rect 4050 230 4150 250
rect 4220 410 4320 430
rect 4220 350 4240 410
rect 4300 350 4320 410
rect 4220 310 4320 350
rect 4220 250 4240 310
rect 4300 250 4320 310
rect 4220 230 4320 250
rect 4520 410 4620 430
rect 4520 350 4540 410
rect 4600 350 4620 410
rect 4520 310 4620 350
rect 4520 250 4540 310
rect 4600 250 4620 310
rect 4520 230 4620 250
rect 4690 410 4790 430
rect 4690 350 4710 410
rect 4770 350 4790 410
rect 4690 310 4790 350
rect 4690 250 4710 310
rect 4770 250 4790 310
rect 4690 230 4790 250
rect 4860 410 4960 430
rect 4860 350 4880 410
rect 4940 350 4960 410
rect 4860 310 4960 350
rect 4860 250 4880 310
rect 4940 250 4960 310
rect 4860 230 4960 250
rect 5030 410 5130 430
rect 5030 350 5050 410
rect 5110 350 5130 410
rect 5030 310 5130 350
rect 5030 250 5050 310
rect 5110 250 5130 310
rect 5030 230 5130 250
rect 5200 410 5300 430
rect 5200 350 5220 410
rect 5280 350 5300 410
rect 5200 310 5300 350
rect 5200 250 5220 310
rect 5280 250 5300 310
rect 5200 230 5300 250
rect 5370 410 5470 430
rect 5370 350 5390 410
rect 5450 350 5470 410
rect 5370 310 5470 350
rect 5370 250 5390 310
rect 5450 250 5470 310
rect 5370 230 5470 250
rect 5540 410 5640 430
rect 5540 350 5560 410
rect 5620 350 5640 410
rect 5540 310 5640 350
rect 5540 250 5560 310
rect 5620 250 5640 310
rect 5540 230 5640 250
rect 5710 410 5810 430
rect 5710 350 5730 410
rect 5790 350 5810 410
rect 5710 310 5810 350
rect 5710 250 5730 310
rect 5790 250 5810 310
rect 5710 230 5810 250
rect 5880 410 5980 430
rect 5880 350 5900 410
rect 5960 350 5980 410
rect 5880 310 5980 350
rect 5880 250 5900 310
rect 5960 250 5980 310
rect 5880 230 5980 250
rect 6050 410 6150 430
rect 6050 350 6070 410
rect 6130 350 6150 410
rect 6050 310 6150 350
rect 6050 250 6070 310
rect 6130 250 6150 310
rect 6050 230 6150 250
rect 6220 410 6320 430
rect 6220 350 6240 410
rect 6300 350 6320 410
rect 6220 310 6320 350
rect 6220 250 6240 310
rect 6300 250 6320 310
rect 6220 230 6320 250
rect 6390 410 6490 430
rect 6390 350 6410 410
rect 6470 350 6490 410
rect 6390 310 6490 350
rect 6390 250 6410 310
rect 6470 250 6490 310
rect 6390 230 6490 250
rect 6560 410 6660 430
rect 6560 350 6580 410
rect 6640 350 6660 410
rect 6560 310 6660 350
rect 6560 250 6580 310
rect 6640 250 6660 310
rect 6560 230 6660 250
rect 6730 410 6830 430
rect 6730 350 6750 410
rect 6810 350 6830 410
rect 6730 310 6830 350
rect 6730 250 6750 310
rect 6810 250 6830 310
rect 6730 230 6830 250
rect 6900 410 7000 430
rect 6900 350 6920 410
rect 6980 350 7000 410
rect 6900 310 7000 350
rect 6900 250 6920 310
rect 6980 250 7000 310
rect 6900 230 7000 250
rect 7070 410 7170 430
rect 7070 350 7090 410
rect 7150 350 7170 410
rect 7070 310 7170 350
rect 7070 250 7090 310
rect 7150 250 7170 310
rect 7070 230 7170 250
rect 7240 410 7340 430
rect 7240 350 7260 410
rect 7320 350 7340 410
rect 7240 310 7340 350
rect 7240 250 7260 310
rect 7320 250 7340 310
rect 7240 230 7340 250
rect 7410 410 7510 430
rect 7410 350 7430 410
rect 7490 350 7510 410
rect 7410 310 7510 350
rect 7410 250 7430 310
rect 7490 250 7510 310
rect 7410 230 7510 250
rect 7580 410 7680 430
rect 7580 350 7600 410
rect 7660 350 7680 410
rect 7580 310 7680 350
rect 7580 250 7600 310
rect 7660 250 7680 310
rect 7580 230 7680 250
rect 7750 410 7850 430
rect 7750 350 7770 410
rect 7830 350 7850 410
rect 7750 310 7850 350
rect 7750 250 7770 310
rect 7830 250 7850 310
rect 7750 230 7850 250
rect 7920 410 8020 430
rect 7920 350 7940 410
rect 8000 350 8020 410
rect 7920 310 8020 350
rect 7920 250 7940 310
rect 8000 250 8020 310
rect 7920 230 8020 250
rect 8090 410 8190 430
rect 8090 350 8110 410
rect 8170 350 8190 410
rect 8090 310 8190 350
rect 8090 250 8110 310
rect 8170 250 8190 310
rect 8090 230 8190 250
rect 8260 410 8360 430
rect 8260 350 8280 410
rect 8340 350 8360 410
rect 8260 310 8360 350
rect 8260 250 8280 310
rect 8340 250 8360 310
rect 8260 230 8360 250
rect 8430 410 8530 430
rect 8430 350 8450 410
rect 8510 350 8530 410
rect 8430 310 8530 350
rect 8430 250 8450 310
rect 8510 250 8530 310
rect 8430 230 8530 250
rect 8600 410 8700 430
rect 8600 350 8620 410
rect 8680 350 8700 410
rect 8600 310 8700 350
rect 8600 250 8620 310
rect 8680 250 8700 310
rect 8600 230 8700 250
rect 8770 410 8870 430
rect 8770 350 8790 410
rect 8850 350 8870 410
rect 8770 310 8870 350
rect 8770 250 8790 310
rect 8850 250 8870 310
rect 8770 230 8870 250
rect 8940 410 9040 430
rect 8940 350 8960 410
rect 9020 350 9040 410
rect 8940 310 9040 350
rect 8940 250 8960 310
rect 9020 250 9040 310
rect 8940 230 9040 250
rect 9110 410 9210 430
rect 9110 350 9130 410
rect 9190 350 9210 410
rect 9110 310 9210 350
rect 9110 250 9130 310
rect 9190 250 9210 310
rect 9110 230 9210 250
rect 9280 410 9380 430
rect 9280 350 9300 410
rect 9360 350 9380 410
rect 9280 310 9380 350
rect 9280 250 9300 310
rect 9360 250 9380 310
rect 9280 230 9380 250
rect 9450 410 9550 430
rect 9450 350 9470 410
rect 9530 350 9550 410
rect 9450 310 9550 350
rect 9450 250 9470 310
rect 9530 250 9550 310
rect 9450 230 9550 250
rect 9620 410 9720 430
rect 9620 350 9640 410
rect 9700 350 9720 410
rect 9620 310 9720 350
rect 9620 250 9640 310
rect 9700 250 9720 310
rect 9620 230 9720 250
rect 9790 410 9890 430
rect 9790 350 9810 410
rect 9870 350 9890 410
rect 9790 310 9890 350
rect 9790 250 9810 310
rect 9870 250 9890 310
rect 9790 230 9890 250
rect 9960 410 10060 430
rect 9960 350 9980 410
rect 10040 350 10060 410
rect 9960 310 10060 350
rect 9960 250 9980 310
rect 10040 250 10060 310
rect 9960 230 10060 250
rect 10130 410 10230 430
rect 10130 350 10150 410
rect 10210 350 10230 410
rect 10130 310 10230 350
rect 10130 250 10150 310
rect 10210 250 10230 310
rect 10130 230 10230 250
rect 10300 410 10400 430
rect 10300 350 10320 410
rect 10380 350 10400 410
rect 10300 310 10400 350
rect 10300 250 10320 310
rect 10380 250 10400 310
rect 10300 230 10400 250
rect 10470 410 10570 430
rect 10470 350 10490 410
rect 10550 350 10570 410
rect 10470 310 10570 350
rect 10470 250 10490 310
rect 10550 250 10570 310
rect 10470 230 10570 250
rect 10640 410 10740 430
rect 10640 350 10660 410
rect 10720 350 10740 410
rect 10640 310 10740 350
rect 10640 250 10660 310
rect 10720 250 10740 310
rect 10640 230 10740 250
rect 10810 410 10910 430
rect 10810 350 10830 410
rect 10890 350 10910 410
rect 10810 310 10910 350
rect 10810 250 10830 310
rect 10890 250 10910 310
rect 10810 230 10910 250
rect 10980 410 11080 430
rect 10980 350 11000 410
rect 11060 350 11080 410
rect 10980 310 11080 350
rect 10980 250 11000 310
rect 11060 250 11080 310
rect 10980 230 11080 250
rect 11150 410 11250 430
rect 11150 350 11170 410
rect 11230 350 11250 410
rect 11150 310 11250 350
rect 11150 250 11170 310
rect 11230 250 11250 310
rect 11150 230 11250 250
rect 11320 410 11420 430
rect 11320 350 11340 410
rect 11400 350 11420 410
rect 11320 310 11420 350
rect 11320 250 11340 310
rect 11400 250 11420 310
rect 11320 230 11420 250
rect 11490 410 11590 430
rect 11490 350 11510 410
rect 11570 350 11590 410
rect 11490 310 11590 350
rect 11490 250 11510 310
rect 11570 250 11590 310
rect 11490 230 11590 250
rect 11660 410 11760 430
rect 11660 350 11680 410
rect 11740 350 11760 410
rect 11660 310 11760 350
rect 11660 250 11680 310
rect 11740 250 11760 310
rect 11660 230 11760 250
rect 11830 410 11930 430
rect 11830 350 11850 410
rect 11910 350 11930 410
rect 11830 310 11930 350
rect 11830 250 11850 310
rect 11910 250 11930 310
rect 11830 230 11930 250
rect 12000 410 12100 430
rect 12000 350 12020 410
rect 12080 350 12100 410
rect 12000 310 12100 350
rect 12000 250 12020 310
rect 12080 250 12100 310
rect 12000 230 12100 250
rect 12170 410 12270 430
rect 12170 350 12190 410
rect 12250 350 12270 410
rect 12170 310 12270 350
rect 12170 250 12190 310
rect 12250 250 12270 310
rect 12170 230 12270 250
rect 12340 410 12440 430
rect 12340 350 12360 410
rect 12420 350 12440 410
rect 12340 310 12440 350
rect 12340 250 12360 310
rect 12420 250 12440 310
rect 12340 230 12440 250
rect 12510 410 12610 430
rect 12510 350 12530 410
rect 12590 350 12610 410
rect 12510 310 12610 350
rect 12510 250 12530 310
rect 12590 250 12610 310
rect 12510 230 12610 250
rect 12680 410 12780 430
rect 12680 350 12700 410
rect 12760 350 12780 410
rect 12680 310 12780 350
rect 12680 250 12700 310
rect 12760 250 12780 310
rect 12680 230 12780 250
rect 12850 410 12950 430
rect 12850 350 12870 410
rect 12930 350 12950 410
rect 12850 310 12950 350
rect 12850 250 12870 310
rect 12930 250 12950 310
rect 12850 230 12950 250
rect 13020 410 13120 430
rect 13020 350 13040 410
rect 13100 350 13120 410
rect 13020 310 13120 350
rect 13020 250 13040 310
rect 13100 250 13120 310
rect 13020 230 13120 250
rect 13190 410 13290 430
rect 13190 350 13210 410
rect 13270 350 13290 410
rect 13190 310 13290 350
rect 13190 250 13210 310
rect 13270 250 13290 310
rect 13190 230 13290 250
rect 13360 410 13460 430
rect 13360 350 13380 410
rect 13440 350 13460 410
rect 13360 310 13460 350
rect 13360 250 13380 310
rect 13440 250 13460 310
rect 13360 230 13460 250
rect 13530 410 13630 430
rect 13530 350 13550 410
rect 13610 350 13630 410
rect 13530 310 13630 350
rect 13530 250 13550 310
rect 13610 250 13630 310
rect 13530 230 13630 250
rect 13700 410 13800 430
rect 13700 350 13720 410
rect 13780 350 13800 410
rect 13700 310 13800 350
rect 13700 250 13720 310
rect 13780 250 13800 310
rect 13700 230 13800 250
rect 13870 410 13970 430
rect 13870 350 13890 410
rect 13950 350 13970 410
rect 13870 310 13970 350
rect 13870 250 13890 310
rect 13950 250 13970 310
rect 13870 230 13970 250
rect 14040 410 14140 430
rect 14040 350 14060 410
rect 14120 350 14140 410
rect 14040 310 14140 350
rect 14040 250 14060 310
rect 14120 250 14140 310
rect 14040 230 14140 250
rect 14210 410 14310 430
rect 14210 350 14230 410
rect 14290 350 14310 410
rect 14210 310 14310 350
rect 14210 250 14230 310
rect 14290 250 14310 310
rect 14210 230 14310 250
rect 14380 410 14480 430
rect 14380 350 14400 410
rect 14460 350 14480 410
rect 14380 310 14480 350
rect 14380 250 14400 310
rect 14460 250 14480 310
rect 14380 230 14480 250
rect 14550 410 14650 430
rect 14550 350 14570 410
rect 14630 350 14650 410
rect 14550 310 14650 350
rect 14550 250 14570 310
rect 14630 250 14650 310
rect 14550 230 14650 250
rect 14720 410 14820 430
rect 14720 350 14740 410
rect 14800 350 14820 410
rect 14720 310 14820 350
rect 14720 250 14740 310
rect 14800 250 14820 310
rect 14720 230 14820 250
rect 14890 410 14990 430
rect 14890 350 14910 410
rect 14970 350 14990 410
rect 14890 310 14990 350
rect 14890 250 14910 310
rect 14970 250 14990 310
rect 14890 230 14990 250
rect 15060 410 15160 430
rect 15060 350 15080 410
rect 15140 350 15160 410
rect 15060 310 15160 350
rect 15060 250 15080 310
rect 15140 250 15160 310
rect 15060 230 15160 250
rect 15230 410 15330 430
rect 15230 350 15250 410
rect 15310 350 15330 410
rect 15230 310 15330 350
rect 15230 250 15250 310
rect 15310 250 15330 310
rect 15230 230 15330 250
rect 15400 410 15500 430
rect 15400 350 15420 410
rect 15480 350 15500 410
rect 15400 310 15500 350
rect 15400 250 15420 310
rect 15480 250 15500 310
rect 15400 230 15500 250
rect 15700 410 15800 430
rect 15700 350 15720 410
rect 15780 350 15800 410
rect 15700 310 15800 350
rect 15700 250 15720 310
rect 15780 250 15800 310
rect 15700 230 15800 250
rect 15870 410 15970 430
rect 15870 350 15890 410
rect 15950 350 15970 410
rect 15870 310 15970 350
rect 15870 250 15890 310
rect 15950 250 15970 310
rect 15870 230 15970 250
rect 16040 410 16140 430
rect 16040 350 16060 410
rect 16120 350 16140 410
rect 16040 310 16140 350
rect 16040 250 16060 310
rect 16120 250 16140 310
rect 16040 230 16140 250
rect 16210 410 16310 430
rect 16210 350 16230 410
rect 16290 350 16310 410
rect 16210 310 16310 350
rect 16210 250 16230 310
rect 16290 250 16310 310
rect 16210 230 16310 250
rect 16380 410 16480 430
rect 16380 350 16400 410
rect 16460 350 16480 410
rect 16380 310 16480 350
rect 16380 250 16400 310
rect 16460 250 16480 310
rect 16380 230 16480 250
rect 16550 410 16650 430
rect 16550 350 16570 410
rect 16630 350 16650 410
rect 16550 310 16650 350
rect 16550 250 16570 310
rect 16630 250 16650 310
rect 16550 230 16650 250
rect 16720 410 16820 430
rect 16720 350 16740 410
rect 16800 350 16820 410
rect 16720 310 16820 350
rect 16720 250 16740 310
rect 16800 250 16820 310
rect 16720 230 16820 250
rect 16890 410 16990 430
rect 16890 350 16910 410
rect 16970 350 16990 410
rect 16890 310 16990 350
rect 16890 250 16910 310
rect 16970 250 16990 310
rect 16890 230 16990 250
rect 17060 410 17160 430
rect 17060 350 17080 410
rect 17140 350 17160 410
rect 17060 310 17160 350
rect 17060 250 17080 310
rect 17140 250 17160 310
rect 17060 230 17160 250
rect 17230 410 17330 430
rect 17230 350 17250 410
rect 17310 350 17330 410
rect 17230 310 17330 350
rect 17230 250 17250 310
rect 17310 250 17330 310
rect 17230 230 17330 250
rect 17400 410 17500 430
rect 17400 350 17420 410
rect 17480 350 17500 410
rect 17400 310 17500 350
rect 17400 250 17420 310
rect 17480 250 17500 310
rect 17400 230 17500 250
rect 17570 410 17670 430
rect 17570 350 17590 410
rect 17650 350 17670 410
rect 17570 310 17670 350
rect 17570 250 17590 310
rect 17650 250 17670 310
rect 17570 230 17670 250
rect 17740 410 17840 430
rect 17740 350 17760 410
rect 17820 350 17840 410
rect 17740 310 17840 350
rect 17740 250 17760 310
rect 17820 250 17840 310
rect 17740 230 17840 250
rect 17910 410 18010 430
rect 17910 350 17930 410
rect 17990 350 18010 410
rect 17910 310 18010 350
rect 17910 250 17930 310
rect 17990 250 18010 310
rect 17910 230 18010 250
rect 18080 410 18180 430
rect 18080 350 18100 410
rect 18160 350 18180 410
rect 18080 310 18180 350
rect 18080 250 18100 310
rect 18160 250 18180 310
rect 18080 230 18180 250
rect 18250 410 18350 430
rect 18250 350 18270 410
rect 18330 350 18350 410
rect 18250 310 18350 350
rect 18250 250 18270 310
rect 18330 250 18350 310
rect 18250 230 18350 250
rect 18420 410 18520 430
rect 18420 350 18440 410
rect 18500 350 18520 410
rect 18420 310 18520 350
rect 18420 250 18440 310
rect 18500 250 18520 310
rect 18420 230 18520 250
rect 18590 410 18690 430
rect 18590 350 18610 410
rect 18670 350 18690 410
rect 18590 310 18690 350
rect 18590 250 18610 310
rect 18670 250 18690 310
rect 18590 230 18690 250
rect 18760 410 18860 430
rect 18760 350 18780 410
rect 18840 350 18860 410
rect 18760 310 18860 350
rect 18760 250 18780 310
rect 18840 250 18860 310
rect 18760 230 18860 250
rect 18930 410 19030 430
rect 18930 350 18950 410
rect 19010 350 19030 410
rect 18930 310 19030 350
rect 18930 250 18950 310
rect 19010 250 19030 310
rect 18930 230 19030 250
rect 19100 410 19200 430
rect 19100 350 19120 410
rect 19180 350 19200 410
rect 19100 310 19200 350
rect 19100 250 19120 310
rect 19180 250 19200 310
rect 19100 230 19200 250
rect 19270 410 19370 430
rect 19270 350 19290 410
rect 19350 350 19370 410
rect 19270 310 19370 350
rect 19270 250 19290 310
rect 19350 250 19370 310
rect 19270 230 19370 250
rect 19440 410 19540 430
rect 19440 350 19460 410
rect 19520 350 19540 410
rect 19440 310 19540 350
rect 19440 250 19460 310
rect 19520 250 19540 310
rect 19440 230 19540 250
rect 19610 410 19710 430
rect 19610 350 19630 410
rect 19690 350 19710 410
rect 19610 310 19710 350
rect 19610 250 19630 310
rect 19690 250 19710 310
rect 19610 230 19710 250
rect 19780 410 19880 430
rect 19780 350 19800 410
rect 19860 350 19880 410
rect 19780 310 19880 350
rect 19780 250 19800 310
rect 19860 250 19880 310
rect 19780 230 19880 250
rect 19950 410 20050 430
rect 19950 350 19970 410
rect 20030 350 20050 410
rect 19950 310 20050 350
rect 19950 250 19970 310
rect 20030 250 20050 310
rect 19950 230 20050 250
rect 20120 410 20220 430
rect 20120 350 20140 410
rect 20200 350 20220 410
rect 20120 310 20220 350
rect 20120 250 20140 310
rect 20200 250 20220 310
rect 20120 230 20220 250
rect 20290 410 20390 430
rect 20290 350 20310 410
rect 20370 350 20390 410
rect 20290 310 20390 350
rect 20290 250 20310 310
rect 20370 250 20390 310
rect 20290 230 20390 250
rect 20460 410 20560 430
rect 20460 350 20480 410
rect 20540 350 20560 410
rect 20460 310 20560 350
rect 20460 250 20480 310
rect 20540 250 20560 310
rect 20460 230 20560 250
rect 20630 410 20730 430
rect 20630 350 20650 410
rect 20710 350 20730 410
rect 20630 310 20730 350
rect 20630 250 20650 310
rect 20710 250 20730 310
rect 20630 230 20730 250
rect 20800 410 20900 430
rect 20800 350 20820 410
rect 20880 350 20900 410
rect 20800 310 20900 350
rect 20800 250 20820 310
rect 20880 250 20900 310
rect 20800 230 20900 250
rect 20970 410 21070 430
rect 20970 350 20990 410
rect 21050 350 21070 410
rect 20970 310 21070 350
rect 20970 250 20990 310
rect 21050 250 21070 310
rect 20970 230 21070 250
rect 21140 410 21240 430
rect 21140 350 21160 410
rect 21220 350 21240 410
rect 21140 310 21240 350
rect 21140 250 21160 310
rect 21220 250 21240 310
rect 21140 230 21240 250
rect 21310 410 21410 430
rect 21310 350 21330 410
rect 21390 350 21410 410
rect 21310 310 21410 350
rect 21310 250 21330 310
rect 21390 250 21410 310
rect 21310 230 21410 250
rect 21480 410 21580 430
rect 21480 350 21500 410
rect 21560 350 21580 410
rect 21480 310 21580 350
rect 21480 250 21500 310
rect 21560 250 21580 310
rect 21480 230 21580 250
rect 21650 410 21750 430
rect 21650 350 21670 410
rect 21730 350 21750 410
rect 21650 310 21750 350
rect 21650 250 21670 310
rect 21730 250 21750 310
rect 21650 230 21750 250
rect 21820 410 21920 430
rect 21820 350 21840 410
rect 21900 350 21920 410
rect 21820 310 21920 350
rect 21820 250 21840 310
rect 21900 250 21920 310
rect 21820 230 21920 250
rect 21990 410 22090 430
rect 21990 350 22010 410
rect 22070 350 22090 410
rect 21990 310 22090 350
rect 21990 250 22010 310
rect 22070 250 22090 310
rect 21990 230 22090 250
rect 22160 410 22260 430
rect 22160 350 22180 410
rect 22240 350 22260 410
rect 22160 310 22260 350
rect 22160 250 22180 310
rect 22240 250 22260 310
rect 22160 230 22260 250
rect 22330 410 22430 430
rect 22330 350 22350 410
rect 22410 350 22430 410
rect 22330 310 22430 350
rect 22330 250 22350 310
rect 22410 250 22430 310
rect 22330 230 22430 250
rect 22500 410 22600 430
rect 22500 350 22520 410
rect 22580 350 22600 410
rect 22500 310 22600 350
rect 22500 250 22520 310
rect 22580 250 22600 310
rect 22500 230 22600 250
rect 22670 410 22770 430
rect 22670 350 22690 410
rect 22750 350 22770 410
rect 22670 310 22770 350
rect 22670 250 22690 310
rect 22750 250 22770 310
rect 22670 230 22770 250
rect 22840 410 22940 430
rect 22840 350 22860 410
rect 22920 350 22940 410
rect 22840 310 22940 350
rect 22840 250 22860 310
rect 22920 250 22940 310
rect 22840 230 22940 250
rect 23010 410 23110 430
rect 23010 350 23030 410
rect 23090 350 23110 410
rect 23010 310 23110 350
rect 23010 250 23030 310
rect 23090 250 23110 310
rect 23010 230 23110 250
rect 23180 410 23280 430
rect 23180 350 23200 410
rect 23260 350 23280 410
rect 23180 310 23280 350
rect 23180 250 23200 310
rect 23260 250 23280 310
rect 23180 230 23280 250
rect 23350 410 23450 430
rect 23350 350 23370 410
rect 23430 350 23450 410
rect 23350 310 23450 350
rect 23350 250 23370 310
rect 23430 250 23450 310
rect 23350 230 23450 250
rect 23520 410 23620 430
rect 23520 350 23540 410
rect 23600 350 23620 410
rect 23520 310 23620 350
rect 23520 250 23540 310
rect 23600 250 23620 310
rect 23520 230 23620 250
rect 23690 410 23790 430
rect 23690 350 23710 410
rect 23770 350 23790 410
rect 23690 310 23790 350
rect 23690 250 23710 310
rect 23770 250 23790 310
rect 23690 230 23790 250
rect 23860 410 23960 430
rect 23860 350 23880 410
rect 23940 350 23960 410
rect 23860 310 23960 350
rect 23860 250 23880 310
rect 23940 250 23960 310
rect 23860 230 23960 250
rect 24030 410 24130 430
rect 24030 350 24050 410
rect 24110 350 24130 410
rect 24030 310 24130 350
rect 24030 250 24050 310
rect 24110 250 24130 310
rect 24030 230 24130 250
rect 24200 410 24300 430
rect 24200 350 24220 410
rect 24280 350 24300 410
rect 24200 310 24300 350
rect 24200 250 24220 310
rect 24280 250 24300 310
rect 24200 230 24300 250
rect 24370 410 24470 430
rect 24370 350 24390 410
rect 24450 350 24470 410
rect 24370 310 24470 350
rect 24370 250 24390 310
rect 24450 250 24470 310
rect 24370 230 24470 250
rect 24540 410 24640 430
rect 24540 350 24560 410
rect 24620 350 24640 410
rect 24540 310 24640 350
rect 24540 250 24560 310
rect 24620 250 24640 310
rect 24540 230 24640 250
rect 24710 410 24810 430
rect 24710 350 24730 410
rect 24790 350 24810 410
rect 24710 310 24810 350
rect 24710 250 24730 310
rect 24790 250 24810 310
rect 24710 230 24810 250
rect 24880 410 24980 430
rect 24880 350 24900 410
rect 24960 350 24980 410
rect 24880 310 24980 350
rect 24880 250 24900 310
rect 24960 250 24980 310
rect 24880 230 24980 250
rect 25050 410 25150 430
rect 25050 350 25070 410
rect 25130 350 25150 410
rect 25050 310 25150 350
rect 25050 250 25070 310
rect 25130 250 25150 310
rect 25050 230 25150 250
rect 25220 410 25320 430
rect 25220 350 25240 410
rect 25300 350 25320 410
rect 25220 310 25320 350
rect 25220 250 25240 310
rect 25300 250 25320 310
rect 25220 230 25320 250
rect 25390 410 25490 430
rect 25390 350 25410 410
rect 25470 350 25490 410
rect 25390 310 25490 350
rect 25390 250 25410 310
rect 25470 250 25490 310
rect 25390 230 25490 250
rect 25560 410 25660 430
rect 25560 350 25580 410
rect 25640 350 25660 410
rect 25560 310 25660 350
rect 25560 250 25580 310
rect 25640 250 25660 310
rect 25560 230 25660 250
rect 25730 410 25830 430
rect 25730 350 25750 410
rect 25810 350 25830 410
rect 25730 310 25830 350
rect 25730 250 25750 310
rect 25810 250 25830 310
rect 25730 230 25830 250
rect 25900 410 26000 430
rect 25900 350 25920 410
rect 25980 350 26000 410
rect 25900 310 26000 350
rect 25900 250 25920 310
rect 25980 250 26000 310
rect 25900 230 26000 250
rect 26070 410 26170 430
rect 26070 350 26090 410
rect 26150 350 26170 410
rect 26070 310 26170 350
rect 26070 250 26090 310
rect 26150 250 26170 310
rect 26070 230 26170 250
rect 26240 410 26340 430
rect 26240 350 26260 410
rect 26320 350 26340 410
rect 26240 310 26340 350
rect 26240 250 26260 310
rect 26320 250 26340 310
rect 26240 230 26340 250
rect 26410 410 26510 430
rect 26410 350 26430 410
rect 26490 350 26510 410
rect 26410 310 26510 350
rect 26410 250 26430 310
rect 26490 250 26510 310
rect 26410 230 26510 250
rect 26580 410 26680 430
rect 26580 350 26600 410
rect 26660 350 26680 410
rect 26580 310 26680 350
rect 26580 250 26600 310
rect 26660 250 26680 310
rect 26580 230 26680 250
rect 26750 410 26850 430
rect 26750 350 26770 410
rect 26830 350 26850 410
rect 26750 310 26850 350
rect 26750 250 26770 310
rect 26830 250 26850 310
rect 26750 230 26850 250
rect 26920 410 27020 430
rect 26920 350 26940 410
rect 27000 350 27020 410
rect 26920 310 27020 350
rect 26920 250 26940 310
rect 27000 250 27020 310
rect 26920 230 27020 250
rect 27090 410 27190 430
rect 27090 350 27110 410
rect 27170 350 27190 410
rect 27090 310 27190 350
rect 27090 250 27110 310
rect 27170 250 27190 310
rect 27090 230 27190 250
rect 27260 410 27360 430
rect 27260 350 27280 410
rect 27340 350 27360 410
rect 27260 310 27360 350
rect 27260 250 27280 310
rect 27340 250 27360 310
rect 27260 230 27360 250
rect 27430 410 27530 430
rect 27430 350 27450 410
rect 27510 350 27530 410
rect 27430 310 27530 350
rect 27430 250 27450 310
rect 27510 250 27530 310
rect 27430 230 27530 250
rect 27600 410 27700 430
rect 27600 350 27620 410
rect 27680 350 27700 410
rect 27600 310 27700 350
rect 27600 250 27620 310
rect 27680 250 27700 310
rect 27600 230 27700 250
rect 27770 410 27870 430
rect 27770 350 27790 410
rect 27850 350 27870 410
rect 27770 310 27870 350
rect 27770 250 27790 310
rect 27850 250 27870 310
rect 27770 230 27870 250
rect 27940 410 28040 430
rect 27940 350 27960 410
rect 28020 350 28040 410
rect 27940 310 28040 350
rect 27940 250 27960 310
rect 28020 250 28040 310
rect 27940 230 28040 250
rect 28110 410 28210 430
rect 28110 350 28130 410
rect 28190 350 28210 410
rect 28110 310 28210 350
rect 28110 250 28130 310
rect 28190 250 28210 310
rect 28110 230 28210 250
rect 28280 410 28380 430
rect 28280 350 28300 410
rect 28360 350 28380 410
rect 28280 310 28380 350
rect 28280 250 28300 310
rect 28360 250 28380 310
rect 28280 230 28380 250
rect 28450 410 28550 430
rect 28450 350 28470 410
rect 28530 350 28550 410
rect 28450 310 28550 350
rect 28450 250 28470 310
rect 28530 250 28550 310
rect 28450 230 28550 250
rect 28620 410 28720 430
rect 28620 350 28640 410
rect 28700 350 28720 410
rect 28620 310 28720 350
rect 28620 250 28640 310
rect 28700 250 28720 310
rect 28620 230 28720 250
rect 28790 410 28890 430
rect 28790 350 28810 410
rect 28870 350 28890 410
rect 28790 310 28890 350
rect 28790 250 28810 310
rect 28870 250 28890 310
rect 28790 230 28890 250
rect 28960 410 29060 430
rect 28960 350 28980 410
rect 29040 350 29060 410
rect 28960 310 29060 350
rect 28960 250 28980 310
rect 29040 250 29060 310
rect 28960 230 29060 250
rect 29130 410 29230 430
rect 29130 350 29150 410
rect 29210 350 29230 410
rect 29130 310 29230 350
rect 29130 250 29150 310
rect 29210 250 29230 310
rect 29130 230 29230 250
rect 29300 410 29400 430
rect 29300 350 29320 410
rect 29380 350 29400 410
rect 29300 310 29400 350
rect 29300 250 29320 310
rect 29380 250 29400 310
rect 29300 230 29400 250
rect 29470 410 29570 430
rect 29470 350 29490 410
rect 29550 350 29570 410
rect 29470 310 29570 350
rect 29470 250 29490 310
rect 29550 250 29570 310
rect 29470 230 29570 250
rect 29640 410 29740 430
rect 29640 350 29660 410
rect 29720 350 29740 410
rect 29640 310 29740 350
rect 29640 250 29660 310
rect 29720 250 29740 310
rect 29640 230 29740 250
rect 29810 410 29910 430
rect 29810 350 29830 410
rect 29890 350 29910 410
rect 29810 310 29910 350
rect 29810 250 29830 310
rect 29890 250 29910 310
rect 29810 230 29910 250
rect 29980 410 30080 430
rect 29980 350 30000 410
rect 30060 350 30080 410
rect 29980 310 30080 350
rect 29980 250 30000 310
rect 30060 250 30080 310
rect 29980 230 30080 250
rect 30150 410 30250 430
rect 30150 350 30170 410
rect 30230 350 30250 410
rect 30150 310 30250 350
rect 30150 250 30170 310
rect 30230 250 30250 310
rect 30150 230 30250 250
rect 30320 410 30420 430
rect 30320 350 30340 410
rect 30400 350 30420 410
rect 30320 310 30420 350
rect 30320 250 30340 310
rect 30400 250 30420 310
rect 30320 230 30420 250
rect 30490 410 30590 430
rect 30490 350 30510 410
rect 30570 350 30590 410
rect 30490 310 30590 350
rect 30490 250 30510 310
rect 30570 250 30590 310
rect 30490 230 30590 250
rect 30660 410 30760 430
rect 30660 350 30680 410
rect 30740 350 30760 410
rect 30660 310 30760 350
rect 30660 250 30680 310
rect 30740 250 30760 310
rect 30660 230 30760 250
rect 30830 410 30930 430
rect 30830 350 30850 410
rect 30910 350 30930 410
rect 30830 310 30930 350
rect 30830 250 30850 310
rect 30910 250 30930 310
rect 30830 230 30930 250
rect 31000 410 31100 430
rect 31000 350 31020 410
rect 31080 350 31100 410
rect 31000 310 31100 350
rect 31000 250 31020 310
rect 31080 250 31100 310
rect 31000 230 31100 250
rect 31170 410 31270 430
rect 31170 350 31190 410
rect 31250 350 31270 410
rect 31170 310 31270 350
rect 31170 250 31190 310
rect 31250 250 31270 310
rect 31170 230 31270 250
rect 31340 410 31440 430
rect 31340 350 31360 410
rect 31420 350 31440 410
rect 31340 310 31440 350
rect 31340 250 31360 310
rect 31420 250 31440 310
rect 31340 230 31440 250
rect 31510 410 31610 430
rect 31510 350 31530 410
rect 31590 350 31610 410
rect 31510 310 31610 350
rect 31510 250 31530 310
rect 31590 250 31610 310
rect 31510 230 31610 250
rect 31680 410 31780 430
rect 31680 350 31700 410
rect 31760 350 31780 410
rect 31680 310 31780 350
rect 31680 250 31700 310
rect 31760 250 31780 310
rect 31680 230 31780 250
rect 31850 410 31950 430
rect 31850 350 31870 410
rect 31930 350 31950 410
rect 31850 310 31950 350
rect 31850 250 31870 310
rect 31930 250 31950 310
rect 31850 230 31950 250
rect 32020 410 32120 430
rect 32020 350 32040 410
rect 32100 350 32120 410
rect 32020 310 32120 350
rect 32020 250 32040 310
rect 32100 250 32120 310
rect 32020 230 32120 250
rect 32190 410 32290 430
rect 32190 350 32210 410
rect 32270 350 32290 410
rect 32190 310 32290 350
rect 32190 250 32210 310
rect 32270 250 32290 310
rect 32190 230 32290 250
rect 32360 410 32460 430
rect 32360 350 32380 410
rect 32440 350 32460 410
rect 32360 310 32460 350
rect 32360 250 32380 310
rect 32440 250 32460 310
rect 32360 230 32460 250
rect 32530 410 32630 430
rect 32530 350 32550 410
rect 32610 350 32630 410
rect 32530 310 32630 350
rect 32530 250 32550 310
rect 32610 250 32630 310
rect 32530 230 32630 250
rect 32700 410 32800 430
rect 32700 350 32720 410
rect 32780 350 32800 410
rect 32700 310 32800 350
rect 32700 250 32720 310
rect 32780 250 32800 310
rect 32700 230 32800 250
rect 32870 410 32970 430
rect 32870 350 32890 410
rect 32950 350 32970 410
rect 32870 310 32970 350
rect 32870 250 32890 310
rect 32950 250 32970 310
rect 32870 230 32970 250
rect 33040 410 33140 430
rect 33040 350 33060 410
rect 33120 350 33140 410
rect 33040 310 33140 350
rect 33040 250 33060 310
rect 33120 250 33140 310
rect 33040 230 33140 250
rect 33210 410 33310 430
rect 33210 350 33230 410
rect 33290 350 33310 410
rect 33210 310 33310 350
rect 33210 250 33230 310
rect 33290 250 33310 310
rect 33210 230 33310 250
rect 33380 410 33480 430
rect 33380 350 33400 410
rect 33460 350 33480 410
rect 33380 310 33480 350
rect 33380 250 33400 310
rect 33460 250 33480 310
rect 33380 230 33480 250
rect 33550 410 33650 430
rect 33550 350 33570 410
rect 33630 350 33650 410
rect 33550 310 33650 350
rect 33550 250 33570 310
rect 33630 250 33650 310
rect 33550 230 33650 250
rect 33720 410 33820 430
rect 33720 350 33740 410
rect 33800 350 33820 410
rect 33720 310 33820 350
rect 33720 250 33740 310
rect 33800 250 33820 310
rect 33720 230 33820 250
rect 33890 410 33990 430
rect 33890 350 33910 410
rect 33970 350 33990 410
rect 33890 310 33990 350
rect 33890 250 33910 310
rect 33970 250 33990 310
rect 33890 230 33990 250
rect 34060 410 34160 430
rect 34060 350 34080 410
rect 34140 350 34160 410
rect 34060 310 34160 350
rect 34060 250 34080 310
rect 34140 250 34160 310
rect 34060 230 34160 250
rect 34230 410 34330 430
rect 34230 350 34250 410
rect 34310 350 34330 410
rect 34230 310 34330 350
rect 34230 250 34250 310
rect 34310 250 34330 310
rect 34230 230 34330 250
rect 34400 410 34500 430
rect 34400 350 34420 410
rect 34480 350 34500 410
rect 34400 310 34500 350
rect 34400 250 34420 310
rect 34480 250 34500 310
rect 34400 230 34500 250
rect 34570 410 34670 430
rect 34570 350 34590 410
rect 34650 350 34670 410
rect 34570 310 34670 350
rect 34570 250 34590 310
rect 34650 250 34670 310
rect 34570 230 34670 250
rect 34740 410 34840 430
rect 34740 350 34760 410
rect 34820 350 34840 410
rect 34740 310 34840 350
rect 34740 250 34760 310
rect 34820 250 34840 310
rect 34740 230 34840 250
rect 34910 410 35010 430
rect 34910 350 34930 410
rect 34990 350 35010 410
rect 34910 310 35010 350
rect 34910 250 34930 310
rect 34990 250 35010 310
rect 34910 230 35010 250
rect 35080 410 35180 430
rect 35080 350 35100 410
rect 35160 350 35180 410
rect 35080 310 35180 350
rect 35080 250 35100 310
rect 35160 250 35180 310
rect 35080 230 35180 250
rect 35250 410 35350 430
rect 35250 350 35270 410
rect 35330 350 35350 410
rect 35250 310 35350 350
rect 35250 250 35270 310
rect 35330 250 35350 310
rect 35250 230 35350 250
rect 35420 410 35520 430
rect 35420 350 35440 410
rect 35500 350 35520 410
rect 35420 310 35520 350
rect 35420 250 35440 310
rect 35500 250 35520 310
rect 35420 230 35520 250
rect 35590 410 35690 430
rect 35590 350 35610 410
rect 35670 350 35690 410
rect 35590 310 35690 350
rect 35590 250 35610 310
rect 35670 250 35690 310
rect 35590 230 35690 250
rect 35760 410 35860 430
rect 35760 350 35780 410
rect 35840 350 35860 410
rect 35760 310 35860 350
rect 35760 250 35780 310
rect 35840 250 35860 310
rect 35760 230 35860 250
rect 35930 410 36030 430
rect 35930 350 35950 410
rect 36010 350 36030 410
rect 35930 310 36030 350
rect 35930 250 35950 310
rect 36010 250 36030 310
rect 35930 230 36030 250
rect 36100 410 36200 430
rect 36100 350 36120 410
rect 36180 350 36200 410
rect 36100 310 36200 350
rect 36100 250 36120 310
rect 36180 250 36200 310
rect 36100 230 36200 250
rect 36270 410 36370 430
rect 36270 350 36290 410
rect 36350 350 36370 410
rect 36270 310 36370 350
rect 36270 250 36290 310
rect 36350 250 36370 310
rect 36270 230 36370 250
rect 36440 410 36540 430
rect 36440 350 36460 410
rect 36520 350 36540 410
rect 36440 310 36540 350
rect 36440 250 36460 310
rect 36520 250 36540 310
rect 36440 230 36540 250
rect 36610 410 36710 430
rect 36610 350 36630 410
rect 36690 350 36710 410
rect 36610 310 36710 350
rect 36610 250 36630 310
rect 36690 250 36710 310
rect 36610 230 36710 250
rect 36780 410 36880 430
rect 36780 350 36800 410
rect 36860 350 36880 410
rect 36780 310 36880 350
rect 36780 250 36800 310
rect 36860 250 36880 310
rect 36780 230 36880 250
rect 36950 410 37050 430
rect 36950 350 36970 410
rect 37030 350 37050 410
rect 36950 310 37050 350
rect 36950 250 36970 310
rect 37030 250 37050 310
rect 36950 230 37050 250
rect 37120 410 37220 430
rect 37120 350 37140 410
rect 37200 350 37220 410
rect 37120 310 37220 350
rect 37120 250 37140 310
rect 37200 250 37220 310
rect 37120 230 37220 250
rect 37290 410 37390 430
rect 37290 350 37310 410
rect 37370 350 37390 410
rect 37290 310 37390 350
rect 37290 250 37310 310
rect 37370 250 37390 310
rect 37290 230 37390 250
rect 37460 410 37560 430
rect 37460 350 37480 410
rect 37540 350 37560 410
rect 37460 310 37560 350
rect 37460 250 37480 310
rect 37540 250 37560 310
rect 37460 230 37560 250
rect 37630 410 37730 430
rect 37630 350 37650 410
rect 37710 350 37730 410
rect 37630 310 37730 350
rect 37630 250 37650 310
rect 37710 250 37730 310
rect 37630 230 37730 250
rect 37800 410 37900 430
rect 37800 350 37820 410
rect 37880 350 37900 410
rect 37800 310 37900 350
rect 37800 250 37820 310
rect 37880 250 37900 310
rect 37800 230 37900 250
rect 37970 410 38070 430
rect 37970 350 37990 410
rect 38050 350 38070 410
rect 37970 310 38070 350
rect 37970 250 37990 310
rect 38050 250 38070 310
rect 37970 230 38070 250
rect 38140 410 38240 430
rect 38140 350 38160 410
rect 38220 350 38240 410
rect 38140 310 38240 350
rect 38140 250 38160 310
rect 38220 250 38240 310
rect 38140 230 38240 250
rect 38310 410 38410 430
rect 38310 350 38330 410
rect 38390 350 38410 410
rect 38310 310 38410 350
rect 38310 250 38330 310
rect 38390 250 38410 310
rect 38310 230 38410 250
rect 38480 410 38580 430
rect 38480 350 38500 410
rect 38560 350 38580 410
rect 38480 310 38580 350
rect 38480 250 38500 310
rect 38560 250 38580 310
rect 38480 230 38580 250
rect 38650 410 38750 430
rect 38650 350 38670 410
rect 38730 350 38750 410
rect 38650 310 38750 350
rect 38650 250 38670 310
rect 38730 250 38750 310
rect 38650 230 38750 250
rect 38820 410 38920 430
rect 38820 350 38840 410
rect 38900 350 38920 410
rect 38820 310 38920 350
rect 38820 250 38840 310
rect 38900 250 38920 310
rect 38820 230 38920 250
rect 38990 410 39090 430
rect 38990 350 39010 410
rect 39070 350 39090 410
rect 38990 310 39090 350
rect 38990 250 39010 310
rect 39070 250 39090 310
rect 38990 230 39090 250
rect 39160 410 39260 430
rect 39160 350 39180 410
rect 39240 350 39260 410
rect 39160 310 39260 350
rect 39160 250 39180 310
rect 39240 250 39260 310
rect 39160 230 39260 250
rect 39330 410 39430 430
rect 39330 350 39350 410
rect 39410 350 39430 410
rect 39330 310 39430 350
rect 39330 250 39350 310
rect 39410 250 39430 310
rect 39330 230 39430 250
rect 39500 410 39600 430
rect 39500 350 39520 410
rect 39580 350 39600 410
rect 39500 310 39600 350
rect 39500 250 39520 310
rect 39580 250 39600 310
rect 39500 230 39600 250
rect 39670 410 39770 430
rect 39670 350 39690 410
rect 39750 350 39770 410
rect 39670 310 39770 350
rect 39670 250 39690 310
rect 39750 250 39770 310
rect 39670 230 39770 250
rect 39840 410 39940 430
rect 39840 350 39860 410
rect 39920 350 39940 410
rect 39840 310 39940 350
rect 39840 250 39860 310
rect 39920 250 39940 310
rect 39840 230 39940 250
rect 40010 410 40110 430
rect 40010 350 40030 410
rect 40090 350 40110 410
rect 40010 310 40110 350
rect 40010 250 40030 310
rect 40090 250 40110 310
rect 40010 230 40110 250
rect 40180 410 40280 430
rect 40180 350 40200 410
rect 40260 350 40280 410
rect 40180 310 40280 350
rect 40180 250 40200 310
rect 40260 250 40280 310
rect 40180 230 40280 250
rect 40350 410 40450 430
rect 40350 350 40370 410
rect 40430 350 40450 410
rect 40350 310 40450 350
rect 40350 250 40370 310
rect 40430 250 40450 310
rect 40350 230 40450 250
rect 40520 410 40620 430
rect 40520 350 40540 410
rect 40600 350 40620 410
rect 40520 310 40620 350
rect 40520 250 40540 310
rect 40600 250 40620 310
rect 40520 230 40620 250
rect 40690 410 40790 430
rect 40690 350 40710 410
rect 40770 350 40790 410
rect 40690 310 40790 350
rect 40690 250 40710 310
rect 40770 250 40790 310
rect 40690 230 40790 250
rect 40860 410 40960 430
rect 40860 350 40880 410
rect 40940 350 40960 410
rect 40860 310 40960 350
rect 40860 250 40880 310
rect 40940 250 40960 310
rect 40860 230 40960 250
rect 41030 410 41130 430
rect 41030 350 41050 410
rect 41110 350 41130 410
rect 41030 310 41130 350
rect 41030 250 41050 310
rect 41110 250 41130 310
rect 41030 230 41130 250
rect 41200 410 41300 430
rect 41200 350 41220 410
rect 41280 350 41300 410
rect 41200 310 41300 350
rect 41200 250 41220 310
rect 41280 250 41300 310
rect 41200 230 41300 250
rect 41370 410 41470 430
rect 41370 350 41390 410
rect 41450 350 41470 410
rect 41370 310 41470 350
rect 41370 250 41390 310
rect 41450 250 41470 310
rect 41370 230 41470 250
rect 41540 410 41640 430
rect 41540 350 41560 410
rect 41620 350 41640 410
rect 41540 310 41640 350
rect 41540 250 41560 310
rect 41620 250 41640 310
rect 41540 230 41640 250
rect 41710 410 41810 430
rect 41710 350 41730 410
rect 41790 350 41810 410
rect 41710 310 41810 350
rect 41710 250 41730 310
rect 41790 250 41810 310
rect 41710 230 41810 250
rect 41880 410 41980 430
rect 41880 350 41900 410
rect 41960 350 41980 410
rect 41880 310 41980 350
rect 41880 250 41900 310
rect 41960 250 41980 310
rect 41880 230 41980 250
rect 42050 410 42150 430
rect 42050 350 42070 410
rect 42130 350 42150 410
rect 42050 310 42150 350
rect 42050 250 42070 310
rect 42130 250 42150 310
rect 42050 230 42150 250
rect 42220 410 42320 430
rect 42220 350 42240 410
rect 42300 350 42320 410
rect 42220 310 42320 350
rect 42220 250 42240 310
rect 42300 250 42320 310
rect 42220 230 42320 250
rect 42390 410 42490 430
rect 42390 350 42410 410
rect 42470 350 42490 410
rect 42390 310 42490 350
rect 42390 250 42410 310
rect 42470 250 42490 310
rect 42390 230 42490 250
rect 42560 410 42660 430
rect 42560 350 42580 410
rect 42640 350 42660 410
rect 42560 310 42660 350
rect 42560 250 42580 310
rect 42640 250 42660 310
rect 42560 230 42660 250
rect 42730 410 42830 430
rect 42730 350 42750 410
rect 42810 350 42830 410
rect 42730 310 42830 350
rect 42730 250 42750 310
rect 42810 250 42830 310
rect 42730 230 42830 250
rect 42900 410 43000 430
rect 42900 350 42920 410
rect 42980 350 43000 410
rect 42900 310 43000 350
rect 42900 250 42920 310
rect 42980 250 43000 310
rect 42900 230 43000 250
rect 43070 410 43170 430
rect 43070 350 43090 410
rect 43150 350 43170 410
rect 43070 310 43170 350
rect 43070 250 43090 310
rect 43150 250 43170 310
rect 43070 230 43170 250
rect 43240 410 43340 430
rect 43240 350 43260 410
rect 43320 350 43340 410
rect 43240 310 43340 350
rect 43240 250 43260 310
rect 43320 250 43340 310
rect 43240 230 43340 250
rect 43410 410 43510 430
rect 43410 350 43430 410
rect 43490 350 43510 410
rect 43410 310 43510 350
rect 43410 250 43430 310
rect 43490 250 43510 310
rect 43410 230 43510 250
rect 43580 410 43680 430
rect 43580 350 43600 410
rect 43660 350 43680 410
rect 43580 310 43680 350
rect 43580 250 43600 310
rect 43660 250 43680 310
rect 43580 230 43680 250
rect 43750 410 43850 430
rect 43750 350 43770 410
rect 43830 350 43850 410
rect 43750 310 43850 350
rect 43750 250 43770 310
rect 43830 250 43850 310
rect 43750 230 43850 250
rect 43920 410 44020 430
rect 43920 350 43940 410
rect 44000 350 44020 410
rect 43920 310 44020 350
rect 43920 250 43940 310
rect 44000 250 44020 310
rect 43920 230 44020 250
rect 44090 410 44190 430
rect 44090 350 44110 410
rect 44170 350 44190 410
rect 44090 310 44190 350
rect 44090 250 44110 310
rect 44170 250 44190 310
rect 44090 230 44190 250
rect 44260 410 44360 430
rect 44260 350 44280 410
rect 44340 350 44360 410
rect 44260 310 44360 350
rect 44260 250 44280 310
rect 44340 250 44360 310
rect 44260 230 44360 250
rect 44430 410 44530 430
rect 44430 350 44450 410
rect 44510 350 44530 410
rect 44430 310 44530 350
rect 44430 250 44450 310
rect 44510 250 44530 310
rect 44430 230 44530 250
rect 44600 410 44700 430
rect 44600 350 44620 410
rect 44680 350 44700 410
rect 44600 310 44700 350
rect 44600 250 44620 310
rect 44680 250 44700 310
rect 44600 230 44700 250
rect 44770 410 44870 430
rect 44770 350 44790 410
rect 44850 350 44870 410
rect 44770 310 44870 350
rect 44770 250 44790 310
rect 44850 250 44870 310
rect 44770 230 44870 250
rect 44940 410 45040 430
rect 44940 350 44960 410
rect 45020 350 45040 410
rect 44940 310 45040 350
rect 44940 250 44960 310
rect 45020 250 45040 310
rect 44940 230 45040 250
rect 45110 410 45210 430
rect 45110 350 45130 410
rect 45190 350 45210 410
rect 45110 310 45210 350
rect 45110 250 45130 310
rect 45190 250 45210 310
rect 45110 230 45210 250
rect 45280 410 45380 430
rect 45280 350 45300 410
rect 45360 350 45380 410
rect 45280 310 45380 350
rect 45280 250 45300 310
rect 45360 250 45380 310
rect 45280 230 45380 250
rect 45450 410 45550 430
rect 45450 350 45470 410
rect 45530 350 45550 410
rect 45450 310 45550 350
rect 45450 250 45470 310
rect 45530 250 45550 310
rect 45450 230 45550 250
rect 45620 410 45720 430
rect 45620 350 45640 410
rect 45700 350 45720 410
rect 45620 310 45720 350
rect 45620 250 45640 310
rect 45700 250 45720 310
rect 45620 230 45720 250
rect 45790 410 45890 430
rect 45790 350 45810 410
rect 45870 350 45890 410
rect 45790 310 45890 350
rect 45790 250 45810 310
rect 45870 250 45890 310
rect 45790 230 45890 250
rect 45960 410 46060 430
rect 45960 350 45980 410
rect 46040 350 46060 410
rect 45960 310 46060 350
rect 45960 250 45980 310
rect 46040 250 46060 310
rect 45960 230 46060 250
rect 46130 410 46230 430
rect 46130 350 46150 410
rect 46210 350 46230 410
rect 46130 310 46230 350
rect 46130 250 46150 310
rect 46210 250 46230 310
rect 46130 230 46230 250
rect 46300 410 46400 430
rect 46300 350 46320 410
rect 46380 350 46400 410
rect 46300 310 46400 350
rect 46300 250 46320 310
rect 46380 250 46400 310
rect 46300 230 46400 250
rect 46470 410 46570 430
rect 46470 350 46490 410
rect 46550 350 46570 410
rect 46470 310 46570 350
rect 46470 250 46490 310
rect 46550 250 46570 310
rect 46470 230 46570 250
rect 46640 410 46740 430
rect 46640 350 46660 410
rect 46720 350 46740 410
rect 46640 310 46740 350
rect 46640 250 46660 310
rect 46720 250 46740 310
rect 46640 230 46740 250
rect 46810 410 46910 430
rect 46810 350 46830 410
rect 46890 350 46910 410
rect 46810 310 46910 350
rect 46810 250 46830 310
rect 46890 250 46910 310
rect 46810 230 46910 250
rect 46980 410 47080 430
rect 46980 350 47000 410
rect 47060 350 47080 410
rect 46980 310 47080 350
rect 46980 250 47000 310
rect 47060 250 47080 310
rect 46980 230 47080 250
rect 47150 410 47250 430
rect 47150 350 47170 410
rect 47230 350 47250 410
rect 47150 310 47250 350
rect 47150 250 47170 310
rect 47230 250 47250 310
rect 47150 230 47250 250
rect 47320 410 47420 430
rect 47320 350 47340 410
rect 47400 350 47420 410
rect 47320 310 47420 350
rect 47320 250 47340 310
rect 47400 250 47420 310
rect 47320 230 47420 250
rect 47490 410 47590 430
rect 47490 350 47510 410
rect 47570 350 47590 410
rect 47490 310 47590 350
rect 47490 250 47510 310
rect 47570 250 47590 310
rect 47490 230 47590 250
rect 47660 410 47760 430
rect 47660 350 47680 410
rect 47740 350 47760 410
rect 47660 310 47760 350
rect 47660 250 47680 310
rect 47740 250 47760 310
rect 47660 230 47760 250
rect 47830 410 47930 430
rect 47830 350 47850 410
rect 47910 350 47930 410
rect 47830 310 47930 350
rect 47830 250 47850 310
rect 47910 250 47930 310
rect 47830 230 47930 250
rect 48000 410 48100 430
rect 48000 350 48020 410
rect 48080 350 48100 410
rect 48000 310 48100 350
rect 48000 250 48020 310
rect 48080 250 48100 310
rect 48000 230 48100 250
rect 48170 410 48270 430
rect 48170 350 48190 410
rect 48250 350 48270 410
rect 48170 310 48270 350
rect 48170 250 48190 310
rect 48250 250 48270 310
rect 48170 230 48270 250
rect 48340 410 48440 430
rect 48340 350 48360 410
rect 48420 350 48440 410
rect 48340 310 48440 350
rect 48340 250 48360 310
rect 48420 250 48440 310
rect 48340 230 48440 250
rect 48510 410 48610 430
rect 48510 350 48530 410
rect 48590 350 48610 410
rect 48510 310 48610 350
rect 48510 250 48530 310
rect 48590 250 48610 310
rect 48510 230 48610 250
rect 48680 410 48780 430
rect 48680 350 48700 410
rect 48760 350 48780 410
rect 48680 310 48780 350
rect 48680 250 48700 310
rect 48760 250 48780 310
rect 48680 230 48780 250
rect 48850 410 48950 430
rect 48850 350 48870 410
rect 48930 350 48950 410
rect 48850 310 48950 350
rect 48850 250 48870 310
rect 48930 250 48950 310
rect 48850 230 48950 250
rect 49020 410 49120 430
rect 49020 350 49040 410
rect 49100 350 49120 410
rect 49020 310 49120 350
rect 49020 250 49040 310
rect 49100 250 49120 310
rect 49020 230 49120 250
rect 49190 410 49290 430
rect 49190 350 49210 410
rect 49270 350 49290 410
rect 49190 310 49290 350
rect 49190 250 49210 310
rect 49270 250 49290 310
rect 49190 230 49290 250
rect 49360 410 49460 430
rect 49360 350 49380 410
rect 49440 350 49460 410
rect 49360 310 49460 350
rect 49360 250 49380 310
rect 49440 250 49460 310
rect 49360 230 49460 250
rect 49530 410 49630 430
rect 49530 350 49550 410
rect 49610 350 49630 410
rect 49530 310 49630 350
rect 49530 250 49550 310
rect 49610 250 49630 310
rect 49530 230 49630 250
rect 49700 410 49800 430
rect 49700 350 49720 410
rect 49780 350 49800 410
rect 49700 310 49800 350
rect 49700 250 49720 310
rect 49780 250 49800 310
rect 49700 230 49800 250
rect 49870 410 49970 430
rect 49870 350 49890 410
rect 49950 350 49970 410
rect 49870 310 49970 350
rect 49870 250 49890 310
rect 49950 250 49970 310
rect 49870 230 49970 250
rect 50040 410 50140 430
rect 50040 350 50060 410
rect 50120 350 50140 410
rect 50040 310 50140 350
rect 50040 250 50060 310
rect 50120 250 50140 310
rect 50040 230 50140 250
rect 50210 410 50310 430
rect 50210 350 50230 410
rect 50290 350 50310 410
rect 50210 310 50310 350
rect 50210 250 50230 310
rect 50290 250 50310 310
rect 50210 230 50310 250
rect 50380 410 50480 430
rect 50380 350 50400 410
rect 50460 350 50480 410
rect 50380 310 50480 350
rect 50380 250 50400 310
rect 50460 250 50480 310
rect 50380 230 50480 250
rect 50550 410 50650 430
rect 50550 350 50570 410
rect 50630 350 50650 410
rect 50550 310 50650 350
rect 50550 250 50570 310
rect 50630 250 50650 310
rect 50550 230 50650 250
rect 50720 410 50820 430
rect 50720 350 50740 410
rect 50800 350 50820 410
rect 50720 310 50820 350
rect 50720 250 50740 310
rect 50800 250 50820 310
rect 50720 230 50820 250
rect 50890 410 50990 430
rect 50890 350 50910 410
rect 50970 350 50990 410
rect 50890 310 50990 350
rect 50890 250 50910 310
rect 50970 250 50990 310
rect 50890 230 50990 250
rect 51060 410 51160 430
rect 51060 350 51080 410
rect 51140 350 51160 410
rect 51060 310 51160 350
rect 51060 250 51080 310
rect 51140 250 51160 310
rect 51060 230 51160 250
rect 51230 410 51330 430
rect 51230 350 51250 410
rect 51310 350 51330 410
rect 51230 310 51330 350
rect 51230 250 51250 310
rect 51310 250 51330 310
rect 51230 230 51330 250
rect 51400 410 51500 430
rect 51400 350 51420 410
rect 51480 350 51500 410
rect 51400 310 51500 350
rect 51400 250 51420 310
rect 51480 250 51500 310
rect 51400 230 51500 250
rect 51570 410 51670 430
rect 51570 350 51590 410
rect 51650 350 51670 410
rect 51570 310 51670 350
rect 51570 250 51590 310
rect 51650 250 51670 310
rect 51570 230 51670 250
rect 51740 410 51840 430
rect 51740 350 51760 410
rect 51820 350 51840 410
rect 51740 310 51840 350
rect 51740 250 51760 310
rect 51820 250 51840 310
rect 51740 230 51840 250
rect 51910 410 52010 430
rect 51910 350 51930 410
rect 51990 350 52010 410
rect 51910 310 52010 350
rect 51910 250 51930 310
rect 51990 250 52010 310
rect 51910 230 52010 250
rect 52080 410 52180 430
rect 52080 350 52100 410
rect 52160 350 52180 410
rect 52080 310 52180 350
rect 52080 250 52100 310
rect 52160 250 52180 310
rect 52080 230 52180 250
rect 52250 410 52350 430
rect 52250 350 52270 410
rect 52330 350 52350 410
rect 52250 310 52350 350
rect 52250 250 52270 310
rect 52330 250 52350 310
rect 52250 230 52350 250
rect 52420 410 52520 430
rect 52420 350 52440 410
rect 52500 350 52520 410
rect 52420 310 52520 350
rect 52420 250 52440 310
rect 52500 250 52520 310
rect 52420 230 52520 250
rect 52590 410 52690 430
rect 52590 350 52610 410
rect 52670 350 52690 410
rect 52590 310 52690 350
rect 52590 250 52610 310
rect 52670 250 52690 310
rect 52590 230 52690 250
rect 52760 410 52860 430
rect 52760 350 52780 410
rect 52840 350 52860 410
rect 52760 310 52860 350
rect 52760 250 52780 310
rect 52840 250 52860 310
rect 52760 230 52860 250
rect 52930 410 53030 430
rect 52930 350 52950 410
rect 53010 350 53030 410
rect 52930 310 53030 350
rect 52930 250 52950 310
rect 53010 250 53030 310
rect 52930 230 53030 250
rect 53100 410 53200 430
rect 53100 350 53120 410
rect 53180 350 53200 410
rect 53100 310 53200 350
rect 53100 250 53120 310
rect 53180 250 53200 310
rect 53100 230 53200 250
rect 53270 410 53370 430
rect 53270 350 53290 410
rect 53350 350 53370 410
rect 53270 310 53370 350
rect 53270 250 53290 310
rect 53350 250 53370 310
rect 53270 230 53370 250
rect 53440 410 53540 430
rect 53440 350 53460 410
rect 53520 350 53540 410
rect 53440 310 53540 350
rect 53440 250 53460 310
rect 53520 250 53540 310
rect 53440 230 53540 250
rect 53610 410 53710 430
rect 53610 350 53630 410
rect 53690 350 53710 410
rect 53610 310 53710 350
rect 53610 250 53630 310
rect 53690 250 53710 310
rect 53610 230 53710 250
rect 53780 410 53880 430
rect 53780 350 53800 410
rect 53860 350 53880 410
rect 53780 310 53880 350
rect 53780 250 53800 310
rect 53860 250 53880 310
rect 53780 230 53880 250
rect 53950 410 54050 430
rect 53950 350 53970 410
rect 54030 350 54050 410
rect 53950 310 54050 350
rect 53950 250 53970 310
rect 54030 250 54050 310
rect 53950 230 54050 250
rect 54120 410 54220 430
rect 54120 350 54140 410
rect 54200 350 54220 410
rect 54120 310 54220 350
rect 54120 250 54140 310
rect 54200 250 54220 310
rect 54120 230 54220 250
rect 54290 410 54390 430
rect 54290 350 54310 410
rect 54370 350 54390 410
rect 54290 310 54390 350
rect 54290 250 54310 310
rect 54370 250 54390 310
rect 54290 230 54390 250
rect 54460 410 54560 430
rect 54460 350 54480 410
rect 54540 350 54560 410
rect 54460 310 54560 350
rect 54460 250 54480 310
rect 54540 250 54560 310
rect 54460 230 54560 250
rect 54630 410 54730 430
rect 54630 350 54650 410
rect 54710 350 54730 410
rect 54630 310 54730 350
rect 54630 250 54650 310
rect 54710 250 54730 310
rect 54630 230 54730 250
rect 54800 410 54900 430
rect 54800 350 54820 410
rect 54880 350 54900 410
rect 54800 310 54900 350
rect 54800 250 54820 310
rect 54880 250 54900 310
rect 54800 230 54900 250
rect 54970 410 55070 430
rect 54970 350 54990 410
rect 55050 350 55070 410
rect 54970 310 55070 350
rect 54970 250 54990 310
rect 55050 250 55070 310
rect 54970 230 55070 250
rect 55140 410 55240 430
rect 55140 350 55160 410
rect 55220 350 55240 410
rect 55140 310 55240 350
rect 55140 250 55160 310
rect 55220 250 55240 310
rect 55140 230 55240 250
rect 55310 410 55410 430
rect 55310 350 55330 410
rect 55390 350 55410 410
rect 55310 310 55410 350
rect 55310 250 55330 310
rect 55390 250 55410 310
rect 55310 230 55410 250
rect 55480 410 55580 430
rect 55480 350 55500 410
rect 55560 350 55580 410
rect 55480 310 55580 350
rect 55480 250 55500 310
rect 55560 250 55580 310
rect 55480 230 55580 250
rect 55650 410 55750 430
rect 55650 350 55670 410
rect 55730 350 55750 410
rect 55650 310 55750 350
rect 55650 250 55670 310
rect 55730 250 55750 310
rect 55650 230 55750 250
rect 55820 410 55920 430
rect 55820 350 55840 410
rect 55900 350 55920 410
rect 55820 310 55920 350
rect 55820 250 55840 310
rect 55900 250 55920 310
rect 55820 230 55920 250
rect 55990 410 56090 430
rect 55990 350 56010 410
rect 56070 350 56090 410
rect 55990 310 56090 350
rect 55990 250 56010 310
rect 56070 250 56090 310
rect 55990 230 56090 250
rect 56160 410 56260 430
rect 56160 350 56180 410
rect 56240 350 56260 410
rect 56160 310 56260 350
rect 56160 250 56180 310
rect 56240 250 56260 310
rect 56160 230 56260 250
rect 56330 410 56430 430
rect 56330 350 56350 410
rect 56410 350 56430 410
rect 56330 310 56430 350
rect 56330 250 56350 310
rect 56410 250 56430 310
rect 56330 230 56430 250
rect 56500 410 56600 430
rect 56500 350 56520 410
rect 56580 350 56600 410
rect 56500 310 56600 350
rect 56500 250 56520 310
rect 56580 250 56600 310
rect 56500 230 56600 250
rect 56670 410 56770 430
rect 56670 350 56690 410
rect 56750 350 56770 410
rect 56670 310 56770 350
rect 56670 250 56690 310
rect 56750 250 56770 310
rect 56670 230 56770 250
rect 56840 410 56940 430
rect 56840 350 56860 410
rect 56920 350 56940 410
rect 56840 310 56940 350
rect 56840 250 56860 310
rect 56920 250 56940 310
rect 56840 230 56940 250
rect 57010 410 57110 430
rect 57010 350 57030 410
rect 57090 350 57110 410
rect 57010 310 57110 350
rect 57010 250 57030 310
rect 57090 250 57110 310
rect 57010 230 57110 250
rect 57180 410 57280 430
rect 57180 350 57200 410
rect 57260 350 57280 410
rect 57180 310 57280 350
rect 57180 250 57200 310
rect 57260 250 57280 310
rect 57180 230 57280 250
rect 57350 410 57450 430
rect 57350 350 57370 410
rect 57430 350 57450 410
rect 57350 310 57450 350
rect 57350 250 57370 310
rect 57430 250 57450 310
rect 57350 230 57450 250
rect 57520 410 57620 430
rect 57520 350 57540 410
rect 57600 350 57620 410
rect 57520 310 57620 350
rect 57520 250 57540 310
rect 57600 250 57620 310
rect 57520 230 57620 250
rect 57690 410 57790 430
rect 57690 350 57710 410
rect 57770 350 57790 410
rect 57690 310 57790 350
rect 57690 250 57710 310
rect 57770 250 57790 310
rect 57690 230 57790 250
rect 57860 410 57960 430
rect 57860 350 57880 410
rect 57940 350 57960 410
rect 57860 310 57960 350
rect 57860 250 57880 310
rect 57940 250 57960 310
rect 57860 230 57960 250
rect 58030 410 58130 430
rect 58030 350 58050 410
rect 58110 350 58130 410
rect 58030 310 58130 350
rect 58030 250 58050 310
rect 58110 250 58130 310
rect 58030 230 58130 250
rect 58200 410 58300 430
rect 58200 350 58220 410
rect 58280 350 58300 410
rect 58200 310 58300 350
rect 58200 250 58220 310
rect 58280 250 58300 310
rect 58200 230 58300 250
rect 58370 410 58470 430
rect 58370 350 58390 410
rect 58450 350 58470 410
rect 58370 310 58470 350
rect 58370 250 58390 310
rect 58450 250 58470 310
rect 58370 230 58470 250
rect 58540 410 58640 430
rect 58540 350 58560 410
rect 58620 350 58640 410
rect 58540 310 58640 350
rect 58540 250 58560 310
rect 58620 250 58640 310
rect 58540 230 58640 250
rect 58710 410 58810 430
rect 58710 350 58730 410
rect 58790 350 58810 410
rect 58710 310 58810 350
rect 58710 250 58730 310
rect 58790 250 58810 310
rect 58710 230 58810 250
rect 58880 410 58980 430
rect 58880 350 58900 410
rect 58960 350 58980 410
rect 58880 310 58980 350
rect 58880 250 58900 310
rect 58960 250 58980 310
rect 58880 230 58980 250
rect 59050 410 59150 430
rect 59050 350 59070 410
rect 59130 350 59150 410
rect 59050 310 59150 350
rect 59050 250 59070 310
rect 59130 250 59150 310
rect 59050 230 59150 250
rect 59220 410 59320 430
rect 59220 350 59240 410
rect 59300 350 59320 410
rect 59220 310 59320 350
rect 59220 250 59240 310
rect 59300 250 59320 310
rect 59220 230 59320 250
rect 50 110 150 130
rect 50 30 70 110
rect 130 30 150 110
rect 50 10 150 30
rect 430 80 530 100
rect 430 20 450 80
rect 510 20 530 80
rect 430 0 530 20
rect 600 80 700 100
rect 600 20 620 80
rect 680 20 700 80
rect 600 0 700 20
rect 770 80 870 100
rect 770 20 790 80
rect 850 20 870 80
rect 770 0 870 20
rect 940 80 1040 100
rect 940 20 960 80
rect 1020 20 1040 80
rect 940 0 1040 20
rect 1110 80 1210 100
rect 1110 20 1130 80
rect 1190 20 1210 80
rect 1110 0 1210 20
rect 1500 80 1600 100
rect 1500 20 1520 80
rect 1580 20 1600 80
rect 1500 0 1600 20
rect 1670 80 1770 100
rect 1670 20 1690 80
rect 1750 20 1770 80
rect 1670 0 1770 20
rect 1840 80 1940 100
rect 1840 20 1860 80
rect 1920 20 1940 80
rect 1840 0 1940 20
rect 2010 80 2110 100
rect 2010 20 2030 80
rect 2090 20 2110 80
rect 2010 0 2110 20
rect 2180 80 2280 100
rect 2180 20 2200 80
rect 2260 20 2280 80
rect 2180 0 2280 20
rect 2350 80 2450 100
rect 2350 20 2370 80
rect 2430 20 2450 80
rect 2350 0 2450 20
rect 2520 80 2620 100
rect 2520 20 2540 80
rect 2600 20 2620 80
rect 2520 0 2620 20
rect 2690 80 2790 100
rect 2690 20 2710 80
rect 2770 20 2790 80
rect 2690 0 2790 20
rect 2860 80 2960 100
rect 2860 20 2880 80
rect 2940 20 2960 80
rect 2860 0 2960 20
rect 3030 80 3130 100
rect 3030 20 3050 80
rect 3110 20 3130 80
rect 3030 0 3130 20
rect 3200 80 3300 100
rect 3200 20 3220 80
rect 3280 20 3300 80
rect 3200 0 3300 20
rect 3370 80 3470 100
rect 3370 20 3390 80
rect 3450 20 3470 80
rect 3370 0 3470 20
rect 3540 80 3640 100
rect 3540 20 3560 80
rect 3620 20 3640 80
rect 3540 0 3640 20
rect 3710 80 3810 100
rect 3710 20 3730 80
rect 3790 20 3810 80
rect 3710 0 3810 20
rect 3880 80 3980 100
rect 3880 20 3900 80
rect 3960 20 3980 80
rect 3880 0 3980 20
rect 4050 80 4150 100
rect 4050 20 4070 80
rect 4130 20 4150 80
rect 4050 0 4150 20
rect 4220 80 4320 100
rect 4220 20 4240 80
rect 4300 20 4320 80
rect 4220 0 4320 20
rect 4520 80 4620 100
rect 4520 20 4540 80
rect 4600 20 4620 80
rect 4520 0 4620 20
rect 4690 80 4790 100
rect 4690 20 4710 80
rect 4770 20 4790 80
rect 4690 0 4790 20
rect 4860 80 4960 100
rect 4860 20 4880 80
rect 4940 20 4960 80
rect 4860 0 4960 20
rect 5030 80 5130 100
rect 5030 20 5050 80
rect 5110 20 5130 80
rect 5030 0 5130 20
rect 5200 80 5300 100
rect 5200 20 5220 80
rect 5280 20 5300 80
rect 5200 0 5300 20
rect 5370 80 5470 100
rect 5370 20 5390 80
rect 5450 20 5470 80
rect 5370 0 5470 20
rect 5540 80 5640 100
rect 5540 20 5560 80
rect 5620 20 5640 80
rect 5540 0 5640 20
rect 5710 80 5810 100
rect 5710 20 5730 80
rect 5790 20 5810 80
rect 5710 0 5810 20
rect 5880 80 5980 100
rect 5880 20 5900 80
rect 5960 20 5980 80
rect 5880 0 5980 20
rect 6050 80 6150 100
rect 6050 20 6070 80
rect 6130 20 6150 80
rect 6050 0 6150 20
rect 6220 80 6320 100
rect 6220 20 6240 80
rect 6300 20 6320 80
rect 6220 0 6320 20
rect 6390 80 6490 100
rect 6390 20 6410 80
rect 6470 20 6490 80
rect 6390 0 6490 20
rect 6560 80 6660 100
rect 6560 20 6580 80
rect 6640 20 6660 80
rect 6560 0 6660 20
rect 6730 80 6830 100
rect 6730 20 6750 80
rect 6810 20 6830 80
rect 6730 0 6830 20
rect 6900 80 7000 100
rect 6900 20 6920 80
rect 6980 20 7000 80
rect 6900 0 7000 20
rect 7070 80 7170 100
rect 7070 20 7090 80
rect 7150 20 7170 80
rect 7070 0 7170 20
rect 7240 80 7340 100
rect 7240 20 7260 80
rect 7320 20 7340 80
rect 7240 0 7340 20
rect 7410 80 7510 100
rect 7410 20 7430 80
rect 7490 20 7510 80
rect 7410 0 7510 20
rect 7580 80 7680 100
rect 7580 20 7600 80
rect 7660 20 7680 80
rect 7580 0 7680 20
rect 7750 80 7850 100
rect 7750 20 7770 80
rect 7830 20 7850 80
rect 7750 0 7850 20
rect 7920 80 8020 100
rect 7920 20 7940 80
rect 8000 20 8020 80
rect 7920 0 8020 20
rect 8090 80 8190 100
rect 8090 20 8110 80
rect 8170 20 8190 80
rect 8090 0 8190 20
rect 8260 80 8360 100
rect 8260 20 8280 80
rect 8340 20 8360 80
rect 8260 0 8360 20
rect 8430 80 8530 100
rect 8430 20 8450 80
rect 8510 20 8530 80
rect 8430 0 8530 20
rect 8600 80 8700 100
rect 8600 20 8620 80
rect 8680 20 8700 80
rect 8600 0 8700 20
rect 8770 80 8870 100
rect 8770 20 8790 80
rect 8850 20 8870 80
rect 8770 0 8870 20
rect 8940 80 9040 100
rect 8940 20 8960 80
rect 9020 20 9040 80
rect 8940 0 9040 20
rect 9110 80 9210 100
rect 9110 20 9130 80
rect 9190 20 9210 80
rect 9110 0 9210 20
rect 9280 80 9380 100
rect 9280 20 9300 80
rect 9360 20 9380 80
rect 9280 0 9380 20
rect 9450 80 9550 100
rect 9450 20 9470 80
rect 9530 20 9550 80
rect 9450 0 9550 20
rect 9620 80 9720 100
rect 9620 20 9640 80
rect 9700 20 9720 80
rect 9620 0 9720 20
rect 9790 80 9890 100
rect 9790 20 9810 80
rect 9870 20 9890 80
rect 9790 0 9890 20
rect 9960 80 10060 100
rect 9960 20 9980 80
rect 10040 20 10060 80
rect 9960 0 10060 20
rect 10130 80 10230 100
rect 10130 20 10150 80
rect 10210 20 10230 80
rect 10130 0 10230 20
rect 10300 80 10400 100
rect 10300 20 10320 80
rect 10380 20 10400 80
rect 10300 0 10400 20
rect 10470 80 10570 100
rect 10470 20 10490 80
rect 10550 20 10570 80
rect 10470 0 10570 20
rect 10640 80 10740 100
rect 10640 20 10660 80
rect 10720 20 10740 80
rect 10640 0 10740 20
rect 10810 80 10910 100
rect 10810 20 10830 80
rect 10890 20 10910 80
rect 10810 0 10910 20
rect 10980 80 11080 100
rect 10980 20 11000 80
rect 11060 20 11080 80
rect 10980 0 11080 20
rect 11150 80 11250 100
rect 11150 20 11170 80
rect 11230 20 11250 80
rect 11150 0 11250 20
rect 11320 80 11420 100
rect 11320 20 11340 80
rect 11400 20 11420 80
rect 11320 0 11420 20
rect 11490 80 11590 100
rect 11490 20 11510 80
rect 11570 20 11590 80
rect 11490 0 11590 20
rect 11660 80 11760 100
rect 11660 20 11680 80
rect 11740 20 11760 80
rect 11660 0 11760 20
rect 11830 80 11930 100
rect 11830 20 11850 80
rect 11910 20 11930 80
rect 11830 0 11930 20
rect 12000 80 12100 100
rect 12000 20 12020 80
rect 12080 20 12100 80
rect 12000 0 12100 20
rect 12170 80 12270 100
rect 12170 20 12190 80
rect 12250 20 12270 80
rect 12170 0 12270 20
rect 12340 80 12440 100
rect 12340 20 12360 80
rect 12420 20 12440 80
rect 12340 0 12440 20
rect 12510 80 12610 100
rect 12510 20 12530 80
rect 12590 20 12610 80
rect 12510 0 12610 20
rect 12680 80 12780 100
rect 12680 20 12700 80
rect 12760 20 12780 80
rect 12680 0 12780 20
rect 12850 80 12950 100
rect 12850 20 12870 80
rect 12930 20 12950 80
rect 12850 0 12950 20
rect 13020 80 13120 100
rect 13020 20 13040 80
rect 13100 20 13120 80
rect 13020 0 13120 20
rect 13190 80 13290 100
rect 13190 20 13210 80
rect 13270 20 13290 80
rect 13190 0 13290 20
rect 13360 80 13460 100
rect 13360 20 13380 80
rect 13440 20 13460 80
rect 13360 0 13460 20
rect 13530 80 13630 100
rect 13530 20 13550 80
rect 13610 20 13630 80
rect 13530 0 13630 20
rect 13700 80 13800 100
rect 13700 20 13720 80
rect 13780 20 13800 80
rect 13700 0 13800 20
rect 13870 80 13970 100
rect 13870 20 13890 80
rect 13950 20 13970 80
rect 13870 0 13970 20
rect 14040 80 14140 100
rect 14040 20 14060 80
rect 14120 20 14140 80
rect 14040 0 14140 20
rect 14210 80 14310 100
rect 14210 20 14230 80
rect 14290 20 14310 80
rect 14210 0 14310 20
rect 14380 80 14480 100
rect 14380 20 14400 80
rect 14460 20 14480 80
rect 14380 0 14480 20
rect 14550 80 14650 100
rect 14550 20 14570 80
rect 14630 20 14650 80
rect 14550 0 14650 20
rect 14720 80 14820 100
rect 14720 20 14740 80
rect 14800 20 14820 80
rect 14720 0 14820 20
rect 14890 80 14990 100
rect 14890 20 14910 80
rect 14970 20 14990 80
rect 14890 0 14990 20
rect 15060 80 15160 100
rect 15060 20 15080 80
rect 15140 20 15160 80
rect 15060 0 15160 20
rect 15230 80 15330 100
rect 15230 20 15250 80
rect 15310 20 15330 80
rect 15230 0 15330 20
rect 15400 80 15500 100
rect 15400 20 15420 80
rect 15480 20 15500 80
rect 15400 0 15500 20
rect 15700 80 15800 100
rect 15700 20 15720 80
rect 15780 20 15800 80
rect 15700 0 15800 20
rect 15870 80 15970 100
rect 15870 20 15890 80
rect 15950 20 15970 80
rect 15870 0 15970 20
rect 16040 80 16140 100
rect 16040 20 16060 80
rect 16120 20 16140 80
rect 16040 0 16140 20
rect 16210 80 16310 100
rect 16210 20 16230 80
rect 16290 20 16310 80
rect 16210 0 16310 20
rect 16380 80 16480 100
rect 16380 20 16400 80
rect 16460 20 16480 80
rect 16380 0 16480 20
rect 16550 80 16650 100
rect 16550 20 16570 80
rect 16630 20 16650 80
rect 16550 0 16650 20
rect 16720 80 16820 100
rect 16720 20 16740 80
rect 16800 20 16820 80
rect 16720 0 16820 20
rect 16890 80 16990 100
rect 16890 20 16910 80
rect 16970 20 16990 80
rect 16890 0 16990 20
rect 17060 80 17160 100
rect 17060 20 17080 80
rect 17140 20 17160 80
rect 17060 0 17160 20
rect 17230 80 17330 100
rect 17230 20 17250 80
rect 17310 20 17330 80
rect 17230 0 17330 20
rect 17400 80 17500 100
rect 17400 20 17420 80
rect 17480 20 17500 80
rect 17400 0 17500 20
rect 17570 80 17670 100
rect 17570 20 17590 80
rect 17650 20 17670 80
rect 17570 0 17670 20
rect 17740 80 17840 100
rect 17740 20 17760 80
rect 17820 20 17840 80
rect 17740 0 17840 20
rect 17910 80 18010 100
rect 17910 20 17930 80
rect 17990 20 18010 80
rect 17910 0 18010 20
rect 18080 80 18180 100
rect 18080 20 18100 80
rect 18160 20 18180 80
rect 18080 0 18180 20
rect 18250 80 18350 100
rect 18250 20 18270 80
rect 18330 20 18350 80
rect 18250 0 18350 20
rect 18420 80 18520 100
rect 18420 20 18440 80
rect 18500 20 18520 80
rect 18420 0 18520 20
rect 18590 80 18690 100
rect 18590 20 18610 80
rect 18670 20 18690 80
rect 18590 0 18690 20
rect 18760 80 18860 100
rect 18760 20 18780 80
rect 18840 20 18860 80
rect 18760 0 18860 20
rect 18930 80 19030 100
rect 18930 20 18950 80
rect 19010 20 19030 80
rect 18930 0 19030 20
rect 19100 80 19200 100
rect 19100 20 19120 80
rect 19180 20 19200 80
rect 19100 0 19200 20
rect 19270 80 19370 100
rect 19270 20 19290 80
rect 19350 20 19370 80
rect 19270 0 19370 20
rect 19440 80 19540 100
rect 19440 20 19460 80
rect 19520 20 19540 80
rect 19440 0 19540 20
rect 19610 80 19710 100
rect 19610 20 19630 80
rect 19690 20 19710 80
rect 19610 0 19710 20
rect 19780 80 19880 100
rect 19780 20 19800 80
rect 19860 20 19880 80
rect 19780 0 19880 20
rect 19950 80 20050 100
rect 19950 20 19970 80
rect 20030 20 20050 80
rect 19950 0 20050 20
rect 20120 80 20220 100
rect 20120 20 20140 80
rect 20200 20 20220 80
rect 20120 0 20220 20
rect 20290 80 20390 100
rect 20290 20 20310 80
rect 20370 20 20390 80
rect 20290 0 20390 20
rect 20460 80 20560 100
rect 20460 20 20480 80
rect 20540 20 20560 80
rect 20460 0 20560 20
rect 20630 80 20730 100
rect 20630 20 20650 80
rect 20710 20 20730 80
rect 20630 0 20730 20
rect 20800 80 20900 100
rect 20800 20 20820 80
rect 20880 20 20900 80
rect 20800 0 20900 20
rect 20970 80 21070 100
rect 20970 20 20990 80
rect 21050 20 21070 80
rect 20970 0 21070 20
rect 21140 80 21240 100
rect 21140 20 21160 80
rect 21220 20 21240 80
rect 21140 0 21240 20
rect 21310 80 21410 100
rect 21310 20 21330 80
rect 21390 20 21410 80
rect 21310 0 21410 20
rect 21480 80 21580 100
rect 21480 20 21500 80
rect 21560 20 21580 80
rect 21480 0 21580 20
rect 21650 80 21750 100
rect 21650 20 21670 80
rect 21730 20 21750 80
rect 21650 0 21750 20
rect 21820 80 21920 100
rect 21820 20 21840 80
rect 21900 20 21920 80
rect 21820 0 21920 20
rect 21990 80 22090 100
rect 21990 20 22010 80
rect 22070 20 22090 80
rect 21990 0 22090 20
rect 22160 80 22260 100
rect 22160 20 22180 80
rect 22240 20 22260 80
rect 22160 0 22260 20
rect 22330 80 22430 100
rect 22330 20 22350 80
rect 22410 20 22430 80
rect 22330 0 22430 20
rect 22500 80 22600 100
rect 22500 20 22520 80
rect 22580 20 22600 80
rect 22500 0 22600 20
rect 22670 80 22770 100
rect 22670 20 22690 80
rect 22750 20 22770 80
rect 22670 0 22770 20
rect 22840 80 22940 100
rect 22840 20 22860 80
rect 22920 20 22940 80
rect 22840 0 22940 20
rect 23010 80 23110 100
rect 23010 20 23030 80
rect 23090 20 23110 80
rect 23010 0 23110 20
rect 23180 80 23280 100
rect 23180 20 23200 80
rect 23260 20 23280 80
rect 23180 0 23280 20
rect 23350 80 23450 100
rect 23350 20 23370 80
rect 23430 20 23450 80
rect 23350 0 23450 20
rect 23520 80 23620 100
rect 23520 20 23540 80
rect 23600 20 23620 80
rect 23520 0 23620 20
rect 23690 80 23790 100
rect 23690 20 23710 80
rect 23770 20 23790 80
rect 23690 0 23790 20
rect 23860 80 23960 100
rect 23860 20 23880 80
rect 23940 20 23960 80
rect 23860 0 23960 20
rect 24030 80 24130 100
rect 24030 20 24050 80
rect 24110 20 24130 80
rect 24030 0 24130 20
rect 24200 80 24300 100
rect 24200 20 24220 80
rect 24280 20 24300 80
rect 24200 0 24300 20
rect 24370 80 24470 100
rect 24370 20 24390 80
rect 24450 20 24470 80
rect 24370 0 24470 20
rect 24540 80 24640 100
rect 24540 20 24560 80
rect 24620 20 24640 80
rect 24540 0 24640 20
rect 24710 80 24810 100
rect 24710 20 24730 80
rect 24790 20 24810 80
rect 24710 0 24810 20
rect 24880 80 24980 100
rect 24880 20 24900 80
rect 24960 20 24980 80
rect 24880 0 24980 20
rect 25050 80 25150 100
rect 25050 20 25070 80
rect 25130 20 25150 80
rect 25050 0 25150 20
rect 25220 80 25320 100
rect 25220 20 25240 80
rect 25300 20 25320 80
rect 25220 0 25320 20
rect 25390 80 25490 100
rect 25390 20 25410 80
rect 25470 20 25490 80
rect 25390 0 25490 20
rect 25560 80 25660 100
rect 25560 20 25580 80
rect 25640 20 25660 80
rect 25560 0 25660 20
rect 25730 80 25830 100
rect 25730 20 25750 80
rect 25810 20 25830 80
rect 25730 0 25830 20
rect 25900 80 26000 100
rect 25900 20 25920 80
rect 25980 20 26000 80
rect 25900 0 26000 20
rect 26070 80 26170 100
rect 26070 20 26090 80
rect 26150 20 26170 80
rect 26070 0 26170 20
rect 26240 80 26340 100
rect 26240 20 26260 80
rect 26320 20 26340 80
rect 26240 0 26340 20
rect 26410 80 26510 100
rect 26410 20 26430 80
rect 26490 20 26510 80
rect 26410 0 26510 20
rect 26580 80 26680 100
rect 26580 20 26600 80
rect 26660 20 26680 80
rect 26580 0 26680 20
rect 26750 80 26850 100
rect 26750 20 26770 80
rect 26830 20 26850 80
rect 26750 0 26850 20
rect 26920 80 27020 100
rect 26920 20 26940 80
rect 27000 20 27020 80
rect 26920 0 27020 20
rect 27090 80 27190 100
rect 27090 20 27110 80
rect 27170 20 27190 80
rect 27090 0 27190 20
rect 27260 80 27360 100
rect 27260 20 27280 80
rect 27340 20 27360 80
rect 27260 0 27360 20
rect 27430 80 27530 100
rect 27430 20 27450 80
rect 27510 20 27530 80
rect 27430 0 27530 20
rect 27600 80 27700 100
rect 27600 20 27620 80
rect 27680 20 27700 80
rect 27600 0 27700 20
rect 27770 80 27870 100
rect 27770 20 27790 80
rect 27850 20 27870 80
rect 27770 0 27870 20
rect 27940 80 28040 100
rect 27940 20 27960 80
rect 28020 20 28040 80
rect 27940 0 28040 20
rect 28110 80 28210 100
rect 28110 20 28130 80
rect 28190 20 28210 80
rect 28110 0 28210 20
rect 28280 80 28380 100
rect 28280 20 28300 80
rect 28360 20 28380 80
rect 28280 0 28380 20
rect 28450 80 28550 100
rect 28450 20 28470 80
rect 28530 20 28550 80
rect 28450 0 28550 20
rect 28620 80 28720 100
rect 28620 20 28640 80
rect 28700 20 28720 80
rect 28620 0 28720 20
rect 28790 80 28890 100
rect 28790 20 28810 80
rect 28870 20 28890 80
rect 28790 0 28890 20
rect 28960 80 29060 100
rect 28960 20 28980 80
rect 29040 20 29060 80
rect 28960 0 29060 20
rect 29130 80 29230 100
rect 29130 20 29150 80
rect 29210 20 29230 80
rect 29130 0 29230 20
rect 29300 80 29400 100
rect 29300 20 29320 80
rect 29380 20 29400 80
rect 29300 0 29400 20
rect 29470 80 29570 100
rect 29470 20 29490 80
rect 29550 20 29570 80
rect 29470 0 29570 20
rect 29640 80 29740 100
rect 29640 20 29660 80
rect 29720 20 29740 80
rect 29640 0 29740 20
rect 29810 80 29910 100
rect 29810 20 29830 80
rect 29890 20 29910 80
rect 29810 0 29910 20
rect 29980 80 30080 100
rect 29980 20 30000 80
rect 30060 20 30080 80
rect 29980 0 30080 20
rect 30150 80 30250 100
rect 30150 20 30170 80
rect 30230 20 30250 80
rect 30150 0 30250 20
rect 30320 80 30420 100
rect 30320 20 30340 80
rect 30400 20 30420 80
rect 30320 0 30420 20
rect 30490 80 30590 100
rect 30490 20 30510 80
rect 30570 20 30590 80
rect 30490 0 30590 20
rect 30660 80 30760 100
rect 30660 20 30680 80
rect 30740 20 30760 80
rect 30660 0 30760 20
rect 30830 80 30930 100
rect 30830 20 30850 80
rect 30910 20 30930 80
rect 30830 0 30930 20
rect 31000 80 31100 100
rect 31000 20 31020 80
rect 31080 20 31100 80
rect 31000 0 31100 20
rect 31170 80 31270 100
rect 31170 20 31190 80
rect 31250 20 31270 80
rect 31170 0 31270 20
rect 31340 80 31440 100
rect 31340 20 31360 80
rect 31420 20 31440 80
rect 31340 0 31440 20
rect 31510 80 31610 100
rect 31510 20 31530 80
rect 31590 20 31610 80
rect 31510 0 31610 20
rect 31680 80 31780 100
rect 31680 20 31700 80
rect 31760 20 31780 80
rect 31680 0 31780 20
rect 31850 80 31950 100
rect 31850 20 31870 80
rect 31930 20 31950 80
rect 31850 0 31950 20
rect 32020 80 32120 100
rect 32020 20 32040 80
rect 32100 20 32120 80
rect 32020 0 32120 20
rect 32190 80 32290 100
rect 32190 20 32210 80
rect 32270 20 32290 80
rect 32190 0 32290 20
rect 32360 80 32460 100
rect 32360 20 32380 80
rect 32440 20 32460 80
rect 32360 0 32460 20
rect 32530 80 32630 100
rect 32530 20 32550 80
rect 32610 20 32630 80
rect 32530 0 32630 20
rect 32700 80 32800 100
rect 32700 20 32720 80
rect 32780 20 32800 80
rect 32700 0 32800 20
rect 32870 80 32970 100
rect 32870 20 32890 80
rect 32950 20 32970 80
rect 32870 0 32970 20
rect 33040 80 33140 100
rect 33040 20 33060 80
rect 33120 20 33140 80
rect 33040 0 33140 20
rect 33210 80 33310 100
rect 33210 20 33230 80
rect 33290 20 33310 80
rect 33210 0 33310 20
rect 33380 80 33480 100
rect 33380 20 33400 80
rect 33460 20 33480 80
rect 33380 0 33480 20
rect 33550 80 33650 100
rect 33550 20 33570 80
rect 33630 20 33650 80
rect 33550 0 33650 20
rect 33720 80 33820 100
rect 33720 20 33740 80
rect 33800 20 33820 80
rect 33720 0 33820 20
rect 33890 80 33990 100
rect 33890 20 33910 80
rect 33970 20 33990 80
rect 33890 0 33990 20
rect 34060 80 34160 100
rect 34060 20 34080 80
rect 34140 20 34160 80
rect 34060 0 34160 20
rect 34230 80 34330 100
rect 34230 20 34250 80
rect 34310 20 34330 80
rect 34230 0 34330 20
rect 34400 80 34500 100
rect 34400 20 34420 80
rect 34480 20 34500 80
rect 34400 0 34500 20
rect 34570 80 34670 100
rect 34570 20 34590 80
rect 34650 20 34670 80
rect 34570 0 34670 20
rect 34740 80 34840 100
rect 34740 20 34760 80
rect 34820 20 34840 80
rect 34740 0 34840 20
rect 34910 80 35010 100
rect 34910 20 34930 80
rect 34990 20 35010 80
rect 34910 0 35010 20
rect 35080 80 35180 100
rect 35080 20 35100 80
rect 35160 20 35180 80
rect 35080 0 35180 20
rect 35250 80 35350 100
rect 35250 20 35270 80
rect 35330 20 35350 80
rect 35250 0 35350 20
rect 35420 80 35520 100
rect 35420 20 35440 80
rect 35500 20 35520 80
rect 35420 0 35520 20
rect 35590 80 35690 100
rect 35590 20 35610 80
rect 35670 20 35690 80
rect 35590 0 35690 20
rect 35760 80 35860 100
rect 35760 20 35780 80
rect 35840 20 35860 80
rect 35760 0 35860 20
rect 35930 80 36030 100
rect 35930 20 35950 80
rect 36010 20 36030 80
rect 35930 0 36030 20
rect 36100 80 36200 100
rect 36100 20 36120 80
rect 36180 20 36200 80
rect 36100 0 36200 20
rect 36270 80 36370 100
rect 36270 20 36290 80
rect 36350 20 36370 80
rect 36270 0 36370 20
rect 36440 80 36540 100
rect 36440 20 36460 80
rect 36520 20 36540 80
rect 36440 0 36540 20
rect 36610 80 36710 100
rect 36610 20 36630 80
rect 36690 20 36710 80
rect 36610 0 36710 20
rect 36780 80 36880 100
rect 36780 20 36800 80
rect 36860 20 36880 80
rect 36780 0 36880 20
rect 36950 80 37050 100
rect 36950 20 36970 80
rect 37030 20 37050 80
rect 36950 0 37050 20
rect 37120 80 37220 100
rect 37120 20 37140 80
rect 37200 20 37220 80
rect 37120 0 37220 20
rect 37290 80 37390 100
rect 37290 20 37310 80
rect 37370 20 37390 80
rect 37290 0 37390 20
rect 37460 80 37560 100
rect 37460 20 37480 80
rect 37540 20 37560 80
rect 37460 0 37560 20
rect 37630 80 37730 100
rect 37630 20 37650 80
rect 37710 20 37730 80
rect 37630 0 37730 20
rect 37800 80 37900 100
rect 37800 20 37820 80
rect 37880 20 37900 80
rect 37800 0 37900 20
rect 37970 80 38070 100
rect 37970 20 37990 80
rect 38050 20 38070 80
rect 37970 0 38070 20
rect 38140 80 38240 100
rect 38140 20 38160 80
rect 38220 20 38240 80
rect 38140 0 38240 20
rect 38310 80 38410 100
rect 38310 20 38330 80
rect 38390 20 38410 80
rect 38310 0 38410 20
rect 38480 80 38580 100
rect 38480 20 38500 80
rect 38560 20 38580 80
rect 38480 0 38580 20
rect 38650 80 38750 100
rect 38650 20 38670 80
rect 38730 20 38750 80
rect 38650 0 38750 20
rect 38820 80 38920 100
rect 38820 20 38840 80
rect 38900 20 38920 80
rect 38820 0 38920 20
rect 38990 80 39090 100
rect 38990 20 39010 80
rect 39070 20 39090 80
rect 38990 0 39090 20
rect 39160 80 39260 100
rect 39160 20 39180 80
rect 39240 20 39260 80
rect 39160 0 39260 20
rect 39330 80 39430 100
rect 39330 20 39350 80
rect 39410 20 39430 80
rect 39330 0 39430 20
rect 39500 80 39600 100
rect 39500 20 39520 80
rect 39580 20 39600 80
rect 39500 0 39600 20
rect 39670 80 39770 100
rect 39670 20 39690 80
rect 39750 20 39770 80
rect 39670 0 39770 20
rect 39840 80 39940 100
rect 39840 20 39860 80
rect 39920 20 39940 80
rect 39840 0 39940 20
rect 40010 80 40110 100
rect 40010 20 40030 80
rect 40090 20 40110 80
rect 40010 0 40110 20
rect 40180 80 40280 100
rect 40180 20 40200 80
rect 40260 20 40280 80
rect 40180 0 40280 20
rect 40350 80 40450 100
rect 40350 20 40370 80
rect 40430 20 40450 80
rect 40350 0 40450 20
rect 40520 80 40620 100
rect 40520 20 40540 80
rect 40600 20 40620 80
rect 40520 0 40620 20
rect 40690 80 40790 100
rect 40690 20 40710 80
rect 40770 20 40790 80
rect 40690 0 40790 20
rect 40860 80 40960 100
rect 40860 20 40880 80
rect 40940 20 40960 80
rect 40860 0 40960 20
rect 41030 80 41130 100
rect 41030 20 41050 80
rect 41110 20 41130 80
rect 41030 0 41130 20
rect 41200 80 41300 100
rect 41200 20 41220 80
rect 41280 20 41300 80
rect 41200 0 41300 20
rect 41370 80 41470 100
rect 41370 20 41390 80
rect 41450 20 41470 80
rect 41370 0 41470 20
rect 41540 80 41640 100
rect 41540 20 41560 80
rect 41620 20 41640 80
rect 41540 0 41640 20
rect 41710 80 41810 100
rect 41710 20 41730 80
rect 41790 20 41810 80
rect 41710 0 41810 20
rect 41880 80 41980 100
rect 41880 20 41900 80
rect 41960 20 41980 80
rect 41880 0 41980 20
rect 42050 80 42150 100
rect 42050 20 42070 80
rect 42130 20 42150 80
rect 42050 0 42150 20
rect 42220 80 42320 100
rect 42220 20 42240 80
rect 42300 20 42320 80
rect 42220 0 42320 20
rect 42390 80 42490 100
rect 42390 20 42410 80
rect 42470 20 42490 80
rect 42390 0 42490 20
rect 42560 80 42660 100
rect 42560 20 42580 80
rect 42640 20 42660 80
rect 42560 0 42660 20
rect 42730 80 42830 100
rect 42730 20 42750 80
rect 42810 20 42830 80
rect 42730 0 42830 20
rect 42900 80 43000 100
rect 42900 20 42920 80
rect 42980 20 43000 80
rect 42900 0 43000 20
rect 43070 80 43170 100
rect 43070 20 43090 80
rect 43150 20 43170 80
rect 43070 0 43170 20
rect 43240 80 43340 100
rect 43240 20 43260 80
rect 43320 20 43340 80
rect 43240 0 43340 20
rect 43410 80 43510 100
rect 43410 20 43430 80
rect 43490 20 43510 80
rect 43410 0 43510 20
rect 43580 80 43680 100
rect 43580 20 43600 80
rect 43660 20 43680 80
rect 43580 0 43680 20
rect 43750 80 43850 100
rect 43750 20 43770 80
rect 43830 20 43850 80
rect 43750 0 43850 20
rect 43920 80 44020 100
rect 43920 20 43940 80
rect 44000 20 44020 80
rect 43920 0 44020 20
rect 44090 80 44190 100
rect 44090 20 44110 80
rect 44170 20 44190 80
rect 44090 0 44190 20
rect 44260 80 44360 100
rect 44260 20 44280 80
rect 44340 20 44360 80
rect 44260 0 44360 20
rect 44430 80 44530 100
rect 44430 20 44450 80
rect 44510 20 44530 80
rect 44430 0 44530 20
rect 44600 80 44700 100
rect 44600 20 44620 80
rect 44680 20 44700 80
rect 44600 0 44700 20
rect 44770 80 44870 100
rect 44770 20 44790 80
rect 44850 20 44870 80
rect 44770 0 44870 20
rect 44940 80 45040 100
rect 44940 20 44960 80
rect 45020 20 45040 80
rect 44940 0 45040 20
rect 45110 80 45210 100
rect 45110 20 45130 80
rect 45190 20 45210 80
rect 45110 0 45210 20
rect 45280 80 45380 100
rect 45280 20 45300 80
rect 45360 20 45380 80
rect 45280 0 45380 20
rect 45450 80 45550 100
rect 45450 20 45470 80
rect 45530 20 45550 80
rect 45450 0 45550 20
rect 45620 80 45720 100
rect 45620 20 45640 80
rect 45700 20 45720 80
rect 45620 0 45720 20
rect 45790 80 45890 100
rect 45790 20 45810 80
rect 45870 20 45890 80
rect 45790 0 45890 20
rect 45960 80 46060 100
rect 45960 20 45980 80
rect 46040 20 46060 80
rect 45960 0 46060 20
rect 46130 80 46230 100
rect 46130 20 46150 80
rect 46210 20 46230 80
rect 46130 0 46230 20
rect 46300 80 46400 100
rect 46300 20 46320 80
rect 46380 20 46400 80
rect 46300 0 46400 20
rect 46470 80 46570 100
rect 46470 20 46490 80
rect 46550 20 46570 80
rect 46470 0 46570 20
rect 46640 80 46740 100
rect 46640 20 46660 80
rect 46720 20 46740 80
rect 46640 0 46740 20
rect 46810 80 46910 100
rect 46810 20 46830 80
rect 46890 20 46910 80
rect 46810 0 46910 20
rect 46980 80 47080 100
rect 46980 20 47000 80
rect 47060 20 47080 80
rect 46980 0 47080 20
rect 47150 80 47250 100
rect 47150 20 47170 80
rect 47230 20 47250 80
rect 47150 0 47250 20
rect 47320 80 47420 100
rect 47320 20 47340 80
rect 47400 20 47420 80
rect 47320 0 47420 20
rect 47490 80 47590 100
rect 47490 20 47510 80
rect 47570 20 47590 80
rect 47490 0 47590 20
rect 47660 80 47760 100
rect 47660 20 47680 80
rect 47740 20 47760 80
rect 47660 0 47760 20
rect 47830 80 47930 100
rect 47830 20 47850 80
rect 47910 20 47930 80
rect 47830 0 47930 20
rect 48000 80 48100 100
rect 48000 20 48020 80
rect 48080 20 48100 80
rect 48000 0 48100 20
rect 48170 80 48270 100
rect 48170 20 48190 80
rect 48250 20 48270 80
rect 48170 0 48270 20
rect 48340 80 48440 100
rect 48340 20 48360 80
rect 48420 20 48440 80
rect 48340 0 48440 20
rect 48510 80 48610 100
rect 48510 20 48530 80
rect 48590 20 48610 80
rect 48510 0 48610 20
rect 48680 80 48780 100
rect 48680 20 48700 80
rect 48760 20 48780 80
rect 48680 0 48780 20
rect 48850 80 48950 100
rect 48850 20 48870 80
rect 48930 20 48950 80
rect 48850 0 48950 20
rect 49020 80 49120 100
rect 49020 20 49040 80
rect 49100 20 49120 80
rect 49020 0 49120 20
rect 49190 80 49290 100
rect 49190 20 49210 80
rect 49270 20 49290 80
rect 49190 0 49290 20
rect 49360 80 49460 100
rect 49360 20 49380 80
rect 49440 20 49460 80
rect 49360 0 49460 20
rect 49530 80 49630 100
rect 49530 20 49550 80
rect 49610 20 49630 80
rect 49530 0 49630 20
rect 49700 80 49800 100
rect 49700 20 49720 80
rect 49780 20 49800 80
rect 49700 0 49800 20
rect 49870 80 49970 100
rect 49870 20 49890 80
rect 49950 20 49970 80
rect 49870 0 49970 20
rect 50040 80 50140 100
rect 50040 20 50060 80
rect 50120 20 50140 80
rect 50040 0 50140 20
rect 50210 80 50310 100
rect 50210 20 50230 80
rect 50290 20 50310 80
rect 50210 0 50310 20
rect 50380 80 50480 100
rect 50380 20 50400 80
rect 50460 20 50480 80
rect 50380 0 50480 20
rect 50550 80 50650 100
rect 50550 20 50570 80
rect 50630 20 50650 80
rect 50550 0 50650 20
rect 50720 80 50820 100
rect 50720 20 50740 80
rect 50800 20 50820 80
rect 50720 0 50820 20
rect 50890 80 50990 100
rect 50890 20 50910 80
rect 50970 20 50990 80
rect 50890 0 50990 20
rect 51060 80 51160 100
rect 51060 20 51080 80
rect 51140 20 51160 80
rect 51060 0 51160 20
rect 51230 80 51330 100
rect 51230 20 51250 80
rect 51310 20 51330 80
rect 51230 0 51330 20
rect 51400 80 51500 100
rect 51400 20 51420 80
rect 51480 20 51500 80
rect 51400 0 51500 20
rect 51570 80 51670 100
rect 51570 20 51590 80
rect 51650 20 51670 80
rect 51570 0 51670 20
rect 51740 80 51840 100
rect 51740 20 51760 80
rect 51820 20 51840 80
rect 51740 0 51840 20
rect 51910 80 52010 100
rect 51910 20 51930 80
rect 51990 20 52010 80
rect 51910 0 52010 20
rect 52080 80 52180 100
rect 52080 20 52100 80
rect 52160 20 52180 80
rect 52080 0 52180 20
rect 52250 80 52350 100
rect 52250 20 52270 80
rect 52330 20 52350 80
rect 52250 0 52350 20
rect 52420 80 52520 100
rect 52420 20 52440 80
rect 52500 20 52520 80
rect 52420 0 52520 20
rect 52590 80 52690 100
rect 52590 20 52610 80
rect 52670 20 52690 80
rect 52590 0 52690 20
rect 52760 80 52860 100
rect 52760 20 52780 80
rect 52840 20 52860 80
rect 52760 0 52860 20
rect 52930 80 53030 100
rect 52930 20 52950 80
rect 53010 20 53030 80
rect 52930 0 53030 20
rect 53100 80 53200 100
rect 53100 20 53120 80
rect 53180 20 53200 80
rect 53100 0 53200 20
rect 53270 80 53370 100
rect 53270 20 53290 80
rect 53350 20 53370 80
rect 53270 0 53370 20
rect 53440 80 53540 100
rect 53440 20 53460 80
rect 53520 20 53540 80
rect 53440 0 53540 20
rect 53610 80 53710 100
rect 53610 20 53630 80
rect 53690 20 53710 80
rect 53610 0 53710 20
rect 53780 80 53880 100
rect 53780 20 53800 80
rect 53860 20 53880 80
rect 53780 0 53880 20
rect 53950 80 54050 100
rect 53950 20 53970 80
rect 54030 20 54050 80
rect 53950 0 54050 20
rect 54120 80 54220 100
rect 54120 20 54140 80
rect 54200 20 54220 80
rect 54120 0 54220 20
rect 54290 80 54390 100
rect 54290 20 54310 80
rect 54370 20 54390 80
rect 54290 0 54390 20
rect 54460 80 54560 100
rect 54460 20 54480 80
rect 54540 20 54560 80
rect 54460 0 54560 20
rect 54630 80 54730 100
rect 54630 20 54650 80
rect 54710 20 54730 80
rect 54630 0 54730 20
rect 54800 80 54900 100
rect 54800 20 54820 80
rect 54880 20 54900 80
rect 54800 0 54900 20
rect 54970 80 55070 100
rect 54970 20 54990 80
rect 55050 20 55070 80
rect 54970 0 55070 20
rect 55140 80 55240 100
rect 55140 20 55160 80
rect 55220 20 55240 80
rect 55140 0 55240 20
rect 55310 80 55410 100
rect 55310 20 55330 80
rect 55390 20 55410 80
rect 55310 0 55410 20
rect 55480 80 55580 100
rect 55480 20 55500 80
rect 55560 20 55580 80
rect 55480 0 55580 20
rect 55650 80 55750 100
rect 55650 20 55670 80
rect 55730 20 55750 80
rect 55650 0 55750 20
rect 55820 80 55920 100
rect 55820 20 55840 80
rect 55900 20 55920 80
rect 55820 0 55920 20
rect 55990 80 56090 100
rect 55990 20 56010 80
rect 56070 20 56090 80
rect 55990 0 56090 20
rect 56160 80 56260 100
rect 56160 20 56180 80
rect 56240 20 56260 80
rect 56160 0 56260 20
rect 56330 80 56430 100
rect 56330 20 56350 80
rect 56410 20 56430 80
rect 56330 0 56430 20
rect 56500 80 56600 100
rect 56500 20 56520 80
rect 56580 20 56600 80
rect 56500 0 56600 20
rect 56670 80 56770 100
rect 56670 20 56690 80
rect 56750 20 56770 80
rect 56670 0 56770 20
rect 56840 80 56940 100
rect 56840 20 56860 80
rect 56920 20 56940 80
rect 56840 0 56940 20
rect 57010 80 57110 100
rect 57010 20 57030 80
rect 57090 20 57110 80
rect 57010 0 57110 20
rect 57180 80 57280 100
rect 57180 20 57200 80
rect 57260 20 57280 80
rect 57180 0 57280 20
rect 57350 80 57450 100
rect 57350 20 57370 80
rect 57430 20 57450 80
rect 57350 0 57450 20
rect 57520 80 57620 100
rect 57520 20 57540 80
rect 57600 20 57620 80
rect 57520 0 57620 20
rect 57690 80 57790 100
rect 57690 20 57710 80
rect 57770 20 57790 80
rect 57690 0 57790 20
rect 57860 80 57960 100
rect 57860 20 57880 80
rect 57940 20 57960 80
rect 57860 0 57960 20
rect 58030 80 58130 100
rect 58030 20 58050 80
rect 58110 20 58130 80
rect 58030 0 58130 20
rect 58200 80 58300 100
rect 58200 20 58220 80
rect 58280 20 58300 80
rect 58200 0 58300 20
rect 58370 80 58470 100
rect 58370 20 58390 80
rect 58450 20 58470 80
rect 58370 0 58470 20
rect 58540 80 58640 100
rect 58540 20 58560 80
rect 58620 20 58640 80
rect 58540 0 58640 20
rect 58710 80 58810 100
rect 58710 20 58730 80
rect 58790 20 58810 80
rect 58710 0 58810 20
rect 58880 80 58980 100
rect 58880 20 58900 80
rect 58960 20 58980 80
rect 58880 0 58980 20
rect 59050 80 59150 100
rect 59050 20 59070 80
rect 59130 20 59150 80
rect 59050 0 59150 20
rect 59220 80 59320 100
rect 59220 20 59240 80
rect 59300 20 59320 80
rect 59220 0 59320 20
rect 10 -60 110 -40
rect 10 -120 30 -60
rect 90 -120 110 -60
rect 10 -140 110 -120
rect 180 -60 280 -40
rect 180 -120 200 -60
rect 260 -120 280 -60
rect 180 -140 280 -120
rect 510 -60 620 -40
rect 510 -120 530 -60
rect 600 -120 620 -60
rect 510 -140 620 -120
rect 680 -60 790 -40
rect 680 -120 700 -60
rect 770 -120 790 -60
rect 680 -140 790 -120
rect 850 -60 960 -40
rect 850 -120 870 -60
rect 940 -120 960 -60
rect 850 -140 960 -120
rect 1020 -60 1130 -40
rect 1020 -120 1040 -60
rect 1110 -120 1130 -60
rect 1020 -140 1130 -120
rect 1580 -60 1690 -40
rect 1580 -120 1600 -60
rect 1670 -120 1690 -60
rect 1580 -140 1690 -120
rect 1750 -60 1860 -40
rect 1750 -120 1770 -60
rect 1840 -120 1860 -60
rect 1750 -140 1860 -120
rect 1920 -60 2030 -40
rect 1920 -120 1940 -60
rect 2010 -120 2030 -60
rect 1920 -140 2030 -120
rect 2090 -60 2200 -40
rect 2090 -120 2110 -60
rect 2180 -120 2200 -60
rect 2090 -140 2200 -120
rect 2260 -60 2370 -40
rect 2260 -120 2280 -60
rect 2350 -120 2370 -60
rect 2260 -140 2370 -120
rect 2430 -60 2540 -40
rect 2430 -120 2450 -60
rect 2520 -120 2540 -60
rect 2430 -140 2540 -120
rect 2600 -60 2710 -40
rect 2600 -120 2620 -60
rect 2690 -120 2710 -60
rect 2600 -140 2710 -120
rect 2770 -60 2880 -40
rect 2770 -120 2790 -60
rect 2860 -120 2880 -60
rect 2770 -140 2880 -120
rect 2940 -60 3050 -40
rect 2940 -120 2960 -60
rect 3030 -120 3050 -60
rect 2940 -140 3050 -120
rect 3110 -60 3220 -40
rect 3110 -120 3130 -60
rect 3200 -120 3220 -60
rect 3110 -140 3220 -120
rect 3280 -60 3390 -40
rect 3280 -120 3300 -60
rect 3370 -120 3390 -60
rect 3280 -140 3390 -120
rect 3450 -60 3560 -40
rect 3450 -120 3470 -60
rect 3540 -120 3560 -60
rect 3450 -140 3560 -120
rect 3620 -60 3730 -40
rect 3620 -120 3640 -60
rect 3710 -120 3730 -60
rect 3620 -140 3730 -120
rect 3790 -60 3900 -40
rect 3790 -120 3810 -60
rect 3880 -120 3900 -60
rect 3790 -140 3900 -120
rect 3960 -60 4070 -40
rect 3960 -120 3980 -60
rect 4050 -120 4070 -60
rect 3960 -140 4070 -120
rect 4130 -60 4240 -40
rect 4130 -120 4150 -60
rect 4220 -120 4240 -60
rect 4130 -140 4240 -120
rect 4600 -60 4710 -40
rect 4600 -120 4620 -60
rect 4690 -120 4710 -60
rect 4600 -140 4710 -120
rect 4770 -60 4880 -40
rect 4770 -120 4790 -60
rect 4860 -120 4880 -60
rect 4770 -140 4880 -120
rect 4940 -60 5050 -40
rect 4940 -120 4960 -60
rect 5030 -120 5050 -60
rect 4940 -140 5050 -120
rect 5110 -60 5220 -40
rect 5110 -120 5130 -60
rect 5200 -120 5220 -60
rect 5110 -140 5220 -120
rect 5280 -60 5390 -40
rect 5280 -120 5300 -60
rect 5370 -120 5390 -60
rect 5280 -140 5390 -120
rect 5450 -60 5560 -40
rect 5450 -120 5470 -60
rect 5540 -120 5560 -60
rect 5450 -140 5560 -120
rect 5620 -60 5730 -40
rect 5620 -120 5640 -60
rect 5710 -120 5730 -60
rect 5620 -140 5730 -120
rect 5790 -60 5900 -40
rect 5790 -120 5810 -60
rect 5880 -120 5900 -60
rect 5790 -140 5900 -120
rect 5960 -60 6070 -40
rect 5960 -120 5980 -60
rect 6050 -120 6070 -60
rect 5960 -140 6070 -120
rect 6130 -60 6240 -40
rect 6130 -120 6150 -60
rect 6220 -120 6240 -60
rect 6130 -140 6240 -120
rect 6300 -60 6410 -40
rect 6300 -120 6320 -60
rect 6390 -120 6410 -60
rect 6300 -140 6410 -120
rect 6470 -60 6580 -40
rect 6470 -120 6490 -60
rect 6560 -120 6580 -60
rect 6470 -140 6580 -120
rect 6640 -60 6750 -40
rect 6640 -120 6660 -60
rect 6730 -120 6750 -60
rect 6640 -140 6750 -120
rect 6810 -60 6920 -40
rect 6810 -120 6830 -60
rect 6900 -120 6920 -60
rect 6810 -140 6920 -120
rect 6980 -60 7090 -40
rect 6980 -120 7000 -60
rect 7070 -120 7090 -60
rect 6980 -140 7090 -120
rect 7150 -60 7260 -40
rect 7150 -120 7170 -60
rect 7240 -120 7260 -60
rect 7150 -140 7260 -120
rect 7320 -60 7430 -40
rect 7320 -120 7340 -60
rect 7410 -120 7430 -60
rect 7320 -140 7430 -120
rect 7490 -60 7600 -40
rect 7490 -120 7510 -60
rect 7580 -120 7600 -60
rect 7490 -140 7600 -120
rect 7660 -60 7770 -40
rect 7660 -120 7680 -60
rect 7750 -120 7770 -60
rect 7660 -140 7770 -120
rect 7830 -60 7940 -40
rect 7830 -120 7850 -60
rect 7920 -120 7940 -60
rect 7830 -140 7940 -120
rect 8000 -60 8110 -40
rect 8000 -120 8020 -60
rect 8090 -120 8110 -60
rect 8000 -140 8110 -120
rect 8170 -60 8280 -40
rect 8170 -120 8190 -60
rect 8260 -120 8280 -60
rect 8170 -140 8280 -120
rect 8340 -60 8450 -40
rect 8340 -120 8360 -60
rect 8430 -120 8450 -60
rect 8340 -140 8450 -120
rect 8510 -60 8620 -40
rect 8510 -120 8530 -60
rect 8600 -120 8620 -60
rect 8510 -140 8620 -120
rect 8680 -60 8790 -40
rect 8680 -120 8700 -60
rect 8770 -120 8790 -60
rect 8680 -140 8790 -120
rect 8850 -60 8960 -40
rect 8850 -120 8870 -60
rect 8940 -120 8960 -60
rect 8850 -140 8960 -120
rect 9020 -60 9130 -40
rect 9020 -120 9040 -60
rect 9110 -120 9130 -60
rect 9020 -140 9130 -120
rect 9190 -60 9300 -40
rect 9190 -120 9210 -60
rect 9280 -120 9300 -60
rect 9190 -140 9300 -120
rect 9360 -60 9470 -40
rect 9360 -120 9380 -60
rect 9450 -120 9470 -60
rect 9360 -140 9470 -120
rect 9530 -60 9640 -40
rect 9530 -120 9550 -60
rect 9620 -120 9640 -60
rect 9530 -140 9640 -120
rect 9700 -60 9810 -40
rect 9700 -120 9720 -60
rect 9790 -120 9810 -60
rect 9700 -140 9810 -120
rect 9870 -60 9980 -40
rect 9870 -120 9890 -60
rect 9960 -120 9980 -60
rect 9870 -140 9980 -120
rect 10040 -60 10150 -40
rect 10040 -120 10060 -60
rect 10130 -120 10150 -60
rect 10040 -140 10150 -120
rect 10210 -60 10320 -40
rect 10210 -120 10230 -60
rect 10300 -120 10320 -60
rect 10210 -140 10320 -120
rect 10380 -60 10490 -40
rect 10380 -120 10400 -60
rect 10470 -120 10490 -60
rect 10380 -140 10490 -120
rect 10550 -60 10660 -40
rect 10550 -120 10570 -60
rect 10640 -120 10660 -60
rect 10550 -140 10660 -120
rect 10720 -60 10830 -40
rect 10720 -120 10740 -60
rect 10810 -120 10830 -60
rect 10720 -140 10830 -120
rect 10890 -60 11000 -40
rect 10890 -120 10910 -60
rect 10980 -120 11000 -60
rect 10890 -140 11000 -120
rect 11060 -60 11170 -40
rect 11060 -120 11080 -60
rect 11150 -120 11170 -60
rect 11060 -140 11170 -120
rect 11230 -60 11340 -40
rect 11230 -120 11250 -60
rect 11320 -120 11340 -60
rect 11230 -140 11340 -120
rect 11400 -60 11510 -40
rect 11400 -120 11420 -60
rect 11490 -120 11510 -60
rect 11400 -140 11510 -120
rect 11570 -60 11680 -40
rect 11570 -120 11590 -60
rect 11660 -120 11680 -60
rect 11570 -140 11680 -120
rect 11740 -60 11850 -40
rect 11740 -120 11760 -60
rect 11830 -120 11850 -60
rect 11740 -140 11850 -120
rect 11910 -60 12020 -40
rect 11910 -120 11930 -60
rect 12000 -120 12020 -60
rect 11910 -140 12020 -120
rect 12080 -60 12190 -40
rect 12080 -120 12100 -60
rect 12170 -120 12190 -60
rect 12080 -140 12190 -120
rect 12250 -60 12360 -40
rect 12250 -120 12270 -60
rect 12340 -120 12360 -60
rect 12250 -140 12360 -120
rect 12420 -60 12530 -40
rect 12420 -120 12440 -60
rect 12510 -120 12530 -60
rect 12420 -140 12530 -120
rect 12590 -60 12700 -40
rect 12590 -120 12610 -60
rect 12680 -120 12700 -60
rect 12590 -140 12700 -120
rect 12760 -60 12870 -40
rect 12760 -120 12780 -60
rect 12850 -120 12870 -60
rect 12760 -140 12870 -120
rect 12930 -60 13040 -40
rect 12930 -120 12950 -60
rect 13020 -120 13040 -60
rect 12930 -140 13040 -120
rect 13100 -60 13210 -40
rect 13100 -120 13120 -60
rect 13190 -120 13210 -60
rect 13100 -140 13210 -120
rect 13270 -60 13380 -40
rect 13270 -120 13290 -60
rect 13360 -120 13380 -60
rect 13270 -140 13380 -120
rect 13440 -60 13550 -40
rect 13440 -120 13460 -60
rect 13530 -120 13550 -60
rect 13440 -140 13550 -120
rect 13610 -60 13720 -40
rect 13610 -120 13630 -60
rect 13700 -120 13720 -60
rect 13610 -140 13720 -120
rect 13780 -60 13890 -40
rect 13780 -120 13800 -60
rect 13870 -120 13890 -60
rect 13780 -140 13890 -120
rect 13950 -60 14060 -40
rect 13950 -120 13970 -60
rect 14040 -120 14060 -60
rect 13950 -140 14060 -120
rect 14120 -60 14230 -40
rect 14120 -120 14140 -60
rect 14210 -120 14230 -60
rect 14120 -140 14230 -120
rect 14290 -60 14400 -40
rect 14290 -120 14310 -60
rect 14380 -120 14400 -60
rect 14290 -140 14400 -120
rect 14460 -60 14570 -40
rect 14460 -120 14480 -60
rect 14550 -120 14570 -60
rect 14460 -140 14570 -120
rect 14630 -60 14740 -40
rect 14630 -120 14650 -60
rect 14720 -120 14740 -60
rect 14630 -140 14740 -120
rect 14800 -60 14910 -40
rect 14800 -120 14820 -60
rect 14890 -120 14910 -60
rect 14800 -140 14910 -120
rect 14970 -60 15080 -40
rect 14970 -120 14990 -60
rect 15060 -120 15080 -60
rect 14970 -140 15080 -120
rect 15140 -60 15250 -40
rect 15140 -120 15160 -60
rect 15230 -120 15250 -60
rect 15140 -140 15250 -120
rect 15310 -60 15420 -40
rect 15310 -120 15330 -60
rect 15400 -120 15420 -60
rect 15310 -140 15420 -120
rect 15780 -60 15890 -40
rect 15780 -120 15800 -60
rect 15870 -120 15890 -60
rect 15780 -140 15890 -120
rect 15950 -60 16060 -40
rect 15950 -120 15970 -60
rect 16040 -120 16060 -60
rect 15950 -140 16060 -120
rect 16120 -60 16230 -40
rect 16120 -120 16140 -60
rect 16210 -120 16230 -60
rect 16120 -140 16230 -120
rect 16290 -60 16400 -40
rect 16290 -120 16310 -60
rect 16380 -120 16400 -60
rect 16290 -140 16400 -120
rect 16460 -60 16570 -40
rect 16460 -120 16480 -60
rect 16550 -120 16570 -60
rect 16460 -140 16570 -120
rect 16630 -60 16740 -40
rect 16630 -120 16650 -60
rect 16720 -120 16740 -60
rect 16630 -140 16740 -120
rect 16800 -60 16910 -40
rect 16800 -120 16820 -60
rect 16890 -120 16910 -60
rect 16800 -140 16910 -120
rect 16970 -60 17080 -40
rect 16970 -120 16990 -60
rect 17060 -120 17080 -60
rect 16970 -140 17080 -120
rect 17140 -60 17250 -40
rect 17140 -120 17160 -60
rect 17230 -120 17250 -60
rect 17140 -140 17250 -120
rect 17310 -60 17420 -40
rect 17310 -120 17330 -60
rect 17400 -120 17420 -60
rect 17310 -140 17420 -120
rect 17480 -60 17590 -40
rect 17480 -120 17500 -60
rect 17570 -120 17590 -60
rect 17480 -140 17590 -120
rect 17650 -60 17760 -40
rect 17650 -120 17670 -60
rect 17740 -120 17760 -60
rect 17650 -140 17760 -120
rect 17820 -60 17930 -40
rect 17820 -120 17840 -60
rect 17910 -120 17930 -60
rect 17820 -140 17930 -120
rect 17990 -60 18100 -40
rect 17990 -120 18010 -60
rect 18080 -120 18100 -60
rect 17990 -140 18100 -120
rect 18160 -60 18270 -40
rect 18160 -120 18180 -60
rect 18250 -120 18270 -60
rect 18160 -140 18270 -120
rect 18330 -60 18440 -40
rect 18330 -120 18350 -60
rect 18420 -120 18440 -60
rect 18330 -140 18440 -120
rect 18500 -60 18610 -40
rect 18500 -120 18520 -60
rect 18590 -120 18610 -60
rect 18500 -140 18610 -120
rect 18670 -60 18780 -40
rect 18670 -120 18690 -60
rect 18760 -120 18780 -60
rect 18670 -140 18780 -120
rect 18840 -60 18950 -40
rect 18840 -120 18860 -60
rect 18930 -120 18950 -60
rect 18840 -140 18950 -120
rect 19010 -60 19120 -40
rect 19010 -120 19030 -60
rect 19100 -120 19120 -60
rect 19010 -140 19120 -120
rect 19180 -60 19290 -40
rect 19180 -120 19200 -60
rect 19270 -120 19290 -60
rect 19180 -140 19290 -120
rect 19350 -60 19460 -40
rect 19350 -120 19370 -60
rect 19440 -120 19460 -60
rect 19350 -140 19460 -120
rect 19520 -60 19630 -40
rect 19520 -120 19540 -60
rect 19610 -120 19630 -60
rect 19520 -140 19630 -120
rect 19690 -60 19800 -40
rect 19690 -120 19710 -60
rect 19780 -120 19800 -60
rect 19690 -140 19800 -120
rect 19860 -60 19970 -40
rect 19860 -120 19880 -60
rect 19950 -120 19970 -60
rect 19860 -140 19970 -120
rect 20030 -60 20140 -40
rect 20030 -120 20050 -60
rect 20120 -120 20140 -60
rect 20030 -140 20140 -120
rect 20200 -60 20310 -40
rect 20200 -120 20220 -60
rect 20290 -120 20310 -60
rect 20200 -140 20310 -120
rect 20370 -60 20480 -40
rect 20370 -120 20390 -60
rect 20460 -120 20480 -60
rect 20370 -140 20480 -120
rect 20540 -60 20650 -40
rect 20540 -120 20560 -60
rect 20630 -120 20650 -60
rect 20540 -140 20650 -120
rect 20710 -60 20820 -40
rect 20710 -120 20730 -60
rect 20800 -120 20820 -60
rect 20710 -140 20820 -120
rect 20880 -60 20990 -40
rect 20880 -120 20900 -60
rect 20970 -120 20990 -60
rect 20880 -140 20990 -120
rect 21050 -60 21160 -40
rect 21050 -120 21070 -60
rect 21140 -120 21160 -60
rect 21050 -140 21160 -120
rect 21220 -60 21330 -40
rect 21220 -120 21240 -60
rect 21310 -120 21330 -60
rect 21220 -140 21330 -120
rect 21390 -60 21500 -40
rect 21390 -120 21410 -60
rect 21480 -120 21500 -60
rect 21390 -140 21500 -120
rect 21560 -60 21670 -40
rect 21560 -120 21580 -60
rect 21650 -120 21670 -60
rect 21560 -140 21670 -120
rect 21730 -60 21840 -40
rect 21730 -120 21750 -60
rect 21820 -120 21840 -60
rect 21730 -140 21840 -120
rect 21900 -60 22010 -40
rect 21900 -120 21920 -60
rect 21990 -120 22010 -60
rect 21900 -140 22010 -120
rect 22070 -60 22180 -40
rect 22070 -120 22090 -60
rect 22160 -120 22180 -60
rect 22070 -140 22180 -120
rect 22240 -60 22350 -40
rect 22240 -120 22260 -60
rect 22330 -120 22350 -60
rect 22240 -140 22350 -120
rect 22410 -60 22520 -40
rect 22410 -120 22430 -60
rect 22500 -120 22520 -60
rect 22410 -140 22520 -120
rect 22580 -60 22690 -40
rect 22580 -120 22600 -60
rect 22670 -120 22690 -60
rect 22580 -140 22690 -120
rect 22750 -60 22860 -40
rect 22750 -120 22770 -60
rect 22840 -120 22860 -60
rect 22750 -140 22860 -120
rect 22920 -60 23030 -40
rect 22920 -120 22940 -60
rect 23010 -120 23030 -60
rect 22920 -140 23030 -120
rect 23090 -60 23200 -40
rect 23090 -120 23110 -60
rect 23180 -120 23200 -60
rect 23090 -140 23200 -120
rect 23260 -60 23370 -40
rect 23260 -120 23280 -60
rect 23350 -120 23370 -60
rect 23260 -140 23370 -120
rect 23430 -60 23540 -40
rect 23430 -120 23450 -60
rect 23520 -120 23540 -60
rect 23430 -140 23540 -120
rect 23600 -60 23710 -40
rect 23600 -120 23620 -60
rect 23690 -120 23710 -60
rect 23600 -140 23710 -120
rect 23770 -60 23880 -40
rect 23770 -120 23790 -60
rect 23860 -120 23880 -60
rect 23770 -140 23880 -120
rect 23940 -60 24050 -40
rect 23940 -120 23960 -60
rect 24030 -120 24050 -60
rect 23940 -140 24050 -120
rect 24110 -60 24220 -40
rect 24110 -120 24130 -60
rect 24200 -120 24220 -60
rect 24110 -140 24220 -120
rect 24280 -60 24390 -40
rect 24280 -120 24300 -60
rect 24370 -120 24390 -60
rect 24280 -140 24390 -120
rect 24450 -60 24560 -40
rect 24450 -120 24470 -60
rect 24540 -120 24560 -60
rect 24450 -140 24560 -120
rect 24620 -60 24730 -40
rect 24620 -120 24640 -60
rect 24710 -120 24730 -60
rect 24620 -140 24730 -120
rect 24790 -60 24900 -40
rect 24790 -120 24810 -60
rect 24880 -120 24900 -60
rect 24790 -140 24900 -120
rect 24960 -60 25070 -40
rect 24960 -120 24980 -60
rect 25050 -120 25070 -60
rect 24960 -140 25070 -120
rect 25130 -60 25240 -40
rect 25130 -120 25150 -60
rect 25220 -120 25240 -60
rect 25130 -140 25240 -120
rect 25300 -60 25410 -40
rect 25300 -120 25320 -60
rect 25390 -120 25410 -60
rect 25300 -140 25410 -120
rect 25470 -60 25580 -40
rect 25470 -120 25490 -60
rect 25560 -120 25580 -60
rect 25470 -140 25580 -120
rect 25640 -60 25750 -40
rect 25640 -120 25660 -60
rect 25730 -120 25750 -60
rect 25640 -140 25750 -120
rect 25810 -60 25920 -40
rect 25810 -120 25830 -60
rect 25900 -120 25920 -60
rect 25810 -140 25920 -120
rect 25980 -60 26090 -40
rect 25980 -120 26000 -60
rect 26070 -120 26090 -60
rect 25980 -140 26090 -120
rect 26150 -60 26260 -40
rect 26150 -120 26170 -60
rect 26240 -120 26260 -60
rect 26150 -140 26260 -120
rect 26320 -60 26430 -40
rect 26320 -120 26340 -60
rect 26410 -120 26430 -60
rect 26320 -140 26430 -120
rect 26490 -60 26600 -40
rect 26490 -120 26510 -60
rect 26580 -120 26600 -60
rect 26490 -140 26600 -120
rect 26660 -60 26770 -40
rect 26660 -120 26680 -60
rect 26750 -120 26770 -60
rect 26660 -140 26770 -120
rect 26830 -60 26940 -40
rect 26830 -120 26850 -60
rect 26920 -120 26940 -60
rect 26830 -140 26940 -120
rect 27000 -60 27110 -40
rect 27000 -120 27020 -60
rect 27090 -120 27110 -60
rect 27000 -140 27110 -120
rect 27170 -60 27280 -40
rect 27170 -120 27190 -60
rect 27260 -120 27280 -60
rect 27170 -140 27280 -120
rect 27340 -60 27450 -40
rect 27340 -120 27360 -60
rect 27430 -120 27450 -60
rect 27340 -140 27450 -120
rect 27510 -60 27620 -40
rect 27510 -120 27530 -60
rect 27600 -120 27620 -60
rect 27510 -140 27620 -120
rect 27680 -60 27790 -40
rect 27680 -120 27700 -60
rect 27770 -120 27790 -60
rect 27680 -140 27790 -120
rect 27850 -60 27960 -40
rect 27850 -120 27870 -60
rect 27940 -120 27960 -60
rect 27850 -140 27960 -120
rect 28020 -60 28130 -40
rect 28020 -120 28040 -60
rect 28110 -120 28130 -60
rect 28020 -140 28130 -120
rect 28190 -60 28300 -40
rect 28190 -120 28210 -60
rect 28280 -120 28300 -60
rect 28190 -140 28300 -120
rect 28360 -60 28470 -40
rect 28360 -120 28380 -60
rect 28450 -120 28470 -60
rect 28360 -140 28470 -120
rect 28530 -60 28640 -40
rect 28530 -120 28550 -60
rect 28620 -120 28640 -60
rect 28530 -140 28640 -120
rect 28700 -60 28810 -40
rect 28700 -120 28720 -60
rect 28790 -120 28810 -60
rect 28700 -140 28810 -120
rect 28870 -60 28980 -40
rect 28870 -120 28890 -60
rect 28960 -120 28980 -60
rect 28870 -140 28980 -120
rect 29040 -60 29150 -40
rect 29040 -120 29060 -60
rect 29130 -120 29150 -60
rect 29040 -140 29150 -120
rect 29210 -60 29320 -40
rect 29210 -120 29230 -60
rect 29300 -120 29320 -60
rect 29210 -140 29320 -120
rect 29380 -60 29490 -40
rect 29380 -120 29400 -60
rect 29470 -120 29490 -60
rect 29380 -140 29490 -120
rect 29550 -60 29660 -40
rect 29550 -120 29570 -60
rect 29640 -120 29660 -60
rect 29550 -140 29660 -120
rect 29720 -60 29830 -40
rect 29720 -120 29740 -60
rect 29810 -120 29830 -60
rect 29720 -140 29830 -120
rect 29890 -60 30000 -40
rect 29890 -120 29910 -60
rect 29980 -120 30000 -60
rect 29890 -140 30000 -120
rect 30060 -60 30170 -40
rect 30060 -120 30080 -60
rect 30150 -120 30170 -60
rect 30060 -140 30170 -120
rect 30230 -60 30340 -40
rect 30230 -120 30250 -60
rect 30320 -120 30340 -60
rect 30230 -140 30340 -120
rect 30400 -60 30510 -40
rect 30400 -120 30420 -60
rect 30490 -120 30510 -60
rect 30400 -140 30510 -120
rect 30570 -60 30680 -40
rect 30570 -120 30590 -60
rect 30660 -120 30680 -60
rect 30570 -140 30680 -120
rect 30740 -60 30850 -40
rect 30740 -120 30760 -60
rect 30830 -120 30850 -60
rect 30740 -140 30850 -120
rect 30910 -60 31020 -40
rect 30910 -120 30930 -60
rect 31000 -120 31020 -60
rect 30910 -140 31020 -120
rect 31080 -60 31190 -40
rect 31080 -120 31100 -60
rect 31170 -120 31190 -60
rect 31080 -140 31190 -120
rect 31250 -60 31360 -40
rect 31250 -120 31270 -60
rect 31340 -120 31360 -60
rect 31250 -140 31360 -120
rect 31420 -60 31530 -40
rect 31420 -120 31440 -60
rect 31510 -120 31530 -60
rect 31420 -140 31530 -120
rect 31590 -60 31700 -40
rect 31590 -120 31610 -60
rect 31680 -120 31700 -60
rect 31590 -140 31700 -120
rect 31760 -60 31870 -40
rect 31760 -120 31780 -60
rect 31850 -120 31870 -60
rect 31760 -140 31870 -120
rect 31930 -60 32040 -40
rect 31930 -120 31950 -60
rect 32020 -120 32040 -60
rect 31930 -140 32040 -120
rect 32100 -60 32210 -40
rect 32100 -120 32120 -60
rect 32190 -120 32210 -60
rect 32100 -140 32210 -120
rect 32270 -60 32380 -40
rect 32270 -120 32290 -60
rect 32360 -120 32380 -60
rect 32270 -140 32380 -120
rect 32440 -60 32550 -40
rect 32440 -120 32460 -60
rect 32530 -120 32550 -60
rect 32440 -140 32550 -120
rect 32610 -60 32720 -40
rect 32610 -120 32630 -60
rect 32700 -120 32720 -60
rect 32610 -140 32720 -120
rect 32780 -60 32890 -40
rect 32780 -120 32800 -60
rect 32870 -120 32890 -60
rect 32780 -140 32890 -120
rect 32950 -60 33060 -40
rect 32950 -120 32970 -60
rect 33040 -120 33060 -60
rect 32950 -140 33060 -120
rect 33120 -60 33230 -40
rect 33120 -120 33140 -60
rect 33210 -120 33230 -60
rect 33120 -140 33230 -120
rect 33290 -60 33400 -40
rect 33290 -120 33310 -60
rect 33380 -120 33400 -60
rect 33290 -140 33400 -120
rect 33460 -60 33570 -40
rect 33460 -120 33480 -60
rect 33550 -120 33570 -60
rect 33460 -140 33570 -120
rect 33630 -60 33740 -40
rect 33630 -120 33650 -60
rect 33720 -120 33740 -60
rect 33630 -140 33740 -120
rect 33800 -60 33910 -40
rect 33800 -120 33820 -60
rect 33890 -120 33910 -60
rect 33800 -140 33910 -120
rect 33970 -60 34080 -40
rect 33970 -120 33990 -60
rect 34060 -120 34080 -60
rect 33970 -140 34080 -120
rect 34140 -60 34250 -40
rect 34140 -120 34160 -60
rect 34230 -120 34250 -60
rect 34140 -140 34250 -120
rect 34310 -60 34420 -40
rect 34310 -120 34330 -60
rect 34400 -120 34420 -60
rect 34310 -140 34420 -120
rect 34480 -60 34590 -40
rect 34480 -120 34500 -60
rect 34570 -120 34590 -60
rect 34480 -140 34590 -120
rect 34650 -60 34760 -40
rect 34650 -120 34670 -60
rect 34740 -120 34760 -60
rect 34650 -140 34760 -120
rect 34820 -60 34930 -40
rect 34820 -120 34840 -60
rect 34910 -120 34930 -60
rect 34820 -140 34930 -120
rect 34990 -60 35100 -40
rect 34990 -120 35010 -60
rect 35080 -120 35100 -60
rect 34990 -140 35100 -120
rect 35160 -60 35270 -40
rect 35160 -120 35180 -60
rect 35250 -120 35270 -60
rect 35160 -140 35270 -120
rect 35330 -60 35440 -40
rect 35330 -120 35350 -60
rect 35420 -120 35440 -60
rect 35330 -140 35440 -120
rect 35500 -60 35610 -40
rect 35500 -120 35520 -60
rect 35590 -120 35610 -60
rect 35500 -140 35610 -120
rect 35670 -60 35780 -40
rect 35670 -120 35690 -60
rect 35760 -120 35780 -60
rect 35670 -140 35780 -120
rect 35840 -60 35950 -40
rect 35840 -120 35860 -60
rect 35930 -120 35950 -60
rect 35840 -140 35950 -120
rect 36010 -60 36120 -40
rect 36010 -120 36030 -60
rect 36100 -120 36120 -60
rect 36010 -140 36120 -120
rect 36180 -60 36290 -40
rect 36180 -120 36200 -60
rect 36270 -120 36290 -60
rect 36180 -140 36290 -120
rect 36350 -60 36460 -40
rect 36350 -120 36370 -60
rect 36440 -120 36460 -60
rect 36350 -140 36460 -120
rect 36520 -60 36630 -40
rect 36520 -120 36540 -60
rect 36610 -120 36630 -60
rect 36520 -140 36630 -120
rect 36690 -60 36800 -40
rect 36690 -120 36710 -60
rect 36780 -120 36800 -60
rect 36690 -140 36800 -120
rect 36860 -60 36970 -40
rect 36860 -120 36880 -60
rect 36950 -120 36970 -60
rect 36860 -140 36970 -120
rect 37030 -60 37140 -40
rect 37030 -120 37050 -60
rect 37120 -120 37140 -60
rect 37030 -140 37140 -120
rect 37200 -60 37310 -40
rect 37200 -120 37220 -60
rect 37290 -120 37310 -60
rect 37200 -140 37310 -120
rect 37370 -60 37480 -40
rect 37370 -120 37390 -60
rect 37460 -120 37480 -60
rect 37370 -140 37480 -120
rect 37540 -60 37650 -40
rect 37540 -120 37560 -60
rect 37630 -120 37650 -60
rect 37540 -140 37650 -120
rect 37710 -60 37820 -40
rect 37710 -120 37730 -60
rect 37800 -120 37820 -60
rect 37710 -140 37820 -120
rect 37880 -60 37990 -40
rect 37880 -120 37900 -60
rect 37970 -120 37990 -60
rect 37880 -140 37990 -120
rect 38050 -60 38160 -40
rect 38050 -120 38070 -60
rect 38140 -120 38160 -60
rect 38050 -140 38160 -120
rect 38220 -60 38330 -40
rect 38220 -120 38240 -60
rect 38310 -120 38330 -60
rect 38220 -140 38330 -120
rect 38390 -60 38500 -40
rect 38390 -120 38410 -60
rect 38480 -120 38500 -60
rect 38390 -140 38500 -120
rect 38560 -60 38670 -40
rect 38560 -120 38580 -60
rect 38650 -120 38670 -60
rect 38560 -140 38670 -120
rect 38730 -60 38840 -40
rect 38730 -120 38750 -60
rect 38820 -120 38840 -60
rect 38730 -140 38840 -120
rect 38900 -60 39010 -40
rect 38900 -120 38920 -60
rect 38990 -120 39010 -60
rect 38900 -140 39010 -120
rect 39070 -60 39180 -40
rect 39070 -120 39090 -60
rect 39160 -120 39180 -60
rect 39070 -140 39180 -120
rect 39240 -60 39350 -40
rect 39240 -120 39260 -60
rect 39330 -120 39350 -60
rect 39240 -140 39350 -120
rect 39410 -60 39520 -40
rect 39410 -120 39430 -60
rect 39500 -120 39520 -60
rect 39410 -140 39520 -120
rect 39580 -60 39690 -40
rect 39580 -120 39600 -60
rect 39670 -120 39690 -60
rect 39580 -140 39690 -120
rect 39750 -60 39860 -40
rect 39750 -120 39770 -60
rect 39840 -120 39860 -60
rect 39750 -140 39860 -120
rect 39920 -60 40030 -40
rect 39920 -120 39940 -60
rect 40010 -120 40030 -60
rect 39920 -140 40030 -120
rect 40090 -60 40200 -40
rect 40090 -120 40110 -60
rect 40180 -120 40200 -60
rect 40090 -140 40200 -120
rect 40260 -60 40370 -40
rect 40260 -120 40280 -60
rect 40350 -120 40370 -60
rect 40260 -140 40370 -120
rect 40430 -60 40540 -40
rect 40430 -120 40450 -60
rect 40520 -120 40540 -60
rect 40430 -140 40540 -120
rect 40600 -60 40710 -40
rect 40600 -120 40620 -60
rect 40690 -120 40710 -60
rect 40600 -140 40710 -120
rect 40770 -60 40880 -40
rect 40770 -120 40790 -60
rect 40860 -120 40880 -60
rect 40770 -140 40880 -120
rect 40940 -60 41050 -40
rect 40940 -120 40960 -60
rect 41030 -120 41050 -60
rect 40940 -140 41050 -120
rect 41110 -60 41220 -40
rect 41110 -120 41130 -60
rect 41200 -120 41220 -60
rect 41110 -140 41220 -120
rect 41280 -60 41390 -40
rect 41280 -120 41300 -60
rect 41370 -120 41390 -60
rect 41280 -140 41390 -120
rect 41450 -60 41560 -40
rect 41450 -120 41470 -60
rect 41540 -120 41560 -60
rect 41450 -140 41560 -120
rect 41620 -60 41730 -40
rect 41620 -120 41640 -60
rect 41710 -120 41730 -60
rect 41620 -140 41730 -120
rect 41790 -60 41900 -40
rect 41790 -120 41810 -60
rect 41880 -120 41900 -60
rect 41790 -140 41900 -120
rect 41960 -60 42070 -40
rect 41960 -120 41980 -60
rect 42050 -120 42070 -60
rect 41960 -140 42070 -120
rect 42130 -60 42240 -40
rect 42130 -120 42150 -60
rect 42220 -120 42240 -60
rect 42130 -140 42240 -120
rect 42300 -60 42410 -40
rect 42300 -120 42320 -60
rect 42390 -120 42410 -60
rect 42300 -140 42410 -120
rect 42470 -60 42580 -40
rect 42470 -120 42490 -60
rect 42560 -120 42580 -60
rect 42470 -140 42580 -120
rect 42640 -60 42750 -40
rect 42640 -120 42660 -60
rect 42730 -120 42750 -60
rect 42640 -140 42750 -120
rect 42810 -60 42920 -40
rect 42810 -120 42830 -60
rect 42900 -120 42920 -60
rect 42810 -140 42920 -120
rect 42980 -60 43090 -40
rect 42980 -120 43000 -60
rect 43070 -120 43090 -60
rect 42980 -140 43090 -120
rect 43150 -60 43260 -40
rect 43150 -120 43170 -60
rect 43240 -120 43260 -60
rect 43150 -140 43260 -120
rect 43320 -60 43430 -40
rect 43320 -120 43340 -60
rect 43410 -120 43430 -60
rect 43320 -140 43430 -120
rect 43490 -60 43600 -40
rect 43490 -120 43510 -60
rect 43580 -120 43600 -60
rect 43490 -140 43600 -120
rect 43660 -60 43770 -40
rect 43660 -120 43680 -60
rect 43750 -120 43770 -60
rect 43660 -140 43770 -120
rect 43830 -60 43940 -40
rect 43830 -120 43850 -60
rect 43920 -120 43940 -60
rect 43830 -140 43940 -120
rect 44000 -60 44110 -40
rect 44000 -120 44020 -60
rect 44090 -120 44110 -60
rect 44000 -140 44110 -120
rect 44170 -60 44280 -40
rect 44170 -120 44190 -60
rect 44260 -120 44280 -60
rect 44170 -140 44280 -120
rect 44340 -60 44450 -40
rect 44340 -120 44360 -60
rect 44430 -120 44450 -60
rect 44340 -140 44450 -120
rect 44510 -60 44620 -40
rect 44510 -120 44530 -60
rect 44600 -120 44620 -60
rect 44510 -140 44620 -120
rect 44680 -60 44790 -40
rect 44680 -120 44700 -60
rect 44770 -120 44790 -60
rect 44680 -140 44790 -120
rect 44850 -60 44960 -40
rect 44850 -120 44870 -60
rect 44940 -120 44960 -60
rect 44850 -140 44960 -120
rect 45020 -60 45130 -40
rect 45020 -120 45040 -60
rect 45110 -120 45130 -60
rect 45020 -140 45130 -120
rect 45190 -60 45300 -40
rect 45190 -120 45210 -60
rect 45280 -120 45300 -60
rect 45190 -140 45300 -120
rect 45360 -60 45470 -40
rect 45360 -120 45380 -60
rect 45450 -120 45470 -60
rect 45360 -140 45470 -120
rect 45530 -60 45640 -40
rect 45530 -120 45550 -60
rect 45620 -120 45640 -60
rect 45530 -140 45640 -120
rect 45700 -60 45810 -40
rect 45700 -120 45720 -60
rect 45790 -120 45810 -60
rect 45700 -140 45810 -120
rect 45870 -60 45980 -40
rect 45870 -120 45890 -60
rect 45960 -120 45980 -60
rect 45870 -140 45980 -120
rect 46040 -60 46150 -40
rect 46040 -120 46060 -60
rect 46130 -120 46150 -60
rect 46040 -140 46150 -120
rect 46210 -60 46320 -40
rect 46210 -120 46230 -60
rect 46300 -120 46320 -60
rect 46210 -140 46320 -120
rect 46380 -60 46490 -40
rect 46380 -120 46400 -60
rect 46470 -120 46490 -60
rect 46380 -140 46490 -120
rect 46550 -60 46660 -40
rect 46550 -120 46570 -60
rect 46640 -120 46660 -60
rect 46550 -140 46660 -120
rect 46720 -60 46830 -40
rect 46720 -120 46740 -60
rect 46810 -120 46830 -60
rect 46720 -140 46830 -120
rect 46890 -60 47000 -40
rect 46890 -120 46910 -60
rect 46980 -120 47000 -60
rect 46890 -140 47000 -120
rect 47060 -60 47170 -40
rect 47060 -120 47080 -60
rect 47150 -120 47170 -60
rect 47060 -140 47170 -120
rect 47230 -60 47340 -40
rect 47230 -120 47250 -60
rect 47320 -120 47340 -60
rect 47230 -140 47340 -120
rect 47400 -60 47510 -40
rect 47400 -120 47420 -60
rect 47490 -120 47510 -60
rect 47400 -140 47510 -120
rect 47570 -60 47680 -40
rect 47570 -120 47590 -60
rect 47660 -120 47680 -60
rect 47570 -140 47680 -120
rect 47740 -60 47850 -40
rect 47740 -120 47760 -60
rect 47830 -120 47850 -60
rect 47740 -140 47850 -120
rect 47910 -60 48020 -40
rect 47910 -120 47930 -60
rect 48000 -120 48020 -60
rect 47910 -140 48020 -120
rect 48080 -60 48190 -40
rect 48080 -120 48100 -60
rect 48170 -120 48190 -60
rect 48080 -140 48190 -120
rect 48250 -60 48360 -40
rect 48250 -120 48270 -60
rect 48340 -120 48360 -60
rect 48250 -140 48360 -120
rect 48420 -60 48530 -40
rect 48420 -120 48440 -60
rect 48510 -120 48530 -60
rect 48420 -140 48530 -120
rect 48590 -60 48700 -40
rect 48590 -120 48610 -60
rect 48680 -120 48700 -60
rect 48590 -140 48700 -120
rect 48760 -60 48870 -40
rect 48760 -120 48780 -60
rect 48850 -120 48870 -60
rect 48760 -140 48870 -120
rect 48930 -60 49040 -40
rect 48930 -120 48950 -60
rect 49020 -120 49040 -60
rect 48930 -140 49040 -120
rect 49100 -60 49210 -40
rect 49100 -120 49120 -60
rect 49190 -120 49210 -60
rect 49100 -140 49210 -120
rect 49270 -60 49380 -40
rect 49270 -120 49290 -60
rect 49360 -120 49380 -60
rect 49270 -140 49380 -120
rect 49440 -60 49550 -40
rect 49440 -120 49460 -60
rect 49530 -120 49550 -60
rect 49440 -140 49550 -120
rect 49610 -60 49720 -40
rect 49610 -120 49630 -60
rect 49700 -120 49720 -60
rect 49610 -140 49720 -120
rect 49780 -60 49890 -40
rect 49780 -120 49800 -60
rect 49870 -120 49890 -60
rect 49780 -140 49890 -120
rect 49950 -60 50060 -40
rect 49950 -120 49970 -60
rect 50040 -120 50060 -60
rect 49950 -140 50060 -120
rect 50120 -60 50230 -40
rect 50120 -120 50140 -60
rect 50210 -120 50230 -60
rect 50120 -140 50230 -120
rect 50290 -60 50400 -40
rect 50290 -120 50310 -60
rect 50380 -120 50400 -60
rect 50290 -140 50400 -120
rect 50460 -60 50570 -40
rect 50460 -120 50480 -60
rect 50550 -120 50570 -60
rect 50460 -140 50570 -120
rect 50630 -60 50740 -40
rect 50630 -120 50650 -60
rect 50720 -120 50740 -60
rect 50630 -140 50740 -120
rect 50800 -60 50910 -40
rect 50800 -120 50820 -60
rect 50890 -120 50910 -60
rect 50800 -140 50910 -120
rect 50970 -60 51080 -40
rect 50970 -120 50990 -60
rect 51060 -120 51080 -60
rect 50970 -140 51080 -120
rect 51140 -60 51250 -40
rect 51140 -120 51160 -60
rect 51230 -120 51250 -60
rect 51140 -140 51250 -120
rect 51310 -60 51420 -40
rect 51310 -120 51330 -60
rect 51400 -120 51420 -60
rect 51310 -140 51420 -120
rect 51480 -60 51590 -40
rect 51480 -120 51500 -60
rect 51570 -120 51590 -60
rect 51480 -140 51590 -120
rect 51650 -60 51760 -40
rect 51650 -120 51670 -60
rect 51740 -120 51760 -60
rect 51650 -140 51760 -120
rect 51820 -60 51930 -40
rect 51820 -120 51840 -60
rect 51910 -120 51930 -60
rect 51820 -140 51930 -120
rect 51990 -60 52100 -40
rect 51990 -120 52010 -60
rect 52080 -120 52100 -60
rect 51990 -140 52100 -120
rect 52160 -60 52270 -40
rect 52160 -120 52180 -60
rect 52250 -120 52270 -60
rect 52160 -140 52270 -120
rect 52330 -60 52440 -40
rect 52330 -120 52350 -60
rect 52420 -120 52440 -60
rect 52330 -140 52440 -120
rect 52500 -60 52610 -40
rect 52500 -120 52520 -60
rect 52590 -120 52610 -60
rect 52500 -140 52610 -120
rect 52670 -60 52780 -40
rect 52670 -120 52690 -60
rect 52760 -120 52780 -60
rect 52670 -140 52780 -120
rect 52840 -60 52950 -40
rect 52840 -120 52860 -60
rect 52930 -120 52950 -60
rect 52840 -140 52950 -120
rect 53010 -60 53120 -40
rect 53010 -120 53030 -60
rect 53100 -120 53120 -60
rect 53010 -140 53120 -120
rect 53180 -60 53290 -40
rect 53180 -120 53200 -60
rect 53270 -120 53290 -60
rect 53180 -140 53290 -120
rect 53350 -60 53460 -40
rect 53350 -120 53370 -60
rect 53440 -120 53460 -60
rect 53350 -140 53460 -120
rect 53520 -60 53630 -40
rect 53520 -120 53540 -60
rect 53610 -120 53630 -60
rect 53520 -140 53630 -120
rect 53690 -60 53800 -40
rect 53690 -120 53710 -60
rect 53780 -120 53800 -60
rect 53690 -140 53800 -120
rect 53860 -60 53970 -40
rect 53860 -120 53880 -60
rect 53950 -120 53970 -60
rect 53860 -140 53970 -120
rect 54030 -60 54140 -40
rect 54030 -120 54050 -60
rect 54120 -120 54140 -60
rect 54030 -140 54140 -120
rect 54200 -60 54310 -40
rect 54200 -120 54220 -60
rect 54290 -120 54310 -60
rect 54200 -140 54310 -120
rect 54370 -60 54480 -40
rect 54370 -120 54390 -60
rect 54460 -120 54480 -60
rect 54370 -140 54480 -120
rect 54540 -60 54650 -40
rect 54540 -120 54560 -60
rect 54630 -120 54650 -60
rect 54540 -140 54650 -120
rect 54710 -60 54820 -40
rect 54710 -120 54730 -60
rect 54800 -120 54820 -60
rect 54710 -140 54820 -120
rect 54880 -60 54990 -40
rect 54880 -120 54900 -60
rect 54970 -120 54990 -60
rect 54880 -140 54990 -120
rect 55050 -60 55160 -40
rect 55050 -120 55070 -60
rect 55140 -120 55160 -60
rect 55050 -140 55160 -120
rect 55220 -60 55330 -40
rect 55220 -120 55240 -60
rect 55310 -120 55330 -60
rect 55220 -140 55330 -120
rect 55390 -60 55500 -40
rect 55390 -120 55410 -60
rect 55480 -120 55500 -60
rect 55390 -140 55500 -120
rect 55560 -60 55670 -40
rect 55560 -120 55580 -60
rect 55650 -120 55670 -60
rect 55560 -140 55670 -120
rect 55730 -60 55840 -40
rect 55730 -120 55750 -60
rect 55820 -120 55840 -60
rect 55730 -140 55840 -120
rect 55900 -60 56010 -40
rect 55900 -120 55920 -60
rect 55990 -120 56010 -60
rect 55900 -140 56010 -120
rect 56070 -60 56180 -40
rect 56070 -120 56090 -60
rect 56160 -120 56180 -60
rect 56070 -140 56180 -120
rect 56240 -60 56350 -40
rect 56240 -120 56260 -60
rect 56330 -120 56350 -60
rect 56240 -140 56350 -120
rect 56410 -60 56520 -40
rect 56410 -120 56430 -60
rect 56500 -120 56520 -60
rect 56410 -140 56520 -120
rect 56580 -60 56690 -40
rect 56580 -120 56600 -60
rect 56670 -120 56690 -60
rect 56580 -140 56690 -120
rect 56750 -60 56860 -40
rect 56750 -120 56770 -60
rect 56840 -120 56860 -60
rect 56750 -140 56860 -120
rect 56920 -60 57030 -40
rect 56920 -120 56940 -60
rect 57010 -120 57030 -60
rect 56920 -140 57030 -120
rect 57090 -60 57200 -40
rect 57090 -120 57110 -60
rect 57180 -120 57200 -60
rect 57090 -140 57200 -120
rect 57260 -60 57370 -40
rect 57260 -120 57280 -60
rect 57350 -120 57370 -60
rect 57260 -140 57370 -120
rect 57430 -60 57540 -40
rect 57430 -120 57450 -60
rect 57520 -120 57540 -60
rect 57430 -140 57540 -120
rect 57600 -60 57710 -40
rect 57600 -120 57620 -60
rect 57690 -120 57710 -60
rect 57600 -140 57710 -120
rect 57770 -60 57880 -40
rect 57770 -120 57790 -60
rect 57860 -120 57880 -60
rect 57770 -140 57880 -120
rect 57940 -60 58050 -40
rect 57940 -120 57960 -60
rect 58030 -120 58050 -60
rect 57940 -140 58050 -120
rect 58110 -60 58220 -40
rect 58110 -120 58130 -60
rect 58200 -120 58220 -60
rect 58110 -140 58220 -120
rect 58280 -60 58390 -40
rect 58280 -120 58300 -60
rect 58370 -120 58390 -60
rect 58280 -140 58390 -120
rect 58450 -60 58560 -40
rect 58450 -120 58470 -60
rect 58540 -120 58560 -60
rect 58450 -140 58560 -120
rect 58620 -60 58730 -40
rect 58620 -120 58640 -60
rect 58710 -120 58730 -60
rect 58620 -140 58730 -120
rect 58790 -60 58900 -40
rect 58790 -120 58810 -60
rect 58880 -120 58900 -60
rect 58790 -140 58900 -120
rect 58960 -60 59070 -40
rect 58960 -120 58980 -60
rect 59050 -120 59070 -60
rect 58960 -140 59070 -120
rect 59130 -60 59240 -40
rect 59130 -120 59150 -60
rect 59220 -120 59240 -60
rect 59130 -140 59240 -120
rect 2070 -260 2400 -240
rect 2070 -390 2120 -260
rect 2350 -390 2400 -260
rect 2070 -410 2400 -390
rect 5088 -268 5418 -248
rect 5088 -398 5138 -268
rect 5368 -398 5418 -268
rect 5088 -418 5418 -398
rect 7574 -268 7904 -248
rect 7574 -398 7624 -268
rect 7854 -398 7904 -268
rect 7574 -418 7904 -398
rect 8994 -268 9324 -248
rect 8994 -398 9044 -268
rect 9274 -398 9324 -268
rect 8994 -418 9324 -398
rect 13618 -264 13948 -244
rect 13618 -394 13668 -264
rect 13898 -394 13948 -264
rect 13618 -414 13948 -394
rect 16818 -264 17148 -244
rect 16818 -394 16868 -264
rect 17098 -394 17148 -264
rect 16818 -414 17148 -394
rect 20374 -264 20704 -244
rect 20374 -394 20424 -264
rect 20654 -394 20704 -264
rect 20374 -414 20704 -394
rect 25708 -264 26038 -244
rect 25708 -394 25758 -264
rect 25988 -394 26038 -264
rect 25708 -414 26038 -394
rect 28552 -264 28882 -244
rect 28552 -394 28602 -264
rect 28832 -394 28882 -264
rect 28552 -414 28882 -394
rect 32464 -264 32794 -244
rect 32464 -394 32514 -264
rect 32744 -394 32794 -264
rect 32464 -414 32794 -394
rect 34620 -264 34950 -244
rect 34620 -394 34670 -264
rect 34900 -394 34950 -264
rect 34620 -414 34950 -394
rect 37442 -264 37772 -244
rect 37442 -394 37492 -264
rect 37722 -394 37772 -264
rect 37442 -414 37772 -394
rect 40642 -264 40972 -244
rect 40642 -394 40692 -264
rect 40922 -394 40972 -264
rect 40642 -414 40972 -394
rect 45618 -264 45948 -244
rect 45618 -394 45668 -264
rect 45898 -394 45948 -264
rect 45618 -414 45948 -394
rect 48818 -264 49148 -244
rect 48818 -394 48868 -264
rect 49098 -394 49148 -264
rect 48818 -414 49148 -394
rect 50952 -264 51282 -244
rect 50952 -394 51002 -264
rect 51232 -394 51282 -264
rect 50952 -414 51282 -394
rect 54508 -264 54838 -244
rect 54508 -394 54558 -264
rect 54788 -394 54838 -264
rect 54508 -414 54838 -394
rect 57352 -264 57682 -244
rect 57352 -394 57402 -264
rect 57632 -394 57682 -264
rect 57352 -414 57682 -394
rect 61264 -264 61594 -244
rect 61264 -394 61314 -264
rect 61544 -394 61594 -264
rect 61264 -414 61594 -394
rect 64108 -264 64438 -244
rect 64108 -394 64158 -264
rect 64388 -394 64438 -264
rect 64108 -414 64438 -394
rect 67664 -264 67994 -244
rect 67664 -394 67714 -264
rect 67944 -394 67994 -264
rect 67664 -414 67994 -394
rect 70508 -264 70838 -244
rect 70508 -394 70558 -264
rect 70788 -394 70838 -264
rect 70508 -414 70838 -394
rect 74418 -264 74748 -244
rect 74418 -394 74468 -264
rect 74698 -394 74748 -264
rect 74418 -414 74748 -394
rect 78330 -264 78660 -244
rect 78330 -394 78380 -264
rect 78610 -394 78660 -264
rect 78330 -414 78660 -394
rect 82242 -264 82572 -244
rect 82242 -394 82292 -264
rect 82522 -394 82572 -264
rect 82242 -414 82572 -394
rect 86152 -264 86482 -244
rect 86152 -394 86202 -264
rect 86432 -394 86482 -264
rect 86152 -414 86482 -394
rect 210 -530 320 -510
rect 210 -590 230 -530
rect 300 -590 320 -530
rect 210 -610 320 -590
rect 380 -530 490 -510
rect 380 -590 400 -530
rect 470 -590 490 -530
rect 380 -610 490 -590
rect 550 -530 660 -510
rect 550 -590 570 -530
rect 640 -590 660 -530
rect 550 -610 660 -590
rect 720 -530 830 -510
rect 720 -590 740 -530
rect 810 -590 830 -530
rect 720 -610 830 -590
rect 890 -530 1000 -510
rect 890 -590 910 -530
rect 980 -590 1000 -530
rect 890 -610 1000 -590
rect 1060 -530 1170 -510
rect 1060 -590 1080 -530
rect 1150 -590 1170 -530
rect 1060 -610 1170 -590
rect 1230 -530 1340 -510
rect 1230 -590 1250 -530
rect 1320 -590 1340 -530
rect 1230 -610 1340 -590
rect 1400 -530 1510 -510
rect 1400 -590 1420 -530
rect 1490 -590 1510 -530
rect 1400 -610 1510 -590
rect 1570 -530 1680 -510
rect 1570 -590 1590 -530
rect 1660 -590 1680 -530
rect 1570 -610 1680 -590
rect 1740 -530 1850 -510
rect 1740 -590 1760 -530
rect 1830 -590 1850 -530
rect 1740 -610 1850 -590
rect 1910 -530 2020 -510
rect 1910 -590 1930 -530
rect 2000 -590 2020 -530
rect 1910 -610 2020 -590
rect 2080 -530 2190 -510
rect 2080 -590 2100 -530
rect 2170 -590 2190 -530
rect 2080 -610 2190 -590
rect 2250 -530 2360 -510
rect 2250 -590 2270 -530
rect 2340 -590 2360 -530
rect 2250 -610 2360 -590
rect 2420 -530 2530 -510
rect 2420 -590 2440 -530
rect 2510 -590 2530 -530
rect 2420 -610 2530 -590
rect 2590 -530 2700 -510
rect 2590 -590 2610 -530
rect 2680 -590 2700 -530
rect 2590 -610 2700 -590
rect 2760 -530 2870 -510
rect 2760 -590 2780 -530
rect 2850 -590 2870 -530
rect 2760 -610 2870 -590
rect 2930 -530 3040 -510
rect 2930 -590 2950 -530
rect 3020 -590 3040 -530
rect 2930 -610 3040 -590
rect 3100 -530 3210 -510
rect 3100 -590 3120 -530
rect 3190 -590 3210 -530
rect 3100 -610 3210 -590
rect 3270 -530 3380 -510
rect 3270 -590 3290 -530
rect 3360 -590 3380 -530
rect 3270 -610 3380 -590
rect 3440 -530 3550 -510
rect 3440 -590 3460 -530
rect 3530 -590 3550 -530
rect 3440 -610 3550 -590
rect 3610 -530 3720 -510
rect 3610 -590 3630 -530
rect 3700 -590 3720 -530
rect 3610 -610 3720 -590
rect 3780 -530 3890 -510
rect 3780 -590 3800 -530
rect 3870 -590 3890 -530
rect 3780 -610 3890 -590
rect 3950 -530 4060 -510
rect 3950 -590 3970 -530
rect 4040 -590 4060 -530
rect 3950 -610 4060 -590
rect 4120 -530 4230 -510
rect 4120 -590 4140 -530
rect 4210 -590 4230 -530
rect 4120 -610 4230 -590
rect 4290 -530 4400 -510
rect 4290 -590 4310 -530
rect 4380 -590 4400 -530
rect 4290 -610 4400 -590
rect 4460 -530 4570 -510
rect 4460 -590 4480 -530
rect 4550 -590 4570 -530
rect 4460 -610 4570 -590
rect 4630 -530 4740 -510
rect 4630 -590 4650 -530
rect 4720 -590 4740 -530
rect 4630 -610 4740 -590
rect 4800 -530 4910 -510
rect 4800 -590 4820 -530
rect 4890 -590 4910 -530
rect 4800 -610 4910 -590
rect 4970 -530 5080 -510
rect 4970 -590 4990 -530
rect 5060 -590 5080 -530
rect 4970 -610 5080 -590
rect 5140 -530 5250 -510
rect 5140 -590 5160 -530
rect 5230 -590 5250 -530
rect 5140 -610 5250 -590
rect 5310 -530 5420 -510
rect 5310 -590 5330 -530
rect 5400 -590 5420 -530
rect 5310 -610 5420 -590
rect 5480 -530 5590 -510
rect 5480 -590 5500 -530
rect 5570 -590 5590 -530
rect 5480 -610 5590 -590
rect 5650 -530 5760 -510
rect 5650 -590 5670 -530
rect 5740 -590 5760 -530
rect 5650 -610 5760 -590
rect 5820 -530 5930 -510
rect 5820 -590 5840 -530
rect 5910 -590 5930 -530
rect 5820 -610 5930 -590
rect 5990 -530 6100 -510
rect 5990 -590 6010 -530
rect 6080 -590 6100 -530
rect 5990 -610 6100 -590
rect 6160 -530 6270 -510
rect 6160 -590 6180 -530
rect 6250 -590 6270 -530
rect 6160 -610 6270 -590
rect 6330 -530 6440 -510
rect 6330 -590 6350 -530
rect 6420 -590 6440 -530
rect 6330 -610 6440 -590
rect 6500 -530 6610 -510
rect 6500 -590 6520 -530
rect 6590 -590 6610 -530
rect 6500 -610 6610 -590
rect 6670 -530 6780 -510
rect 6670 -590 6690 -530
rect 6760 -590 6780 -530
rect 6670 -610 6780 -590
rect 6840 -530 6950 -510
rect 6840 -590 6860 -530
rect 6930 -590 6950 -530
rect 6840 -610 6950 -590
rect 7010 -530 7120 -510
rect 7010 -590 7030 -530
rect 7100 -590 7120 -530
rect 7010 -610 7120 -590
rect 7180 -530 7290 -510
rect 7180 -590 7200 -530
rect 7270 -590 7290 -530
rect 7180 -610 7290 -590
rect 7350 -530 7460 -510
rect 7350 -590 7370 -530
rect 7440 -590 7460 -530
rect 7350 -610 7460 -590
rect 7520 -530 7630 -510
rect 7520 -590 7540 -530
rect 7610 -590 7630 -530
rect 7520 -610 7630 -590
rect 7690 -530 7800 -510
rect 7690 -590 7710 -530
rect 7780 -590 7800 -530
rect 7690 -610 7800 -590
rect 7860 -530 7970 -510
rect 7860 -590 7880 -530
rect 7950 -590 7970 -530
rect 7860 -610 7970 -590
rect 8030 -530 8140 -510
rect 8030 -590 8050 -530
rect 8120 -590 8140 -530
rect 8030 -610 8140 -590
rect 8200 -530 8310 -510
rect 8200 -590 8220 -530
rect 8290 -590 8310 -530
rect 8200 -610 8310 -590
rect 8370 -530 8480 -510
rect 8370 -590 8390 -530
rect 8460 -590 8480 -530
rect 8370 -610 8480 -590
rect 8540 -530 8650 -510
rect 8540 -590 8560 -530
rect 8630 -590 8650 -530
rect 8540 -610 8650 -590
rect 8710 -530 8820 -510
rect 8710 -590 8730 -530
rect 8800 -590 8820 -530
rect 8710 -610 8820 -590
rect 8880 -530 8990 -510
rect 8880 -590 8900 -530
rect 8970 -590 8990 -530
rect 8880 -610 8990 -590
rect 9050 -530 9160 -510
rect 9050 -590 9070 -530
rect 9140 -590 9160 -530
rect 9050 -610 9160 -590
rect 9220 -530 9330 -510
rect 9220 -590 9240 -530
rect 9310 -590 9330 -530
rect 9220 -610 9330 -590
rect 9390 -530 9500 -510
rect 9390 -590 9410 -530
rect 9480 -590 9500 -530
rect 9390 -610 9500 -590
rect 9560 -530 9670 -510
rect 9560 -590 9580 -530
rect 9650 -590 9670 -530
rect 9560 -610 9670 -590
rect 9730 -530 9840 -510
rect 9730 -590 9750 -530
rect 9820 -590 9840 -530
rect 9730 -610 9840 -590
rect 9900 -530 10010 -510
rect 9900 -590 9920 -530
rect 9990 -590 10010 -530
rect 9900 -610 10010 -590
rect 10070 -530 10180 -510
rect 10070 -590 10090 -530
rect 10160 -590 10180 -530
rect 10070 -610 10180 -590
rect 10240 -530 10350 -510
rect 10240 -590 10260 -530
rect 10330 -590 10350 -530
rect 10240 -610 10350 -590
rect 10410 -530 10520 -510
rect 10410 -590 10430 -530
rect 10500 -590 10520 -530
rect 10410 -610 10520 -590
rect 10580 -530 10690 -510
rect 10580 -590 10600 -530
rect 10670 -590 10690 -530
rect 10580 -610 10690 -590
rect 10750 -530 10860 -510
rect 10750 -590 10770 -530
rect 10840 -590 10860 -530
rect 10750 -610 10860 -590
rect 10920 -530 11030 -510
rect 10920 -590 10940 -530
rect 11010 -590 11030 -530
rect 10920 -610 11030 -590
rect 11090 -530 11200 -510
rect 11090 -590 11110 -530
rect 11180 -590 11200 -530
rect 11090 -610 11200 -590
rect 11260 -530 11370 -510
rect 11260 -590 11280 -530
rect 11350 -590 11370 -530
rect 11260 -610 11370 -590
rect 11430 -530 11540 -510
rect 11430 -590 11450 -530
rect 11520 -590 11540 -530
rect 11430 -610 11540 -590
rect 11600 -530 11710 -510
rect 11600 -590 11620 -530
rect 11690 -590 11710 -530
rect 11600 -610 11710 -590
rect 11770 -530 11880 -510
rect 11770 -590 11790 -530
rect 11860 -590 11880 -530
rect 11770 -610 11880 -590
rect 11940 -530 12050 -510
rect 11940 -590 11960 -530
rect 12030 -590 12050 -530
rect 11940 -610 12050 -590
rect 12110 -530 12220 -510
rect 12110 -590 12130 -530
rect 12200 -590 12220 -530
rect 12110 -610 12220 -590
rect 12280 -530 12390 -510
rect 12280 -590 12300 -530
rect 12370 -590 12390 -530
rect 12280 -610 12390 -590
rect 12450 -530 12560 -510
rect 12450 -590 12470 -530
rect 12540 -590 12560 -530
rect 12450 -610 12560 -590
rect 12620 -530 12730 -510
rect 12620 -590 12640 -530
rect 12710 -590 12730 -530
rect 12620 -610 12730 -590
rect 12790 -530 12900 -510
rect 12790 -590 12810 -530
rect 12880 -590 12900 -530
rect 12790 -610 12900 -590
rect 12960 -530 13070 -510
rect 12960 -590 12980 -530
rect 13050 -590 13070 -530
rect 12960 -610 13070 -590
rect 13130 -530 13240 -510
rect 13130 -590 13150 -530
rect 13220 -590 13240 -530
rect 13130 -610 13240 -590
rect 13300 -530 13410 -510
rect 13300 -590 13320 -530
rect 13390 -590 13410 -530
rect 13300 -610 13410 -590
rect 13470 -530 13580 -510
rect 13470 -590 13490 -530
rect 13560 -590 13580 -530
rect 13470 -610 13580 -590
rect 13640 -530 13750 -510
rect 13640 -590 13660 -530
rect 13730 -590 13750 -530
rect 13640 -610 13750 -590
rect 13810 -530 13920 -510
rect 13810 -590 13830 -530
rect 13900 -590 13920 -530
rect 13810 -610 13920 -590
rect 13980 -530 14090 -510
rect 13980 -590 14000 -530
rect 14070 -590 14090 -530
rect 13980 -610 14090 -590
rect 14150 -530 14260 -510
rect 14150 -590 14170 -530
rect 14240 -590 14260 -530
rect 14150 -610 14260 -590
rect 14320 -530 14430 -510
rect 14320 -590 14340 -530
rect 14410 -590 14430 -530
rect 14320 -610 14430 -590
rect 14490 -530 14600 -510
rect 14490 -590 14510 -530
rect 14580 -590 14600 -530
rect 14490 -610 14600 -590
rect 14660 -530 14770 -510
rect 14660 -590 14680 -530
rect 14750 -590 14770 -530
rect 14660 -610 14770 -590
rect 14830 -530 14940 -510
rect 14830 -590 14850 -530
rect 14920 -590 14940 -530
rect 14830 -610 14940 -590
rect 15000 -530 15110 -510
rect 15000 -590 15020 -530
rect 15090 -590 15110 -530
rect 15000 -610 15110 -590
rect 15170 -530 15280 -510
rect 15170 -590 15190 -530
rect 15260 -590 15280 -530
rect 15170 -610 15280 -590
rect 15340 -530 15450 -510
rect 15340 -590 15360 -530
rect 15430 -590 15450 -530
rect 15340 -610 15450 -590
rect 15510 -530 15620 -510
rect 15510 -590 15530 -530
rect 15600 -590 15620 -530
rect 15510 -610 15620 -590
rect 15680 -530 15790 -510
rect 15680 -590 15700 -530
rect 15770 -590 15790 -530
rect 15680 -610 15790 -590
rect 15850 -530 15960 -510
rect 15850 -590 15870 -530
rect 15940 -590 15960 -530
rect 15850 -610 15960 -590
rect 16020 -530 16130 -510
rect 16020 -590 16040 -530
rect 16110 -590 16130 -530
rect 16020 -610 16130 -590
rect 16190 -530 16300 -510
rect 16190 -590 16210 -530
rect 16280 -590 16300 -530
rect 16190 -610 16300 -590
rect 16360 -530 16470 -510
rect 16360 -590 16380 -530
rect 16450 -590 16470 -530
rect 16360 -610 16470 -590
rect 16530 -530 16640 -510
rect 16530 -590 16550 -530
rect 16620 -590 16640 -530
rect 16530 -610 16640 -590
rect 16700 -530 16810 -510
rect 16700 -590 16720 -530
rect 16790 -590 16810 -530
rect 16700 -610 16810 -590
rect 16870 -530 16980 -510
rect 16870 -590 16890 -530
rect 16960 -590 16980 -530
rect 16870 -610 16980 -590
rect 17040 -530 17150 -510
rect 17040 -590 17060 -530
rect 17130 -590 17150 -530
rect 17040 -610 17150 -590
rect 17210 -530 17320 -510
rect 17210 -590 17230 -530
rect 17300 -590 17320 -530
rect 17210 -610 17320 -590
rect 17380 -530 17490 -510
rect 17380 -590 17400 -530
rect 17470 -590 17490 -530
rect 17380 -610 17490 -590
rect 17550 -530 17660 -510
rect 17550 -590 17570 -530
rect 17640 -590 17660 -530
rect 17550 -610 17660 -590
rect 17720 -530 17830 -510
rect 17720 -590 17740 -530
rect 17810 -590 17830 -530
rect 17720 -610 17830 -590
rect 17890 -530 18000 -510
rect 17890 -590 17910 -530
rect 17980 -590 18000 -530
rect 17890 -610 18000 -590
rect 18060 -530 18170 -510
rect 18060 -590 18080 -530
rect 18150 -590 18170 -530
rect 18060 -610 18170 -590
rect 18230 -530 18340 -510
rect 18230 -590 18250 -530
rect 18320 -590 18340 -530
rect 18230 -610 18340 -590
rect 18400 -530 18510 -510
rect 18400 -590 18420 -530
rect 18490 -590 18510 -530
rect 18400 -610 18510 -590
rect 18570 -530 18680 -510
rect 18570 -590 18590 -530
rect 18660 -590 18680 -530
rect 18570 -610 18680 -590
rect 18740 -530 18850 -510
rect 18740 -590 18760 -530
rect 18830 -590 18850 -530
rect 18740 -610 18850 -590
rect 18910 -530 19020 -510
rect 18910 -590 18930 -530
rect 19000 -590 19020 -530
rect 18910 -610 19020 -590
rect 19080 -530 19190 -510
rect 19080 -590 19100 -530
rect 19170 -590 19190 -530
rect 19080 -610 19190 -590
rect 19250 -530 19360 -510
rect 19250 -590 19270 -530
rect 19340 -590 19360 -530
rect 19250 -610 19360 -590
rect 19420 -530 19530 -510
rect 19420 -590 19440 -530
rect 19510 -590 19530 -530
rect 19420 -610 19530 -590
rect 19590 -530 19700 -510
rect 19590 -590 19610 -530
rect 19680 -590 19700 -530
rect 19590 -610 19700 -590
rect 19760 -530 19870 -510
rect 19760 -590 19780 -530
rect 19850 -590 19870 -530
rect 19760 -610 19870 -590
rect 19930 -530 20040 -510
rect 19930 -590 19950 -530
rect 20020 -590 20040 -530
rect 19930 -610 20040 -590
rect 20100 -530 20210 -510
rect 20100 -590 20120 -530
rect 20190 -590 20210 -530
rect 20100 -610 20210 -590
rect 20270 -530 20380 -510
rect 20270 -590 20290 -530
rect 20360 -590 20380 -530
rect 20270 -610 20380 -590
rect 20440 -530 20550 -510
rect 20440 -590 20460 -530
rect 20530 -590 20550 -530
rect 20440 -610 20550 -590
rect 20610 -530 20720 -510
rect 20610 -590 20630 -530
rect 20700 -590 20720 -530
rect 20610 -610 20720 -590
rect 20780 -530 20890 -510
rect 20780 -590 20800 -530
rect 20870 -590 20890 -530
rect 20780 -610 20890 -590
rect 20950 -530 21060 -510
rect 20950 -590 20970 -530
rect 21040 -590 21060 -530
rect 20950 -610 21060 -590
rect 21120 -530 21230 -510
rect 21120 -590 21140 -530
rect 21210 -590 21230 -530
rect 21120 -610 21230 -590
rect 21290 -530 21400 -510
rect 21290 -590 21310 -530
rect 21380 -590 21400 -530
rect 21290 -610 21400 -590
rect 21460 -530 21570 -510
rect 21460 -590 21480 -530
rect 21550 -590 21570 -530
rect 21460 -610 21570 -590
rect 21630 -530 21740 -510
rect 21630 -590 21650 -530
rect 21720 -590 21740 -530
rect 21630 -610 21740 -590
rect 21800 -530 21910 -510
rect 21800 -590 21820 -530
rect 21890 -590 21910 -530
rect 21800 -610 21910 -590
rect 21970 -530 22080 -510
rect 21970 -590 21990 -530
rect 22060 -590 22080 -530
rect 21970 -610 22080 -590
rect 22140 -530 22250 -510
rect 22140 -590 22160 -530
rect 22230 -590 22250 -530
rect 22140 -610 22250 -590
rect 22310 -530 22420 -510
rect 22310 -590 22330 -530
rect 22400 -590 22420 -530
rect 22310 -610 22420 -590
rect 22480 -530 22590 -510
rect 22480 -590 22500 -530
rect 22570 -590 22590 -530
rect 22480 -610 22590 -590
rect 22650 -530 22760 -510
rect 22650 -590 22670 -530
rect 22740 -590 22760 -530
rect 22650 -610 22760 -590
rect 22820 -530 22930 -510
rect 22820 -590 22840 -530
rect 22910 -590 22930 -530
rect 22820 -610 22930 -590
rect 22990 -530 23100 -510
rect 22990 -590 23010 -530
rect 23080 -590 23100 -530
rect 22990 -610 23100 -590
rect 23160 -530 23270 -510
rect 23160 -590 23180 -530
rect 23250 -590 23270 -530
rect 23160 -610 23270 -590
rect 23330 -530 23440 -510
rect 23330 -590 23350 -530
rect 23420 -590 23440 -530
rect 23330 -610 23440 -590
rect 23500 -530 23610 -510
rect 23500 -590 23520 -530
rect 23590 -590 23610 -530
rect 23500 -610 23610 -590
rect 23670 -530 23780 -510
rect 23670 -590 23690 -530
rect 23760 -590 23780 -530
rect 23670 -610 23780 -590
rect 23840 -530 23950 -510
rect 23840 -590 23860 -530
rect 23930 -590 23950 -530
rect 23840 -610 23950 -590
rect 24010 -530 24120 -510
rect 24010 -590 24030 -530
rect 24100 -590 24120 -530
rect 24010 -610 24120 -590
rect 24180 -530 24290 -510
rect 24180 -590 24200 -530
rect 24270 -590 24290 -530
rect 24180 -610 24290 -590
rect 24350 -530 24460 -510
rect 24350 -590 24370 -530
rect 24440 -590 24460 -530
rect 24350 -610 24460 -590
rect 24520 -530 24630 -510
rect 24520 -590 24540 -530
rect 24610 -590 24630 -530
rect 24520 -610 24630 -590
rect 24690 -530 24800 -510
rect 24690 -590 24710 -530
rect 24780 -590 24800 -530
rect 24690 -610 24800 -590
rect 24860 -530 24970 -510
rect 24860 -590 24880 -530
rect 24950 -590 24970 -530
rect 24860 -610 24970 -590
rect 25030 -530 25140 -510
rect 25030 -590 25050 -530
rect 25120 -590 25140 -530
rect 25030 -610 25140 -590
rect 25200 -530 25310 -510
rect 25200 -590 25220 -530
rect 25290 -590 25310 -530
rect 25200 -610 25310 -590
rect 25370 -530 25480 -510
rect 25370 -590 25390 -530
rect 25460 -590 25480 -530
rect 25370 -610 25480 -590
rect 25540 -530 25650 -510
rect 25540 -590 25560 -530
rect 25630 -590 25650 -530
rect 25540 -610 25650 -590
rect 25710 -530 25820 -510
rect 25710 -590 25730 -530
rect 25800 -590 25820 -530
rect 25710 -610 25820 -590
rect 25880 -530 25990 -510
rect 25880 -590 25900 -530
rect 25970 -590 25990 -530
rect 25880 -610 25990 -590
rect 26050 -530 26160 -510
rect 26050 -590 26070 -530
rect 26140 -590 26160 -530
rect 26050 -610 26160 -590
rect 26220 -530 26330 -510
rect 26220 -590 26240 -530
rect 26310 -590 26330 -530
rect 26220 -610 26330 -590
rect 26390 -530 26500 -510
rect 26390 -590 26410 -530
rect 26480 -590 26500 -530
rect 26390 -610 26500 -590
rect 26560 -530 26670 -510
rect 26560 -590 26580 -530
rect 26650 -590 26670 -530
rect 26560 -610 26670 -590
rect 26730 -530 26840 -510
rect 26730 -590 26750 -530
rect 26820 -590 26840 -530
rect 26730 -610 26840 -590
rect 26900 -530 27010 -510
rect 26900 -590 26920 -530
rect 26990 -590 27010 -530
rect 26900 -610 27010 -590
rect 27070 -530 27180 -510
rect 27070 -590 27090 -530
rect 27160 -590 27180 -530
rect 27070 -610 27180 -590
rect 27240 -530 27350 -510
rect 27240 -590 27260 -530
rect 27330 -590 27350 -530
rect 27240 -610 27350 -590
rect 27410 -530 27520 -510
rect 27410 -590 27430 -530
rect 27500 -590 27520 -530
rect 27410 -610 27520 -590
rect 27580 -530 27690 -510
rect 27580 -590 27600 -530
rect 27670 -590 27690 -530
rect 27580 -610 27690 -590
rect 27750 -530 27860 -510
rect 27750 -590 27770 -530
rect 27840 -590 27860 -530
rect 27750 -610 27860 -590
rect 27920 -530 28030 -510
rect 27920 -590 27940 -530
rect 28010 -590 28030 -530
rect 27920 -610 28030 -590
rect 28090 -530 28200 -510
rect 28090 -590 28110 -530
rect 28180 -590 28200 -530
rect 28090 -610 28200 -590
rect 28260 -530 28370 -510
rect 28260 -590 28280 -530
rect 28350 -590 28370 -530
rect 28260 -610 28370 -590
rect 28430 -530 28540 -510
rect 28430 -590 28450 -530
rect 28520 -590 28540 -530
rect 28430 -610 28540 -590
rect 28600 -530 28710 -510
rect 28600 -590 28620 -530
rect 28690 -590 28710 -530
rect 28600 -610 28710 -590
rect 28770 -530 28880 -510
rect 28770 -590 28790 -530
rect 28860 -590 28880 -530
rect 28770 -610 28880 -590
rect 28940 -530 29050 -510
rect 28940 -590 28960 -530
rect 29030 -590 29050 -530
rect 28940 -610 29050 -590
rect 29110 -530 29220 -510
rect 29110 -590 29130 -530
rect 29200 -590 29220 -530
rect 29110 -610 29220 -590
rect 29280 -530 29390 -510
rect 29280 -590 29300 -530
rect 29370 -590 29390 -530
rect 29280 -610 29390 -590
rect 29450 -530 29560 -510
rect 29450 -590 29470 -530
rect 29540 -590 29560 -530
rect 29450 -610 29560 -590
rect 29620 -530 29730 -510
rect 29620 -590 29640 -530
rect 29710 -590 29730 -530
rect 29620 -610 29730 -590
rect 29790 -530 29900 -510
rect 29790 -590 29810 -530
rect 29880 -590 29900 -530
rect 29790 -610 29900 -590
rect 29960 -530 30070 -510
rect 29960 -590 29980 -530
rect 30050 -590 30070 -530
rect 29960 -610 30070 -590
rect 30130 -530 30240 -510
rect 30130 -590 30150 -530
rect 30220 -590 30240 -530
rect 30130 -610 30240 -590
rect 30300 -530 30410 -510
rect 30300 -590 30320 -530
rect 30390 -590 30410 -530
rect 30300 -610 30410 -590
rect 30470 -530 30580 -510
rect 30470 -590 30490 -530
rect 30560 -590 30580 -530
rect 30470 -610 30580 -590
rect 30640 -530 30750 -510
rect 30640 -590 30660 -530
rect 30730 -590 30750 -530
rect 30640 -610 30750 -590
rect 30810 -530 30920 -510
rect 30810 -590 30830 -530
rect 30900 -590 30920 -530
rect 30810 -610 30920 -590
rect 30980 -530 31090 -510
rect 30980 -590 31000 -530
rect 31070 -590 31090 -530
rect 30980 -610 31090 -590
rect 31150 -530 31260 -510
rect 31150 -590 31170 -530
rect 31240 -590 31260 -530
rect 31150 -610 31260 -590
rect 31320 -530 31430 -510
rect 31320 -590 31340 -530
rect 31410 -590 31430 -530
rect 31320 -610 31430 -590
rect 31490 -530 31600 -510
rect 31490 -590 31510 -530
rect 31580 -590 31600 -530
rect 31490 -610 31600 -590
rect 31660 -530 31770 -510
rect 31660 -590 31680 -530
rect 31750 -590 31770 -530
rect 31660 -610 31770 -590
rect 31830 -530 31940 -510
rect 31830 -590 31850 -530
rect 31920 -590 31940 -530
rect 31830 -610 31940 -590
rect 32000 -530 32110 -510
rect 32000 -590 32020 -530
rect 32090 -590 32110 -530
rect 32000 -610 32110 -590
rect 32170 -530 32280 -510
rect 32170 -590 32190 -530
rect 32260 -590 32280 -530
rect 32170 -610 32280 -590
rect 32340 -530 32450 -510
rect 32340 -590 32360 -530
rect 32430 -590 32450 -530
rect 32340 -610 32450 -590
rect 32510 -530 32620 -510
rect 32510 -590 32530 -530
rect 32600 -590 32620 -530
rect 32510 -610 32620 -590
rect 32680 -530 32790 -510
rect 32680 -590 32700 -530
rect 32770 -590 32790 -530
rect 32680 -610 32790 -590
rect 32850 -530 32960 -510
rect 32850 -590 32870 -530
rect 32940 -590 32960 -530
rect 32850 -610 32960 -590
rect 33020 -530 33130 -510
rect 33020 -590 33040 -530
rect 33110 -590 33130 -530
rect 33020 -610 33130 -590
rect 33190 -530 33300 -510
rect 33190 -590 33210 -530
rect 33280 -590 33300 -530
rect 33190 -610 33300 -590
rect 33360 -530 33470 -510
rect 33360 -590 33380 -530
rect 33450 -590 33470 -530
rect 33360 -610 33470 -590
rect 33530 -530 33640 -510
rect 33530 -590 33550 -530
rect 33620 -590 33640 -530
rect 33530 -610 33640 -590
rect 33700 -530 33810 -510
rect 33700 -590 33720 -530
rect 33790 -590 33810 -530
rect 33700 -610 33810 -590
rect 33870 -530 33980 -510
rect 33870 -590 33890 -530
rect 33960 -590 33980 -530
rect 33870 -610 33980 -590
rect 34040 -530 34150 -510
rect 34040 -590 34060 -530
rect 34130 -590 34150 -530
rect 34040 -610 34150 -590
rect 34210 -530 34320 -510
rect 34210 -590 34230 -530
rect 34300 -590 34320 -530
rect 34210 -610 34320 -590
rect 34380 -530 34490 -510
rect 34380 -590 34400 -530
rect 34470 -590 34490 -530
rect 34380 -610 34490 -590
rect 34550 -530 34660 -510
rect 34550 -590 34570 -530
rect 34640 -590 34660 -530
rect 34550 -610 34660 -590
rect 34720 -530 34830 -510
rect 34720 -590 34740 -530
rect 34810 -590 34830 -530
rect 34720 -610 34830 -590
rect 34890 -530 35000 -510
rect 34890 -590 34910 -530
rect 34980 -590 35000 -530
rect 34890 -610 35000 -590
rect 35060 -530 35170 -510
rect 35060 -590 35080 -530
rect 35150 -590 35170 -530
rect 35060 -610 35170 -590
rect 35230 -530 35340 -510
rect 35230 -590 35250 -530
rect 35320 -590 35340 -530
rect 35230 -610 35340 -590
rect 35400 -530 35510 -510
rect 35400 -590 35420 -530
rect 35490 -590 35510 -530
rect 35400 -610 35510 -590
rect 35570 -530 35680 -510
rect 35570 -590 35590 -530
rect 35660 -590 35680 -530
rect 35570 -610 35680 -590
rect 35740 -530 35850 -510
rect 35740 -590 35760 -530
rect 35830 -590 35850 -530
rect 35740 -610 35850 -590
rect 35910 -530 36020 -510
rect 35910 -590 35930 -530
rect 36000 -590 36020 -530
rect 35910 -610 36020 -590
rect 36080 -530 36190 -510
rect 36080 -590 36100 -530
rect 36170 -590 36190 -530
rect 36080 -610 36190 -590
rect 36250 -530 36360 -510
rect 36250 -590 36270 -530
rect 36340 -590 36360 -530
rect 36250 -610 36360 -590
rect 36420 -530 36530 -510
rect 36420 -590 36440 -530
rect 36510 -590 36530 -530
rect 36420 -610 36530 -590
rect 36590 -530 36700 -510
rect 36590 -590 36610 -530
rect 36680 -590 36700 -530
rect 36590 -610 36700 -590
rect 36760 -530 36870 -510
rect 36760 -590 36780 -530
rect 36850 -590 36870 -530
rect 36760 -610 36870 -590
rect 36930 -530 37040 -510
rect 36930 -590 36950 -530
rect 37020 -590 37040 -530
rect 36930 -610 37040 -590
rect 37100 -530 37210 -510
rect 37100 -590 37120 -530
rect 37190 -590 37210 -530
rect 37100 -610 37210 -590
rect 37270 -530 37380 -510
rect 37270 -590 37290 -530
rect 37360 -590 37380 -530
rect 37270 -610 37380 -590
rect 37440 -530 37550 -510
rect 37440 -590 37460 -530
rect 37530 -590 37550 -530
rect 37440 -610 37550 -590
rect 37610 -530 37720 -510
rect 37610 -590 37630 -530
rect 37700 -590 37720 -530
rect 37610 -610 37720 -590
rect 37780 -530 37890 -510
rect 37780 -590 37800 -530
rect 37870 -590 37890 -530
rect 37780 -610 37890 -590
rect 37950 -530 38060 -510
rect 37950 -590 37970 -530
rect 38040 -590 38060 -530
rect 37950 -610 38060 -590
rect 38120 -530 38230 -510
rect 38120 -590 38140 -530
rect 38210 -590 38230 -530
rect 38120 -610 38230 -590
rect 38290 -530 38400 -510
rect 38290 -590 38310 -530
rect 38380 -590 38400 -530
rect 38290 -610 38400 -590
rect 38460 -530 38570 -510
rect 38460 -590 38480 -530
rect 38550 -590 38570 -530
rect 38460 -610 38570 -590
rect 38630 -530 38740 -510
rect 38630 -590 38650 -530
rect 38720 -590 38740 -530
rect 38630 -610 38740 -590
rect 38800 -530 38910 -510
rect 38800 -590 38820 -530
rect 38890 -590 38910 -530
rect 38800 -610 38910 -590
rect 38970 -530 39080 -510
rect 38970 -590 38990 -530
rect 39060 -590 39080 -530
rect 38970 -610 39080 -590
rect 39140 -530 39250 -510
rect 39140 -590 39160 -530
rect 39230 -590 39250 -530
rect 39140 -610 39250 -590
rect 39310 -530 39420 -510
rect 39310 -590 39330 -530
rect 39400 -590 39420 -530
rect 39310 -610 39420 -590
rect 39480 -530 39590 -510
rect 39480 -590 39500 -530
rect 39570 -590 39590 -530
rect 39480 -610 39590 -590
rect 39650 -530 39760 -510
rect 39650 -590 39670 -530
rect 39740 -590 39760 -530
rect 39650 -610 39760 -590
rect 39820 -530 39930 -510
rect 39820 -590 39840 -530
rect 39910 -590 39930 -530
rect 39820 -610 39930 -590
rect 39990 -530 40100 -510
rect 39990 -590 40010 -530
rect 40080 -590 40100 -530
rect 39990 -610 40100 -590
rect 40160 -530 40270 -510
rect 40160 -590 40180 -530
rect 40250 -590 40270 -530
rect 40160 -610 40270 -590
rect 40330 -530 40440 -510
rect 40330 -590 40350 -530
rect 40420 -590 40440 -530
rect 40330 -610 40440 -590
rect 40500 -530 40610 -510
rect 40500 -590 40520 -530
rect 40590 -590 40610 -530
rect 40500 -610 40610 -590
rect 40670 -530 40780 -510
rect 40670 -590 40690 -530
rect 40760 -590 40780 -530
rect 40670 -610 40780 -590
rect 40840 -530 40950 -510
rect 40840 -590 40860 -530
rect 40930 -590 40950 -530
rect 40840 -610 40950 -590
rect 41010 -530 41120 -510
rect 41010 -590 41030 -530
rect 41100 -590 41120 -530
rect 41010 -610 41120 -590
rect 41180 -530 41290 -510
rect 41180 -590 41200 -530
rect 41270 -590 41290 -530
rect 41180 -610 41290 -590
rect 41350 -530 41460 -510
rect 41350 -590 41370 -530
rect 41440 -590 41460 -530
rect 41350 -610 41460 -590
rect 41520 -530 41630 -510
rect 41520 -590 41540 -530
rect 41610 -590 41630 -530
rect 41520 -610 41630 -590
rect 41690 -530 41800 -510
rect 41690 -590 41710 -530
rect 41780 -590 41800 -530
rect 41690 -610 41800 -590
rect 41860 -530 41970 -510
rect 41860 -590 41880 -530
rect 41950 -590 41970 -530
rect 41860 -610 41970 -590
rect 42030 -530 42140 -510
rect 42030 -590 42050 -530
rect 42120 -590 42140 -530
rect 42030 -610 42140 -590
rect 42200 -530 42310 -510
rect 42200 -590 42220 -530
rect 42290 -590 42310 -530
rect 42200 -610 42310 -590
rect 42370 -530 42480 -510
rect 42370 -590 42390 -530
rect 42460 -590 42480 -530
rect 42370 -610 42480 -590
rect 42540 -530 42650 -510
rect 42540 -590 42560 -530
rect 42630 -590 42650 -530
rect 42540 -610 42650 -590
rect 42710 -530 42820 -510
rect 42710 -590 42730 -530
rect 42800 -590 42820 -530
rect 42710 -610 42820 -590
rect 42880 -530 42990 -510
rect 42880 -590 42900 -530
rect 42970 -590 42990 -530
rect 42880 -610 42990 -590
rect 43050 -530 43160 -510
rect 43050 -590 43070 -530
rect 43140 -590 43160 -530
rect 43050 -610 43160 -590
rect 43220 -530 43330 -510
rect 43220 -590 43240 -530
rect 43310 -590 43330 -530
rect 43220 -610 43330 -590
rect 43390 -530 43500 -510
rect 43390 -590 43410 -530
rect 43480 -590 43500 -530
rect 43390 -610 43500 -590
rect 43560 -530 43670 -510
rect 43560 -590 43580 -530
rect 43650 -590 43670 -530
rect 43560 -610 43670 -590
rect 43730 -530 43840 -510
rect 43730 -590 43750 -530
rect 43820 -590 43840 -530
rect 43730 -610 43840 -590
rect 43900 -530 44010 -510
rect 43900 -590 43920 -530
rect 43990 -590 44010 -530
rect 43900 -610 44010 -590
rect 44070 -530 44180 -510
rect 44070 -590 44090 -530
rect 44160 -590 44180 -530
rect 44070 -610 44180 -590
rect 44240 -530 44350 -510
rect 44240 -590 44260 -530
rect 44330 -590 44350 -530
rect 44240 -610 44350 -590
rect 44410 -530 44520 -510
rect 44410 -590 44430 -530
rect 44500 -590 44520 -530
rect 44410 -610 44520 -590
rect 44580 -530 44690 -510
rect 44580 -590 44600 -530
rect 44670 -590 44690 -530
rect 44580 -610 44690 -590
rect 44750 -530 44860 -510
rect 44750 -590 44770 -530
rect 44840 -590 44860 -530
rect 44750 -610 44860 -590
rect 44920 -530 45030 -510
rect 44920 -590 44940 -530
rect 45010 -590 45030 -530
rect 44920 -610 45030 -590
rect 45090 -530 45200 -510
rect 45090 -590 45110 -530
rect 45180 -590 45200 -530
rect 45090 -610 45200 -590
rect 45260 -530 45370 -510
rect 45260 -590 45280 -530
rect 45350 -590 45370 -530
rect 45260 -610 45370 -590
rect 45430 -530 45540 -510
rect 45430 -590 45450 -530
rect 45520 -590 45540 -530
rect 45430 -610 45540 -590
rect 45600 -530 45710 -510
rect 45600 -590 45620 -530
rect 45690 -590 45710 -530
rect 45600 -610 45710 -590
rect 45770 -530 45880 -510
rect 45770 -590 45790 -530
rect 45860 -590 45880 -530
rect 45770 -610 45880 -590
rect 45940 -530 46050 -510
rect 45940 -590 45960 -530
rect 46030 -590 46050 -530
rect 45940 -610 46050 -590
rect 46110 -530 46220 -510
rect 46110 -590 46130 -530
rect 46200 -590 46220 -530
rect 46110 -610 46220 -590
rect 46280 -530 46390 -510
rect 46280 -590 46300 -530
rect 46370 -590 46390 -530
rect 46280 -610 46390 -590
rect 46450 -530 46560 -510
rect 46450 -590 46470 -530
rect 46540 -590 46560 -530
rect 46450 -610 46560 -590
rect 46620 -530 46730 -510
rect 46620 -590 46640 -530
rect 46710 -590 46730 -530
rect 46620 -610 46730 -590
rect 46790 -530 46900 -510
rect 46790 -590 46810 -530
rect 46880 -590 46900 -530
rect 46790 -610 46900 -590
rect 46960 -530 47070 -510
rect 46960 -590 46980 -530
rect 47050 -590 47070 -530
rect 46960 -610 47070 -590
rect 47130 -530 47240 -510
rect 47130 -590 47150 -530
rect 47220 -590 47240 -530
rect 47130 -610 47240 -590
rect 47300 -530 47410 -510
rect 47300 -590 47320 -530
rect 47390 -590 47410 -530
rect 47300 -610 47410 -590
rect 47470 -530 47580 -510
rect 47470 -590 47490 -530
rect 47560 -590 47580 -530
rect 47470 -610 47580 -590
rect 47640 -530 47750 -510
rect 47640 -590 47660 -530
rect 47730 -590 47750 -530
rect 47640 -610 47750 -590
rect 47810 -530 47920 -510
rect 47810 -590 47830 -530
rect 47900 -590 47920 -530
rect 47810 -610 47920 -590
rect 47980 -530 48090 -510
rect 47980 -590 48000 -530
rect 48070 -590 48090 -530
rect 47980 -610 48090 -590
rect 48150 -530 48260 -510
rect 48150 -590 48170 -530
rect 48240 -590 48260 -530
rect 48150 -610 48260 -590
rect 48320 -530 48430 -510
rect 48320 -590 48340 -530
rect 48410 -590 48430 -530
rect 48320 -610 48430 -590
rect 48490 -530 48600 -510
rect 48490 -590 48510 -530
rect 48580 -590 48600 -530
rect 48490 -610 48600 -590
rect 48660 -530 48770 -510
rect 48660 -590 48680 -530
rect 48750 -590 48770 -530
rect 48660 -610 48770 -590
rect 48830 -530 48940 -510
rect 48830 -590 48850 -530
rect 48920 -590 48940 -530
rect 48830 -610 48940 -590
rect 49000 -530 49110 -510
rect 49000 -590 49020 -530
rect 49090 -590 49110 -530
rect 49000 -610 49110 -590
rect 49170 -530 49280 -510
rect 49170 -590 49190 -530
rect 49260 -590 49280 -530
rect 49170 -610 49280 -590
rect 49340 -530 49450 -510
rect 49340 -590 49360 -530
rect 49430 -590 49450 -530
rect 49340 -610 49450 -590
rect 49510 -530 49620 -510
rect 49510 -590 49530 -530
rect 49600 -590 49620 -530
rect 49510 -610 49620 -590
rect 49680 -530 49790 -510
rect 49680 -590 49700 -530
rect 49770 -590 49790 -530
rect 49680 -610 49790 -590
rect 49850 -530 49960 -510
rect 49850 -590 49870 -530
rect 49940 -590 49960 -530
rect 49850 -610 49960 -590
rect 50020 -530 50130 -510
rect 50020 -590 50040 -530
rect 50110 -590 50130 -530
rect 50020 -610 50130 -590
rect 50190 -530 50300 -510
rect 50190 -590 50210 -530
rect 50280 -590 50300 -530
rect 50190 -610 50300 -590
rect 50360 -530 50470 -510
rect 50360 -590 50380 -530
rect 50450 -590 50470 -530
rect 50360 -610 50470 -590
rect 50530 -530 50640 -510
rect 50530 -590 50550 -530
rect 50620 -590 50640 -530
rect 50530 -610 50640 -590
rect 50700 -530 50810 -510
rect 50700 -590 50720 -530
rect 50790 -590 50810 -530
rect 50700 -610 50810 -590
rect 50870 -530 50980 -510
rect 50870 -590 50890 -530
rect 50960 -590 50980 -530
rect 50870 -610 50980 -590
rect 51040 -530 51150 -510
rect 51040 -590 51060 -530
rect 51130 -590 51150 -530
rect 51040 -610 51150 -590
rect 51210 -530 51320 -510
rect 51210 -590 51230 -530
rect 51300 -590 51320 -530
rect 51210 -610 51320 -590
rect 51380 -530 51490 -510
rect 51380 -590 51400 -530
rect 51470 -590 51490 -530
rect 51380 -610 51490 -590
rect 51550 -530 51660 -510
rect 51550 -590 51570 -530
rect 51640 -590 51660 -530
rect 51550 -610 51660 -590
rect 51720 -530 51830 -510
rect 51720 -590 51740 -530
rect 51810 -590 51830 -530
rect 51720 -610 51830 -590
rect 51890 -530 52000 -510
rect 51890 -590 51910 -530
rect 51980 -590 52000 -530
rect 51890 -610 52000 -590
rect 52060 -530 52170 -510
rect 52060 -590 52080 -530
rect 52150 -590 52170 -530
rect 52060 -610 52170 -590
rect 52230 -530 52340 -510
rect 52230 -590 52250 -530
rect 52320 -590 52340 -530
rect 52230 -610 52340 -590
rect 52400 -530 52510 -510
rect 52400 -590 52420 -530
rect 52490 -590 52510 -530
rect 52400 -610 52510 -590
rect 52570 -530 52680 -510
rect 52570 -590 52590 -530
rect 52660 -590 52680 -530
rect 52570 -610 52680 -590
rect 52740 -530 52850 -510
rect 52740 -590 52760 -530
rect 52830 -590 52850 -530
rect 52740 -610 52850 -590
rect 52910 -530 53020 -510
rect 52910 -590 52930 -530
rect 53000 -590 53020 -530
rect 52910 -610 53020 -590
rect 53080 -530 53190 -510
rect 53080 -590 53100 -530
rect 53170 -590 53190 -530
rect 53080 -610 53190 -590
rect 53250 -530 53360 -510
rect 53250 -590 53270 -530
rect 53340 -590 53360 -530
rect 53250 -610 53360 -590
rect 53420 -530 53530 -510
rect 53420 -590 53440 -530
rect 53510 -590 53530 -530
rect 53420 -610 53530 -590
rect 53590 -530 53700 -510
rect 53590 -590 53610 -530
rect 53680 -590 53700 -530
rect 53590 -610 53700 -590
rect 53760 -530 53870 -510
rect 53760 -590 53780 -530
rect 53850 -590 53870 -530
rect 53760 -610 53870 -590
rect 53930 -530 54040 -510
rect 53930 -590 53950 -530
rect 54020 -590 54040 -530
rect 53930 -610 54040 -590
rect 54100 -530 54210 -510
rect 54100 -590 54120 -530
rect 54190 -590 54210 -530
rect 54100 -610 54210 -590
rect 54270 -530 54380 -510
rect 54270 -590 54290 -530
rect 54360 -590 54380 -530
rect 54270 -610 54380 -590
rect 54440 -530 54550 -510
rect 54440 -590 54460 -530
rect 54530 -590 54550 -530
rect 54440 -610 54550 -590
rect 54610 -530 54720 -510
rect 54610 -590 54630 -530
rect 54700 -590 54720 -530
rect 54610 -610 54720 -590
rect 54780 -530 54890 -510
rect 54780 -590 54800 -530
rect 54870 -590 54890 -530
rect 54780 -610 54890 -590
rect 54950 -530 55060 -510
rect 54950 -590 54970 -530
rect 55040 -590 55060 -530
rect 54950 -610 55060 -590
rect 55120 -530 55230 -510
rect 55120 -590 55140 -530
rect 55210 -590 55230 -530
rect 55120 -610 55230 -590
rect 55290 -530 55400 -510
rect 55290 -590 55310 -530
rect 55380 -590 55400 -530
rect 55290 -610 55400 -590
rect 55460 -530 55570 -510
rect 55460 -590 55480 -530
rect 55550 -590 55570 -530
rect 55460 -610 55570 -590
rect 55630 -530 55740 -510
rect 55630 -590 55650 -530
rect 55720 -590 55740 -530
rect 55630 -610 55740 -590
rect 55800 -530 55910 -510
rect 55800 -590 55820 -530
rect 55890 -590 55910 -530
rect 55800 -610 55910 -590
rect 55970 -530 56080 -510
rect 55970 -590 55990 -530
rect 56060 -590 56080 -530
rect 55970 -610 56080 -590
rect 56140 -530 56250 -510
rect 56140 -590 56160 -530
rect 56230 -590 56250 -530
rect 56140 -610 56250 -590
rect 56310 -530 56420 -510
rect 56310 -590 56330 -530
rect 56400 -590 56420 -530
rect 56310 -610 56420 -590
rect 56480 -530 56590 -510
rect 56480 -590 56500 -530
rect 56570 -590 56590 -530
rect 56480 -610 56590 -590
rect 56650 -530 56760 -510
rect 56650 -590 56670 -530
rect 56740 -590 56760 -530
rect 56650 -610 56760 -590
rect 56820 -530 56930 -510
rect 56820 -590 56840 -530
rect 56910 -590 56930 -530
rect 56820 -610 56930 -590
rect 56990 -530 57100 -510
rect 56990 -590 57010 -530
rect 57080 -590 57100 -530
rect 56990 -610 57100 -590
rect 57160 -530 57270 -510
rect 57160 -590 57180 -530
rect 57250 -590 57270 -530
rect 57160 -610 57270 -590
rect 57330 -530 57440 -510
rect 57330 -590 57350 -530
rect 57420 -590 57440 -530
rect 57330 -610 57440 -590
rect 57500 -530 57610 -510
rect 57500 -590 57520 -530
rect 57590 -590 57610 -530
rect 57500 -610 57610 -590
rect 57670 -530 57780 -510
rect 57670 -590 57690 -530
rect 57760 -590 57780 -530
rect 57670 -610 57780 -590
rect 57840 -530 57950 -510
rect 57840 -590 57860 -530
rect 57930 -590 57950 -530
rect 57840 -610 57950 -590
rect 58010 -530 58120 -510
rect 58010 -590 58030 -530
rect 58100 -590 58120 -530
rect 58010 -610 58120 -590
rect 58180 -530 58290 -510
rect 58180 -590 58200 -530
rect 58270 -590 58290 -530
rect 58180 -610 58290 -590
rect 58350 -530 58460 -510
rect 58350 -590 58370 -530
rect 58440 -590 58460 -530
rect 58350 -610 58460 -590
rect 58520 -530 58630 -510
rect 58520 -590 58540 -530
rect 58610 -590 58630 -530
rect 58520 -610 58630 -590
rect 58690 -530 58800 -510
rect 58690 -590 58710 -530
rect 58780 -590 58800 -530
rect 58690 -610 58800 -590
rect 58860 -530 58970 -510
rect 58860 -590 58880 -530
rect 58950 -590 58970 -530
rect 58860 -610 58970 -590
rect 59030 -530 59140 -510
rect 59030 -590 59050 -530
rect 59120 -590 59140 -530
rect 59030 -610 59140 -590
rect 59200 -530 59310 -510
rect 59200 -590 59220 -530
rect 59290 -590 59310 -530
rect 59200 -610 59310 -590
rect 59370 -530 59480 -510
rect 59370 -590 59390 -530
rect 59460 -590 59480 -530
rect 59370 -610 59480 -590
rect 59540 -530 59650 -510
rect 59540 -590 59560 -530
rect 59630 -590 59650 -530
rect 59540 -610 59650 -590
rect 59710 -530 59820 -510
rect 59710 -590 59730 -530
rect 59800 -590 59820 -530
rect 59710 -610 59820 -590
rect 59880 -530 59990 -510
rect 59880 -590 59900 -530
rect 59970 -590 59990 -530
rect 59880 -610 59990 -590
rect 60050 -530 60160 -510
rect 60050 -590 60070 -530
rect 60140 -590 60160 -530
rect 60050 -610 60160 -590
rect 60220 -530 60330 -510
rect 60220 -590 60240 -530
rect 60310 -590 60330 -530
rect 60220 -610 60330 -590
rect 60390 -530 60500 -510
rect 60390 -590 60410 -530
rect 60480 -590 60500 -530
rect 60390 -610 60500 -590
rect 60560 -530 60670 -510
rect 60560 -590 60580 -530
rect 60650 -590 60670 -530
rect 60560 -610 60670 -590
rect 60730 -530 60840 -510
rect 60730 -590 60750 -530
rect 60820 -590 60840 -530
rect 60730 -610 60840 -590
rect 60900 -530 61010 -510
rect 60900 -590 60920 -530
rect 60990 -590 61010 -530
rect 60900 -610 61010 -590
rect 61070 -530 61180 -510
rect 61070 -590 61090 -530
rect 61160 -590 61180 -530
rect 61070 -610 61180 -590
rect 61240 -530 61350 -510
rect 61240 -590 61260 -530
rect 61330 -590 61350 -530
rect 61240 -610 61350 -590
rect 61410 -530 61520 -510
rect 61410 -590 61430 -530
rect 61500 -590 61520 -530
rect 61410 -610 61520 -590
rect 61580 -530 61690 -510
rect 61580 -590 61600 -530
rect 61670 -590 61690 -530
rect 61580 -610 61690 -590
rect 61750 -530 61860 -510
rect 61750 -590 61770 -530
rect 61840 -590 61860 -530
rect 61750 -610 61860 -590
rect 61920 -530 62030 -510
rect 61920 -590 61940 -530
rect 62010 -590 62030 -530
rect 61920 -610 62030 -590
rect 62090 -530 62200 -510
rect 62090 -590 62110 -530
rect 62180 -590 62200 -530
rect 62090 -610 62200 -590
rect 62260 -530 62370 -510
rect 62260 -590 62280 -530
rect 62350 -590 62370 -530
rect 62260 -610 62370 -590
rect 62430 -530 62540 -510
rect 62430 -590 62450 -530
rect 62520 -590 62540 -530
rect 62430 -610 62540 -590
rect 62600 -530 62710 -510
rect 62600 -590 62620 -530
rect 62690 -590 62710 -530
rect 62600 -610 62710 -590
rect 62770 -530 62880 -510
rect 62770 -590 62790 -530
rect 62860 -590 62880 -530
rect 62770 -610 62880 -590
rect 62940 -530 63050 -510
rect 62940 -590 62960 -530
rect 63030 -590 63050 -530
rect 62940 -610 63050 -590
rect 63110 -530 63220 -510
rect 63110 -590 63130 -530
rect 63200 -590 63220 -530
rect 63110 -610 63220 -590
rect 63280 -530 63390 -510
rect 63280 -590 63300 -530
rect 63370 -590 63390 -530
rect 63280 -610 63390 -590
rect 63450 -530 63560 -510
rect 63450 -590 63470 -530
rect 63540 -590 63560 -530
rect 63450 -610 63560 -590
rect 63620 -530 63730 -510
rect 63620 -590 63640 -530
rect 63710 -590 63730 -530
rect 63620 -610 63730 -590
rect 63790 -530 63900 -510
rect 63790 -590 63810 -530
rect 63880 -590 63900 -530
rect 63790 -610 63900 -590
rect 63960 -530 64070 -510
rect 63960 -590 63980 -530
rect 64050 -590 64070 -530
rect 63960 -610 64070 -590
rect 64130 -530 64240 -510
rect 64130 -590 64150 -530
rect 64220 -590 64240 -530
rect 64130 -610 64240 -590
rect 64300 -530 64410 -510
rect 64300 -590 64320 -530
rect 64390 -590 64410 -530
rect 64300 -610 64410 -590
rect 64470 -530 64580 -510
rect 64470 -590 64490 -530
rect 64560 -590 64580 -530
rect 64470 -610 64580 -590
rect 64640 -530 64750 -510
rect 64640 -590 64660 -530
rect 64730 -590 64750 -530
rect 64640 -610 64750 -590
rect 64810 -530 64920 -510
rect 64810 -590 64830 -530
rect 64900 -590 64920 -530
rect 64810 -610 64920 -590
rect 64980 -530 65090 -510
rect 64980 -590 65000 -530
rect 65070 -590 65090 -530
rect 64980 -610 65090 -590
rect 65150 -530 65260 -510
rect 65150 -590 65170 -530
rect 65240 -590 65260 -530
rect 65150 -610 65260 -590
rect 65320 -530 65430 -510
rect 65320 -590 65340 -530
rect 65410 -590 65430 -530
rect 65320 -610 65430 -590
rect 65490 -530 65600 -510
rect 65490 -590 65510 -530
rect 65580 -590 65600 -530
rect 65490 -610 65600 -590
rect 65660 -530 65770 -510
rect 65660 -590 65680 -530
rect 65750 -590 65770 -530
rect 65660 -610 65770 -590
rect 65830 -530 65940 -510
rect 65830 -590 65850 -530
rect 65920 -590 65940 -530
rect 65830 -610 65940 -590
rect 66000 -530 66110 -510
rect 66000 -590 66020 -530
rect 66090 -590 66110 -530
rect 66000 -610 66110 -590
rect 66170 -530 66280 -510
rect 66170 -590 66190 -530
rect 66260 -590 66280 -530
rect 66170 -610 66280 -590
rect 66340 -530 66450 -510
rect 66340 -590 66360 -530
rect 66430 -590 66450 -530
rect 66340 -610 66450 -590
rect 66510 -530 66620 -510
rect 66510 -590 66530 -530
rect 66600 -590 66620 -530
rect 66510 -610 66620 -590
rect 66680 -530 66790 -510
rect 66680 -590 66700 -530
rect 66770 -590 66790 -530
rect 66680 -610 66790 -590
rect 66850 -530 66960 -510
rect 66850 -590 66870 -530
rect 66940 -590 66960 -530
rect 66850 -610 66960 -590
rect 67020 -530 67130 -510
rect 67020 -590 67040 -530
rect 67110 -590 67130 -530
rect 67020 -610 67130 -590
rect 67190 -530 67300 -510
rect 67190 -590 67210 -530
rect 67280 -590 67300 -530
rect 67190 -610 67300 -590
rect 67360 -530 67470 -510
rect 67360 -590 67380 -530
rect 67450 -590 67470 -530
rect 67360 -610 67470 -590
rect 67530 -530 67640 -510
rect 67530 -590 67550 -530
rect 67620 -590 67640 -530
rect 67530 -610 67640 -590
rect 67700 -530 67810 -510
rect 67700 -590 67720 -530
rect 67790 -590 67810 -530
rect 67700 -610 67810 -590
rect 67870 -530 67980 -510
rect 67870 -590 67890 -530
rect 67960 -590 67980 -530
rect 67870 -610 67980 -590
rect 68040 -530 68150 -510
rect 68040 -590 68060 -530
rect 68130 -590 68150 -530
rect 68040 -610 68150 -590
rect 68210 -530 68320 -510
rect 68210 -590 68230 -530
rect 68300 -590 68320 -530
rect 68210 -610 68320 -590
rect 68380 -530 68490 -510
rect 68380 -590 68400 -530
rect 68470 -590 68490 -530
rect 68380 -610 68490 -590
rect 68550 -530 68660 -510
rect 68550 -590 68570 -530
rect 68640 -590 68660 -530
rect 68550 -610 68660 -590
rect 68720 -530 68830 -510
rect 68720 -590 68740 -530
rect 68810 -590 68830 -530
rect 68720 -610 68830 -590
rect 68890 -530 69000 -510
rect 68890 -590 68910 -530
rect 68980 -590 69000 -530
rect 68890 -610 69000 -590
rect 69060 -530 69170 -510
rect 69060 -590 69080 -530
rect 69150 -590 69170 -530
rect 69060 -610 69170 -590
rect 69230 -530 69340 -510
rect 69230 -590 69250 -530
rect 69320 -590 69340 -530
rect 69230 -610 69340 -590
rect 69400 -530 69510 -510
rect 69400 -590 69420 -530
rect 69490 -590 69510 -530
rect 69400 -610 69510 -590
rect 69570 -530 69680 -510
rect 69570 -590 69590 -530
rect 69660 -590 69680 -530
rect 69570 -610 69680 -590
rect 69740 -530 69850 -510
rect 69740 -590 69760 -530
rect 69830 -590 69850 -530
rect 69740 -610 69850 -590
rect 69910 -530 70020 -510
rect 69910 -590 69930 -530
rect 70000 -590 70020 -530
rect 69910 -610 70020 -590
rect 70080 -530 70190 -510
rect 70080 -590 70100 -530
rect 70170 -590 70190 -530
rect 70080 -610 70190 -590
rect 70250 -530 70360 -510
rect 70250 -590 70270 -530
rect 70340 -590 70360 -530
rect 70250 -610 70360 -590
rect 70420 -530 70530 -510
rect 70420 -590 70440 -530
rect 70510 -590 70530 -530
rect 70420 -610 70530 -590
rect 70590 -530 70700 -510
rect 70590 -590 70610 -530
rect 70680 -590 70700 -530
rect 70590 -610 70700 -590
rect 70760 -530 70870 -510
rect 70760 -590 70780 -530
rect 70850 -590 70870 -530
rect 70760 -610 70870 -590
rect 70930 -530 71040 -510
rect 70930 -590 70950 -530
rect 71020 -590 71040 -530
rect 70930 -610 71040 -590
rect 71100 -530 71210 -510
rect 71100 -590 71120 -530
rect 71190 -590 71210 -530
rect 71100 -610 71210 -590
rect 71270 -530 71380 -510
rect 71270 -590 71290 -530
rect 71360 -590 71380 -530
rect 71270 -610 71380 -590
rect 71440 -530 71550 -510
rect 71440 -590 71460 -530
rect 71530 -590 71550 -530
rect 71440 -610 71550 -590
rect 71610 -530 71720 -510
rect 71610 -590 71630 -530
rect 71700 -590 71720 -530
rect 71610 -610 71720 -590
rect 71780 -530 71890 -510
rect 71780 -590 71800 -530
rect 71870 -590 71890 -530
rect 71780 -610 71890 -590
rect 71950 -530 72060 -510
rect 71950 -590 71970 -530
rect 72040 -590 72060 -530
rect 71950 -610 72060 -590
rect 72120 -530 72230 -510
rect 72120 -590 72140 -530
rect 72210 -590 72230 -530
rect 72120 -610 72230 -590
rect 72290 -530 72400 -510
rect 72290 -590 72310 -530
rect 72380 -590 72400 -530
rect 72290 -610 72400 -590
rect 72460 -530 72570 -510
rect 72460 -590 72480 -530
rect 72550 -590 72570 -530
rect 72460 -610 72570 -590
rect 72630 -530 72740 -510
rect 72630 -590 72650 -530
rect 72720 -590 72740 -530
rect 72630 -610 72740 -590
rect 72800 -530 72910 -510
rect 72800 -590 72820 -530
rect 72890 -590 72910 -530
rect 72800 -610 72910 -590
rect 72970 -530 73080 -510
rect 72970 -590 72990 -530
rect 73060 -590 73080 -530
rect 72970 -610 73080 -590
rect 73140 -530 73250 -510
rect 73140 -590 73160 -530
rect 73230 -590 73250 -530
rect 73140 -610 73250 -590
rect 73310 -530 73420 -510
rect 73310 -590 73330 -530
rect 73400 -590 73420 -530
rect 73310 -610 73420 -590
rect 73480 -530 73590 -510
rect 73480 -590 73500 -530
rect 73570 -590 73590 -530
rect 73480 -610 73590 -590
rect 73650 -530 73760 -510
rect 73650 -590 73670 -530
rect 73740 -590 73760 -530
rect 73650 -610 73760 -590
rect 73820 -530 73930 -510
rect 73820 -590 73840 -530
rect 73910 -590 73930 -530
rect 73820 -610 73930 -590
rect 73990 -530 74100 -510
rect 73990 -590 74010 -530
rect 74080 -590 74100 -530
rect 73990 -610 74100 -590
rect 74160 -530 74270 -510
rect 74160 -590 74180 -530
rect 74250 -590 74270 -530
rect 74160 -610 74270 -590
rect 74330 -530 74440 -510
rect 74330 -590 74350 -530
rect 74420 -590 74440 -530
rect 74330 -610 74440 -590
rect 74500 -530 74610 -510
rect 74500 -590 74520 -530
rect 74590 -590 74610 -530
rect 74500 -610 74610 -590
rect 74670 -530 74780 -510
rect 74670 -590 74690 -530
rect 74760 -590 74780 -530
rect 74670 -610 74780 -590
rect 74840 -530 74950 -510
rect 74840 -590 74860 -530
rect 74930 -590 74950 -530
rect 74840 -610 74950 -590
rect 75010 -530 75120 -510
rect 75010 -590 75030 -530
rect 75100 -590 75120 -530
rect 75010 -610 75120 -590
rect 75180 -530 75290 -510
rect 75180 -590 75200 -530
rect 75270 -590 75290 -530
rect 75180 -610 75290 -590
rect 75350 -530 75460 -510
rect 75350 -590 75370 -530
rect 75440 -590 75460 -530
rect 75350 -610 75460 -590
rect 75520 -530 75630 -510
rect 75520 -590 75540 -530
rect 75610 -590 75630 -530
rect 75520 -610 75630 -590
rect 75690 -530 75800 -510
rect 75690 -590 75710 -530
rect 75780 -590 75800 -530
rect 75690 -610 75800 -590
rect 75860 -530 75970 -510
rect 75860 -590 75880 -530
rect 75950 -590 75970 -530
rect 75860 -610 75970 -590
rect 76030 -530 76140 -510
rect 76030 -590 76050 -530
rect 76120 -590 76140 -530
rect 76030 -610 76140 -590
rect 76200 -530 76310 -510
rect 76200 -590 76220 -530
rect 76290 -590 76310 -530
rect 76200 -610 76310 -590
rect 76370 -530 76480 -510
rect 76370 -590 76390 -530
rect 76460 -590 76480 -530
rect 76370 -610 76480 -590
rect 76540 -530 76650 -510
rect 76540 -590 76560 -530
rect 76630 -590 76650 -530
rect 76540 -610 76650 -590
rect 76710 -530 76820 -510
rect 76710 -590 76730 -530
rect 76800 -590 76820 -530
rect 76710 -610 76820 -590
rect 76880 -530 76990 -510
rect 76880 -590 76900 -530
rect 76970 -590 76990 -530
rect 76880 -610 76990 -590
rect 77050 -530 77160 -510
rect 77050 -590 77070 -530
rect 77140 -590 77160 -530
rect 77050 -610 77160 -590
rect 77220 -530 77330 -510
rect 77220 -590 77240 -530
rect 77310 -590 77330 -530
rect 77220 -610 77330 -590
rect 77390 -530 77500 -510
rect 77390 -590 77410 -530
rect 77480 -590 77500 -530
rect 77390 -610 77500 -590
rect 77560 -530 77670 -510
rect 77560 -590 77580 -530
rect 77650 -590 77670 -530
rect 77560 -610 77670 -590
rect 77730 -530 77840 -510
rect 77730 -590 77750 -530
rect 77820 -590 77840 -530
rect 77730 -610 77840 -590
rect 77900 -530 78010 -510
rect 77900 -590 77920 -530
rect 77990 -590 78010 -530
rect 77900 -610 78010 -590
rect 78070 -530 78180 -510
rect 78070 -590 78090 -530
rect 78160 -590 78180 -530
rect 78070 -610 78180 -590
rect 78240 -530 78350 -510
rect 78240 -590 78260 -530
rect 78330 -590 78350 -530
rect 78240 -610 78350 -590
rect 78410 -530 78520 -510
rect 78410 -590 78430 -530
rect 78500 -590 78520 -530
rect 78410 -610 78520 -590
rect 78580 -530 78690 -510
rect 78580 -590 78600 -530
rect 78670 -590 78690 -530
rect 78580 -610 78690 -590
rect 78750 -530 78860 -510
rect 78750 -590 78770 -530
rect 78840 -590 78860 -530
rect 78750 -610 78860 -590
rect 78920 -530 79030 -510
rect 78920 -590 78940 -530
rect 79010 -590 79030 -530
rect 78920 -610 79030 -590
rect 79090 -530 79200 -510
rect 79090 -590 79110 -530
rect 79180 -590 79200 -530
rect 79090 -610 79200 -590
rect 79260 -530 79370 -510
rect 79260 -590 79280 -530
rect 79350 -590 79370 -530
rect 79260 -610 79370 -590
rect 79430 -530 79540 -510
rect 79430 -590 79450 -530
rect 79520 -590 79540 -530
rect 79430 -610 79540 -590
rect 79600 -530 79710 -510
rect 79600 -590 79620 -530
rect 79690 -590 79710 -530
rect 79600 -610 79710 -590
rect 79770 -530 79880 -510
rect 79770 -590 79790 -530
rect 79860 -590 79880 -530
rect 79770 -610 79880 -590
rect 79940 -530 80050 -510
rect 79940 -590 79960 -530
rect 80030 -590 80050 -530
rect 79940 -610 80050 -590
rect 80110 -530 80220 -510
rect 80110 -590 80130 -530
rect 80200 -590 80220 -530
rect 80110 -610 80220 -590
rect 80280 -530 80390 -510
rect 80280 -590 80300 -530
rect 80370 -590 80390 -530
rect 80280 -610 80390 -590
rect 80450 -530 80560 -510
rect 80450 -590 80470 -530
rect 80540 -590 80560 -530
rect 80450 -610 80560 -590
rect 80620 -530 80730 -510
rect 80620 -590 80640 -530
rect 80710 -590 80730 -530
rect 80620 -610 80730 -590
rect 80790 -530 80900 -510
rect 80790 -590 80810 -530
rect 80880 -590 80900 -530
rect 80790 -610 80900 -590
rect 80960 -530 81070 -510
rect 80960 -590 80980 -530
rect 81050 -590 81070 -530
rect 80960 -610 81070 -590
rect 81130 -530 81240 -510
rect 81130 -590 81150 -530
rect 81220 -590 81240 -530
rect 81130 -610 81240 -590
rect 81300 -530 81410 -510
rect 81300 -590 81320 -530
rect 81390 -590 81410 -530
rect 81300 -610 81410 -590
rect 81470 -530 81580 -510
rect 81470 -590 81490 -530
rect 81560 -590 81580 -530
rect 81470 -610 81580 -590
rect 81640 -530 81750 -510
rect 81640 -590 81660 -530
rect 81730 -590 81750 -530
rect 81640 -610 81750 -590
rect 81810 -530 81920 -510
rect 81810 -590 81830 -530
rect 81900 -590 81920 -530
rect 81810 -610 81920 -590
rect 81980 -530 82090 -510
rect 81980 -590 82000 -530
rect 82070 -590 82090 -530
rect 81980 -610 82090 -590
rect 82150 -530 82260 -510
rect 82150 -590 82170 -530
rect 82240 -590 82260 -530
rect 82150 -610 82260 -590
rect 82320 -530 82430 -510
rect 82320 -590 82340 -530
rect 82410 -590 82430 -530
rect 82320 -610 82430 -590
rect 82490 -530 82600 -510
rect 82490 -590 82510 -530
rect 82580 -590 82600 -530
rect 82490 -610 82600 -590
rect 82660 -530 82770 -510
rect 82660 -590 82680 -530
rect 82750 -590 82770 -530
rect 82660 -610 82770 -590
rect 82830 -530 82940 -510
rect 82830 -590 82850 -530
rect 82920 -590 82940 -530
rect 82830 -610 82940 -590
rect 83000 -530 83110 -510
rect 83000 -590 83020 -530
rect 83090 -590 83110 -530
rect 83000 -610 83110 -590
rect 83170 -530 83280 -510
rect 83170 -590 83190 -530
rect 83260 -590 83280 -530
rect 83170 -610 83280 -590
rect 83340 -530 83450 -510
rect 83340 -590 83360 -530
rect 83430 -590 83450 -530
rect 83340 -610 83450 -590
rect 83510 -530 83620 -510
rect 83510 -590 83530 -530
rect 83600 -590 83620 -530
rect 83510 -610 83620 -590
rect 83680 -530 83790 -510
rect 83680 -590 83700 -530
rect 83770 -590 83790 -530
rect 83680 -610 83790 -590
rect 83850 -530 83960 -510
rect 83850 -590 83870 -530
rect 83940 -590 83960 -530
rect 83850 -610 83960 -590
rect 84020 -530 84130 -510
rect 84020 -590 84040 -530
rect 84110 -590 84130 -530
rect 84020 -610 84130 -590
rect 84190 -530 84300 -510
rect 84190 -590 84210 -530
rect 84280 -590 84300 -530
rect 84190 -610 84300 -590
rect 84360 -530 84470 -510
rect 84360 -590 84380 -530
rect 84450 -590 84470 -530
rect 84360 -610 84470 -590
rect 84530 -530 84640 -510
rect 84530 -590 84550 -530
rect 84620 -590 84640 -530
rect 84530 -610 84640 -590
rect 84700 -530 84810 -510
rect 84700 -590 84720 -530
rect 84790 -590 84810 -530
rect 84700 -610 84810 -590
rect 84870 -530 84980 -510
rect 84870 -590 84890 -530
rect 84960 -590 84980 -530
rect 84870 -610 84980 -590
rect 85040 -530 85150 -510
rect 85040 -590 85060 -530
rect 85130 -590 85150 -530
rect 85040 -610 85150 -590
rect 85210 -530 85320 -510
rect 85210 -590 85230 -530
rect 85300 -590 85320 -530
rect 85210 -610 85320 -590
rect 85380 -530 85490 -510
rect 85380 -590 85400 -530
rect 85470 -590 85490 -530
rect 85380 -610 85490 -590
rect 85550 -530 85660 -510
rect 85550 -590 85570 -530
rect 85640 -590 85660 -530
rect 85550 -610 85660 -590
rect 85720 -530 85830 -510
rect 85720 -590 85740 -530
rect 85810 -590 85830 -530
rect 85720 -610 85830 -590
rect 85890 -530 86000 -510
rect 85890 -590 85910 -530
rect 85980 -590 86000 -530
rect 85890 -610 86000 -590
rect 86060 -530 86170 -510
rect 86060 -590 86080 -530
rect 86150 -590 86170 -530
rect 86060 -610 86170 -590
rect 86230 -530 86340 -510
rect 86230 -590 86250 -530
rect 86320 -590 86340 -530
rect 86230 -610 86340 -590
rect 86400 -530 86510 -510
rect 86400 -590 86420 -530
rect 86490 -590 86510 -530
rect 86400 -610 86510 -590
rect 86570 -530 86680 -510
rect 86570 -590 86590 -530
rect 86660 -590 86680 -530
rect 86570 -610 86680 -590
rect 86740 -530 86850 -510
rect 86740 -590 86760 -530
rect 86830 -590 86850 -530
rect 86740 -610 86850 -590
rect 86910 -530 87020 -510
rect 86910 -590 86930 -530
rect 87000 -590 87020 -530
rect 86910 -610 87020 -590
rect 87080 -530 87190 -510
rect 87080 -590 87100 -530
rect 87170 -590 87190 -530
rect 87080 -610 87190 -590
rect 130 -670 230 -650
rect 130 -730 150 -670
rect 210 -730 230 -670
rect 130 -770 230 -730
rect 130 -830 150 -770
rect 210 -830 230 -770
rect 130 -850 230 -830
rect 300 -670 400 -650
rect 300 -730 320 -670
rect 380 -730 400 -670
rect 300 -770 400 -730
rect 300 -830 320 -770
rect 380 -830 400 -770
rect 300 -850 400 -830
rect 470 -670 570 -650
rect 470 -730 490 -670
rect 550 -730 570 -670
rect 470 -770 570 -730
rect 470 -830 490 -770
rect 550 -830 570 -770
rect 470 -850 570 -830
rect 640 -670 740 -650
rect 640 -730 660 -670
rect 720 -730 740 -670
rect 640 -770 740 -730
rect 640 -830 660 -770
rect 720 -830 740 -770
rect 640 -850 740 -830
rect 810 -670 910 -650
rect 810 -730 830 -670
rect 890 -730 910 -670
rect 810 -770 910 -730
rect 810 -830 830 -770
rect 890 -830 910 -770
rect 810 -850 910 -830
rect 980 -670 1080 -650
rect 980 -730 1000 -670
rect 1060 -730 1080 -670
rect 980 -770 1080 -730
rect 980 -830 1000 -770
rect 1060 -830 1080 -770
rect 980 -850 1080 -830
rect 1150 -670 1250 -650
rect 1150 -730 1170 -670
rect 1230 -730 1250 -670
rect 1150 -770 1250 -730
rect 1150 -830 1170 -770
rect 1230 -830 1250 -770
rect 1150 -850 1250 -830
rect 1320 -670 1420 -650
rect 1320 -730 1340 -670
rect 1400 -730 1420 -670
rect 1320 -770 1420 -730
rect 1320 -830 1340 -770
rect 1400 -830 1420 -770
rect 1320 -850 1420 -830
rect 1490 -670 1590 -650
rect 1490 -730 1510 -670
rect 1570 -730 1590 -670
rect 1490 -770 1590 -730
rect 1490 -830 1510 -770
rect 1570 -830 1590 -770
rect 1490 -850 1590 -830
rect 1660 -670 1760 -650
rect 1660 -730 1680 -670
rect 1740 -730 1760 -670
rect 1660 -770 1760 -730
rect 1660 -830 1680 -770
rect 1740 -830 1760 -770
rect 1660 -850 1760 -830
rect 1830 -670 1930 -650
rect 1830 -730 1850 -670
rect 1910 -730 1930 -670
rect 1830 -770 1930 -730
rect 1830 -830 1850 -770
rect 1910 -830 1930 -770
rect 1830 -850 1930 -830
rect 2000 -670 2100 -650
rect 2000 -730 2020 -670
rect 2080 -730 2100 -670
rect 2000 -770 2100 -730
rect 2000 -830 2020 -770
rect 2080 -830 2100 -770
rect 2000 -850 2100 -830
rect 2170 -670 2270 -650
rect 2170 -730 2190 -670
rect 2250 -730 2270 -670
rect 2170 -770 2270 -730
rect 2170 -830 2190 -770
rect 2250 -830 2270 -770
rect 2170 -850 2270 -830
rect 2340 -670 2440 -650
rect 2340 -730 2360 -670
rect 2420 -730 2440 -670
rect 2340 -770 2440 -730
rect 2340 -830 2360 -770
rect 2420 -830 2440 -770
rect 2340 -850 2440 -830
rect 2510 -670 2610 -650
rect 2510 -730 2530 -670
rect 2590 -730 2610 -670
rect 2510 -770 2610 -730
rect 2510 -830 2530 -770
rect 2590 -830 2610 -770
rect 2510 -850 2610 -830
rect 2680 -670 2780 -650
rect 2680 -730 2700 -670
rect 2760 -730 2780 -670
rect 2680 -770 2780 -730
rect 2680 -830 2700 -770
rect 2760 -830 2780 -770
rect 2680 -850 2780 -830
rect 2850 -670 2950 -650
rect 2850 -730 2870 -670
rect 2930 -730 2950 -670
rect 2850 -770 2950 -730
rect 2850 -830 2870 -770
rect 2930 -830 2950 -770
rect 2850 -850 2950 -830
rect 3020 -670 3120 -650
rect 3020 -730 3040 -670
rect 3100 -730 3120 -670
rect 3020 -770 3120 -730
rect 3020 -830 3040 -770
rect 3100 -830 3120 -770
rect 3020 -850 3120 -830
rect 3190 -670 3290 -650
rect 3190 -730 3210 -670
rect 3270 -730 3290 -670
rect 3190 -770 3290 -730
rect 3190 -830 3210 -770
rect 3270 -830 3290 -770
rect 3190 -850 3290 -830
rect 3360 -670 3460 -650
rect 3360 -730 3380 -670
rect 3440 -730 3460 -670
rect 3360 -770 3460 -730
rect 3360 -830 3380 -770
rect 3440 -830 3460 -770
rect 3360 -850 3460 -830
rect 3530 -670 3630 -650
rect 3530 -730 3550 -670
rect 3610 -730 3630 -670
rect 3530 -770 3630 -730
rect 3530 -830 3550 -770
rect 3610 -830 3630 -770
rect 3530 -850 3630 -830
rect 3700 -670 3800 -650
rect 3700 -730 3720 -670
rect 3780 -730 3800 -670
rect 3700 -770 3800 -730
rect 3700 -830 3720 -770
rect 3780 -830 3800 -770
rect 3700 -850 3800 -830
rect 3870 -670 3970 -650
rect 3870 -730 3890 -670
rect 3950 -730 3970 -670
rect 3870 -770 3970 -730
rect 3870 -830 3890 -770
rect 3950 -830 3970 -770
rect 3870 -850 3970 -830
rect 4040 -670 4140 -650
rect 4040 -730 4060 -670
rect 4120 -730 4140 -670
rect 4040 -770 4140 -730
rect 4040 -830 4060 -770
rect 4120 -830 4140 -770
rect 4040 -850 4140 -830
rect 4210 -670 4310 -650
rect 4210 -730 4230 -670
rect 4290 -730 4310 -670
rect 4210 -770 4310 -730
rect 4210 -830 4230 -770
rect 4290 -830 4310 -770
rect 4210 -850 4310 -830
rect 4380 -670 4480 -650
rect 4380 -730 4400 -670
rect 4460 -730 4480 -670
rect 4380 -770 4480 -730
rect 4380 -830 4400 -770
rect 4460 -830 4480 -770
rect 4380 -850 4480 -830
rect 4550 -670 4650 -650
rect 4550 -730 4570 -670
rect 4630 -730 4650 -670
rect 4550 -770 4650 -730
rect 4550 -830 4570 -770
rect 4630 -830 4650 -770
rect 4550 -850 4650 -830
rect 4720 -670 4820 -650
rect 4720 -730 4740 -670
rect 4800 -730 4820 -670
rect 4720 -770 4820 -730
rect 4720 -830 4740 -770
rect 4800 -830 4820 -770
rect 4720 -850 4820 -830
rect 4890 -670 4990 -650
rect 4890 -730 4910 -670
rect 4970 -730 4990 -670
rect 4890 -770 4990 -730
rect 4890 -830 4910 -770
rect 4970 -830 4990 -770
rect 4890 -850 4990 -830
rect 5060 -670 5160 -650
rect 5060 -730 5080 -670
rect 5140 -730 5160 -670
rect 5060 -770 5160 -730
rect 5060 -830 5080 -770
rect 5140 -830 5160 -770
rect 5060 -850 5160 -830
rect 5230 -670 5330 -650
rect 5230 -730 5250 -670
rect 5310 -730 5330 -670
rect 5230 -770 5330 -730
rect 5230 -830 5250 -770
rect 5310 -830 5330 -770
rect 5230 -850 5330 -830
rect 5400 -670 5500 -650
rect 5400 -730 5420 -670
rect 5480 -730 5500 -670
rect 5400 -770 5500 -730
rect 5400 -830 5420 -770
rect 5480 -830 5500 -770
rect 5400 -850 5500 -830
rect 5570 -670 5670 -650
rect 5570 -730 5590 -670
rect 5650 -730 5670 -670
rect 5570 -770 5670 -730
rect 5570 -830 5590 -770
rect 5650 -830 5670 -770
rect 5570 -850 5670 -830
rect 5740 -670 5840 -650
rect 5740 -730 5760 -670
rect 5820 -730 5840 -670
rect 5740 -770 5840 -730
rect 5740 -830 5760 -770
rect 5820 -830 5840 -770
rect 5740 -850 5840 -830
rect 5910 -670 6010 -650
rect 5910 -730 5930 -670
rect 5990 -730 6010 -670
rect 5910 -770 6010 -730
rect 5910 -830 5930 -770
rect 5990 -830 6010 -770
rect 5910 -850 6010 -830
rect 6080 -670 6180 -650
rect 6080 -730 6100 -670
rect 6160 -730 6180 -670
rect 6080 -770 6180 -730
rect 6080 -830 6100 -770
rect 6160 -830 6180 -770
rect 6080 -850 6180 -830
rect 6250 -670 6350 -650
rect 6250 -730 6270 -670
rect 6330 -730 6350 -670
rect 6250 -770 6350 -730
rect 6250 -830 6270 -770
rect 6330 -830 6350 -770
rect 6250 -850 6350 -830
rect 6420 -670 6520 -650
rect 6420 -730 6440 -670
rect 6500 -730 6520 -670
rect 6420 -770 6520 -730
rect 6420 -830 6440 -770
rect 6500 -830 6520 -770
rect 6420 -850 6520 -830
rect 6590 -670 6690 -650
rect 6590 -730 6610 -670
rect 6670 -730 6690 -670
rect 6590 -770 6690 -730
rect 6590 -830 6610 -770
rect 6670 -830 6690 -770
rect 6590 -850 6690 -830
rect 6760 -670 6860 -650
rect 6760 -730 6780 -670
rect 6840 -730 6860 -670
rect 6760 -770 6860 -730
rect 6760 -830 6780 -770
rect 6840 -830 6860 -770
rect 6760 -850 6860 -830
rect 6930 -670 7030 -650
rect 6930 -730 6950 -670
rect 7010 -730 7030 -670
rect 6930 -770 7030 -730
rect 6930 -830 6950 -770
rect 7010 -830 7030 -770
rect 6930 -850 7030 -830
rect 7100 -670 7200 -650
rect 7100 -730 7120 -670
rect 7180 -730 7200 -670
rect 7100 -770 7200 -730
rect 7100 -830 7120 -770
rect 7180 -830 7200 -770
rect 7100 -850 7200 -830
rect 7270 -670 7370 -650
rect 7270 -730 7290 -670
rect 7350 -730 7370 -670
rect 7270 -770 7370 -730
rect 7270 -830 7290 -770
rect 7350 -830 7370 -770
rect 7270 -850 7370 -830
rect 7440 -670 7540 -650
rect 7440 -730 7460 -670
rect 7520 -730 7540 -670
rect 7440 -770 7540 -730
rect 7440 -830 7460 -770
rect 7520 -830 7540 -770
rect 7440 -850 7540 -830
rect 7610 -670 7710 -650
rect 7610 -730 7630 -670
rect 7690 -730 7710 -670
rect 7610 -770 7710 -730
rect 7610 -830 7630 -770
rect 7690 -830 7710 -770
rect 7610 -850 7710 -830
rect 7780 -670 7880 -650
rect 7780 -730 7800 -670
rect 7860 -730 7880 -670
rect 7780 -770 7880 -730
rect 7780 -830 7800 -770
rect 7860 -830 7880 -770
rect 7780 -850 7880 -830
rect 7950 -670 8050 -650
rect 7950 -730 7970 -670
rect 8030 -730 8050 -670
rect 7950 -770 8050 -730
rect 7950 -830 7970 -770
rect 8030 -830 8050 -770
rect 7950 -850 8050 -830
rect 8120 -670 8220 -650
rect 8120 -730 8140 -670
rect 8200 -730 8220 -670
rect 8120 -770 8220 -730
rect 8120 -830 8140 -770
rect 8200 -830 8220 -770
rect 8120 -850 8220 -830
rect 8290 -670 8390 -650
rect 8290 -730 8310 -670
rect 8370 -730 8390 -670
rect 8290 -770 8390 -730
rect 8290 -830 8310 -770
rect 8370 -830 8390 -770
rect 8290 -850 8390 -830
rect 8460 -670 8560 -650
rect 8460 -730 8480 -670
rect 8540 -730 8560 -670
rect 8460 -770 8560 -730
rect 8460 -830 8480 -770
rect 8540 -830 8560 -770
rect 8460 -850 8560 -830
rect 8630 -670 8730 -650
rect 8630 -730 8650 -670
rect 8710 -730 8730 -670
rect 8630 -770 8730 -730
rect 8630 -830 8650 -770
rect 8710 -830 8730 -770
rect 8630 -850 8730 -830
rect 8800 -670 8900 -650
rect 8800 -730 8820 -670
rect 8880 -730 8900 -670
rect 8800 -770 8900 -730
rect 8800 -830 8820 -770
rect 8880 -830 8900 -770
rect 8800 -850 8900 -830
rect 8970 -670 9070 -650
rect 8970 -730 8990 -670
rect 9050 -730 9070 -670
rect 8970 -770 9070 -730
rect 8970 -830 8990 -770
rect 9050 -830 9070 -770
rect 8970 -850 9070 -830
rect 9140 -670 9240 -650
rect 9140 -730 9160 -670
rect 9220 -730 9240 -670
rect 9140 -770 9240 -730
rect 9140 -830 9160 -770
rect 9220 -830 9240 -770
rect 9140 -850 9240 -830
rect 9310 -670 9410 -650
rect 9310 -730 9330 -670
rect 9390 -730 9410 -670
rect 9310 -770 9410 -730
rect 9310 -830 9330 -770
rect 9390 -830 9410 -770
rect 9310 -850 9410 -830
rect 9480 -670 9580 -650
rect 9480 -730 9500 -670
rect 9560 -730 9580 -670
rect 9480 -770 9580 -730
rect 9480 -830 9500 -770
rect 9560 -830 9580 -770
rect 9480 -850 9580 -830
rect 9650 -670 9750 -650
rect 9650 -730 9670 -670
rect 9730 -730 9750 -670
rect 9650 -770 9750 -730
rect 9650 -830 9670 -770
rect 9730 -830 9750 -770
rect 9650 -850 9750 -830
rect 9820 -670 9920 -650
rect 9820 -730 9840 -670
rect 9900 -730 9920 -670
rect 9820 -770 9920 -730
rect 9820 -830 9840 -770
rect 9900 -830 9920 -770
rect 9820 -850 9920 -830
rect 9990 -670 10090 -650
rect 9990 -730 10010 -670
rect 10070 -730 10090 -670
rect 9990 -770 10090 -730
rect 9990 -830 10010 -770
rect 10070 -830 10090 -770
rect 9990 -850 10090 -830
rect 10160 -670 10260 -650
rect 10160 -730 10180 -670
rect 10240 -730 10260 -670
rect 10160 -770 10260 -730
rect 10160 -830 10180 -770
rect 10240 -830 10260 -770
rect 10160 -850 10260 -830
rect 10330 -670 10430 -650
rect 10330 -730 10350 -670
rect 10410 -730 10430 -670
rect 10330 -770 10430 -730
rect 10330 -830 10350 -770
rect 10410 -830 10430 -770
rect 10330 -850 10430 -830
rect 10500 -670 10600 -650
rect 10500 -730 10520 -670
rect 10580 -730 10600 -670
rect 10500 -770 10600 -730
rect 10500 -830 10520 -770
rect 10580 -830 10600 -770
rect 10500 -850 10600 -830
rect 10670 -670 10770 -650
rect 10670 -730 10690 -670
rect 10750 -730 10770 -670
rect 10670 -770 10770 -730
rect 10670 -830 10690 -770
rect 10750 -830 10770 -770
rect 10670 -850 10770 -830
rect 10840 -670 10940 -650
rect 10840 -730 10860 -670
rect 10920 -730 10940 -670
rect 10840 -770 10940 -730
rect 10840 -830 10860 -770
rect 10920 -830 10940 -770
rect 10840 -850 10940 -830
rect 11010 -670 11110 -650
rect 11010 -730 11030 -670
rect 11090 -730 11110 -670
rect 11010 -770 11110 -730
rect 11010 -830 11030 -770
rect 11090 -830 11110 -770
rect 11010 -850 11110 -830
rect 11180 -670 11280 -650
rect 11180 -730 11200 -670
rect 11260 -730 11280 -670
rect 11180 -770 11280 -730
rect 11180 -830 11200 -770
rect 11260 -830 11280 -770
rect 11180 -850 11280 -830
rect 11350 -670 11450 -650
rect 11350 -730 11370 -670
rect 11430 -730 11450 -670
rect 11350 -770 11450 -730
rect 11350 -830 11370 -770
rect 11430 -830 11450 -770
rect 11350 -850 11450 -830
rect 11520 -670 11620 -650
rect 11520 -730 11540 -670
rect 11600 -730 11620 -670
rect 11520 -770 11620 -730
rect 11520 -830 11540 -770
rect 11600 -830 11620 -770
rect 11520 -850 11620 -830
rect 11690 -670 11790 -650
rect 11690 -730 11710 -670
rect 11770 -730 11790 -670
rect 11690 -770 11790 -730
rect 11690 -830 11710 -770
rect 11770 -830 11790 -770
rect 11690 -850 11790 -830
rect 11860 -670 11960 -650
rect 11860 -730 11880 -670
rect 11940 -730 11960 -670
rect 11860 -770 11960 -730
rect 11860 -830 11880 -770
rect 11940 -830 11960 -770
rect 11860 -850 11960 -830
rect 12030 -670 12130 -650
rect 12030 -730 12050 -670
rect 12110 -730 12130 -670
rect 12030 -770 12130 -730
rect 12030 -830 12050 -770
rect 12110 -830 12130 -770
rect 12030 -850 12130 -830
rect 12200 -670 12300 -650
rect 12200 -730 12220 -670
rect 12280 -730 12300 -670
rect 12200 -770 12300 -730
rect 12200 -830 12220 -770
rect 12280 -830 12300 -770
rect 12200 -850 12300 -830
rect 12370 -670 12470 -650
rect 12370 -730 12390 -670
rect 12450 -730 12470 -670
rect 12370 -770 12470 -730
rect 12370 -830 12390 -770
rect 12450 -830 12470 -770
rect 12370 -850 12470 -830
rect 12540 -670 12640 -650
rect 12540 -730 12560 -670
rect 12620 -730 12640 -670
rect 12540 -770 12640 -730
rect 12540 -830 12560 -770
rect 12620 -830 12640 -770
rect 12540 -850 12640 -830
rect 12710 -670 12810 -650
rect 12710 -730 12730 -670
rect 12790 -730 12810 -670
rect 12710 -770 12810 -730
rect 12710 -830 12730 -770
rect 12790 -830 12810 -770
rect 12710 -850 12810 -830
rect 12880 -670 12980 -650
rect 12880 -730 12900 -670
rect 12960 -730 12980 -670
rect 12880 -770 12980 -730
rect 12880 -830 12900 -770
rect 12960 -830 12980 -770
rect 12880 -850 12980 -830
rect 13050 -670 13150 -650
rect 13050 -730 13070 -670
rect 13130 -730 13150 -670
rect 13050 -770 13150 -730
rect 13050 -830 13070 -770
rect 13130 -830 13150 -770
rect 13050 -850 13150 -830
rect 13220 -670 13320 -650
rect 13220 -730 13240 -670
rect 13300 -730 13320 -670
rect 13220 -770 13320 -730
rect 13220 -830 13240 -770
rect 13300 -830 13320 -770
rect 13220 -850 13320 -830
rect 13390 -670 13490 -650
rect 13390 -730 13410 -670
rect 13470 -730 13490 -670
rect 13390 -770 13490 -730
rect 13390 -830 13410 -770
rect 13470 -830 13490 -770
rect 13390 -850 13490 -830
rect 13560 -670 13660 -650
rect 13560 -730 13580 -670
rect 13640 -730 13660 -670
rect 13560 -770 13660 -730
rect 13560 -830 13580 -770
rect 13640 -830 13660 -770
rect 13560 -850 13660 -830
rect 13730 -670 13830 -650
rect 13730 -730 13750 -670
rect 13810 -730 13830 -670
rect 13730 -770 13830 -730
rect 13730 -830 13750 -770
rect 13810 -830 13830 -770
rect 13730 -850 13830 -830
rect 13900 -670 14000 -650
rect 13900 -730 13920 -670
rect 13980 -730 14000 -670
rect 13900 -770 14000 -730
rect 13900 -830 13920 -770
rect 13980 -830 14000 -770
rect 13900 -850 14000 -830
rect 14070 -670 14170 -650
rect 14070 -730 14090 -670
rect 14150 -730 14170 -670
rect 14070 -770 14170 -730
rect 14070 -830 14090 -770
rect 14150 -830 14170 -770
rect 14070 -850 14170 -830
rect 14240 -670 14340 -650
rect 14240 -730 14260 -670
rect 14320 -730 14340 -670
rect 14240 -770 14340 -730
rect 14240 -830 14260 -770
rect 14320 -830 14340 -770
rect 14240 -850 14340 -830
rect 14410 -670 14510 -650
rect 14410 -730 14430 -670
rect 14490 -730 14510 -670
rect 14410 -770 14510 -730
rect 14410 -830 14430 -770
rect 14490 -830 14510 -770
rect 14410 -850 14510 -830
rect 14580 -670 14680 -650
rect 14580 -730 14600 -670
rect 14660 -730 14680 -670
rect 14580 -770 14680 -730
rect 14580 -830 14600 -770
rect 14660 -830 14680 -770
rect 14580 -850 14680 -830
rect 14750 -670 14850 -650
rect 14750 -730 14770 -670
rect 14830 -730 14850 -670
rect 14750 -770 14850 -730
rect 14750 -830 14770 -770
rect 14830 -830 14850 -770
rect 14750 -850 14850 -830
rect 14920 -670 15020 -650
rect 14920 -730 14940 -670
rect 15000 -730 15020 -670
rect 14920 -770 15020 -730
rect 14920 -830 14940 -770
rect 15000 -830 15020 -770
rect 14920 -850 15020 -830
rect 15090 -670 15190 -650
rect 15090 -730 15110 -670
rect 15170 -730 15190 -670
rect 15090 -770 15190 -730
rect 15090 -830 15110 -770
rect 15170 -830 15190 -770
rect 15090 -850 15190 -830
rect 15260 -670 15360 -650
rect 15260 -730 15280 -670
rect 15340 -730 15360 -670
rect 15260 -770 15360 -730
rect 15260 -830 15280 -770
rect 15340 -830 15360 -770
rect 15260 -850 15360 -830
rect 15430 -670 15530 -650
rect 15430 -730 15450 -670
rect 15510 -730 15530 -670
rect 15430 -770 15530 -730
rect 15430 -830 15450 -770
rect 15510 -830 15530 -770
rect 15430 -850 15530 -830
rect 15600 -670 15700 -650
rect 15600 -730 15620 -670
rect 15680 -730 15700 -670
rect 15600 -770 15700 -730
rect 15600 -830 15620 -770
rect 15680 -830 15700 -770
rect 15600 -850 15700 -830
rect 15770 -670 15870 -650
rect 15770 -730 15790 -670
rect 15850 -730 15870 -670
rect 15770 -770 15870 -730
rect 15770 -830 15790 -770
rect 15850 -830 15870 -770
rect 15770 -850 15870 -830
rect 15940 -670 16040 -650
rect 15940 -730 15960 -670
rect 16020 -730 16040 -670
rect 15940 -770 16040 -730
rect 15940 -830 15960 -770
rect 16020 -830 16040 -770
rect 15940 -850 16040 -830
rect 16110 -670 16210 -650
rect 16110 -730 16130 -670
rect 16190 -730 16210 -670
rect 16110 -770 16210 -730
rect 16110 -830 16130 -770
rect 16190 -830 16210 -770
rect 16110 -850 16210 -830
rect 16280 -670 16380 -650
rect 16280 -730 16300 -670
rect 16360 -730 16380 -670
rect 16280 -770 16380 -730
rect 16280 -830 16300 -770
rect 16360 -830 16380 -770
rect 16280 -850 16380 -830
rect 16450 -670 16550 -650
rect 16450 -730 16470 -670
rect 16530 -730 16550 -670
rect 16450 -770 16550 -730
rect 16450 -830 16470 -770
rect 16530 -830 16550 -770
rect 16450 -850 16550 -830
rect 16620 -670 16720 -650
rect 16620 -730 16640 -670
rect 16700 -730 16720 -670
rect 16620 -770 16720 -730
rect 16620 -830 16640 -770
rect 16700 -830 16720 -770
rect 16620 -850 16720 -830
rect 16790 -670 16890 -650
rect 16790 -730 16810 -670
rect 16870 -730 16890 -670
rect 16790 -770 16890 -730
rect 16790 -830 16810 -770
rect 16870 -830 16890 -770
rect 16790 -850 16890 -830
rect 16960 -670 17060 -650
rect 16960 -730 16980 -670
rect 17040 -730 17060 -670
rect 16960 -770 17060 -730
rect 16960 -830 16980 -770
rect 17040 -830 17060 -770
rect 16960 -850 17060 -830
rect 17130 -670 17230 -650
rect 17130 -730 17150 -670
rect 17210 -730 17230 -670
rect 17130 -770 17230 -730
rect 17130 -830 17150 -770
rect 17210 -830 17230 -770
rect 17130 -850 17230 -830
rect 17300 -670 17400 -650
rect 17300 -730 17320 -670
rect 17380 -730 17400 -670
rect 17300 -770 17400 -730
rect 17300 -830 17320 -770
rect 17380 -830 17400 -770
rect 17300 -850 17400 -830
rect 17470 -670 17570 -650
rect 17470 -730 17490 -670
rect 17550 -730 17570 -670
rect 17470 -770 17570 -730
rect 17470 -830 17490 -770
rect 17550 -830 17570 -770
rect 17470 -850 17570 -830
rect 17640 -670 17740 -650
rect 17640 -730 17660 -670
rect 17720 -730 17740 -670
rect 17640 -770 17740 -730
rect 17640 -830 17660 -770
rect 17720 -830 17740 -770
rect 17640 -850 17740 -830
rect 17810 -670 17910 -650
rect 17810 -730 17830 -670
rect 17890 -730 17910 -670
rect 17810 -770 17910 -730
rect 17810 -830 17830 -770
rect 17890 -830 17910 -770
rect 17810 -850 17910 -830
rect 17980 -670 18080 -650
rect 17980 -730 18000 -670
rect 18060 -730 18080 -670
rect 17980 -770 18080 -730
rect 17980 -830 18000 -770
rect 18060 -830 18080 -770
rect 17980 -850 18080 -830
rect 18150 -670 18250 -650
rect 18150 -730 18170 -670
rect 18230 -730 18250 -670
rect 18150 -770 18250 -730
rect 18150 -830 18170 -770
rect 18230 -830 18250 -770
rect 18150 -850 18250 -830
rect 18320 -670 18420 -650
rect 18320 -730 18340 -670
rect 18400 -730 18420 -670
rect 18320 -770 18420 -730
rect 18320 -830 18340 -770
rect 18400 -830 18420 -770
rect 18320 -850 18420 -830
rect 18490 -670 18590 -650
rect 18490 -730 18510 -670
rect 18570 -730 18590 -670
rect 18490 -770 18590 -730
rect 18490 -830 18510 -770
rect 18570 -830 18590 -770
rect 18490 -850 18590 -830
rect 18660 -670 18760 -650
rect 18660 -730 18680 -670
rect 18740 -730 18760 -670
rect 18660 -770 18760 -730
rect 18660 -830 18680 -770
rect 18740 -830 18760 -770
rect 18660 -850 18760 -830
rect 18830 -670 18930 -650
rect 18830 -730 18850 -670
rect 18910 -730 18930 -670
rect 18830 -770 18930 -730
rect 18830 -830 18850 -770
rect 18910 -830 18930 -770
rect 18830 -850 18930 -830
rect 19000 -670 19100 -650
rect 19000 -730 19020 -670
rect 19080 -730 19100 -670
rect 19000 -770 19100 -730
rect 19000 -830 19020 -770
rect 19080 -830 19100 -770
rect 19000 -850 19100 -830
rect 19170 -670 19270 -650
rect 19170 -730 19190 -670
rect 19250 -730 19270 -670
rect 19170 -770 19270 -730
rect 19170 -830 19190 -770
rect 19250 -830 19270 -770
rect 19170 -850 19270 -830
rect 19340 -670 19440 -650
rect 19340 -730 19360 -670
rect 19420 -730 19440 -670
rect 19340 -770 19440 -730
rect 19340 -830 19360 -770
rect 19420 -830 19440 -770
rect 19340 -850 19440 -830
rect 19510 -670 19610 -650
rect 19510 -730 19530 -670
rect 19590 -730 19610 -670
rect 19510 -770 19610 -730
rect 19510 -830 19530 -770
rect 19590 -830 19610 -770
rect 19510 -850 19610 -830
rect 19680 -670 19780 -650
rect 19680 -730 19700 -670
rect 19760 -730 19780 -670
rect 19680 -770 19780 -730
rect 19680 -830 19700 -770
rect 19760 -830 19780 -770
rect 19680 -850 19780 -830
rect 19850 -670 19950 -650
rect 19850 -730 19870 -670
rect 19930 -730 19950 -670
rect 19850 -770 19950 -730
rect 19850 -830 19870 -770
rect 19930 -830 19950 -770
rect 19850 -850 19950 -830
rect 20020 -670 20120 -650
rect 20020 -730 20040 -670
rect 20100 -730 20120 -670
rect 20020 -770 20120 -730
rect 20020 -830 20040 -770
rect 20100 -830 20120 -770
rect 20020 -850 20120 -830
rect 20190 -670 20290 -650
rect 20190 -730 20210 -670
rect 20270 -730 20290 -670
rect 20190 -770 20290 -730
rect 20190 -830 20210 -770
rect 20270 -830 20290 -770
rect 20190 -850 20290 -830
rect 20360 -670 20460 -650
rect 20360 -730 20380 -670
rect 20440 -730 20460 -670
rect 20360 -770 20460 -730
rect 20360 -830 20380 -770
rect 20440 -830 20460 -770
rect 20360 -850 20460 -830
rect 20530 -670 20630 -650
rect 20530 -730 20550 -670
rect 20610 -730 20630 -670
rect 20530 -770 20630 -730
rect 20530 -830 20550 -770
rect 20610 -830 20630 -770
rect 20530 -850 20630 -830
rect 20700 -670 20800 -650
rect 20700 -730 20720 -670
rect 20780 -730 20800 -670
rect 20700 -770 20800 -730
rect 20700 -830 20720 -770
rect 20780 -830 20800 -770
rect 20700 -850 20800 -830
rect 20870 -670 20970 -650
rect 20870 -730 20890 -670
rect 20950 -730 20970 -670
rect 20870 -770 20970 -730
rect 20870 -830 20890 -770
rect 20950 -830 20970 -770
rect 20870 -850 20970 -830
rect 21040 -670 21140 -650
rect 21040 -730 21060 -670
rect 21120 -730 21140 -670
rect 21040 -770 21140 -730
rect 21040 -830 21060 -770
rect 21120 -830 21140 -770
rect 21040 -850 21140 -830
rect 21210 -670 21310 -650
rect 21210 -730 21230 -670
rect 21290 -730 21310 -670
rect 21210 -770 21310 -730
rect 21210 -830 21230 -770
rect 21290 -830 21310 -770
rect 21210 -850 21310 -830
rect 21380 -670 21480 -650
rect 21380 -730 21400 -670
rect 21460 -730 21480 -670
rect 21380 -770 21480 -730
rect 21380 -830 21400 -770
rect 21460 -830 21480 -770
rect 21380 -850 21480 -830
rect 21550 -670 21650 -650
rect 21550 -730 21570 -670
rect 21630 -730 21650 -670
rect 21550 -770 21650 -730
rect 21550 -830 21570 -770
rect 21630 -830 21650 -770
rect 21550 -850 21650 -830
rect 21720 -670 21820 -650
rect 21720 -730 21740 -670
rect 21800 -730 21820 -670
rect 21720 -770 21820 -730
rect 21720 -830 21740 -770
rect 21800 -830 21820 -770
rect 21720 -850 21820 -830
rect 21890 -670 21990 -650
rect 21890 -730 21910 -670
rect 21970 -730 21990 -670
rect 21890 -770 21990 -730
rect 21890 -830 21910 -770
rect 21970 -830 21990 -770
rect 21890 -850 21990 -830
rect 22060 -670 22160 -650
rect 22060 -730 22080 -670
rect 22140 -730 22160 -670
rect 22060 -770 22160 -730
rect 22060 -830 22080 -770
rect 22140 -830 22160 -770
rect 22060 -850 22160 -830
rect 22230 -670 22330 -650
rect 22230 -730 22250 -670
rect 22310 -730 22330 -670
rect 22230 -770 22330 -730
rect 22230 -830 22250 -770
rect 22310 -830 22330 -770
rect 22230 -850 22330 -830
rect 22400 -670 22500 -650
rect 22400 -730 22420 -670
rect 22480 -730 22500 -670
rect 22400 -770 22500 -730
rect 22400 -830 22420 -770
rect 22480 -830 22500 -770
rect 22400 -850 22500 -830
rect 22570 -670 22670 -650
rect 22570 -730 22590 -670
rect 22650 -730 22670 -670
rect 22570 -770 22670 -730
rect 22570 -830 22590 -770
rect 22650 -830 22670 -770
rect 22570 -850 22670 -830
rect 22740 -670 22840 -650
rect 22740 -730 22760 -670
rect 22820 -730 22840 -670
rect 22740 -770 22840 -730
rect 22740 -830 22760 -770
rect 22820 -830 22840 -770
rect 22740 -850 22840 -830
rect 22910 -670 23010 -650
rect 22910 -730 22930 -670
rect 22990 -730 23010 -670
rect 22910 -770 23010 -730
rect 22910 -830 22930 -770
rect 22990 -830 23010 -770
rect 22910 -850 23010 -830
rect 23080 -670 23180 -650
rect 23080 -730 23100 -670
rect 23160 -730 23180 -670
rect 23080 -770 23180 -730
rect 23080 -830 23100 -770
rect 23160 -830 23180 -770
rect 23080 -850 23180 -830
rect 23250 -670 23350 -650
rect 23250 -730 23270 -670
rect 23330 -730 23350 -670
rect 23250 -770 23350 -730
rect 23250 -830 23270 -770
rect 23330 -830 23350 -770
rect 23250 -850 23350 -830
rect 23420 -670 23520 -650
rect 23420 -730 23440 -670
rect 23500 -730 23520 -670
rect 23420 -770 23520 -730
rect 23420 -830 23440 -770
rect 23500 -830 23520 -770
rect 23420 -850 23520 -830
rect 23590 -670 23690 -650
rect 23590 -730 23610 -670
rect 23670 -730 23690 -670
rect 23590 -770 23690 -730
rect 23590 -830 23610 -770
rect 23670 -830 23690 -770
rect 23590 -850 23690 -830
rect 23760 -670 23860 -650
rect 23760 -730 23780 -670
rect 23840 -730 23860 -670
rect 23760 -770 23860 -730
rect 23760 -830 23780 -770
rect 23840 -830 23860 -770
rect 23760 -850 23860 -830
rect 23930 -670 24030 -650
rect 23930 -730 23950 -670
rect 24010 -730 24030 -670
rect 23930 -770 24030 -730
rect 23930 -830 23950 -770
rect 24010 -830 24030 -770
rect 23930 -850 24030 -830
rect 24100 -670 24200 -650
rect 24100 -730 24120 -670
rect 24180 -730 24200 -670
rect 24100 -770 24200 -730
rect 24100 -830 24120 -770
rect 24180 -830 24200 -770
rect 24100 -850 24200 -830
rect 24270 -670 24370 -650
rect 24270 -730 24290 -670
rect 24350 -730 24370 -670
rect 24270 -770 24370 -730
rect 24270 -830 24290 -770
rect 24350 -830 24370 -770
rect 24270 -850 24370 -830
rect 24440 -670 24540 -650
rect 24440 -730 24460 -670
rect 24520 -730 24540 -670
rect 24440 -770 24540 -730
rect 24440 -830 24460 -770
rect 24520 -830 24540 -770
rect 24440 -850 24540 -830
rect 24610 -670 24710 -650
rect 24610 -730 24630 -670
rect 24690 -730 24710 -670
rect 24610 -770 24710 -730
rect 24610 -830 24630 -770
rect 24690 -830 24710 -770
rect 24610 -850 24710 -830
rect 24780 -670 24880 -650
rect 24780 -730 24800 -670
rect 24860 -730 24880 -670
rect 24780 -770 24880 -730
rect 24780 -830 24800 -770
rect 24860 -830 24880 -770
rect 24780 -850 24880 -830
rect 24950 -670 25050 -650
rect 24950 -730 24970 -670
rect 25030 -730 25050 -670
rect 24950 -770 25050 -730
rect 24950 -830 24970 -770
rect 25030 -830 25050 -770
rect 24950 -850 25050 -830
rect 25120 -670 25220 -650
rect 25120 -730 25140 -670
rect 25200 -730 25220 -670
rect 25120 -770 25220 -730
rect 25120 -830 25140 -770
rect 25200 -830 25220 -770
rect 25120 -850 25220 -830
rect 25290 -670 25390 -650
rect 25290 -730 25310 -670
rect 25370 -730 25390 -670
rect 25290 -770 25390 -730
rect 25290 -830 25310 -770
rect 25370 -830 25390 -770
rect 25290 -850 25390 -830
rect 25460 -670 25560 -650
rect 25460 -730 25480 -670
rect 25540 -730 25560 -670
rect 25460 -770 25560 -730
rect 25460 -830 25480 -770
rect 25540 -830 25560 -770
rect 25460 -850 25560 -830
rect 25630 -670 25730 -650
rect 25630 -730 25650 -670
rect 25710 -730 25730 -670
rect 25630 -770 25730 -730
rect 25630 -830 25650 -770
rect 25710 -830 25730 -770
rect 25630 -850 25730 -830
rect 25800 -670 25900 -650
rect 25800 -730 25820 -670
rect 25880 -730 25900 -670
rect 25800 -770 25900 -730
rect 25800 -830 25820 -770
rect 25880 -830 25900 -770
rect 25800 -850 25900 -830
rect 25970 -670 26070 -650
rect 25970 -730 25990 -670
rect 26050 -730 26070 -670
rect 25970 -770 26070 -730
rect 25970 -830 25990 -770
rect 26050 -830 26070 -770
rect 25970 -850 26070 -830
rect 26140 -670 26240 -650
rect 26140 -730 26160 -670
rect 26220 -730 26240 -670
rect 26140 -770 26240 -730
rect 26140 -830 26160 -770
rect 26220 -830 26240 -770
rect 26140 -850 26240 -830
rect 26310 -670 26410 -650
rect 26310 -730 26330 -670
rect 26390 -730 26410 -670
rect 26310 -770 26410 -730
rect 26310 -830 26330 -770
rect 26390 -830 26410 -770
rect 26310 -850 26410 -830
rect 26480 -670 26580 -650
rect 26480 -730 26500 -670
rect 26560 -730 26580 -670
rect 26480 -770 26580 -730
rect 26480 -830 26500 -770
rect 26560 -830 26580 -770
rect 26480 -850 26580 -830
rect 26650 -670 26750 -650
rect 26650 -730 26670 -670
rect 26730 -730 26750 -670
rect 26650 -770 26750 -730
rect 26650 -830 26670 -770
rect 26730 -830 26750 -770
rect 26650 -850 26750 -830
rect 26820 -670 26920 -650
rect 26820 -730 26840 -670
rect 26900 -730 26920 -670
rect 26820 -770 26920 -730
rect 26820 -830 26840 -770
rect 26900 -830 26920 -770
rect 26820 -850 26920 -830
rect 26990 -670 27090 -650
rect 26990 -730 27010 -670
rect 27070 -730 27090 -670
rect 26990 -770 27090 -730
rect 26990 -830 27010 -770
rect 27070 -830 27090 -770
rect 26990 -850 27090 -830
rect 27160 -670 27260 -650
rect 27160 -730 27180 -670
rect 27240 -730 27260 -670
rect 27160 -770 27260 -730
rect 27160 -830 27180 -770
rect 27240 -830 27260 -770
rect 27160 -850 27260 -830
rect 27330 -670 27430 -650
rect 27330 -730 27350 -670
rect 27410 -730 27430 -670
rect 27330 -770 27430 -730
rect 27330 -830 27350 -770
rect 27410 -830 27430 -770
rect 27330 -850 27430 -830
rect 27500 -670 27600 -650
rect 27500 -730 27520 -670
rect 27580 -730 27600 -670
rect 27500 -770 27600 -730
rect 27500 -830 27520 -770
rect 27580 -830 27600 -770
rect 27500 -850 27600 -830
rect 27670 -670 27770 -650
rect 27670 -730 27690 -670
rect 27750 -730 27770 -670
rect 27670 -770 27770 -730
rect 27670 -830 27690 -770
rect 27750 -830 27770 -770
rect 27670 -850 27770 -830
rect 27840 -670 27940 -650
rect 27840 -730 27860 -670
rect 27920 -730 27940 -670
rect 27840 -770 27940 -730
rect 27840 -830 27860 -770
rect 27920 -830 27940 -770
rect 27840 -850 27940 -830
rect 28010 -670 28110 -650
rect 28010 -730 28030 -670
rect 28090 -730 28110 -670
rect 28010 -770 28110 -730
rect 28010 -830 28030 -770
rect 28090 -830 28110 -770
rect 28010 -850 28110 -830
rect 28180 -670 28280 -650
rect 28180 -730 28200 -670
rect 28260 -730 28280 -670
rect 28180 -770 28280 -730
rect 28180 -830 28200 -770
rect 28260 -830 28280 -770
rect 28180 -850 28280 -830
rect 28350 -670 28450 -650
rect 28350 -730 28370 -670
rect 28430 -730 28450 -670
rect 28350 -770 28450 -730
rect 28350 -830 28370 -770
rect 28430 -830 28450 -770
rect 28350 -850 28450 -830
rect 28520 -670 28620 -650
rect 28520 -730 28540 -670
rect 28600 -730 28620 -670
rect 28520 -770 28620 -730
rect 28520 -830 28540 -770
rect 28600 -830 28620 -770
rect 28520 -850 28620 -830
rect 28690 -670 28790 -650
rect 28690 -730 28710 -670
rect 28770 -730 28790 -670
rect 28690 -770 28790 -730
rect 28690 -830 28710 -770
rect 28770 -830 28790 -770
rect 28690 -850 28790 -830
rect 28860 -670 28960 -650
rect 28860 -730 28880 -670
rect 28940 -730 28960 -670
rect 28860 -770 28960 -730
rect 28860 -830 28880 -770
rect 28940 -830 28960 -770
rect 28860 -850 28960 -830
rect 29030 -670 29130 -650
rect 29030 -730 29050 -670
rect 29110 -730 29130 -670
rect 29030 -770 29130 -730
rect 29030 -830 29050 -770
rect 29110 -830 29130 -770
rect 29030 -850 29130 -830
rect 29200 -670 29300 -650
rect 29200 -730 29220 -670
rect 29280 -730 29300 -670
rect 29200 -770 29300 -730
rect 29200 -830 29220 -770
rect 29280 -830 29300 -770
rect 29200 -850 29300 -830
rect 29370 -670 29470 -650
rect 29370 -730 29390 -670
rect 29450 -730 29470 -670
rect 29370 -770 29470 -730
rect 29370 -830 29390 -770
rect 29450 -830 29470 -770
rect 29370 -850 29470 -830
rect 29540 -670 29640 -650
rect 29540 -730 29560 -670
rect 29620 -730 29640 -670
rect 29540 -770 29640 -730
rect 29540 -830 29560 -770
rect 29620 -830 29640 -770
rect 29540 -850 29640 -830
rect 29710 -670 29810 -650
rect 29710 -730 29730 -670
rect 29790 -730 29810 -670
rect 29710 -770 29810 -730
rect 29710 -830 29730 -770
rect 29790 -830 29810 -770
rect 29710 -850 29810 -830
rect 29880 -670 29980 -650
rect 29880 -730 29900 -670
rect 29960 -730 29980 -670
rect 29880 -770 29980 -730
rect 29880 -830 29900 -770
rect 29960 -830 29980 -770
rect 29880 -850 29980 -830
rect 30050 -670 30150 -650
rect 30050 -730 30070 -670
rect 30130 -730 30150 -670
rect 30050 -770 30150 -730
rect 30050 -830 30070 -770
rect 30130 -830 30150 -770
rect 30050 -850 30150 -830
rect 30220 -670 30320 -650
rect 30220 -730 30240 -670
rect 30300 -730 30320 -670
rect 30220 -770 30320 -730
rect 30220 -830 30240 -770
rect 30300 -830 30320 -770
rect 30220 -850 30320 -830
rect 30390 -670 30490 -650
rect 30390 -730 30410 -670
rect 30470 -730 30490 -670
rect 30390 -770 30490 -730
rect 30390 -830 30410 -770
rect 30470 -830 30490 -770
rect 30390 -850 30490 -830
rect 30560 -670 30660 -650
rect 30560 -730 30580 -670
rect 30640 -730 30660 -670
rect 30560 -770 30660 -730
rect 30560 -830 30580 -770
rect 30640 -830 30660 -770
rect 30560 -850 30660 -830
rect 30730 -670 30830 -650
rect 30730 -730 30750 -670
rect 30810 -730 30830 -670
rect 30730 -770 30830 -730
rect 30730 -830 30750 -770
rect 30810 -830 30830 -770
rect 30730 -850 30830 -830
rect 30900 -670 31000 -650
rect 30900 -730 30920 -670
rect 30980 -730 31000 -670
rect 30900 -770 31000 -730
rect 30900 -830 30920 -770
rect 30980 -830 31000 -770
rect 30900 -850 31000 -830
rect 31070 -670 31170 -650
rect 31070 -730 31090 -670
rect 31150 -730 31170 -670
rect 31070 -770 31170 -730
rect 31070 -830 31090 -770
rect 31150 -830 31170 -770
rect 31070 -850 31170 -830
rect 31240 -670 31340 -650
rect 31240 -730 31260 -670
rect 31320 -730 31340 -670
rect 31240 -770 31340 -730
rect 31240 -830 31260 -770
rect 31320 -830 31340 -770
rect 31240 -850 31340 -830
rect 31410 -670 31510 -650
rect 31410 -730 31430 -670
rect 31490 -730 31510 -670
rect 31410 -770 31510 -730
rect 31410 -830 31430 -770
rect 31490 -830 31510 -770
rect 31410 -850 31510 -830
rect 31580 -670 31680 -650
rect 31580 -730 31600 -670
rect 31660 -730 31680 -670
rect 31580 -770 31680 -730
rect 31580 -830 31600 -770
rect 31660 -830 31680 -770
rect 31580 -850 31680 -830
rect 31750 -670 31850 -650
rect 31750 -730 31770 -670
rect 31830 -730 31850 -670
rect 31750 -770 31850 -730
rect 31750 -830 31770 -770
rect 31830 -830 31850 -770
rect 31750 -850 31850 -830
rect 31920 -670 32020 -650
rect 31920 -730 31940 -670
rect 32000 -730 32020 -670
rect 31920 -770 32020 -730
rect 31920 -830 31940 -770
rect 32000 -830 32020 -770
rect 31920 -850 32020 -830
rect 32090 -670 32190 -650
rect 32090 -730 32110 -670
rect 32170 -730 32190 -670
rect 32090 -770 32190 -730
rect 32090 -830 32110 -770
rect 32170 -830 32190 -770
rect 32090 -850 32190 -830
rect 32260 -670 32360 -650
rect 32260 -730 32280 -670
rect 32340 -730 32360 -670
rect 32260 -770 32360 -730
rect 32260 -830 32280 -770
rect 32340 -830 32360 -770
rect 32260 -850 32360 -830
rect 32430 -670 32530 -650
rect 32430 -730 32450 -670
rect 32510 -730 32530 -670
rect 32430 -770 32530 -730
rect 32430 -830 32450 -770
rect 32510 -830 32530 -770
rect 32430 -850 32530 -830
rect 32600 -670 32700 -650
rect 32600 -730 32620 -670
rect 32680 -730 32700 -670
rect 32600 -770 32700 -730
rect 32600 -830 32620 -770
rect 32680 -830 32700 -770
rect 32600 -850 32700 -830
rect 32770 -670 32870 -650
rect 32770 -730 32790 -670
rect 32850 -730 32870 -670
rect 32770 -770 32870 -730
rect 32770 -830 32790 -770
rect 32850 -830 32870 -770
rect 32770 -850 32870 -830
rect 32940 -670 33040 -650
rect 32940 -730 32960 -670
rect 33020 -730 33040 -670
rect 32940 -770 33040 -730
rect 32940 -830 32960 -770
rect 33020 -830 33040 -770
rect 32940 -850 33040 -830
rect 33110 -670 33210 -650
rect 33110 -730 33130 -670
rect 33190 -730 33210 -670
rect 33110 -770 33210 -730
rect 33110 -830 33130 -770
rect 33190 -830 33210 -770
rect 33110 -850 33210 -830
rect 33280 -670 33380 -650
rect 33280 -730 33300 -670
rect 33360 -730 33380 -670
rect 33280 -770 33380 -730
rect 33280 -830 33300 -770
rect 33360 -830 33380 -770
rect 33280 -850 33380 -830
rect 33450 -670 33550 -650
rect 33450 -730 33470 -670
rect 33530 -730 33550 -670
rect 33450 -770 33550 -730
rect 33450 -830 33470 -770
rect 33530 -830 33550 -770
rect 33450 -850 33550 -830
rect 33620 -670 33720 -650
rect 33620 -730 33640 -670
rect 33700 -730 33720 -670
rect 33620 -770 33720 -730
rect 33620 -830 33640 -770
rect 33700 -830 33720 -770
rect 33620 -850 33720 -830
rect 33790 -670 33890 -650
rect 33790 -730 33810 -670
rect 33870 -730 33890 -670
rect 33790 -770 33890 -730
rect 33790 -830 33810 -770
rect 33870 -830 33890 -770
rect 33790 -850 33890 -830
rect 33960 -670 34060 -650
rect 33960 -730 33980 -670
rect 34040 -730 34060 -670
rect 33960 -770 34060 -730
rect 33960 -830 33980 -770
rect 34040 -830 34060 -770
rect 33960 -850 34060 -830
rect 34130 -670 34230 -650
rect 34130 -730 34150 -670
rect 34210 -730 34230 -670
rect 34130 -770 34230 -730
rect 34130 -830 34150 -770
rect 34210 -830 34230 -770
rect 34130 -850 34230 -830
rect 34300 -670 34400 -650
rect 34300 -730 34320 -670
rect 34380 -730 34400 -670
rect 34300 -770 34400 -730
rect 34300 -830 34320 -770
rect 34380 -830 34400 -770
rect 34300 -850 34400 -830
rect 34470 -670 34570 -650
rect 34470 -730 34490 -670
rect 34550 -730 34570 -670
rect 34470 -770 34570 -730
rect 34470 -830 34490 -770
rect 34550 -830 34570 -770
rect 34470 -850 34570 -830
rect 34640 -670 34740 -650
rect 34640 -730 34660 -670
rect 34720 -730 34740 -670
rect 34640 -770 34740 -730
rect 34640 -830 34660 -770
rect 34720 -830 34740 -770
rect 34640 -850 34740 -830
rect 34810 -670 34910 -650
rect 34810 -730 34830 -670
rect 34890 -730 34910 -670
rect 34810 -770 34910 -730
rect 34810 -830 34830 -770
rect 34890 -830 34910 -770
rect 34810 -850 34910 -830
rect 34980 -670 35080 -650
rect 34980 -730 35000 -670
rect 35060 -730 35080 -670
rect 34980 -770 35080 -730
rect 34980 -830 35000 -770
rect 35060 -830 35080 -770
rect 34980 -850 35080 -830
rect 35150 -670 35250 -650
rect 35150 -730 35170 -670
rect 35230 -730 35250 -670
rect 35150 -770 35250 -730
rect 35150 -830 35170 -770
rect 35230 -830 35250 -770
rect 35150 -850 35250 -830
rect 35320 -670 35420 -650
rect 35320 -730 35340 -670
rect 35400 -730 35420 -670
rect 35320 -770 35420 -730
rect 35320 -830 35340 -770
rect 35400 -830 35420 -770
rect 35320 -850 35420 -830
rect 35490 -670 35590 -650
rect 35490 -730 35510 -670
rect 35570 -730 35590 -670
rect 35490 -770 35590 -730
rect 35490 -830 35510 -770
rect 35570 -830 35590 -770
rect 35490 -850 35590 -830
rect 35660 -670 35760 -650
rect 35660 -730 35680 -670
rect 35740 -730 35760 -670
rect 35660 -770 35760 -730
rect 35660 -830 35680 -770
rect 35740 -830 35760 -770
rect 35660 -850 35760 -830
rect 35830 -670 35930 -650
rect 35830 -730 35850 -670
rect 35910 -730 35930 -670
rect 35830 -770 35930 -730
rect 35830 -830 35850 -770
rect 35910 -830 35930 -770
rect 35830 -850 35930 -830
rect 36000 -670 36100 -650
rect 36000 -730 36020 -670
rect 36080 -730 36100 -670
rect 36000 -770 36100 -730
rect 36000 -830 36020 -770
rect 36080 -830 36100 -770
rect 36000 -850 36100 -830
rect 36170 -670 36270 -650
rect 36170 -730 36190 -670
rect 36250 -730 36270 -670
rect 36170 -770 36270 -730
rect 36170 -830 36190 -770
rect 36250 -830 36270 -770
rect 36170 -850 36270 -830
rect 36340 -670 36440 -650
rect 36340 -730 36360 -670
rect 36420 -730 36440 -670
rect 36340 -770 36440 -730
rect 36340 -830 36360 -770
rect 36420 -830 36440 -770
rect 36340 -850 36440 -830
rect 36510 -670 36610 -650
rect 36510 -730 36530 -670
rect 36590 -730 36610 -670
rect 36510 -770 36610 -730
rect 36510 -830 36530 -770
rect 36590 -830 36610 -770
rect 36510 -850 36610 -830
rect 36680 -670 36780 -650
rect 36680 -730 36700 -670
rect 36760 -730 36780 -670
rect 36680 -770 36780 -730
rect 36680 -830 36700 -770
rect 36760 -830 36780 -770
rect 36680 -850 36780 -830
rect 36850 -670 36950 -650
rect 36850 -730 36870 -670
rect 36930 -730 36950 -670
rect 36850 -770 36950 -730
rect 36850 -830 36870 -770
rect 36930 -830 36950 -770
rect 36850 -850 36950 -830
rect 37020 -670 37120 -650
rect 37020 -730 37040 -670
rect 37100 -730 37120 -670
rect 37020 -770 37120 -730
rect 37020 -830 37040 -770
rect 37100 -830 37120 -770
rect 37020 -850 37120 -830
rect 37190 -670 37290 -650
rect 37190 -730 37210 -670
rect 37270 -730 37290 -670
rect 37190 -770 37290 -730
rect 37190 -830 37210 -770
rect 37270 -830 37290 -770
rect 37190 -850 37290 -830
rect 37360 -670 37460 -650
rect 37360 -730 37380 -670
rect 37440 -730 37460 -670
rect 37360 -770 37460 -730
rect 37360 -830 37380 -770
rect 37440 -830 37460 -770
rect 37360 -850 37460 -830
rect 37530 -670 37630 -650
rect 37530 -730 37550 -670
rect 37610 -730 37630 -670
rect 37530 -770 37630 -730
rect 37530 -830 37550 -770
rect 37610 -830 37630 -770
rect 37530 -850 37630 -830
rect 37700 -670 37800 -650
rect 37700 -730 37720 -670
rect 37780 -730 37800 -670
rect 37700 -770 37800 -730
rect 37700 -830 37720 -770
rect 37780 -830 37800 -770
rect 37700 -850 37800 -830
rect 37870 -670 37970 -650
rect 37870 -730 37890 -670
rect 37950 -730 37970 -670
rect 37870 -770 37970 -730
rect 37870 -830 37890 -770
rect 37950 -830 37970 -770
rect 37870 -850 37970 -830
rect 38040 -670 38140 -650
rect 38040 -730 38060 -670
rect 38120 -730 38140 -670
rect 38040 -770 38140 -730
rect 38040 -830 38060 -770
rect 38120 -830 38140 -770
rect 38040 -850 38140 -830
rect 38210 -670 38310 -650
rect 38210 -730 38230 -670
rect 38290 -730 38310 -670
rect 38210 -770 38310 -730
rect 38210 -830 38230 -770
rect 38290 -830 38310 -770
rect 38210 -850 38310 -830
rect 38380 -670 38480 -650
rect 38380 -730 38400 -670
rect 38460 -730 38480 -670
rect 38380 -770 38480 -730
rect 38380 -830 38400 -770
rect 38460 -830 38480 -770
rect 38380 -850 38480 -830
rect 38550 -670 38650 -650
rect 38550 -730 38570 -670
rect 38630 -730 38650 -670
rect 38550 -770 38650 -730
rect 38550 -830 38570 -770
rect 38630 -830 38650 -770
rect 38550 -850 38650 -830
rect 38720 -670 38820 -650
rect 38720 -730 38740 -670
rect 38800 -730 38820 -670
rect 38720 -770 38820 -730
rect 38720 -830 38740 -770
rect 38800 -830 38820 -770
rect 38720 -850 38820 -830
rect 38890 -670 38990 -650
rect 38890 -730 38910 -670
rect 38970 -730 38990 -670
rect 38890 -770 38990 -730
rect 38890 -830 38910 -770
rect 38970 -830 38990 -770
rect 38890 -850 38990 -830
rect 39060 -670 39160 -650
rect 39060 -730 39080 -670
rect 39140 -730 39160 -670
rect 39060 -770 39160 -730
rect 39060 -830 39080 -770
rect 39140 -830 39160 -770
rect 39060 -850 39160 -830
rect 39230 -670 39330 -650
rect 39230 -730 39250 -670
rect 39310 -730 39330 -670
rect 39230 -770 39330 -730
rect 39230 -830 39250 -770
rect 39310 -830 39330 -770
rect 39230 -850 39330 -830
rect 39400 -670 39500 -650
rect 39400 -730 39420 -670
rect 39480 -730 39500 -670
rect 39400 -770 39500 -730
rect 39400 -830 39420 -770
rect 39480 -830 39500 -770
rect 39400 -850 39500 -830
rect 39570 -670 39670 -650
rect 39570 -730 39590 -670
rect 39650 -730 39670 -670
rect 39570 -770 39670 -730
rect 39570 -830 39590 -770
rect 39650 -830 39670 -770
rect 39570 -850 39670 -830
rect 39740 -670 39840 -650
rect 39740 -730 39760 -670
rect 39820 -730 39840 -670
rect 39740 -770 39840 -730
rect 39740 -830 39760 -770
rect 39820 -830 39840 -770
rect 39740 -850 39840 -830
rect 39910 -670 40010 -650
rect 39910 -730 39930 -670
rect 39990 -730 40010 -670
rect 39910 -770 40010 -730
rect 39910 -830 39930 -770
rect 39990 -830 40010 -770
rect 39910 -850 40010 -830
rect 40080 -670 40180 -650
rect 40080 -730 40100 -670
rect 40160 -730 40180 -670
rect 40080 -770 40180 -730
rect 40080 -830 40100 -770
rect 40160 -830 40180 -770
rect 40080 -850 40180 -830
rect 40250 -670 40350 -650
rect 40250 -730 40270 -670
rect 40330 -730 40350 -670
rect 40250 -770 40350 -730
rect 40250 -830 40270 -770
rect 40330 -830 40350 -770
rect 40250 -850 40350 -830
rect 40420 -670 40520 -650
rect 40420 -730 40440 -670
rect 40500 -730 40520 -670
rect 40420 -770 40520 -730
rect 40420 -830 40440 -770
rect 40500 -830 40520 -770
rect 40420 -850 40520 -830
rect 40590 -670 40690 -650
rect 40590 -730 40610 -670
rect 40670 -730 40690 -670
rect 40590 -770 40690 -730
rect 40590 -830 40610 -770
rect 40670 -830 40690 -770
rect 40590 -850 40690 -830
rect 40760 -670 40860 -650
rect 40760 -730 40780 -670
rect 40840 -730 40860 -670
rect 40760 -770 40860 -730
rect 40760 -830 40780 -770
rect 40840 -830 40860 -770
rect 40760 -850 40860 -830
rect 40930 -670 41030 -650
rect 40930 -730 40950 -670
rect 41010 -730 41030 -670
rect 40930 -770 41030 -730
rect 40930 -830 40950 -770
rect 41010 -830 41030 -770
rect 40930 -850 41030 -830
rect 41100 -670 41200 -650
rect 41100 -730 41120 -670
rect 41180 -730 41200 -670
rect 41100 -770 41200 -730
rect 41100 -830 41120 -770
rect 41180 -830 41200 -770
rect 41100 -850 41200 -830
rect 41270 -670 41370 -650
rect 41270 -730 41290 -670
rect 41350 -730 41370 -670
rect 41270 -770 41370 -730
rect 41270 -830 41290 -770
rect 41350 -830 41370 -770
rect 41270 -850 41370 -830
rect 41440 -670 41540 -650
rect 41440 -730 41460 -670
rect 41520 -730 41540 -670
rect 41440 -770 41540 -730
rect 41440 -830 41460 -770
rect 41520 -830 41540 -770
rect 41440 -850 41540 -830
rect 41610 -670 41710 -650
rect 41610 -730 41630 -670
rect 41690 -730 41710 -670
rect 41610 -770 41710 -730
rect 41610 -830 41630 -770
rect 41690 -830 41710 -770
rect 41610 -850 41710 -830
rect 41780 -670 41880 -650
rect 41780 -730 41800 -670
rect 41860 -730 41880 -670
rect 41780 -770 41880 -730
rect 41780 -830 41800 -770
rect 41860 -830 41880 -770
rect 41780 -850 41880 -830
rect 41950 -670 42050 -650
rect 41950 -730 41970 -670
rect 42030 -730 42050 -670
rect 41950 -770 42050 -730
rect 41950 -830 41970 -770
rect 42030 -830 42050 -770
rect 41950 -850 42050 -830
rect 42120 -670 42220 -650
rect 42120 -730 42140 -670
rect 42200 -730 42220 -670
rect 42120 -770 42220 -730
rect 42120 -830 42140 -770
rect 42200 -830 42220 -770
rect 42120 -850 42220 -830
rect 42290 -670 42390 -650
rect 42290 -730 42310 -670
rect 42370 -730 42390 -670
rect 42290 -770 42390 -730
rect 42290 -830 42310 -770
rect 42370 -830 42390 -770
rect 42290 -850 42390 -830
rect 42460 -670 42560 -650
rect 42460 -730 42480 -670
rect 42540 -730 42560 -670
rect 42460 -770 42560 -730
rect 42460 -830 42480 -770
rect 42540 -830 42560 -770
rect 42460 -850 42560 -830
rect 42630 -670 42730 -650
rect 42630 -730 42650 -670
rect 42710 -730 42730 -670
rect 42630 -770 42730 -730
rect 42630 -830 42650 -770
rect 42710 -830 42730 -770
rect 42630 -850 42730 -830
rect 42800 -670 42900 -650
rect 42800 -730 42820 -670
rect 42880 -730 42900 -670
rect 42800 -770 42900 -730
rect 42800 -830 42820 -770
rect 42880 -830 42900 -770
rect 42800 -850 42900 -830
rect 42970 -670 43070 -650
rect 42970 -730 42990 -670
rect 43050 -730 43070 -670
rect 42970 -770 43070 -730
rect 42970 -830 42990 -770
rect 43050 -830 43070 -770
rect 42970 -850 43070 -830
rect 43140 -670 43240 -650
rect 43140 -730 43160 -670
rect 43220 -730 43240 -670
rect 43140 -770 43240 -730
rect 43140 -830 43160 -770
rect 43220 -830 43240 -770
rect 43140 -850 43240 -830
rect 43310 -670 43410 -650
rect 43310 -730 43330 -670
rect 43390 -730 43410 -670
rect 43310 -770 43410 -730
rect 43310 -830 43330 -770
rect 43390 -830 43410 -770
rect 43310 -850 43410 -830
rect 43480 -670 43580 -650
rect 43480 -730 43500 -670
rect 43560 -730 43580 -670
rect 43480 -770 43580 -730
rect 43480 -830 43500 -770
rect 43560 -830 43580 -770
rect 43480 -850 43580 -830
rect 43650 -670 43750 -650
rect 43650 -730 43670 -670
rect 43730 -730 43750 -670
rect 43650 -770 43750 -730
rect 43650 -830 43670 -770
rect 43730 -830 43750 -770
rect 43650 -850 43750 -830
rect 43820 -670 43920 -650
rect 43820 -730 43840 -670
rect 43900 -730 43920 -670
rect 43820 -770 43920 -730
rect 43820 -830 43840 -770
rect 43900 -830 43920 -770
rect 43820 -850 43920 -830
rect 43990 -670 44090 -650
rect 43990 -730 44010 -670
rect 44070 -730 44090 -670
rect 43990 -770 44090 -730
rect 43990 -830 44010 -770
rect 44070 -830 44090 -770
rect 43990 -850 44090 -830
rect 44160 -670 44260 -650
rect 44160 -730 44180 -670
rect 44240 -730 44260 -670
rect 44160 -770 44260 -730
rect 44160 -830 44180 -770
rect 44240 -830 44260 -770
rect 44160 -850 44260 -830
rect 44330 -670 44430 -650
rect 44330 -730 44350 -670
rect 44410 -730 44430 -670
rect 44330 -770 44430 -730
rect 44330 -830 44350 -770
rect 44410 -830 44430 -770
rect 44330 -850 44430 -830
rect 44500 -670 44600 -650
rect 44500 -730 44520 -670
rect 44580 -730 44600 -670
rect 44500 -770 44600 -730
rect 44500 -830 44520 -770
rect 44580 -830 44600 -770
rect 44500 -850 44600 -830
rect 44670 -670 44770 -650
rect 44670 -730 44690 -670
rect 44750 -730 44770 -670
rect 44670 -770 44770 -730
rect 44670 -830 44690 -770
rect 44750 -830 44770 -770
rect 44670 -850 44770 -830
rect 44840 -670 44940 -650
rect 44840 -730 44860 -670
rect 44920 -730 44940 -670
rect 44840 -770 44940 -730
rect 44840 -830 44860 -770
rect 44920 -830 44940 -770
rect 44840 -850 44940 -830
rect 45010 -670 45110 -650
rect 45010 -730 45030 -670
rect 45090 -730 45110 -670
rect 45010 -770 45110 -730
rect 45010 -830 45030 -770
rect 45090 -830 45110 -770
rect 45010 -850 45110 -830
rect 45180 -670 45280 -650
rect 45180 -730 45200 -670
rect 45260 -730 45280 -670
rect 45180 -770 45280 -730
rect 45180 -830 45200 -770
rect 45260 -830 45280 -770
rect 45180 -850 45280 -830
rect 45350 -670 45450 -650
rect 45350 -730 45370 -670
rect 45430 -730 45450 -670
rect 45350 -770 45450 -730
rect 45350 -830 45370 -770
rect 45430 -830 45450 -770
rect 45350 -850 45450 -830
rect 45520 -670 45620 -650
rect 45520 -730 45540 -670
rect 45600 -730 45620 -670
rect 45520 -770 45620 -730
rect 45520 -830 45540 -770
rect 45600 -830 45620 -770
rect 45520 -850 45620 -830
rect 45690 -670 45790 -650
rect 45690 -730 45710 -670
rect 45770 -730 45790 -670
rect 45690 -770 45790 -730
rect 45690 -830 45710 -770
rect 45770 -830 45790 -770
rect 45690 -850 45790 -830
rect 45860 -670 45960 -650
rect 45860 -730 45880 -670
rect 45940 -730 45960 -670
rect 45860 -770 45960 -730
rect 45860 -830 45880 -770
rect 45940 -830 45960 -770
rect 45860 -850 45960 -830
rect 46030 -670 46130 -650
rect 46030 -730 46050 -670
rect 46110 -730 46130 -670
rect 46030 -770 46130 -730
rect 46030 -830 46050 -770
rect 46110 -830 46130 -770
rect 46030 -850 46130 -830
rect 46200 -670 46300 -650
rect 46200 -730 46220 -670
rect 46280 -730 46300 -670
rect 46200 -770 46300 -730
rect 46200 -830 46220 -770
rect 46280 -830 46300 -770
rect 46200 -850 46300 -830
rect 46370 -670 46470 -650
rect 46370 -730 46390 -670
rect 46450 -730 46470 -670
rect 46370 -770 46470 -730
rect 46370 -830 46390 -770
rect 46450 -830 46470 -770
rect 46370 -850 46470 -830
rect 46540 -670 46640 -650
rect 46540 -730 46560 -670
rect 46620 -730 46640 -670
rect 46540 -770 46640 -730
rect 46540 -830 46560 -770
rect 46620 -830 46640 -770
rect 46540 -850 46640 -830
rect 46710 -670 46810 -650
rect 46710 -730 46730 -670
rect 46790 -730 46810 -670
rect 46710 -770 46810 -730
rect 46710 -830 46730 -770
rect 46790 -830 46810 -770
rect 46710 -850 46810 -830
rect 46880 -670 46980 -650
rect 46880 -730 46900 -670
rect 46960 -730 46980 -670
rect 46880 -770 46980 -730
rect 46880 -830 46900 -770
rect 46960 -830 46980 -770
rect 46880 -850 46980 -830
rect 47050 -670 47150 -650
rect 47050 -730 47070 -670
rect 47130 -730 47150 -670
rect 47050 -770 47150 -730
rect 47050 -830 47070 -770
rect 47130 -830 47150 -770
rect 47050 -850 47150 -830
rect 47220 -670 47320 -650
rect 47220 -730 47240 -670
rect 47300 -730 47320 -670
rect 47220 -770 47320 -730
rect 47220 -830 47240 -770
rect 47300 -830 47320 -770
rect 47220 -850 47320 -830
rect 47390 -670 47490 -650
rect 47390 -730 47410 -670
rect 47470 -730 47490 -670
rect 47390 -770 47490 -730
rect 47390 -830 47410 -770
rect 47470 -830 47490 -770
rect 47390 -850 47490 -830
rect 47560 -670 47660 -650
rect 47560 -730 47580 -670
rect 47640 -730 47660 -670
rect 47560 -770 47660 -730
rect 47560 -830 47580 -770
rect 47640 -830 47660 -770
rect 47560 -850 47660 -830
rect 47730 -670 47830 -650
rect 47730 -730 47750 -670
rect 47810 -730 47830 -670
rect 47730 -770 47830 -730
rect 47730 -830 47750 -770
rect 47810 -830 47830 -770
rect 47730 -850 47830 -830
rect 47900 -670 48000 -650
rect 47900 -730 47920 -670
rect 47980 -730 48000 -670
rect 47900 -770 48000 -730
rect 47900 -830 47920 -770
rect 47980 -830 48000 -770
rect 47900 -850 48000 -830
rect 48070 -670 48170 -650
rect 48070 -730 48090 -670
rect 48150 -730 48170 -670
rect 48070 -770 48170 -730
rect 48070 -830 48090 -770
rect 48150 -830 48170 -770
rect 48070 -850 48170 -830
rect 48240 -670 48340 -650
rect 48240 -730 48260 -670
rect 48320 -730 48340 -670
rect 48240 -770 48340 -730
rect 48240 -830 48260 -770
rect 48320 -830 48340 -770
rect 48240 -850 48340 -830
rect 48410 -670 48510 -650
rect 48410 -730 48430 -670
rect 48490 -730 48510 -670
rect 48410 -770 48510 -730
rect 48410 -830 48430 -770
rect 48490 -830 48510 -770
rect 48410 -850 48510 -830
rect 48580 -670 48680 -650
rect 48580 -730 48600 -670
rect 48660 -730 48680 -670
rect 48580 -770 48680 -730
rect 48580 -830 48600 -770
rect 48660 -830 48680 -770
rect 48580 -850 48680 -830
rect 48750 -670 48850 -650
rect 48750 -730 48770 -670
rect 48830 -730 48850 -670
rect 48750 -770 48850 -730
rect 48750 -830 48770 -770
rect 48830 -830 48850 -770
rect 48750 -850 48850 -830
rect 48920 -670 49020 -650
rect 48920 -730 48940 -670
rect 49000 -730 49020 -670
rect 48920 -770 49020 -730
rect 48920 -830 48940 -770
rect 49000 -830 49020 -770
rect 48920 -850 49020 -830
rect 49090 -670 49190 -650
rect 49090 -730 49110 -670
rect 49170 -730 49190 -670
rect 49090 -770 49190 -730
rect 49090 -830 49110 -770
rect 49170 -830 49190 -770
rect 49090 -850 49190 -830
rect 49260 -670 49360 -650
rect 49260 -730 49280 -670
rect 49340 -730 49360 -670
rect 49260 -770 49360 -730
rect 49260 -830 49280 -770
rect 49340 -830 49360 -770
rect 49260 -850 49360 -830
rect 49430 -670 49530 -650
rect 49430 -730 49450 -670
rect 49510 -730 49530 -670
rect 49430 -770 49530 -730
rect 49430 -830 49450 -770
rect 49510 -830 49530 -770
rect 49430 -850 49530 -830
rect 49600 -670 49700 -650
rect 49600 -730 49620 -670
rect 49680 -730 49700 -670
rect 49600 -770 49700 -730
rect 49600 -830 49620 -770
rect 49680 -830 49700 -770
rect 49600 -850 49700 -830
rect 49770 -670 49870 -650
rect 49770 -730 49790 -670
rect 49850 -730 49870 -670
rect 49770 -770 49870 -730
rect 49770 -830 49790 -770
rect 49850 -830 49870 -770
rect 49770 -850 49870 -830
rect 49940 -670 50040 -650
rect 49940 -730 49960 -670
rect 50020 -730 50040 -670
rect 49940 -770 50040 -730
rect 49940 -830 49960 -770
rect 50020 -830 50040 -770
rect 49940 -850 50040 -830
rect 50110 -670 50210 -650
rect 50110 -730 50130 -670
rect 50190 -730 50210 -670
rect 50110 -770 50210 -730
rect 50110 -830 50130 -770
rect 50190 -830 50210 -770
rect 50110 -850 50210 -830
rect 50280 -670 50380 -650
rect 50280 -730 50300 -670
rect 50360 -730 50380 -670
rect 50280 -770 50380 -730
rect 50280 -830 50300 -770
rect 50360 -830 50380 -770
rect 50280 -850 50380 -830
rect 50450 -670 50550 -650
rect 50450 -730 50470 -670
rect 50530 -730 50550 -670
rect 50450 -770 50550 -730
rect 50450 -830 50470 -770
rect 50530 -830 50550 -770
rect 50450 -850 50550 -830
rect 50620 -670 50720 -650
rect 50620 -730 50640 -670
rect 50700 -730 50720 -670
rect 50620 -770 50720 -730
rect 50620 -830 50640 -770
rect 50700 -830 50720 -770
rect 50620 -850 50720 -830
rect 50790 -670 50890 -650
rect 50790 -730 50810 -670
rect 50870 -730 50890 -670
rect 50790 -770 50890 -730
rect 50790 -830 50810 -770
rect 50870 -830 50890 -770
rect 50790 -850 50890 -830
rect 50960 -670 51060 -650
rect 50960 -730 50980 -670
rect 51040 -730 51060 -670
rect 50960 -770 51060 -730
rect 50960 -830 50980 -770
rect 51040 -830 51060 -770
rect 50960 -850 51060 -830
rect 51130 -670 51230 -650
rect 51130 -730 51150 -670
rect 51210 -730 51230 -670
rect 51130 -770 51230 -730
rect 51130 -830 51150 -770
rect 51210 -830 51230 -770
rect 51130 -850 51230 -830
rect 51300 -670 51400 -650
rect 51300 -730 51320 -670
rect 51380 -730 51400 -670
rect 51300 -770 51400 -730
rect 51300 -830 51320 -770
rect 51380 -830 51400 -770
rect 51300 -850 51400 -830
rect 51470 -670 51570 -650
rect 51470 -730 51490 -670
rect 51550 -730 51570 -670
rect 51470 -770 51570 -730
rect 51470 -830 51490 -770
rect 51550 -830 51570 -770
rect 51470 -850 51570 -830
rect 51640 -670 51740 -650
rect 51640 -730 51660 -670
rect 51720 -730 51740 -670
rect 51640 -770 51740 -730
rect 51640 -830 51660 -770
rect 51720 -830 51740 -770
rect 51640 -850 51740 -830
rect 51810 -670 51910 -650
rect 51810 -730 51830 -670
rect 51890 -730 51910 -670
rect 51810 -770 51910 -730
rect 51810 -830 51830 -770
rect 51890 -830 51910 -770
rect 51810 -850 51910 -830
rect 51980 -670 52080 -650
rect 51980 -730 52000 -670
rect 52060 -730 52080 -670
rect 51980 -770 52080 -730
rect 51980 -830 52000 -770
rect 52060 -830 52080 -770
rect 51980 -850 52080 -830
rect 52150 -670 52250 -650
rect 52150 -730 52170 -670
rect 52230 -730 52250 -670
rect 52150 -770 52250 -730
rect 52150 -830 52170 -770
rect 52230 -830 52250 -770
rect 52150 -850 52250 -830
rect 52320 -670 52420 -650
rect 52320 -730 52340 -670
rect 52400 -730 52420 -670
rect 52320 -770 52420 -730
rect 52320 -830 52340 -770
rect 52400 -830 52420 -770
rect 52320 -850 52420 -830
rect 52490 -670 52590 -650
rect 52490 -730 52510 -670
rect 52570 -730 52590 -670
rect 52490 -770 52590 -730
rect 52490 -830 52510 -770
rect 52570 -830 52590 -770
rect 52490 -850 52590 -830
rect 52660 -670 52760 -650
rect 52660 -730 52680 -670
rect 52740 -730 52760 -670
rect 52660 -770 52760 -730
rect 52660 -830 52680 -770
rect 52740 -830 52760 -770
rect 52660 -850 52760 -830
rect 52830 -670 52930 -650
rect 52830 -730 52850 -670
rect 52910 -730 52930 -670
rect 52830 -770 52930 -730
rect 52830 -830 52850 -770
rect 52910 -830 52930 -770
rect 52830 -850 52930 -830
rect 53000 -670 53100 -650
rect 53000 -730 53020 -670
rect 53080 -730 53100 -670
rect 53000 -770 53100 -730
rect 53000 -830 53020 -770
rect 53080 -830 53100 -770
rect 53000 -850 53100 -830
rect 53170 -670 53270 -650
rect 53170 -730 53190 -670
rect 53250 -730 53270 -670
rect 53170 -770 53270 -730
rect 53170 -830 53190 -770
rect 53250 -830 53270 -770
rect 53170 -850 53270 -830
rect 53340 -670 53440 -650
rect 53340 -730 53360 -670
rect 53420 -730 53440 -670
rect 53340 -770 53440 -730
rect 53340 -830 53360 -770
rect 53420 -830 53440 -770
rect 53340 -850 53440 -830
rect 53510 -670 53610 -650
rect 53510 -730 53530 -670
rect 53590 -730 53610 -670
rect 53510 -770 53610 -730
rect 53510 -830 53530 -770
rect 53590 -830 53610 -770
rect 53510 -850 53610 -830
rect 53680 -670 53780 -650
rect 53680 -730 53700 -670
rect 53760 -730 53780 -670
rect 53680 -770 53780 -730
rect 53680 -830 53700 -770
rect 53760 -830 53780 -770
rect 53680 -850 53780 -830
rect 53850 -670 53950 -650
rect 53850 -730 53870 -670
rect 53930 -730 53950 -670
rect 53850 -770 53950 -730
rect 53850 -830 53870 -770
rect 53930 -830 53950 -770
rect 53850 -850 53950 -830
rect 54020 -670 54120 -650
rect 54020 -730 54040 -670
rect 54100 -730 54120 -670
rect 54020 -770 54120 -730
rect 54020 -830 54040 -770
rect 54100 -830 54120 -770
rect 54020 -850 54120 -830
rect 54190 -670 54290 -650
rect 54190 -730 54210 -670
rect 54270 -730 54290 -670
rect 54190 -770 54290 -730
rect 54190 -830 54210 -770
rect 54270 -830 54290 -770
rect 54190 -850 54290 -830
rect 54360 -670 54460 -650
rect 54360 -730 54380 -670
rect 54440 -730 54460 -670
rect 54360 -770 54460 -730
rect 54360 -830 54380 -770
rect 54440 -830 54460 -770
rect 54360 -850 54460 -830
rect 54530 -670 54630 -650
rect 54530 -730 54550 -670
rect 54610 -730 54630 -670
rect 54530 -770 54630 -730
rect 54530 -830 54550 -770
rect 54610 -830 54630 -770
rect 54530 -850 54630 -830
rect 54700 -670 54800 -650
rect 54700 -730 54720 -670
rect 54780 -730 54800 -670
rect 54700 -770 54800 -730
rect 54700 -830 54720 -770
rect 54780 -830 54800 -770
rect 54700 -850 54800 -830
rect 54870 -670 54970 -650
rect 54870 -730 54890 -670
rect 54950 -730 54970 -670
rect 54870 -770 54970 -730
rect 54870 -830 54890 -770
rect 54950 -830 54970 -770
rect 54870 -850 54970 -830
rect 55040 -670 55140 -650
rect 55040 -730 55060 -670
rect 55120 -730 55140 -670
rect 55040 -770 55140 -730
rect 55040 -830 55060 -770
rect 55120 -830 55140 -770
rect 55040 -850 55140 -830
rect 55210 -670 55310 -650
rect 55210 -730 55230 -670
rect 55290 -730 55310 -670
rect 55210 -770 55310 -730
rect 55210 -830 55230 -770
rect 55290 -830 55310 -770
rect 55210 -850 55310 -830
rect 55380 -670 55480 -650
rect 55380 -730 55400 -670
rect 55460 -730 55480 -670
rect 55380 -770 55480 -730
rect 55380 -830 55400 -770
rect 55460 -830 55480 -770
rect 55380 -850 55480 -830
rect 55550 -670 55650 -650
rect 55550 -730 55570 -670
rect 55630 -730 55650 -670
rect 55550 -770 55650 -730
rect 55550 -830 55570 -770
rect 55630 -830 55650 -770
rect 55550 -850 55650 -830
rect 55720 -670 55820 -650
rect 55720 -730 55740 -670
rect 55800 -730 55820 -670
rect 55720 -770 55820 -730
rect 55720 -830 55740 -770
rect 55800 -830 55820 -770
rect 55720 -850 55820 -830
rect 55890 -670 55990 -650
rect 55890 -730 55910 -670
rect 55970 -730 55990 -670
rect 55890 -770 55990 -730
rect 55890 -830 55910 -770
rect 55970 -830 55990 -770
rect 55890 -850 55990 -830
rect 56060 -670 56160 -650
rect 56060 -730 56080 -670
rect 56140 -730 56160 -670
rect 56060 -770 56160 -730
rect 56060 -830 56080 -770
rect 56140 -830 56160 -770
rect 56060 -850 56160 -830
rect 56230 -670 56330 -650
rect 56230 -730 56250 -670
rect 56310 -730 56330 -670
rect 56230 -770 56330 -730
rect 56230 -830 56250 -770
rect 56310 -830 56330 -770
rect 56230 -850 56330 -830
rect 56400 -670 56500 -650
rect 56400 -730 56420 -670
rect 56480 -730 56500 -670
rect 56400 -770 56500 -730
rect 56400 -830 56420 -770
rect 56480 -830 56500 -770
rect 56400 -850 56500 -830
rect 56570 -670 56670 -650
rect 56570 -730 56590 -670
rect 56650 -730 56670 -670
rect 56570 -770 56670 -730
rect 56570 -830 56590 -770
rect 56650 -830 56670 -770
rect 56570 -850 56670 -830
rect 56740 -670 56840 -650
rect 56740 -730 56760 -670
rect 56820 -730 56840 -670
rect 56740 -770 56840 -730
rect 56740 -830 56760 -770
rect 56820 -830 56840 -770
rect 56740 -850 56840 -830
rect 56910 -670 57010 -650
rect 56910 -730 56930 -670
rect 56990 -730 57010 -670
rect 56910 -770 57010 -730
rect 56910 -830 56930 -770
rect 56990 -830 57010 -770
rect 56910 -850 57010 -830
rect 57080 -670 57180 -650
rect 57080 -730 57100 -670
rect 57160 -730 57180 -670
rect 57080 -770 57180 -730
rect 57080 -830 57100 -770
rect 57160 -830 57180 -770
rect 57080 -850 57180 -830
rect 57250 -670 57350 -650
rect 57250 -730 57270 -670
rect 57330 -730 57350 -670
rect 57250 -770 57350 -730
rect 57250 -830 57270 -770
rect 57330 -830 57350 -770
rect 57250 -850 57350 -830
rect 57420 -670 57520 -650
rect 57420 -730 57440 -670
rect 57500 -730 57520 -670
rect 57420 -770 57520 -730
rect 57420 -830 57440 -770
rect 57500 -830 57520 -770
rect 57420 -850 57520 -830
rect 57590 -670 57690 -650
rect 57590 -730 57610 -670
rect 57670 -730 57690 -670
rect 57590 -770 57690 -730
rect 57590 -830 57610 -770
rect 57670 -830 57690 -770
rect 57590 -850 57690 -830
rect 57760 -670 57860 -650
rect 57760 -730 57780 -670
rect 57840 -730 57860 -670
rect 57760 -770 57860 -730
rect 57760 -830 57780 -770
rect 57840 -830 57860 -770
rect 57760 -850 57860 -830
rect 57930 -670 58030 -650
rect 57930 -730 57950 -670
rect 58010 -730 58030 -670
rect 57930 -770 58030 -730
rect 57930 -830 57950 -770
rect 58010 -830 58030 -770
rect 57930 -850 58030 -830
rect 58100 -670 58200 -650
rect 58100 -730 58120 -670
rect 58180 -730 58200 -670
rect 58100 -770 58200 -730
rect 58100 -830 58120 -770
rect 58180 -830 58200 -770
rect 58100 -850 58200 -830
rect 58270 -670 58370 -650
rect 58270 -730 58290 -670
rect 58350 -730 58370 -670
rect 58270 -770 58370 -730
rect 58270 -830 58290 -770
rect 58350 -830 58370 -770
rect 58270 -850 58370 -830
rect 58440 -670 58540 -650
rect 58440 -730 58460 -670
rect 58520 -730 58540 -670
rect 58440 -770 58540 -730
rect 58440 -830 58460 -770
rect 58520 -830 58540 -770
rect 58440 -850 58540 -830
rect 58610 -670 58710 -650
rect 58610 -730 58630 -670
rect 58690 -730 58710 -670
rect 58610 -770 58710 -730
rect 58610 -830 58630 -770
rect 58690 -830 58710 -770
rect 58610 -850 58710 -830
rect 58780 -670 58880 -650
rect 58780 -730 58800 -670
rect 58860 -730 58880 -670
rect 58780 -770 58880 -730
rect 58780 -830 58800 -770
rect 58860 -830 58880 -770
rect 58780 -850 58880 -830
rect 58950 -670 59050 -650
rect 58950 -730 58970 -670
rect 59030 -730 59050 -670
rect 58950 -770 59050 -730
rect 58950 -830 58970 -770
rect 59030 -830 59050 -770
rect 58950 -850 59050 -830
rect 59120 -670 59220 -650
rect 59120 -730 59140 -670
rect 59200 -730 59220 -670
rect 59120 -770 59220 -730
rect 59120 -830 59140 -770
rect 59200 -830 59220 -770
rect 59120 -850 59220 -830
rect 59290 -670 59390 -650
rect 59290 -730 59310 -670
rect 59370 -730 59390 -670
rect 59290 -770 59390 -730
rect 59290 -830 59310 -770
rect 59370 -830 59390 -770
rect 59290 -850 59390 -830
rect 59460 -670 59560 -650
rect 59460 -730 59480 -670
rect 59540 -730 59560 -670
rect 59460 -770 59560 -730
rect 59460 -830 59480 -770
rect 59540 -830 59560 -770
rect 59460 -850 59560 -830
rect 59630 -670 59730 -650
rect 59630 -730 59650 -670
rect 59710 -730 59730 -670
rect 59630 -770 59730 -730
rect 59630 -830 59650 -770
rect 59710 -830 59730 -770
rect 59630 -850 59730 -830
rect 59800 -670 59900 -650
rect 59800 -730 59820 -670
rect 59880 -730 59900 -670
rect 59800 -770 59900 -730
rect 59800 -830 59820 -770
rect 59880 -830 59900 -770
rect 59800 -850 59900 -830
rect 59970 -670 60070 -650
rect 59970 -730 59990 -670
rect 60050 -730 60070 -670
rect 59970 -770 60070 -730
rect 59970 -830 59990 -770
rect 60050 -830 60070 -770
rect 59970 -850 60070 -830
rect 60140 -670 60240 -650
rect 60140 -730 60160 -670
rect 60220 -730 60240 -670
rect 60140 -770 60240 -730
rect 60140 -830 60160 -770
rect 60220 -830 60240 -770
rect 60140 -850 60240 -830
rect 60310 -670 60410 -650
rect 60310 -730 60330 -670
rect 60390 -730 60410 -670
rect 60310 -770 60410 -730
rect 60310 -830 60330 -770
rect 60390 -830 60410 -770
rect 60310 -850 60410 -830
rect 60480 -670 60580 -650
rect 60480 -730 60500 -670
rect 60560 -730 60580 -670
rect 60480 -770 60580 -730
rect 60480 -830 60500 -770
rect 60560 -830 60580 -770
rect 60480 -850 60580 -830
rect 60650 -670 60750 -650
rect 60650 -730 60670 -670
rect 60730 -730 60750 -670
rect 60650 -770 60750 -730
rect 60650 -830 60670 -770
rect 60730 -830 60750 -770
rect 60650 -850 60750 -830
rect 60820 -670 60920 -650
rect 60820 -730 60840 -670
rect 60900 -730 60920 -670
rect 60820 -770 60920 -730
rect 60820 -830 60840 -770
rect 60900 -830 60920 -770
rect 60820 -850 60920 -830
rect 60990 -670 61090 -650
rect 60990 -730 61010 -670
rect 61070 -730 61090 -670
rect 60990 -770 61090 -730
rect 60990 -830 61010 -770
rect 61070 -830 61090 -770
rect 60990 -850 61090 -830
rect 61160 -670 61260 -650
rect 61160 -730 61180 -670
rect 61240 -730 61260 -670
rect 61160 -770 61260 -730
rect 61160 -830 61180 -770
rect 61240 -830 61260 -770
rect 61160 -850 61260 -830
rect 61330 -670 61430 -650
rect 61330 -730 61350 -670
rect 61410 -730 61430 -670
rect 61330 -770 61430 -730
rect 61330 -830 61350 -770
rect 61410 -830 61430 -770
rect 61330 -850 61430 -830
rect 61500 -670 61600 -650
rect 61500 -730 61520 -670
rect 61580 -730 61600 -670
rect 61500 -770 61600 -730
rect 61500 -830 61520 -770
rect 61580 -830 61600 -770
rect 61500 -850 61600 -830
rect 61670 -670 61770 -650
rect 61670 -730 61690 -670
rect 61750 -730 61770 -670
rect 61670 -770 61770 -730
rect 61670 -830 61690 -770
rect 61750 -830 61770 -770
rect 61670 -850 61770 -830
rect 61840 -670 61940 -650
rect 61840 -730 61860 -670
rect 61920 -730 61940 -670
rect 61840 -770 61940 -730
rect 61840 -830 61860 -770
rect 61920 -830 61940 -770
rect 61840 -850 61940 -830
rect 62010 -670 62110 -650
rect 62010 -730 62030 -670
rect 62090 -730 62110 -670
rect 62010 -770 62110 -730
rect 62010 -830 62030 -770
rect 62090 -830 62110 -770
rect 62010 -850 62110 -830
rect 62180 -670 62280 -650
rect 62180 -730 62200 -670
rect 62260 -730 62280 -670
rect 62180 -770 62280 -730
rect 62180 -830 62200 -770
rect 62260 -830 62280 -770
rect 62180 -850 62280 -830
rect 62350 -670 62450 -650
rect 62350 -730 62370 -670
rect 62430 -730 62450 -670
rect 62350 -770 62450 -730
rect 62350 -830 62370 -770
rect 62430 -830 62450 -770
rect 62350 -850 62450 -830
rect 62520 -670 62620 -650
rect 62520 -730 62540 -670
rect 62600 -730 62620 -670
rect 62520 -770 62620 -730
rect 62520 -830 62540 -770
rect 62600 -830 62620 -770
rect 62520 -850 62620 -830
rect 62690 -670 62790 -650
rect 62690 -730 62710 -670
rect 62770 -730 62790 -670
rect 62690 -770 62790 -730
rect 62690 -830 62710 -770
rect 62770 -830 62790 -770
rect 62690 -850 62790 -830
rect 62860 -670 62960 -650
rect 62860 -730 62880 -670
rect 62940 -730 62960 -670
rect 62860 -770 62960 -730
rect 62860 -830 62880 -770
rect 62940 -830 62960 -770
rect 62860 -850 62960 -830
rect 63030 -670 63130 -650
rect 63030 -730 63050 -670
rect 63110 -730 63130 -670
rect 63030 -770 63130 -730
rect 63030 -830 63050 -770
rect 63110 -830 63130 -770
rect 63030 -850 63130 -830
rect 63200 -670 63300 -650
rect 63200 -730 63220 -670
rect 63280 -730 63300 -670
rect 63200 -770 63300 -730
rect 63200 -830 63220 -770
rect 63280 -830 63300 -770
rect 63200 -850 63300 -830
rect 63370 -670 63470 -650
rect 63370 -730 63390 -670
rect 63450 -730 63470 -670
rect 63370 -770 63470 -730
rect 63370 -830 63390 -770
rect 63450 -830 63470 -770
rect 63370 -850 63470 -830
rect 63540 -670 63640 -650
rect 63540 -730 63560 -670
rect 63620 -730 63640 -670
rect 63540 -770 63640 -730
rect 63540 -830 63560 -770
rect 63620 -830 63640 -770
rect 63540 -850 63640 -830
rect 63710 -670 63810 -650
rect 63710 -730 63730 -670
rect 63790 -730 63810 -670
rect 63710 -770 63810 -730
rect 63710 -830 63730 -770
rect 63790 -830 63810 -770
rect 63710 -850 63810 -830
rect 63880 -670 63980 -650
rect 63880 -730 63900 -670
rect 63960 -730 63980 -670
rect 63880 -770 63980 -730
rect 63880 -830 63900 -770
rect 63960 -830 63980 -770
rect 63880 -850 63980 -830
rect 64050 -670 64150 -650
rect 64050 -730 64070 -670
rect 64130 -730 64150 -670
rect 64050 -770 64150 -730
rect 64050 -830 64070 -770
rect 64130 -830 64150 -770
rect 64050 -850 64150 -830
rect 64220 -670 64320 -650
rect 64220 -730 64240 -670
rect 64300 -730 64320 -670
rect 64220 -770 64320 -730
rect 64220 -830 64240 -770
rect 64300 -830 64320 -770
rect 64220 -850 64320 -830
rect 64390 -670 64490 -650
rect 64390 -730 64410 -670
rect 64470 -730 64490 -670
rect 64390 -770 64490 -730
rect 64390 -830 64410 -770
rect 64470 -830 64490 -770
rect 64390 -850 64490 -830
rect 64560 -670 64660 -650
rect 64560 -730 64580 -670
rect 64640 -730 64660 -670
rect 64560 -770 64660 -730
rect 64560 -830 64580 -770
rect 64640 -830 64660 -770
rect 64560 -850 64660 -830
rect 64730 -670 64830 -650
rect 64730 -730 64750 -670
rect 64810 -730 64830 -670
rect 64730 -770 64830 -730
rect 64730 -830 64750 -770
rect 64810 -830 64830 -770
rect 64730 -850 64830 -830
rect 64900 -670 65000 -650
rect 64900 -730 64920 -670
rect 64980 -730 65000 -670
rect 64900 -770 65000 -730
rect 64900 -830 64920 -770
rect 64980 -830 65000 -770
rect 64900 -850 65000 -830
rect 65070 -670 65170 -650
rect 65070 -730 65090 -670
rect 65150 -730 65170 -670
rect 65070 -770 65170 -730
rect 65070 -830 65090 -770
rect 65150 -830 65170 -770
rect 65070 -850 65170 -830
rect 65240 -670 65340 -650
rect 65240 -730 65260 -670
rect 65320 -730 65340 -670
rect 65240 -770 65340 -730
rect 65240 -830 65260 -770
rect 65320 -830 65340 -770
rect 65240 -850 65340 -830
rect 65410 -670 65510 -650
rect 65410 -730 65430 -670
rect 65490 -730 65510 -670
rect 65410 -770 65510 -730
rect 65410 -830 65430 -770
rect 65490 -830 65510 -770
rect 65410 -850 65510 -830
rect 65580 -670 65680 -650
rect 65580 -730 65600 -670
rect 65660 -730 65680 -670
rect 65580 -770 65680 -730
rect 65580 -830 65600 -770
rect 65660 -830 65680 -770
rect 65580 -850 65680 -830
rect 65750 -670 65850 -650
rect 65750 -730 65770 -670
rect 65830 -730 65850 -670
rect 65750 -770 65850 -730
rect 65750 -830 65770 -770
rect 65830 -830 65850 -770
rect 65750 -850 65850 -830
rect 65920 -670 66020 -650
rect 65920 -730 65940 -670
rect 66000 -730 66020 -670
rect 65920 -770 66020 -730
rect 65920 -830 65940 -770
rect 66000 -830 66020 -770
rect 65920 -850 66020 -830
rect 66090 -670 66190 -650
rect 66090 -730 66110 -670
rect 66170 -730 66190 -670
rect 66090 -770 66190 -730
rect 66090 -830 66110 -770
rect 66170 -830 66190 -770
rect 66090 -850 66190 -830
rect 66260 -670 66360 -650
rect 66260 -730 66280 -670
rect 66340 -730 66360 -670
rect 66260 -770 66360 -730
rect 66260 -830 66280 -770
rect 66340 -830 66360 -770
rect 66260 -850 66360 -830
rect 66430 -670 66530 -650
rect 66430 -730 66450 -670
rect 66510 -730 66530 -670
rect 66430 -770 66530 -730
rect 66430 -830 66450 -770
rect 66510 -830 66530 -770
rect 66430 -850 66530 -830
rect 66600 -670 66700 -650
rect 66600 -730 66620 -670
rect 66680 -730 66700 -670
rect 66600 -770 66700 -730
rect 66600 -830 66620 -770
rect 66680 -830 66700 -770
rect 66600 -850 66700 -830
rect 66770 -670 66870 -650
rect 66770 -730 66790 -670
rect 66850 -730 66870 -670
rect 66770 -770 66870 -730
rect 66770 -830 66790 -770
rect 66850 -830 66870 -770
rect 66770 -850 66870 -830
rect 66940 -670 67040 -650
rect 66940 -730 66960 -670
rect 67020 -730 67040 -670
rect 66940 -770 67040 -730
rect 66940 -830 66960 -770
rect 67020 -830 67040 -770
rect 66940 -850 67040 -830
rect 67110 -670 67210 -650
rect 67110 -730 67130 -670
rect 67190 -730 67210 -670
rect 67110 -770 67210 -730
rect 67110 -830 67130 -770
rect 67190 -830 67210 -770
rect 67110 -850 67210 -830
rect 67280 -670 67380 -650
rect 67280 -730 67300 -670
rect 67360 -730 67380 -670
rect 67280 -770 67380 -730
rect 67280 -830 67300 -770
rect 67360 -830 67380 -770
rect 67280 -850 67380 -830
rect 67450 -670 67550 -650
rect 67450 -730 67470 -670
rect 67530 -730 67550 -670
rect 67450 -770 67550 -730
rect 67450 -830 67470 -770
rect 67530 -830 67550 -770
rect 67450 -850 67550 -830
rect 67620 -670 67720 -650
rect 67620 -730 67640 -670
rect 67700 -730 67720 -670
rect 67620 -770 67720 -730
rect 67620 -830 67640 -770
rect 67700 -830 67720 -770
rect 67620 -850 67720 -830
rect 67790 -670 67890 -650
rect 67790 -730 67810 -670
rect 67870 -730 67890 -670
rect 67790 -770 67890 -730
rect 67790 -830 67810 -770
rect 67870 -830 67890 -770
rect 67790 -850 67890 -830
rect 67960 -670 68060 -650
rect 67960 -730 67980 -670
rect 68040 -730 68060 -670
rect 67960 -770 68060 -730
rect 67960 -830 67980 -770
rect 68040 -830 68060 -770
rect 67960 -850 68060 -830
rect 68130 -670 68230 -650
rect 68130 -730 68150 -670
rect 68210 -730 68230 -670
rect 68130 -770 68230 -730
rect 68130 -830 68150 -770
rect 68210 -830 68230 -770
rect 68130 -850 68230 -830
rect 68300 -670 68400 -650
rect 68300 -730 68320 -670
rect 68380 -730 68400 -670
rect 68300 -770 68400 -730
rect 68300 -830 68320 -770
rect 68380 -830 68400 -770
rect 68300 -850 68400 -830
rect 68470 -670 68570 -650
rect 68470 -730 68490 -670
rect 68550 -730 68570 -670
rect 68470 -770 68570 -730
rect 68470 -830 68490 -770
rect 68550 -830 68570 -770
rect 68470 -850 68570 -830
rect 68640 -670 68740 -650
rect 68640 -730 68660 -670
rect 68720 -730 68740 -670
rect 68640 -770 68740 -730
rect 68640 -830 68660 -770
rect 68720 -830 68740 -770
rect 68640 -850 68740 -830
rect 68810 -670 68910 -650
rect 68810 -730 68830 -670
rect 68890 -730 68910 -670
rect 68810 -770 68910 -730
rect 68810 -830 68830 -770
rect 68890 -830 68910 -770
rect 68810 -850 68910 -830
rect 68980 -670 69080 -650
rect 68980 -730 69000 -670
rect 69060 -730 69080 -670
rect 68980 -770 69080 -730
rect 68980 -830 69000 -770
rect 69060 -830 69080 -770
rect 68980 -850 69080 -830
rect 69150 -670 69250 -650
rect 69150 -730 69170 -670
rect 69230 -730 69250 -670
rect 69150 -770 69250 -730
rect 69150 -830 69170 -770
rect 69230 -830 69250 -770
rect 69150 -850 69250 -830
rect 69320 -670 69420 -650
rect 69320 -730 69340 -670
rect 69400 -730 69420 -670
rect 69320 -770 69420 -730
rect 69320 -830 69340 -770
rect 69400 -830 69420 -770
rect 69320 -850 69420 -830
rect 69490 -670 69590 -650
rect 69490 -730 69510 -670
rect 69570 -730 69590 -670
rect 69490 -770 69590 -730
rect 69490 -830 69510 -770
rect 69570 -830 69590 -770
rect 69490 -850 69590 -830
rect 69660 -670 69760 -650
rect 69660 -730 69680 -670
rect 69740 -730 69760 -670
rect 69660 -770 69760 -730
rect 69660 -830 69680 -770
rect 69740 -830 69760 -770
rect 69660 -850 69760 -830
rect 69830 -670 69930 -650
rect 69830 -730 69850 -670
rect 69910 -730 69930 -670
rect 69830 -770 69930 -730
rect 69830 -830 69850 -770
rect 69910 -830 69930 -770
rect 69830 -850 69930 -830
rect 70000 -670 70100 -650
rect 70000 -730 70020 -670
rect 70080 -730 70100 -670
rect 70000 -770 70100 -730
rect 70000 -830 70020 -770
rect 70080 -830 70100 -770
rect 70000 -850 70100 -830
rect 70170 -670 70270 -650
rect 70170 -730 70190 -670
rect 70250 -730 70270 -670
rect 70170 -770 70270 -730
rect 70170 -830 70190 -770
rect 70250 -830 70270 -770
rect 70170 -850 70270 -830
rect 70340 -670 70440 -650
rect 70340 -730 70360 -670
rect 70420 -730 70440 -670
rect 70340 -770 70440 -730
rect 70340 -830 70360 -770
rect 70420 -830 70440 -770
rect 70340 -850 70440 -830
rect 70510 -670 70610 -650
rect 70510 -730 70530 -670
rect 70590 -730 70610 -670
rect 70510 -770 70610 -730
rect 70510 -830 70530 -770
rect 70590 -830 70610 -770
rect 70510 -850 70610 -830
rect 70680 -670 70780 -650
rect 70680 -730 70700 -670
rect 70760 -730 70780 -670
rect 70680 -770 70780 -730
rect 70680 -830 70700 -770
rect 70760 -830 70780 -770
rect 70680 -850 70780 -830
rect 70850 -670 70950 -650
rect 70850 -730 70870 -670
rect 70930 -730 70950 -670
rect 70850 -770 70950 -730
rect 70850 -830 70870 -770
rect 70930 -830 70950 -770
rect 70850 -850 70950 -830
rect 71020 -670 71120 -650
rect 71020 -730 71040 -670
rect 71100 -730 71120 -670
rect 71020 -770 71120 -730
rect 71020 -830 71040 -770
rect 71100 -830 71120 -770
rect 71020 -850 71120 -830
rect 71190 -670 71290 -650
rect 71190 -730 71210 -670
rect 71270 -730 71290 -670
rect 71190 -770 71290 -730
rect 71190 -830 71210 -770
rect 71270 -830 71290 -770
rect 71190 -850 71290 -830
rect 71360 -670 71460 -650
rect 71360 -730 71380 -670
rect 71440 -730 71460 -670
rect 71360 -770 71460 -730
rect 71360 -830 71380 -770
rect 71440 -830 71460 -770
rect 71360 -850 71460 -830
rect 71530 -670 71630 -650
rect 71530 -730 71550 -670
rect 71610 -730 71630 -670
rect 71530 -770 71630 -730
rect 71530 -830 71550 -770
rect 71610 -830 71630 -770
rect 71530 -850 71630 -830
rect 71700 -670 71800 -650
rect 71700 -730 71720 -670
rect 71780 -730 71800 -670
rect 71700 -770 71800 -730
rect 71700 -830 71720 -770
rect 71780 -830 71800 -770
rect 71700 -850 71800 -830
rect 71870 -670 71970 -650
rect 71870 -730 71890 -670
rect 71950 -730 71970 -670
rect 71870 -770 71970 -730
rect 71870 -830 71890 -770
rect 71950 -830 71970 -770
rect 71870 -850 71970 -830
rect 72040 -670 72140 -650
rect 72040 -730 72060 -670
rect 72120 -730 72140 -670
rect 72040 -770 72140 -730
rect 72040 -830 72060 -770
rect 72120 -830 72140 -770
rect 72040 -850 72140 -830
rect 72210 -670 72310 -650
rect 72210 -730 72230 -670
rect 72290 -730 72310 -670
rect 72210 -770 72310 -730
rect 72210 -830 72230 -770
rect 72290 -830 72310 -770
rect 72210 -850 72310 -830
rect 72380 -670 72480 -650
rect 72380 -730 72400 -670
rect 72460 -730 72480 -670
rect 72380 -770 72480 -730
rect 72380 -830 72400 -770
rect 72460 -830 72480 -770
rect 72380 -850 72480 -830
rect 72550 -670 72650 -650
rect 72550 -730 72570 -670
rect 72630 -730 72650 -670
rect 72550 -770 72650 -730
rect 72550 -830 72570 -770
rect 72630 -830 72650 -770
rect 72550 -850 72650 -830
rect 72720 -670 72820 -650
rect 72720 -730 72740 -670
rect 72800 -730 72820 -670
rect 72720 -770 72820 -730
rect 72720 -830 72740 -770
rect 72800 -830 72820 -770
rect 72720 -850 72820 -830
rect 72890 -670 72990 -650
rect 72890 -730 72910 -670
rect 72970 -730 72990 -670
rect 72890 -770 72990 -730
rect 72890 -830 72910 -770
rect 72970 -830 72990 -770
rect 72890 -850 72990 -830
rect 73060 -670 73160 -650
rect 73060 -730 73080 -670
rect 73140 -730 73160 -670
rect 73060 -770 73160 -730
rect 73060 -830 73080 -770
rect 73140 -830 73160 -770
rect 73060 -850 73160 -830
rect 73230 -670 73330 -650
rect 73230 -730 73250 -670
rect 73310 -730 73330 -670
rect 73230 -770 73330 -730
rect 73230 -830 73250 -770
rect 73310 -830 73330 -770
rect 73230 -850 73330 -830
rect 73400 -670 73500 -650
rect 73400 -730 73420 -670
rect 73480 -730 73500 -670
rect 73400 -770 73500 -730
rect 73400 -830 73420 -770
rect 73480 -830 73500 -770
rect 73400 -850 73500 -830
rect 73570 -670 73670 -650
rect 73570 -730 73590 -670
rect 73650 -730 73670 -670
rect 73570 -770 73670 -730
rect 73570 -830 73590 -770
rect 73650 -830 73670 -770
rect 73570 -850 73670 -830
rect 73740 -670 73840 -650
rect 73740 -730 73760 -670
rect 73820 -730 73840 -670
rect 73740 -770 73840 -730
rect 73740 -830 73760 -770
rect 73820 -830 73840 -770
rect 73740 -850 73840 -830
rect 73910 -670 74010 -650
rect 73910 -730 73930 -670
rect 73990 -730 74010 -670
rect 73910 -770 74010 -730
rect 73910 -830 73930 -770
rect 73990 -830 74010 -770
rect 73910 -850 74010 -830
rect 74080 -670 74180 -650
rect 74080 -730 74100 -670
rect 74160 -730 74180 -670
rect 74080 -770 74180 -730
rect 74080 -830 74100 -770
rect 74160 -830 74180 -770
rect 74080 -850 74180 -830
rect 74250 -670 74350 -650
rect 74250 -730 74270 -670
rect 74330 -730 74350 -670
rect 74250 -770 74350 -730
rect 74250 -830 74270 -770
rect 74330 -830 74350 -770
rect 74250 -850 74350 -830
rect 74420 -670 74520 -650
rect 74420 -730 74440 -670
rect 74500 -730 74520 -670
rect 74420 -770 74520 -730
rect 74420 -830 74440 -770
rect 74500 -830 74520 -770
rect 74420 -850 74520 -830
rect 74590 -670 74690 -650
rect 74590 -730 74610 -670
rect 74670 -730 74690 -670
rect 74590 -770 74690 -730
rect 74590 -830 74610 -770
rect 74670 -830 74690 -770
rect 74590 -850 74690 -830
rect 74760 -670 74860 -650
rect 74760 -730 74780 -670
rect 74840 -730 74860 -670
rect 74760 -770 74860 -730
rect 74760 -830 74780 -770
rect 74840 -830 74860 -770
rect 74760 -850 74860 -830
rect 74930 -670 75030 -650
rect 74930 -730 74950 -670
rect 75010 -730 75030 -670
rect 74930 -770 75030 -730
rect 74930 -830 74950 -770
rect 75010 -830 75030 -770
rect 74930 -850 75030 -830
rect 75100 -670 75200 -650
rect 75100 -730 75120 -670
rect 75180 -730 75200 -670
rect 75100 -770 75200 -730
rect 75100 -830 75120 -770
rect 75180 -830 75200 -770
rect 75100 -850 75200 -830
rect 75270 -670 75370 -650
rect 75270 -730 75290 -670
rect 75350 -730 75370 -670
rect 75270 -770 75370 -730
rect 75270 -830 75290 -770
rect 75350 -830 75370 -770
rect 75270 -850 75370 -830
rect 75440 -670 75540 -650
rect 75440 -730 75460 -670
rect 75520 -730 75540 -670
rect 75440 -770 75540 -730
rect 75440 -830 75460 -770
rect 75520 -830 75540 -770
rect 75440 -850 75540 -830
rect 75610 -670 75710 -650
rect 75610 -730 75630 -670
rect 75690 -730 75710 -670
rect 75610 -770 75710 -730
rect 75610 -830 75630 -770
rect 75690 -830 75710 -770
rect 75610 -850 75710 -830
rect 75780 -670 75880 -650
rect 75780 -730 75800 -670
rect 75860 -730 75880 -670
rect 75780 -770 75880 -730
rect 75780 -830 75800 -770
rect 75860 -830 75880 -770
rect 75780 -850 75880 -830
rect 75950 -670 76050 -650
rect 75950 -730 75970 -670
rect 76030 -730 76050 -670
rect 75950 -770 76050 -730
rect 75950 -830 75970 -770
rect 76030 -830 76050 -770
rect 75950 -850 76050 -830
rect 76120 -670 76220 -650
rect 76120 -730 76140 -670
rect 76200 -730 76220 -670
rect 76120 -770 76220 -730
rect 76120 -830 76140 -770
rect 76200 -830 76220 -770
rect 76120 -850 76220 -830
rect 76290 -670 76390 -650
rect 76290 -730 76310 -670
rect 76370 -730 76390 -670
rect 76290 -770 76390 -730
rect 76290 -830 76310 -770
rect 76370 -830 76390 -770
rect 76290 -850 76390 -830
rect 76460 -670 76560 -650
rect 76460 -730 76480 -670
rect 76540 -730 76560 -670
rect 76460 -770 76560 -730
rect 76460 -830 76480 -770
rect 76540 -830 76560 -770
rect 76460 -850 76560 -830
rect 76630 -670 76730 -650
rect 76630 -730 76650 -670
rect 76710 -730 76730 -670
rect 76630 -770 76730 -730
rect 76630 -830 76650 -770
rect 76710 -830 76730 -770
rect 76630 -850 76730 -830
rect 76800 -670 76900 -650
rect 76800 -730 76820 -670
rect 76880 -730 76900 -670
rect 76800 -770 76900 -730
rect 76800 -830 76820 -770
rect 76880 -830 76900 -770
rect 76800 -850 76900 -830
rect 76970 -670 77070 -650
rect 76970 -730 76990 -670
rect 77050 -730 77070 -670
rect 76970 -770 77070 -730
rect 76970 -830 76990 -770
rect 77050 -830 77070 -770
rect 76970 -850 77070 -830
rect 77140 -670 77240 -650
rect 77140 -730 77160 -670
rect 77220 -730 77240 -670
rect 77140 -770 77240 -730
rect 77140 -830 77160 -770
rect 77220 -830 77240 -770
rect 77140 -850 77240 -830
rect 77310 -670 77410 -650
rect 77310 -730 77330 -670
rect 77390 -730 77410 -670
rect 77310 -770 77410 -730
rect 77310 -830 77330 -770
rect 77390 -830 77410 -770
rect 77310 -850 77410 -830
rect 77480 -670 77580 -650
rect 77480 -730 77500 -670
rect 77560 -730 77580 -670
rect 77480 -770 77580 -730
rect 77480 -830 77500 -770
rect 77560 -830 77580 -770
rect 77480 -850 77580 -830
rect 77650 -670 77750 -650
rect 77650 -730 77670 -670
rect 77730 -730 77750 -670
rect 77650 -770 77750 -730
rect 77650 -830 77670 -770
rect 77730 -830 77750 -770
rect 77650 -850 77750 -830
rect 77820 -670 77920 -650
rect 77820 -730 77840 -670
rect 77900 -730 77920 -670
rect 77820 -770 77920 -730
rect 77820 -830 77840 -770
rect 77900 -830 77920 -770
rect 77820 -850 77920 -830
rect 77990 -670 78090 -650
rect 77990 -730 78010 -670
rect 78070 -730 78090 -670
rect 77990 -770 78090 -730
rect 77990 -830 78010 -770
rect 78070 -830 78090 -770
rect 77990 -850 78090 -830
rect 78160 -670 78260 -650
rect 78160 -730 78180 -670
rect 78240 -730 78260 -670
rect 78160 -770 78260 -730
rect 78160 -830 78180 -770
rect 78240 -830 78260 -770
rect 78160 -850 78260 -830
rect 78330 -670 78430 -650
rect 78330 -730 78350 -670
rect 78410 -730 78430 -670
rect 78330 -770 78430 -730
rect 78330 -830 78350 -770
rect 78410 -830 78430 -770
rect 78330 -850 78430 -830
rect 78500 -670 78600 -650
rect 78500 -730 78520 -670
rect 78580 -730 78600 -670
rect 78500 -770 78600 -730
rect 78500 -830 78520 -770
rect 78580 -830 78600 -770
rect 78500 -850 78600 -830
rect 78670 -670 78770 -650
rect 78670 -730 78690 -670
rect 78750 -730 78770 -670
rect 78670 -770 78770 -730
rect 78670 -830 78690 -770
rect 78750 -830 78770 -770
rect 78670 -850 78770 -830
rect 78840 -670 78940 -650
rect 78840 -730 78860 -670
rect 78920 -730 78940 -670
rect 78840 -770 78940 -730
rect 78840 -830 78860 -770
rect 78920 -830 78940 -770
rect 78840 -850 78940 -830
rect 79010 -670 79110 -650
rect 79010 -730 79030 -670
rect 79090 -730 79110 -670
rect 79010 -770 79110 -730
rect 79010 -830 79030 -770
rect 79090 -830 79110 -770
rect 79010 -850 79110 -830
rect 79180 -670 79280 -650
rect 79180 -730 79200 -670
rect 79260 -730 79280 -670
rect 79180 -770 79280 -730
rect 79180 -830 79200 -770
rect 79260 -830 79280 -770
rect 79180 -850 79280 -830
rect 79350 -670 79450 -650
rect 79350 -730 79370 -670
rect 79430 -730 79450 -670
rect 79350 -770 79450 -730
rect 79350 -830 79370 -770
rect 79430 -830 79450 -770
rect 79350 -850 79450 -830
rect 79520 -670 79620 -650
rect 79520 -730 79540 -670
rect 79600 -730 79620 -670
rect 79520 -770 79620 -730
rect 79520 -830 79540 -770
rect 79600 -830 79620 -770
rect 79520 -850 79620 -830
rect 79690 -670 79790 -650
rect 79690 -730 79710 -670
rect 79770 -730 79790 -670
rect 79690 -770 79790 -730
rect 79690 -830 79710 -770
rect 79770 -830 79790 -770
rect 79690 -850 79790 -830
rect 79860 -670 79960 -650
rect 79860 -730 79880 -670
rect 79940 -730 79960 -670
rect 79860 -770 79960 -730
rect 79860 -830 79880 -770
rect 79940 -830 79960 -770
rect 79860 -850 79960 -830
rect 80030 -670 80130 -650
rect 80030 -730 80050 -670
rect 80110 -730 80130 -670
rect 80030 -770 80130 -730
rect 80030 -830 80050 -770
rect 80110 -830 80130 -770
rect 80030 -850 80130 -830
rect 80200 -670 80300 -650
rect 80200 -730 80220 -670
rect 80280 -730 80300 -670
rect 80200 -770 80300 -730
rect 80200 -830 80220 -770
rect 80280 -830 80300 -770
rect 80200 -850 80300 -830
rect 80370 -670 80470 -650
rect 80370 -730 80390 -670
rect 80450 -730 80470 -670
rect 80370 -770 80470 -730
rect 80370 -830 80390 -770
rect 80450 -830 80470 -770
rect 80370 -850 80470 -830
rect 80540 -670 80640 -650
rect 80540 -730 80560 -670
rect 80620 -730 80640 -670
rect 80540 -770 80640 -730
rect 80540 -830 80560 -770
rect 80620 -830 80640 -770
rect 80540 -850 80640 -830
rect 80710 -670 80810 -650
rect 80710 -730 80730 -670
rect 80790 -730 80810 -670
rect 80710 -770 80810 -730
rect 80710 -830 80730 -770
rect 80790 -830 80810 -770
rect 80710 -850 80810 -830
rect 80880 -670 80980 -650
rect 80880 -730 80900 -670
rect 80960 -730 80980 -670
rect 80880 -770 80980 -730
rect 80880 -830 80900 -770
rect 80960 -830 80980 -770
rect 80880 -850 80980 -830
rect 81050 -670 81150 -650
rect 81050 -730 81070 -670
rect 81130 -730 81150 -670
rect 81050 -770 81150 -730
rect 81050 -830 81070 -770
rect 81130 -830 81150 -770
rect 81050 -850 81150 -830
rect 81220 -670 81320 -650
rect 81220 -730 81240 -670
rect 81300 -730 81320 -670
rect 81220 -770 81320 -730
rect 81220 -830 81240 -770
rect 81300 -830 81320 -770
rect 81220 -850 81320 -830
rect 81390 -670 81490 -650
rect 81390 -730 81410 -670
rect 81470 -730 81490 -670
rect 81390 -770 81490 -730
rect 81390 -830 81410 -770
rect 81470 -830 81490 -770
rect 81390 -850 81490 -830
rect 81560 -670 81660 -650
rect 81560 -730 81580 -670
rect 81640 -730 81660 -670
rect 81560 -770 81660 -730
rect 81560 -830 81580 -770
rect 81640 -830 81660 -770
rect 81560 -850 81660 -830
rect 81730 -670 81830 -650
rect 81730 -730 81750 -670
rect 81810 -730 81830 -670
rect 81730 -770 81830 -730
rect 81730 -830 81750 -770
rect 81810 -830 81830 -770
rect 81730 -850 81830 -830
rect 81900 -670 82000 -650
rect 81900 -730 81920 -670
rect 81980 -730 82000 -670
rect 81900 -770 82000 -730
rect 81900 -830 81920 -770
rect 81980 -830 82000 -770
rect 81900 -850 82000 -830
rect 82070 -670 82170 -650
rect 82070 -730 82090 -670
rect 82150 -730 82170 -670
rect 82070 -770 82170 -730
rect 82070 -830 82090 -770
rect 82150 -830 82170 -770
rect 82070 -850 82170 -830
rect 82240 -670 82340 -650
rect 82240 -730 82260 -670
rect 82320 -730 82340 -670
rect 82240 -770 82340 -730
rect 82240 -830 82260 -770
rect 82320 -830 82340 -770
rect 82240 -850 82340 -830
rect 82410 -670 82510 -650
rect 82410 -730 82430 -670
rect 82490 -730 82510 -670
rect 82410 -770 82510 -730
rect 82410 -830 82430 -770
rect 82490 -830 82510 -770
rect 82410 -850 82510 -830
rect 82580 -670 82680 -650
rect 82580 -730 82600 -670
rect 82660 -730 82680 -670
rect 82580 -770 82680 -730
rect 82580 -830 82600 -770
rect 82660 -830 82680 -770
rect 82580 -850 82680 -830
rect 82750 -670 82850 -650
rect 82750 -730 82770 -670
rect 82830 -730 82850 -670
rect 82750 -770 82850 -730
rect 82750 -830 82770 -770
rect 82830 -830 82850 -770
rect 82750 -850 82850 -830
rect 82920 -670 83020 -650
rect 82920 -730 82940 -670
rect 83000 -730 83020 -670
rect 82920 -770 83020 -730
rect 82920 -830 82940 -770
rect 83000 -830 83020 -770
rect 82920 -850 83020 -830
rect 83090 -670 83190 -650
rect 83090 -730 83110 -670
rect 83170 -730 83190 -670
rect 83090 -770 83190 -730
rect 83090 -830 83110 -770
rect 83170 -830 83190 -770
rect 83090 -850 83190 -830
rect 83260 -670 83360 -650
rect 83260 -730 83280 -670
rect 83340 -730 83360 -670
rect 83260 -770 83360 -730
rect 83260 -830 83280 -770
rect 83340 -830 83360 -770
rect 83260 -850 83360 -830
rect 83430 -670 83530 -650
rect 83430 -730 83450 -670
rect 83510 -730 83530 -670
rect 83430 -770 83530 -730
rect 83430 -830 83450 -770
rect 83510 -830 83530 -770
rect 83430 -850 83530 -830
rect 83600 -670 83700 -650
rect 83600 -730 83620 -670
rect 83680 -730 83700 -670
rect 83600 -770 83700 -730
rect 83600 -830 83620 -770
rect 83680 -830 83700 -770
rect 83600 -850 83700 -830
rect 83770 -670 83870 -650
rect 83770 -730 83790 -670
rect 83850 -730 83870 -670
rect 83770 -770 83870 -730
rect 83770 -830 83790 -770
rect 83850 -830 83870 -770
rect 83770 -850 83870 -830
rect 83940 -670 84040 -650
rect 83940 -730 83960 -670
rect 84020 -730 84040 -670
rect 83940 -770 84040 -730
rect 83940 -830 83960 -770
rect 84020 -830 84040 -770
rect 83940 -850 84040 -830
rect 84110 -670 84210 -650
rect 84110 -730 84130 -670
rect 84190 -730 84210 -670
rect 84110 -770 84210 -730
rect 84110 -830 84130 -770
rect 84190 -830 84210 -770
rect 84110 -850 84210 -830
rect 84280 -670 84380 -650
rect 84280 -730 84300 -670
rect 84360 -730 84380 -670
rect 84280 -770 84380 -730
rect 84280 -830 84300 -770
rect 84360 -830 84380 -770
rect 84280 -850 84380 -830
rect 84450 -670 84550 -650
rect 84450 -730 84470 -670
rect 84530 -730 84550 -670
rect 84450 -770 84550 -730
rect 84450 -830 84470 -770
rect 84530 -830 84550 -770
rect 84450 -850 84550 -830
rect 84620 -670 84720 -650
rect 84620 -730 84640 -670
rect 84700 -730 84720 -670
rect 84620 -770 84720 -730
rect 84620 -830 84640 -770
rect 84700 -830 84720 -770
rect 84620 -850 84720 -830
rect 84790 -670 84890 -650
rect 84790 -730 84810 -670
rect 84870 -730 84890 -670
rect 84790 -770 84890 -730
rect 84790 -830 84810 -770
rect 84870 -830 84890 -770
rect 84790 -850 84890 -830
rect 84960 -670 85060 -650
rect 84960 -730 84980 -670
rect 85040 -730 85060 -670
rect 84960 -770 85060 -730
rect 84960 -830 84980 -770
rect 85040 -830 85060 -770
rect 84960 -850 85060 -830
rect 85130 -670 85230 -650
rect 85130 -730 85150 -670
rect 85210 -730 85230 -670
rect 85130 -770 85230 -730
rect 85130 -830 85150 -770
rect 85210 -830 85230 -770
rect 85130 -850 85230 -830
rect 85300 -670 85400 -650
rect 85300 -730 85320 -670
rect 85380 -730 85400 -670
rect 85300 -770 85400 -730
rect 85300 -830 85320 -770
rect 85380 -830 85400 -770
rect 85300 -850 85400 -830
rect 85470 -670 85570 -650
rect 85470 -730 85490 -670
rect 85550 -730 85570 -670
rect 85470 -770 85570 -730
rect 85470 -830 85490 -770
rect 85550 -830 85570 -770
rect 85470 -850 85570 -830
rect 85640 -670 85740 -650
rect 85640 -730 85660 -670
rect 85720 -730 85740 -670
rect 85640 -770 85740 -730
rect 85640 -830 85660 -770
rect 85720 -830 85740 -770
rect 85640 -850 85740 -830
rect 85810 -670 85910 -650
rect 85810 -730 85830 -670
rect 85890 -730 85910 -670
rect 85810 -770 85910 -730
rect 85810 -830 85830 -770
rect 85890 -830 85910 -770
rect 85810 -850 85910 -830
rect 85980 -670 86080 -650
rect 85980 -730 86000 -670
rect 86060 -730 86080 -670
rect 85980 -770 86080 -730
rect 85980 -830 86000 -770
rect 86060 -830 86080 -770
rect 85980 -850 86080 -830
rect 86150 -670 86250 -650
rect 86150 -730 86170 -670
rect 86230 -730 86250 -670
rect 86150 -770 86250 -730
rect 86150 -830 86170 -770
rect 86230 -830 86250 -770
rect 86150 -850 86250 -830
rect 86320 -670 86420 -650
rect 86320 -730 86340 -670
rect 86400 -730 86420 -670
rect 86320 -770 86420 -730
rect 86320 -830 86340 -770
rect 86400 -830 86420 -770
rect 86320 -850 86420 -830
rect 86490 -670 86590 -650
rect 86490 -730 86510 -670
rect 86570 -730 86590 -670
rect 86490 -770 86590 -730
rect 86490 -830 86510 -770
rect 86570 -830 86590 -770
rect 86490 -850 86590 -830
rect 86660 -670 86760 -650
rect 86660 -730 86680 -670
rect 86740 -730 86760 -670
rect 86660 -770 86760 -730
rect 86660 -830 86680 -770
rect 86740 -830 86760 -770
rect 86660 -850 86760 -830
rect 86830 -670 86930 -650
rect 86830 -730 86850 -670
rect 86910 -730 86930 -670
rect 86830 -770 86930 -730
rect 86830 -830 86850 -770
rect 86910 -830 86930 -770
rect 86830 -850 86930 -830
rect 87000 -670 87100 -650
rect 87000 -730 87020 -670
rect 87080 -730 87100 -670
rect 87000 -770 87100 -730
rect 87000 -830 87020 -770
rect 87080 -830 87100 -770
rect 87000 -850 87100 -830
rect 87170 -670 87270 -650
rect 87170 -730 87190 -670
rect 87250 -730 87270 -670
rect 87170 -770 87270 -730
rect 87170 -830 87190 -770
rect 87250 -830 87270 -770
rect 87170 -850 87270 -830
rect 130 -1000 230 -980
rect 130 -1060 150 -1000
rect 210 -1060 230 -1000
rect 130 -1100 230 -1060
rect 130 -1160 150 -1100
rect 210 -1160 230 -1100
rect 130 -1200 230 -1160
rect 130 -1260 150 -1200
rect 210 -1260 230 -1200
rect 130 -1300 230 -1260
rect 130 -1360 150 -1300
rect 210 -1360 230 -1300
rect 130 -1380 230 -1360
rect 300 -1000 400 -980
rect 300 -1060 320 -1000
rect 380 -1060 400 -1000
rect 300 -1100 400 -1060
rect 300 -1160 320 -1100
rect 380 -1160 400 -1100
rect 300 -1200 400 -1160
rect 300 -1260 320 -1200
rect 380 -1260 400 -1200
rect 300 -1300 400 -1260
rect 300 -1360 320 -1300
rect 380 -1360 400 -1300
rect 300 -1380 400 -1360
rect 470 -1000 570 -980
rect 470 -1060 490 -1000
rect 550 -1060 570 -1000
rect 470 -1100 570 -1060
rect 470 -1160 490 -1100
rect 550 -1160 570 -1100
rect 470 -1200 570 -1160
rect 470 -1260 490 -1200
rect 550 -1260 570 -1200
rect 470 -1300 570 -1260
rect 470 -1360 490 -1300
rect 550 -1360 570 -1300
rect 470 -1380 570 -1360
rect 640 -1000 740 -980
rect 640 -1060 660 -1000
rect 720 -1060 740 -1000
rect 640 -1100 740 -1060
rect 640 -1160 660 -1100
rect 720 -1160 740 -1100
rect 640 -1200 740 -1160
rect 640 -1260 660 -1200
rect 720 -1260 740 -1200
rect 640 -1300 740 -1260
rect 640 -1360 660 -1300
rect 720 -1360 740 -1300
rect 640 -1380 740 -1360
rect 810 -1000 910 -980
rect 810 -1060 830 -1000
rect 890 -1060 910 -1000
rect 810 -1100 910 -1060
rect 810 -1160 830 -1100
rect 890 -1160 910 -1100
rect 810 -1200 910 -1160
rect 810 -1260 830 -1200
rect 890 -1260 910 -1200
rect 810 -1300 910 -1260
rect 810 -1360 830 -1300
rect 890 -1360 910 -1300
rect 810 -1380 910 -1360
rect 980 -1000 1080 -980
rect 980 -1060 1000 -1000
rect 1060 -1060 1080 -1000
rect 980 -1100 1080 -1060
rect 980 -1160 1000 -1100
rect 1060 -1160 1080 -1100
rect 980 -1200 1080 -1160
rect 980 -1260 1000 -1200
rect 1060 -1260 1080 -1200
rect 980 -1300 1080 -1260
rect 980 -1360 1000 -1300
rect 1060 -1360 1080 -1300
rect 980 -1380 1080 -1360
rect 1150 -1000 1250 -980
rect 1150 -1060 1170 -1000
rect 1230 -1060 1250 -1000
rect 1150 -1100 1250 -1060
rect 1150 -1160 1170 -1100
rect 1230 -1160 1250 -1100
rect 1150 -1200 1250 -1160
rect 1150 -1260 1170 -1200
rect 1230 -1260 1250 -1200
rect 1150 -1300 1250 -1260
rect 1150 -1360 1170 -1300
rect 1230 -1360 1250 -1300
rect 1150 -1380 1250 -1360
rect 1320 -1000 1420 -980
rect 1320 -1060 1340 -1000
rect 1400 -1060 1420 -1000
rect 1320 -1100 1420 -1060
rect 1320 -1160 1340 -1100
rect 1400 -1160 1420 -1100
rect 1320 -1200 1420 -1160
rect 1320 -1260 1340 -1200
rect 1400 -1260 1420 -1200
rect 1320 -1300 1420 -1260
rect 1320 -1360 1340 -1300
rect 1400 -1360 1420 -1300
rect 1320 -1380 1420 -1360
rect 1490 -1000 1590 -980
rect 1490 -1060 1510 -1000
rect 1570 -1060 1590 -1000
rect 1490 -1100 1590 -1060
rect 1490 -1160 1510 -1100
rect 1570 -1160 1590 -1100
rect 1490 -1200 1590 -1160
rect 1490 -1260 1510 -1200
rect 1570 -1260 1590 -1200
rect 1490 -1300 1590 -1260
rect 1490 -1360 1510 -1300
rect 1570 -1360 1590 -1300
rect 1490 -1380 1590 -1360
rect 1660 -1000 1760 -980
rect 1660 -1060 1680 -1000
rect 1740 -1060 1760 -1000
rect 1660 -1100 1760 -1060
rect 1660 -1160 1680 -1100
rect 1740 -1160 1760 -1100
rect 1660 -1200 1760 -1160
rect 1660 -1260 1680 -1200
rect 1740 -1260 1760 -1200
rect 1660 -1300 1760 -1260
rect 1660 -1360 1680 -1300
rect 1740 -1360 1760 -1300
rect 1660 -1380 1760 -1360
rect 1830 -1000 1930 -980
rect 1830 -1060 1850 -1000
rect 1910 -1060 1930 -1000
rect 1830 -1100 1930 -1060
rect 1830 -1160 1850 -1100
rect 1910 -1160 1930 -1100
rect 1830 -1200 1930 -1160
rect 1830 -1260 1850 -1200
rect 1910 -1260 1930 -1200
rect 1830 -1300 1930 -1260
rect 1830 -1360 1850 -1300
rect 1910 -1360 1930 -1300
rect 1830 -1380 1930 -1360
rect 2000 -1000 2100 -980
rect 2000 -1060 2020 -1000
rect 2080 -1060 2100 -1000
rect 2000 -1100 2100 -1060
rect 2000 -1160 2020 -1100
rect 2080 -1160 2100 -1100
rect 2000 -1200 2100 -1160
rect 2000 -1260 2020 -1200
rect 2080 -1260 2100 -1200
rect 2000 -1300 2100 -1260
rect 2000 -1360 2020 -1300
rect 2080 -1360 2100 -1300
rect 2000 -1380 2100 -1360
rect 2170 -1000 2270 -980
rect 2170 -1060 2190 -1000
rect 2250 -1060 2270 -1000
rect 2170 -1100 2270 -1060
rect 2170 -1160 2190 -1100
rect 2250 -1160 2270 -1100
rect 2170 -1200 2270 -1160
rect 2170 -1260 2190 -1200
rect 2250 -1260 2270 -1200
rect 2170 -1300 2270 -1260
rect 2170 -1360 2190 -1300
rect 2250 -1360 2270 -1300
rect 2170 -1380 2270 -1360
rect 2340 -1000 2440 -980
rect 2340 -1060 2360 -1000
rect 2420 -1060 2440 -1000
rect 2340 -1100 2440 -1060
rect 2340 -1160 2360 -1100
rect 2420 -1160 2440 -1100
rect 2340 -1200 2440 -1160
rect 2340 -1260 2360 -1200
rect 2420 -1260 2440 -1200
rect 2340 -1300 2440 -1260
rect 2340 -1360 2360 -1300
rect 2420 -1360 2440 -1300
rect 2340 -1380 2440 -1360
rect 2510 -1000 2610 -980
rect 2510 -1060 2530 -1000
rect 2590 -1060 2610 -1000
rect 2510 -1100 2610 -1060
rect 2510 -1160 2530 -1100
rect 2590 -1160 2610 -1100
rect 2510 -1200 2610 -1160
rect 2510 -1260 2530 -1200
rect 2590 -1260 2610 -1200
rect 2510 -1300 2610 -1260
rect 2510 -1360 2530 -1300
rect 2590 -1360 2610 -1300
rect 2510 -1380 2610 -1360
rect 2680 -1000 2780 -980
rect 2680 -1060 2700 -1000
rect 2760 -1060 2780 -1000
rect 2680 -1100 2780 -1060
rect 2680 -1160 2700 -1100
rect 2760 -1160 2780 -1100
rect 2680 -1200 2780 -1160
rect 2680 -1260 2700 -1200
rect 2760 -1260 2780 -1200
rect 2680 -1300 2780 -1260
rect 2680 -1360 2700 -1300
rect 2760 -1360 2780 -1300
rect 2680 -1380 2780 -1360
rect 2850 -1000 2950 -980
rect 2850 -1060 2870 -1000
rect 2930 -1060 2950 -1000
rect 2850 -1100 2950 -1060
rect 2850 -1160 2870 -1100
rect 2930 -1160 2950 -1100
rect 2850 -1200 2950 -1160
rect 2850 -1260 2870 -1200
rect 2930 -1260 2950 -1200
rect 2850 -1300 2950 -1260
rect 2850 -1360 2870 -1300
rect 2930 -1360 2950 -1300
rect 2850 -1380 2950 -1360
rect 3020 -1000 3120 -980
rect 3020 -1060 3040 -1000
rect 3100 -1060 3120 -1000
rect 3020 -1100 3120 -1060
rect 3020 -1160 3040 -1100
rect 3100 -1160 3120 -1100
rect 3020 -1200 3120 -1160
rect 3020 -1260 3040 -1200
rect 3100 -1260 3120 -1200
rect 3020 -1300 3120 -1260
rect 3020 -1360 3040 -1300
rect 3100 -1360 3120 -1300
rect 3020 -1380 3120 -1360
rect 3190 -1000 3290 -980
rect 3190 -1060 3210 -1000
rect 3270 -1060 3290 -1000
rect 3190 -1100 3290 -1060
rect 3190 -1160 3210 -1100
rect 3270 -1160 3290 -1100
rect 3190 -1200 3290 -1160
rect 3190 -1260 3210 -1200
rect 3270 -1260 3290 -1200
rect 3190 -1300 3290 -1260
rect 3190 -1360 3210 -1300
rect 3270 -1360 3290 -1300
rect 3190 -1380 3290 -1360
rect 3360 -1000 3460 -980
rect 3360 -1060 3380 -1000
rect 3440 -1060 3460 -1000
rect 3360 -1100 3460 -1060
rect 3360 -1160 3380 -1100
rect 3440 -1160 3460 -1100
rect 3360 -1200 3460 -1160
rect 3360 -1260 3380 -1200
rect 3440 -1260 3460 -1200
rect 3360 -1300 3460 -1260
rect 3360 -1360 3380 -1300
rect 3440 -1360 3460 -1300
rect 3360 -1380 3460 -1360
rect 3530 -1000 3630 -980
rect 3530 -1060 3550 -1000
rect 3610 -1060 3630 -1000
rect 3530 -1100 3630 -1060
rect 3530 -1160 3550 -1100
rect 3610 -1160 3630 -1100
rect 3530 -1200 3630 -1160
rect 3530 -1260 3550 -1200
rect 3610 -1260 3630 -1200
rect 3530 -1300 3630 -1260
rect 3530 -1360 3550 -1300
rect 3610 -1360 3630 -1300
rect 3530 -1380 3630 -1360
rect 3700 -1000 3800 -980
rect 3700 -1060 3720 -1000
rect 3780 -1060 3800 -1000
rect 3700 -1100 3800 -1060
rect 3700 -1160 3720 -1100
rect 3780 -1160 3800 -1100
rect 3700 -1200 3800 -1160
rect 3700 -1260 3720 -1200
rect 3780 -1260 3800 -1200
rect 3700 -1300 3800 -1260
rect 3700 -1360 3720 -1300
rect 3780 -1360 3800 -1300
rect 3700 -1380 3800 -1360
rect 3870 -1000 3970 -980
rect 3870 -1060 3890 -1000
rect 3950 -1060 3970 -1000
rect 3870 -1100 3970 -1060
rect 3870 -1160 3890 -1100
rect 3950 -1160 3970 -1100
rect 3870 -1200 3970 -1160
rect 3870 -1260 3890 -1200
rect 3950 -1260 3970 -1200
rect 3870 -1300 3970 -1260
rect 3870 -1360 3890 -1300
rect 3950 -1360 3970 -1300
rect 3870 -1380 3970 -1360
rect 4040 -1000 4140 -980
rect 4040 -1060 4060 -1000
rect 4120 -1060 4140 -1000
rect 4040 -1100 4140 -1060
rect 4040 -1160 4060 -1100
rect 4120 -1160 4140 -1100
rect 4040 -1200 4140 -1160
rect 4040 -1260 4060 -1200
rect 4120 -1260 4140 -1200
rect 4040 -1300 4140 -1260
rect 4040 -1360 4060 -1300
rect 4120 -1360 4140 -1300
rect 4040 -1380 4140 -1360
rect 4210 -1000 4310 -980
rect 4210 -1060 4230 -1000
rect 4290 -1060 4310 -1000
rect 4210 -1100 4310 -1060
rect 4210 -1160 4230 -1100
rect 4290 -1160 4310 -1100
rect 4210 -1200 4310 -1160
rect 4210 -1260 4230 -1200
rect 4290 -1260 4310 -1200
rect 4210 -1300 4310 -1260
rect 4210 -1360 4230 -1300
rect 4290 -1360 4310 -1300
rect 4210 -1380 4310 -1360
rect 4380 -1000 4480 -980
rect 4380 -1060 4400 -1000
rect 4460 -1060 4480 -1000
rect 4380 -1100 4480 -1060
rect 4380 -1160 4400 -1100
rect 4460 -1160 4480 -1100
rect 4380 -1200 4480 -1160
rect 4380 -1260 4400 -1200
rect 4460 -1260 4480 -1200
rect 4380 -1300 4480 -1260
rect 4380 -1360 4400 -1300
rect 4460 -1360 4480 -1300
rect 4380 -1380 4480 -1360
rect 4550 -1000 4650 -980
rect 4550 -1060 4570 -1000
rect 4630 -1060 4650 -1000
rect 4550 -1100 4650 -1060
rect 4550 -1160 4570 -1100
rect 4630 -1160 4650 -1100
rect 4550 -1200 4650 -1160
rect 4550 -1260 4570 -1200
rect 4630 -1260 4650 -1200
rect 4550 -1300 4650 -1260
rect 4550 -1360 4570 -1300
rect 4630 -1360 4650 -1300
rect 4550 -1380 4650 -1360
rect 4720 -1000 4820 -980
rect 4720 -1060 4740 -1000
rect 4800 -1060 4820 -1000
rect 4720 -1100 4820 -1060
rect 4720 -1160 4740 -1100
rect 4800 -1160 4820 -1100
rect 4720 -1200 4820 -1160
rect 4720 -1260 4740 -1200
rect 4800 -1260 4820 -1200
rect 4720 -1300 4820 -1260
rect 4720 -1360 4740 -1300
rect 4800 -1360 4820 -1300
rect 4720 -1380 4820 -1360
rect 4890 -1000 4990 -980
rect 4890 -1060 4910 -1000
rect 4970 -1060 4990 -1000
rect 4890 -1100 4990 -1060
rect 4890 -1160 4910 -1100
rect 4970 -1160 4990 -1100
rect 4890 -1200 4990 -1160
rect 4890 -1260 4910 -1200
rect 4970 -1260 4990 -1200
rect 4890 -1300 4990 -1260
rect 4890 -1360 4910 -1300
rect 4970 -1360 4990 -1300
rect 4890 -1380 4990 -1360
rect 5060 -1000 5160 -980
rect 5060 -1060 5080 -1000
rect 5140 -1060 5160 -1000
rect 5060 -1100 5160 -1060
rect 5060 -1160 5080 -1100
rect 5140 -1160 5160 -1100
rect 5060 -1200 5160 -1160
rect 5060 -1260 5080 -1200
rect 5140 -1260 5160 -1200
rect 5060 -1300 5160 -1260
rect 5060 -1360 5080 -1300
rect 5140 -1360 5160 -1300
rect 5060 -1380 5160 -1360
rect 5230 -1000 5330 -980
rect 5230 -1060 5250 -1000
rect 5310 -1060 5330 -1000
rect 5230 -1100 5330 -1060
rect 5230 -1160 5250 -1100
rect 5310 -1160 5330 -1100
rect 5230 -1200 5330 -1160
rect 5230 -1260 5250 -1200
rect 5310 -1260 5330 -1200
rect 5230 -1300 5330 -1260
rect 5230 -1360 5250 -1300
rect 5310 -1360 5330 -1300
rect 5230 -1380 5330 -1360
rect 5400 -1000 5500 -980
rect 5400 -1060 5420 -1000
rect 5480 -1060 5500 -1000
rect 5400 -1100 5500 -1060
rect 5400 -1160 5420 -1100
rect 5480 -1160 5500 -1100
rect 5400 -1200 5500 -1160
rect 5400 -1260 5420 -1200
rect 5480 -1260 5500 -1200
rect 5400 -1300 5500 -1260
rect 5400 -1360 5420 -1300
rect 5480 -1360 5500 -1300
rect 5400 -1380 5500 -1360
rect 5570 -1000 5670 -980
rect 5570 -1060 5590 -1000
rect 5650 -1060 5670 -1000
rect 5570 -1100 5670 -1060
rect 5570 -1160 5590 -1100
rect 5650 -1160 5670 -1100
rect 5570 -1200 5670 -1160
rect 5570 -1260 5590 -1200
rect 5650 -1260 5670 -1200
rect 5570 -1300 5670 -1260
rect 5570 -1360 5590 -1300
rect 5650 -1360 5670 -1300
rect 5570 -1380 5670 -1360
rect 5740 -1000 5840 -980
rect 5740 -1060 5760 -1000
rect 5820 -1060 5840 -1000
rect 5740 -1100 5840 -1060
rect 5740 -1160 5760 -1100
rect 5820 -1160 5840 -1100
rect 5740 -1200 5840 -1160
rect 5740 -1260 5760 -1200
rect 5820 -1260 5840 -1200
rect 5740 -1300 5840 -1260
rect 5740 -1360 5760 -1300
rect 5820 -1360 5840 -1300
rect 5740 -1380 5840 -1360
rect 5910 -1000 6010 -980
rect 5910 -1060 5930 -1000
rect 5990 -1060 6010 -1000
rect 5910 -1100 6010 -1060
rect 5910 -1160 5930 -1100
rect 5990 -1160 6010 -1100
rect 5910 -1200 6010 -1160
rect 5910 -1260 5930 -1200
rect 5990 -1260 6010 -1200
rect 5910 -1300 6010 -1260
rect 5910 -1360 5930 -1300
rect 5990 -1360 6010 -1300
rect 5910 -1380 6010 -1360
rect 6080 -1000 6180 -980
rect 6080 -1060 6100 -1000
rect 6160 -1060 6180 -1000
rect 6080 -1100 6180 -1060
rect 6080 -1160 6100 -1100
rect 6160 -1160 6180 -1100
rect 6080 -1200 6180 -1160
rect 6080 -1260 6100 -1200
rect 6160 -1260 6180 -1200
rect 6080 -1300 6180 -1260
rect 6080 -1360 6100 -1300
rect 6160 -1360 6180 -1300
rect 6080 -1380 6180 -1360
rect 6250 -1000 6350 -980
rect 6250 -1060 6270 -1000
rect 6330 -1060 6350 -1000
rect 6250 -1100 6350 -1060
rect 6250 -1160 6270 -1100
rect 6330 -1160 6350 -1100
rect 6250 -1200 6350 -1160
rect 6250 -1260 6270 -1200
rect 6330 -1260 6350 -1200
rect 6250 -1300 6350 -1260
rect 6250 -1360 6270 -1300
rect 6330 -1360 6350 -1300
rect 6250 -1380 6350 -1360
rect 6420 -1000 6520 -980
rect 6420 -1060 6440 -1000
rect 6500 -1060 6520 -1000
rect 6420 -1100 6520 -1060
rect 6420 -1160 6440 -1100
rect 6500 -1160 6520 -1100
rect 6420 -1200 6520 -1160
rect 6420 -1260 6440 -1200
rect 6500 -1260 6520 -1200
rect 6420 -1300 6520 -1260
rect 6420 -1360 6440 -1300
rect 6500 -1360 6520 -1300
rect 6420 -1380 6520 -1360
rect 6590 -1000 6690 -980
rect 6590 -1060 6610 -1000
rect 6670 -1060 6690 -1000
rect 6590 -1100 6690 -1060
rect 6590 -1160 6610 -1100
rect 6670 -1160 6690 -1100
rect 6590 -1200 6690 -1160
rect 6590 -1260 6610 -1200
rect 6670 -1260 6690 -1200
rect 6590 -1300 6690 -1260
rect 6590 -1360 6610 -1300
rect 6670 -1360 6690 -1300
rect 6590 -1380 6690 -1360
rect 6760 -1000 6860 -980
rect 6760 -1060 6780 -1000
rect 6840 -1060 6860 -1000
rect 6760 -1100 6860 -1060
rect 6760 -1160 6780 -1100
rect 6840 -1160 6860 -1100
rect 6760 -1200 6860 -1160
rect 6760 -1260 6780 -1200
rect 6840 -1260 6860 -1200
rect 6760 -1300 6860 -1260
rect 6760 -1360 6780 -1300
rect 6840 -1360 6860 -1300
rect 6760 -1380 6860 -1360
rect 6930 -1000 7030 -980
rect 6930 -1060 6950 -1000
rect 7010 -1060 7030 -1000
rect 6930 -1100 7030 -1060
rect 6930 -1160 6950 -1100
rect 7010 -1160 7030 -1100
rect 6930 -1200 7030 -1160
rect 6930 -1260 6950 -1200
rect 7010 -1260 7030 -1200
rect 6930 -1300 7030 -1260
rect 6930 -1360 6950 -1300
rect 7010 -1360 7030 -1300
rect 6930 -1380 7030 -1360
rect 7100 -1000 7200 -980
rect 7100 -1060 7120 -1000
rect 7180 -1060 7200 -1000
rect 7100 -1100 7200 -1060
rect 7100 -1160 7120 -1100
rect 7180 -1160 7200 -1100
rect 7100 -1200 7200 -1160
rect 7100 -1260 7120 -1200
rect 7180 -1260 7200 -1200
rect 7100 -1300 7200 -1260
rect 7100 -1360 7120 -1300
rect 7180 -1360 7200 -1300
rect 7100 -1380 7200 -1360
rect 7270 -1000 7370 -980
rect 7270 -1060 7290 -1000
rect 7350 -1060 7370 -1000
rect 7270 -1100 7370 -1060
rect 7270 -1160 7290 -1100
rect 7350 -1160 7370 -1100
rect 7270 -1200 7370 -1160
rect 7270 -1260 7290 -1200
rect 7350 -1260 7370 -1200
rect 7270 -1300 7370 -1260
rect 7270 -1360 7290 -1300
rect 7350 -1360 7370 -1300
rect 7270 -1380 7370 -1360
rect 7440 -1000 7540 -980
rect 7440 -1060 7460 -1000
rect 7520 -1060 7540 -1000
rect 7440 -1100 7540 -1060
rect 7440 -1160 7460 -1100
rect 7520 -1160 7540 -1100
rect 7440 -1200 7540 -1160
rect 7440 -1260 7460 -1200
rect 7520 -1260 7540 -1200
rect 7440 -1300 7540 -1260
rect 7440 -1360 7460 -1300
rect 7520 -1360 7540 -1300
rect 7440 -1380 7540 -1360
rect 7610 -1000 7710 -980
rect 7610 -1060 7630 -1000
rect 7690 -1060 7710 -1000
rect 7610 -1100 7710 -1060
rect 7610 -1160 7630 -1100
rect 7690 -1160 7710 -1100
rect 7610 -1200 7710 -1160
rect 7610 -1260 7630 -1200
rect 7690 -1260 7710 -1200
rect 7610 -1300 7710 -1260
rect 7610 -1360 7630 -1300
rect 7690 -1360 7710 -1300
rect 7610 -1380 7710 -1360
rect 7780 -1000 7880 -980
rect 7780 -1060 7800 -1000
rect 7860 -1060 7880 -1000
rect 7780 -1100 7880 -1060
rect 7780 -1160 7800 -1100
rect 7860 -1160 7880 -1100
rect 7780 -1200 7880 -1160
rect 7780 -1260 7800 -1200
rect 7860 -1260 7880 -1200
rect 7780 -1300 7880 -1260
rect 7780 -1360 7800 -1300
rect 7860 -1360 7880 -1300
rect 7780 -1380 7880 -1360
rect 7950 -1000 8050 -980
rect 7950 -1060 7970 -1000
rect 8030 -1060 8050 -1000
rect 7950 -1100 8050 -1060
rect 7950 -1160 7970 -1100
rect 8030 -1160 8050 -1100
rect 7950 -1200 8050 -1160
rect 7950 -1260 7970 -1200
rect 8030 -1260 8050 -1200
rect 7950 -1300 8050 -1260
rect 7950 -1360 7970 -1300
rect 8030 -1360 8050 -1300
rect 7950 -1380 8050 -1360
rect 8120 -1000 8220 -980
rect 8120 -1060 8140 -1000
rect 8200 -1060 8220 -1000
rect 8120 -1100 8220 -1060
rect 8120 -1160 8140 -1100
rect 8200 -1160 8220 -1100
rect 8120 -1200 8220 -1160
rect 8120 -1260 8140 -1200
rect 8200 -1260 8220 -1200
rect 8120 -1300 8220 -1260
rect 8120 -1360 8140 -1300
rect 8200 -1360 8220 -1300
rect 8120 -1380 8220 -1360
rect 8290 -1000 8390 -980
rect 8290 -1060 8310 -1000
rect 8370 -1060 8390 -1000
rect 8290 -1100 8390 -1060
rect 8290 -1160 8310 -1100
rect 8370 -1160 8390 -1100
rect 8290 -1200 8390 -1160
rect 8290 -1260 8310 -1200
rect 8370 -1260 8390 -1200
rect 8290 -1300 8390 -1260
rect 8290 -1360 8310 -1300
rect 8370 -1360 8390 -1300
rect 8290 -1380 8390 -1360
rect 8460 -1000 8560 -980
rect 8460 -1060 8480 -1000
rect 8540 -1060 8560 -1000
rect 8460 -1100 8560 -1060
rect 8460 -1160 8480 -1100
rect 8540 -1160 8560 -1100
rect 8460 -1200 8560 -1160
rect 8460 -1260 8480 -1200
rect 8540 -1260 8560 -1200
rect 8460 -1300 8560 -1260
rect 8460 -1360 8480 -1300
rect 8540 -1360 8560 -1300
rect 8460 -1380 8560 -1360
rect 8630 -1000 8730 -980
rect 8630 -1060 8650 -1000
rect 8710 -1060 8730 -1000
rect 8630 -1100 8730 -1060
rect 8630 -1160 8650 -1100
rect 8710 -1160 8730 -1100
rect 8630 -1200 8730 -1160
rect 8630 -1260 8650 -1200
rect 8710 -1260 8730 -1200
rect 8630 -1300 8730 -1260
rect 8630 -1360 8650 -1300
rect 8710 -1360 8730 -1300
rect 8630 -1380 8730 -1360
rect 8800 -1000 8900 -980
rect 8800 -1060 8820 -1000
rect 8880 -1060 8900 -1000
rect 8800 -1100 8900 -1060
rect 8800 -1160 8820 -1100
rect 8880 -1160 8900 -1100
rect 8800 -1200 8900 -1160
rect 8800 -1260 8820 -1200
rect 8880 -1260 8900 -1200
rect 8800 -1300 8900 -1260
rect 8800 -1360 8820 -1300
rect 8880 -1360 8900 -1300
rect 8800 -1380 8900 -1360
rect 8970 -1000 9070 -980
rect 8970 -1060 8990 -1000
rect 9050 -1060 9070 -1000
rect 8970 -1100 9070 -1060
rect 8970 -1160 8990 -1100
rect 9050 -1160 9070 -1100
rect 8970 -1200 9070 -1160
rect 8970 -1260 8990 -1200
rect 9050 -1260 9070 -1200
rect 8970 -1300 9070 -1260
rect 8970 -1360 8990 -1300
rect 9050 -1360 9070 -1300
rect 8970 -1380 9070 -1360
rect 9140 -1000 9240 -980
rect 9140 -1060 9160 -1000
rect 9220 -1060 9240 -1000
rect 9140 -1100 9240 -1060
rect 9140 -1160 9160 -1100
rect 9220 -1160 9240 -1100
rect 9140 -1200 9240 -1160
rect 9140 -1260 9160 -1200
rect 9220 -1260 9240 -1200
rect 9140 -1300 9240 -1260
rect 9140 -1360 9160 -1300
rect 9220 -1360 9240 -1300
rect 9140 -1380 9240 -1360
rect 9310 -1000 9410 -980
rect 9310 -1060 9330 -1000
rect 9390 -1060 9410 -1000
rect 9310 -1100 9410 -1060
rect 9310 -1160 9330 -1100
rect 9390 -1160 9410 -1100
rect 9310 -1200 9410 -1160
rect 9310 -1260 9330 -1200
rect 9390 -1260 9410 -1200
rect 9310 -1300 9410 -1260
rect 9310 -1360 9330 -1300
rect 9390 -1360 9410 -1300
rect 9310 -1380 9410 -1360
rect 9480 -1000 9580 -980
rect 9480 -1060 9500 -1000
rect 9560 -1060 9580 -1000
rect 9480 -1100 9580 -1060
rect 9480 -1160 9500 -1100
rect 9560 -1160 9580 -1100
rect 9480 -1200 9580 -1160
rect 9480 -1260 9500 -1200
rect 9560 -1260 9580 -1200
rect 9480 -1300 9580 -1260
rect 9480 -1360 9500 -1300
rect 9560 -1360 9580 -1300
rect 9480 -1380 9580 -1360
rect 9650 -1000 9750 -980
rect 9650 -1060 9670 -1000
rect 9730 -1060 9750 -1000
rect 9650 -1100 9750 -1060
rect 9650 -1160 9670 -1100
rect 9730 -1160 9750 -1100
rect 9650 -1200 9750 -1160
rect 9650 -1260 9670 -1200
rect 9730 -1260 9750 -1200
rect 9650 -1300 9750 -1260
rect 9650 -1360 9670 -1300
rect 9730 -1360 9750 -1300
rect 9650 -1380 9750 -1360
rect 9820 -1000 9920 -980
rect 9820 -1060 9840 -1000
rect 9900 -1060 9920 -1000
rect 9820 -1100 9920 -1060
rect 9820 -1160 9840 -1100
rect 9900 -1160 9920 -1100
rect 9820 -1200 9920 -1160
rect 9820 -1260 9840 -1200
rect 9900 -1260 9920 -1200
rect 9820 -1300 9920 -1260
rect 9820 -1360 9840 -1300
rect 9900 -1360 9920 -1300
rect 9820 -1380 9920 -1360
rect 9990 -1000 10090 -980
rect 9990 -1060 10010 -1000
rect 10070 -1060 10090 -1000
rect 9990 -1100 10090 -1060
rect 9990 -1160 10010 -1100
rect 10070 -1160 10090 -1100
rect 9990 -1200 10090 -1160
rect 9990 -1260 10010 -1200
rect 10070 -1260 10090 -1200
rect 9990 -1300 10090 -1260
rect 9990 -1360 10010 -1300
rect 10070 -1360 10090 -1300
rect 9990 -1380 10090 -1360
rect 10160 -1000 10260 -980
rect 10160 -1060 10180 -1000
rect 10240 -1060 10260 -1000
rect 10160 -1100 10260 -1060
rect 10160 -1160 10180 -1100
rect 10240 -1160 10260 -1100
rect 10160 -1200 10260 -1160
rect 10160 -1260 10180 -1200
rect 10240 -1260 10260 -1200
rect 10160 -1300 10260 -1260
rect 10160 -1360 10180 -1300
rect 10240 -1360 10260 -1300
rect 10160 -1380 10260 -1360
rect 10330 -1000 10430 -980
rect 10330 -1060 10350 -1000
rect 10410 -1060 10430 -1000
rect 10330 -1100 10430 -1060
rect 10330 -1160 10350 -1100
rect 10410 -1160 10430 -1100
rect 10330 -1200 10430 -1160
rect 10330 -1260 10350 -1200
rect 10410 -1260 10430 -1200
rect 10330 -1300 10430 -1260
rect 10330 -1360 10350 -1300
rect 10410 -1360 10430 -1300
rect 10330 -1380 10430 -1360
rect 10500 -1000 10600 -980
rect 10500 -1060 10520 -1000
rect 10580 -1060 10600 -1000
rect 10500 -1100 10600 -1060
rect 10500 -1160 10520 -1100
rect 10580 -1160 10600 -1100
rect 10500 -1200 10600 -1160
rect 10500 -1260 10520 -1200
rect 10580 -1260 10600 -1200
rect 10500 -1300 10600 -1260
rect 10500 -1360 10520 -1300
rect 10580 -1360 10600 -1300
rect 10500 -1380 10600 -1360
rect 10670 -1000 10770 -980
rect 10670 -1060 10690 -1000
rect 10750 -1060 10770 -1000
rect 10670 -1100 10770 -1060
rect 10670 -1160 10690 -1100
rect 10750 -1160 10770 -1100
rect 10670 -1200 10770 -1160
rect 10670 -1260 10690 -1200
rect 10750 -1260 10770 -1200
rect 10670 -1300 10770 -1260
rect 10670 -1360 10690 -1300
rect 10750 -1360 10770 -1300
rect 10670 -1380 10770 -1360
rect 10840 -1000 10940 -980
rect 10840 -1060 10860 -1000
rect 10920 -1060 10940 -1000
rect 10840 -1100 10940 -1060
rect 10840 -1160 10860 -1100
rect 10920 -1160 10940 -1100
rect 10840 -1200 10940 -1160
rect 10840 -1260 10860 -1200
rect 10920 -1260 10940 -1200
rect 10840 -1300 10940 -1260
rect 10840 -1360 10860 -1300
rect 10920 -1360 10940 -1300
rect 10840 -1380 10940 -1360
rect 11010 -1000 11110 -980
rect 11010 -1060 11030 -1000
rect 11090 -1060 11110 -1000
rect 11010 -1100 11110 -1060
rect 11010 -1160 11030 -1100
rect 11090 -1160 11110 -1100
rect 11010 -1200 11110 -1160
rect 11010 -1260 11030 -1200
rect 11090 -1260 11110 -1200
rect 11010 -1300 11110 -1260
rect 11010 -1360 11030 -1300
rect 11090 -1360 11110 -1300
rect 11010 -1380 11110 -1360
rect 11180 -1000 11280 -980
rect 11180 -1060 11200 -1000
rect 11260 -1060 11280 -1000
rect 11180 -1100 11280 -1060
rect 11180 -1160 11200 -1100
rect 11260 -1160 11280 -1100
rect 11180 -1200 11280 -1160
rect 11180 -1260 11200 -1200
rect 11260 -1260 11280 -1200
rect 11180 -1300 11280 -1260
rect 11180 -1360 11200 -1300
rect 11260 -1360 11280 -1300
rect 11180 -1380 11280 -1360
rect 11350 -1000 11450 -980
rect 11350 -1060 11370 -1000
rect 11430 -1060 11450 -1000
rect 11350 -1100 11450 -1060
rect 11350 -1160 11370 -1100
rect 11430 -1160 11450 -1100
rect 11350 -1200 11450 -1160
rect 11350 -1260 11370 -1200
rect 11430 -1260 11450 -1200
rect 11350 -1300 11450 -1260
rect 11350 -1360 11370 -1300
rect 11430 -1360 11450 -1300
rect 11350 -1380 11450 -1360
rect 11520 -1000 11620 -980
rect 11520 -1060 11540 -1000
rect 11600 -1060 11620 -1000
rect 11520 -1100 11620 -1060
rect 11520 -1160 11540 -1100
rect 11600 -1160 11620 -1100
rect 11520 -1200 11620 -1160
rect 11520 -1260 11540 -1200
rect 11600 -1260 11620 -1200
rect 11520 -1300 11620 -1260
rect 11520 -1360 11540 -1300
rect 11600 -1360 11620 -1300
rect 11520 -1380 11620 -1360
rect 11690 -1000 11790 -980
rect 11690 -1060 11710 -1000
rect 11770 -1060 11790 -1000
rect 11690 -1100 11790 -1060
rect 11690 -1160 11710 -1100
rect 11770 -1160 11790 -1100
rect 11690 -1200 11790 -1160
rect 11690 -1260 11710 -1200
rect 11770 -1260 11790 -1200
rect 11690 -1300 11790 -1260
rect 11690 -1360 11710 -1300
rect 11770 -1360 11790 -1300
rect 11690 -1380 11790 -1360
rect 11860 -1000 11960 -980
rect 11860 -1060 11880 -1000
rect 11940 -1060 11960 -1000
rect 11860 -1100 11960 -1060
rect 11860 -1160 11880 -1100
rect 11940 -1160 11960 -1100
rect 11860 -1200 11960 -1160
rect 11860 -1260 11880 -1200
rect 11940 -1260 11960 -1200
rect 11860 -1300 11960 -1260
rect 11860 -1360 11880 -1300
rect 11940 -1360 11960 -1300
rect 11860 -1380 11960 -1360
rect 12030 -1000 12130 -980
rect 12030 -1060 12050 -1000
rect 12110 -1060 12130 -1000
rect 12030 -1100 12130 -1060
rect 12030 -1160 12050 -1100
rect 12110 -1160 12130 -1100
rect 12030 -1200 12130 -1160
rect 12030 -1260 12050 -1200
rect 12110 -1260 12130 -1200
rect 12030 -1300 12130 -1260
rect 12030 -1360 12050 -1300
rect 12110 -1360 12130 -1300
rect 12030 -1380 12130 -1360
rect 12200 -1000 12300 -980
rect 12200 -1060 12220 -1000
rect 12280 -1060 12300 -1000
rect 12200 -1100 12300 -1060
rect 12200 -1160 12220 -1100
rect 12280 -1160 12300 -1100
rect 12200 -1200 12300 -1160
rect 12200 -1260 12220 -1200
rect 12280 -1260 12300 -1200
rect 12200 -1300 12300 -1260
rect 12200 -1360 12220 -1300
rect 12280 -1360 12300 -1300
rect 12200 -1380 12300 -1360
rect 12370 -1000 12470 -980
rect 12370 -1060 12390 -1000
rect 12450 -1060 12470 -1000
rect 12370 -1100 12470 -1060
rect 12370 -1160 12390 -1100
rect 12450 -1160 12470 -1100
rect 12370 -1200 12470 -1160
rect 12370 -1260 12390 -1200
rect 12450 -1260 12470 -1200
rect 12370 -1300 12470 -1260
rect 12370 -1360 12390 -1300
rect 12450 -1360 12470 -1300
rect 12370 -1380 12470 -1360
rect 12540 -1000 12640 -980
rect 12540 -1060 12560 -1000
rect 12620 -1060 12640 -1000
rect 12540 -1100 12640 -1060
rect 12540 -1160 12560 -1100
rect 12620 -1160 12640 -1100
rect 12540 -1200 12640 -1160
rect 12540 -1260 12560 -1200
rect 12620 -1260 12640 -1200
rect 12540 -1300 12640 -1260
rect 12540 -1360 12560 -1300
rect 12620 -1360 12640 -1300
rect 12540 -1380 12640 -1360
rect 12710 -1000 12810 -980
rect 12710 -1060 12730 -1000
rect 12790 -1060 12810 -1000
rect 12710 -1100 12810 -1060
rect 12710 -1160 12730 -1100
rect 12790 -1160 12810 -1100
rect 12710 -1200 12810 -1160
rect 12710 -1260 12730 -1200
rect 12790 -1260 12810 -1200
rect 12710 -1300 12810 -1260
rect 12710 -1360 12730 -1300
rect 12790 -1360 12810 -1300
rect 12710 -1380 12810 -1360
rect 12880 -1000 12980 -980
rect 12880 -1060 12900 -1000
rect 12960 -1060 12980 -1000
rect 12880 -1100 12980 -1060
rect 12880 -1160 12900 -1100
rect 12960 -1160 12980 -1100
rect 12880 -1200 12980 -1160
rect 12880 -1260 12900 -1200
rect 12960 -1260 12980 -1200
rect 12880 -1300 12980 -1260
rect 12880 -1360 12900 -1300
rect 12960 -1360 12980 -1300
rect 12880 -1380 12980 -1360
rect 13050 -1000 13150 -980
rect 13050 -1060 13070 -1000
rect 13130 -1060 13150 -1000
rect 13050 -1100 13150 -1060
rect 13050 -1160 13070 -1100
rect 13130 -1160 13150 -1100
rect 13050 -1200 13150 -1160
rect 13050 -1260 13070 -1200
rect 13130 -1260 13150 -1200
rect 13050 -1300 13150 -1260
rect 13050 -1360 13070 -1300
rect 13130 -1360 13150 -1300
rect 13050 -1380 13150 -1360
rect 13220 -1000 13320 -980
rect 13220 -1060 13240 -1000
rect 13300 -1060 13320 -1000
rect 13220 -1100 13320 -1060
rect 13220 -1160 13240 -1100
rect 13300 -1160 13320 -1100
rect 13220 -1200 13320 -1160
rect 13220 -1260 13240 -1200
rect 13300 -1260 13320 -1200
rect 13220 -1300 13320 -1260
rect 13220 -1360 13240 -1300
rect 13300 -1360 13320 -1300
rect 13220 -1380 13320 -1360
rect 13390 -1000 13490 -980
rect 13390 -1060 13410 -1000
rect 13470 -1060 13490 -1000
rect 13390 -1100 13490 -1060
rect 13390 -1160 13410 -1100
rect 13470 -1160 13490 -1100
rect 13390 -1200 13490 -1160
rect 13390 -1260 13410 -1200
rect 13470 -1260 13490 -1200
rect 13390 -1300 13490 -1260
rect 13390 -1360 13410 -1300
rect 13470 -1360 13490 -1300
rect 13390 -1380 13490 -1360
rect 13560 -1000 13660 -980
rect 13560 -1060 13580 -1000
rect 13640 -1060 13660 -1000
rect 13560 -1100 13660 -1060
rect 13560 -1160 13580 -1100
rect 13640 -1160 13660 -1100
rect 13560 -1200 13660 -1160
rect 13560 -1260 13580 -1200
rect 13640 -1260 13660 -1200
rect 13560 -1300 13660 -1260
rect 13560 -1360 13580 -1300
rect 13640 -1360 13660 -1300
rect 13560 -1380 13660 -1360
rect 13730 -1000 13830 -980
rect 13730 -1060 13750 -1000
rect 13810 -1060 13830 -1000
rect 13730 -1100 13830 -1060
rect 13730 -1160 13750 -1100
rect 13810 -1160 13830 -1100
rect 13730 -1200 13830 -1160
rect 13730 -1260 13750 -1200
rect 13810 -1260 13830 -1200
rect 13730 -1300 13830 -1260
rect 13730 -1360 13750 -1300
rect 13810 -1360 13830 -1300
rect 13730 -1380 13830 -1360
rect 13900 -1000 14000 -980
rect 13900 -1060 13920 -1000
rect 13980 -1060 14000 -1000
rect 13900 -1100 14000 -1060
rect 13900 -1160 13920 -1100
rect 13980 -1160 14000 -1100
rect 13900 -1200 14000 -1160
rect 13900 -1260 13920 -1200
rect 13980 -1260 14000 -1200
rect 13900 -1300 14000 -1260
rect 13900 -1360 13920 -1300
rect 13980 -1360 14000 -1300
rect 13900 -1380 14000 -1360
rect 14070 -1000 14170 -980
rect 14070 -1060 14090 -1000
rect 14150 -1060 14170 -1000
rect 14070 -1100 14170 -1060
rect 14070 -1160 14090 -1100
rect 14150 -1160 14170 -1100
rect 14070 -1200 14170 -1160
rect 14070 -1260 14090 -1200
rect 14150 -1260 14170 -1200
rect 14070 -1300 14170 -1260
rect 14070 -1360 14090 -1300
rect 14150 -1360 14170 -1300
rect 14070 -1380 14170 -1360
rect 14240 -1000 14340 -980
rect 14240 -1060 14260 -1000
rect 14320 -1060 14340 -1000
rect 14240 -1100 14340 -1060
rect 14240 -1160 14260 -1100
rect 14320 -1160 14340 -1100
rect 14240 -1200 14340 -1160
rect 14240 -1260 14260 -1200
rect 14320 -1260 14340 -1200
rect 14240 -1300 14340 -1260
rect 14240 -1360 14260 -1300
rect 14320 -1360 14340 -1300
rect 14240 -1380 14340 -1360
rect 14410 -1000 14510 -980
rect 14410 -1060 14430 -1000
rect 14490 -1060 14510 -1000
rect 14410 -1100 14510 -1060
rect 14410 -1160 14430 -1100
rect 14490 -1160 14510 -1100
rect 14410 -1200 14510 -1160
rect 14410 -1260 14430 -1200
rect 14490 -1260 14510 -1200
rect 14410 -1300 14510 -1260
rect 14410 -1360 14430 -1300
rect 14490 -1360 14510 -1300
rect 14410 -1380 14510 -1360
rect 14580 -1000 14680 -980
rect 14580 -1060 14600 -1000
rect 14660 -1060 14680 -1000
rect 14580 -1100 14680 -1060
rect 14580 -1160 14600 -1100
rect 14660 -1160 14680 -1100
rect 14580 -1200 14680 -1160
rect 14580 -1260 14600 -1200
rect 14660 -1260 14680 -1200
rect 14580 -1300 14680 -1260
rect 14580 -1360 14600 -1300
rect 14660 -1360 14680 -1300
rect 14580 -1380 14680 -1360
rect 14750 -1000 14850 -980
rect 14750 -1060 14770 -1000
rect 14830 -1060 14850 -1000
rect 14750 -1100 14850 -1060
rect 14750 -1160 14770 -1100
rect 14830 -1160 14850 -1100
rect 14750 -1200 14850 -1160
rect 14750 -1260 14770 -1200
rect 14830 -1260 14850 -1200
rect 14750 -1300 14850 -1260
rect 14750 -1360 14770 -1300
rect 14830 -1360 14850 -1300
rect 14750 -1380 14850 -1360
rect 14920 -1000 15020 -980
rect 14920 -1060 14940 -1000
rect 15000 -1060 15020 -1000
rect 14920 -1100 15020 -1060
rect 14920 -1160 14940 -1100
rect 15000 -1160 15020 -1100
rect 14920 -1200 15020 -1160
rect 14920 -1260 14940 -1200
rect 15000 -1260 15020 -1200
rect 14920 -1300 15020 -1260
rect 14920 -1360 14940 -1300
rect 15000 -1360 15020 -1300
rect 14920 -1380 15020 -1360
rect 15090 -1000 15190 -980
rect 15090 -1060 15110 -1000
rect 15170 -1060 15190 -1000
rect 15090 -1100 15190 -1060
rect 15090 -1160 15110 -1100
rect 15170 -1160 15190 -1100
rect 15090 -1200 15190 -1160
rect 15090 -1260 15110 -1200
rect 15170 -1260 15190 -1200
rect 15090 -1300 15190 -1260
rect 15090 -1360 15110 -1300
rect 15170 -1360 15190 -1300
rect 15090 -1380 15190 -1360
rect 15260 -1000 15360 -980
rect 15260 -1060 15280 -1000
rect 15340 -1060 15360 -1000
rect 15260 -1100 15360 -1060
rect 15260 -1160 15280 -1100
rect 15340 -1160 15360 -1100
rect 15260 -1200 15360 -1160
rect 15260 -1260 15280 -1200
rect 15340 -1260 15360 -1200
rect 15260 -1300 15360 -1260
rect 15260 -1360 15280 -1300
rect 15340 -1360 15360 -1300
rect 15260 -1380 15360 -1360
rect 15430 -1000 15530 -980
rect 15430 -1060 15450 -1000
rect 15510 -1060 15530 -1000
rect 15430 -1100 15530 -1060
rect 15430 -1160 15450 -1100
rect 15510 -1160 15530 -1100
rect 15430 -1200 15530 -1160
rect 15430 -1260 15450 -1200
rect 15510 -1260 15530 -1200
rect 15430 -1300 15530 -1260
rect 15430 -1360 15450 -1300
rect 15510 -1360 15530 -1300
rect 15430 -1380 15530 -1360
rect 15600 -1000 15700 -980
rect 15600 -1060 15620 -1000
rect 15680 -1060 15700 -1000
rect 15600 -1100 15700 -1060
rect 15600 -1160 15620 -1100
rect 15680 -1160 15700 -1100
rect 15600 -1200 15700 -1160
rect 15600 -1260 15620 -1200
rect 15680 -1260 15700 -1200
rect 15600 -1300 15700 -1260
rect 15600 -1360 15620 -1300
rect 15680 -1360 15700 -1300
rect 15600 -1380 15700 -1360
rect 15770 -1000 15870 -980
rect 15770 -1060 15790 -1000
rect 15850 -1060 15870 -1000
rect 15770 -1100 15870 -1060
rect 15770 -1160 15790 -1100
rect 15850 -1160 15870 -1100
rect 15770 -1200 15870 -1160
rect 15770 -1260 15790 -1200
rect 15850 -1260 15870 -1200
rect 15770 -1300 15870 -1260
rect 15770 -1360 15790 -1300
rect 15850 -1360 15870 -1300
rect 15770 -1380 15870 -1360
rect 15940 -1000 16040 -980
rect 15940 -1060 15960 -1000
rect 16020 -1060 16040 -1000
rect 15940 -1100 16040 -1060
rect 15940 -1160 15960 -1100
rect 16020 -1160 16040 -1100
rect 15940 -1200 16040 -1160
rect 15940 -1260 15960 -1200
rect 16020 -1260 16040 -1200
rect 15940 -1300 16040 -1260
rect 15940 -1360 15960 -1300
rect 16020 -1360 16040 -1300
rect 15940 -1380 16040 -1360
rect 16110 -1000 16210 -980
rect 16110 -1060 16130 -1000
rect 16190 -1060 16210 -1000
rect 16110 -1100 16210 -1060
rect 16110 -1160 16130 -1100
rect 16190 -1160 16210 -1100
rect 16110 -1200 16210 -1160
rect 16110 -1260 16130 -1200
rect 16190 -1260 16210 -1200
rect 16110 -1300 16210 -1260
rect 16110 -1360 16130 -1300
rect 16190 -1360 16210 -1300
rect 16110 -1380 16210 -1360
rect 16280 -1000 16380 -980
rect 16280 -1060 16300 -1000
rect 16360 -1060 16380 -1000
rect 16280 -1100 16380 -1060
rect 16280 -1160 16300 -1100
rect 16360 -1160 16380 -1100
rect 16280 -1200 16380 -1160
rect 16280 -1260 16300 -1200
rect 16360 -1260 16380 -1200
rect 16280 -1300 16380 -1260
rect 16280 -1360 16300 -1300
rect 16360 -1360 16380 -1300
rect 16280 -1380 16380 -1360
rect 16450 -1000 16550 -980
rect 16450 -1060 16470 -1000
rect 16530 -1060 16550 -1000
rect 16450 -1100 16550 -1060
rect 16450 -1160 16470 -1100
rect 16530 -1160 16550 -1100
rect 16450 -1200 16550 -1160
rect 16450 -1260 16470 -1200
rect 16530 -1260 16550 -1200
rect 16450 -1300 16550 -1260
rect 16450 -1360 16470 -1300
rect 16530 -1360 16550 -1300
rect 16450 -1380 16550 -1360
rect 16620 -1000 16720 -980
rect 16620 -1060 16640 -1000
rect 16700 -1060 16720 -1000
rect 16620 -1100 16720 -1060
rect 16620 -1160 16640 -1100
rect 16700 -1160 16720 -1100
rect 16620 -1200 16720 -1160
rect 16620 -1260 16640 -1200
rect 16700 -1260 16720 -1200
rect 16620 -1300 16720 -1260
rect 16620 -1360 16640 -1300
rect 16700 -1360 16720 -1300
rect 16620 -1380 16720 -1360
rect 16790 -1000 16890 -980
rect 16790 -1060 16810 -1000
rect 16870 -1060 16890 -1000
rect 16790 -1100 16890 -1060
rect 16790 -1160 16810 -1100
rect 16870 -1160 16890 -1100
rect 16790 -1200 16890 -1160
rect 16790 -1260 16810 -1200
rect 16870 -1260 16890 -1200
rect 16790 -1300 16890 -1260
rect 16790 -1360 16810 -1300
rect 16870 -1360 16890 -1300
rect 16790 -1380 16890 -1360
rect 16960 -1000 17060 -980
rect 16960 -1060 16980 -1000
rect 17040 -1060 17060 -1000
rect 16960 -1100 17060 -1060
rect 16960 -1160 16980 -1100
rect 17040 -1160 17060 -1100
rect 16960 -1200 17060 -1160
rect 16960 -1260 16980 -1200
rect 17040 -1260 17060 -1200
rect 16960 -1300 17060 -1260
rect 16960 -1360 16980 -1300
rect 17040 -1360 17060 -1300
rect 16960 -1380 17060 -1360
rect 17130 -1000 17230 -980
rect 17130 -1060 17150 -1000
rect 17210 -1060 17230 -1000
rect 17130 -1100 17230 -1060
rect 17130 -1160 17150 -1100
rect 17210 -1160 17230 -1100
rect 17130 -1200 17230 -1160
rect 17130 -1260 17150 -1200
rect 17210 -1260 17230 -1200
rect 17130 -1300 17230 -1260
rect 17130 -1360 17150 -1300
rect 17210 -1360 17230 -1300
rect 17130 -1380 17230 -1360
rect 17300 -1000 17400 -980
rect 17300 -1060 17320 -1000
rect 17380 -1060 17400 -1000
rect 17300 -1100 17400 -1060
rect 17300 -1160 17320 -1100
rect 17380 -1160 17400 -1100
rect 17300 -1200 17400 -1160
rect 17300 -1260 17320 -1200
rect 17380 -1260 17400 -1200
rect 17300 -1300 17400 -1260
rect 17300 -1360 17320 -1300
rect 17380 -1360 17400 -1300
rect 17300 -1380 17400 -1360
rect 17470 -1000 17570 -980
rect 17470 -1060 17490 -1000
rect 17550 -1060 17570 -1000
rect 17470 -1100 17570 -1060
rect 17470 -1160 17490 -1100
rect 17550 -1160 17570 -1100
rect 17470 -1200 17570 -1160
rect 17470 -1260 17490 -1200
rect 17550 -1260 17570 -1200
rect 17470 -1300 17570 -1260
rect 17470 -1360 17490 -1300
rect 17550 -1360 17570 -1300
rect 17470 -1380 17570 -1360
rect 17640 -1000 17740 -980
rect 17640 -1060 17660 -1000
rect 17720 -1060 17740 -1000
rect 17640 -1100 17740 -1060
rect 17640 -1160 17660 -1100
rect 17720 -1160 17740 -1100
rect 17640 -1200 17740 -1160
rect 17640 -1260 17660 -1200
rect 17720 -1260 17740 -1200
rect 17640 -1300 17740 -1260
rect 17640 -1360 17660 -1300
rect 17720 -1360 17740 -1300
rect 17640 -1380 17740 -1360
rect 17810 -1000 17910 -980
rect 17810 -1060 17830 -1000
rect 17890 -1060 17910 -1000
rect 17810 -1100 17910 -1060
rect 17810 -1160 17830 -1100
rect 17890 -1160 17910 -1100
rect 17810 -1200 17910 -1160
rect 17810 -1260 17830 -1200
rect 17890 -1260 17910 -1200
rect 17810 -1300 17910 -1260
rect 17810 -1360 17830 -1300
rect 17890 -1360 17910 -1300
rect 17810 -1380 17910 -1360
rect 17980 -1000 18080 -980
rect 17980 -1060 18000 -1000
rect 18060 -1060 18080 -1000
rect 17980 -1100 18080 -1060
rect 17980 -1160 18000 -1100
rect 18060 -1160 18080 -1100
rect 17980 -1200 18080 -1160
rect 17980 -1260 18000 -1200
rect 18060 -1260 18080 -1200
rect 17980 -1300 18080 -1260
rect 17980 -1360 18000 -1300
rect 18060 -1360 18080 -1300
rect 17980 -1380 18080 -1360
rect 18150 -1000 18250 -980
rect 18150 -1060 18170 -1000
rect 18230 -1060 18250 -1000
rect 18150 -1100 18250 -1060
rect 18150 -1160 18170 -1100
rect 18230 -1160 18250 -1100
rect 18150 -1200 18250 -1160
rect 18150 -1260 18170 -1200
rect 18230 -1260 18250 -1200
rect 18150 -1300 18250 -1260
rect 18150 -1360 18170 -1300
rect 18230 -1360 18250 -1300
rect 18150 -1380 18250 -1360
rect 18320 -1000 18420 -980
rect 18320 -1060 18340 -1000
rect 18400 -1060 18420 -1000
rect 18320 -1100 18420 -1060
rect 18320 -1160 18340 -1100
rect 18400 -1160 18420 -1100
rect 18320 -1200 18420 -1160
rect 18320 -1260 18340 -1200
rect 18400 -1260 18420 -1200
rect 18320 -1300 18420 -1260
rect 18320 -1360 18340 -1300
rect 18400 -1360 18420 -1300
rect 18320 -1380 18420 -1360
rect 18490 -1000 18590 -980
rect 18490 -1060 18510 -1000
rect 18570 -1060 18590 -1000
rect 18490 -1100 18590 -1060
rect 18490 -1160 18510 -1100
rect 18570 -1160 18590 -1100
rect 18490 -1200 18590 -1160
rect 18490 -1260 18510 -1200
rect 18570 -1260 18590 -1200
rect 18490 -1300 18590 -1260
rect 18490 -1360 18510 -1300
rect 18570 -1360 18590 -1300
rect 18490 -1380 18590 -1360
rect 18660 -1000 18760 -980
rect 18660 -1060 18680 -1000
rect 18740 -1060 18760 -1000
rect 18660 -1100 18760 -1060
rect 18660 -1160 18680 -1100
rect 18740 -1160 18760 -1100
rect 18660 -1200 18760 -1160
rect 18660 -1260 18680 -1200
rect 18740 -1260 18760 -1200
rect 18660 -1300 18760 -1260
rect 18660 -1360 18680 -1300
rect 18740 -1360 18760 -1300
rect 18660 -1380 18760 -1360
rect 18830 -1000 18930 -980
rect 18830 -1060 18850 -1000
rect 18910 -1060 18930 -1000
rect 18830 -1100 18930 -1060
rect 18830 -1160 18850 -1100
rect 18910 -1160 18930 -1100
rect 18830 -1200 18930 -1160
rect 18830 -1260 18850 -1200
rect 18910 -1260 18930 -1200
rect 18830 -1300 18930 -1260
rect 18830 -1360 18850 -1300
rect 18910 -1360 18930 -1300
rect 18830 -1380 18930 -1360
rect 19000 -1000 19100 -980
rect 19000 -1060 19020 -1000
rect 19080 -1060 19100 -1000
rect 19000 -1100 19100 -1060
rect 19000 -1160 19020 -1100
rect 19080 -1160 19100 -1100
rect 19000 -1200 19100 -1160
rect 19000 -1260 19020 -1200
rect 19080 -1260 19100 -1200
rect 19000 -1300 19100 -1260
rect 19000 -1360 19020 -1300
rect 19080 -1360 19100 -1300
rect 19000 -1380 19100 -1360
rect 19170 -1000 19270 -980
rect 19170 -1060 19190 -1000
rect 19250 -1060 19270 -1000
rect 19170 -1100 19270 -1060
rect 19170 -1160 19190 -1100
rect 19250 -1160 19270 -1100
rect 19170 -1200 19270 -1160
rect 19170 -1260 19190 -1200
rect 19250 -1260 19270 -1200
rect 19170 -1300 19270 -1260
rect 19170 -1360 19190 -1300
rect 19250 -1360 19270 -1300
rect 19170 -1380 19270 -1360
rect 19340 -1000 19440 -980
rect 19340 -1060 19360 -1000
rect 19420 -1060 19440 -1000
rect 19340 -1100 19440 -1060
rect 19340 -1160 19360 -1100
rect 19420 -1160 19440 -1100
rect 19340 -1200 19440 -1160
rect 19340 -1260 19360 -1200
rect 19420 -1260 19440 -1200
rect 19340 -1300 19440 -1260
rect 19340 -1360 19360 -1300
rect 19420 -1360 19440 -1300
rect 19340 -1380 19440 -1360
rect 19510 -1000 19610 -980
rect 19510 -1060 19530 -1000
rect 19590 -1060 19610 -1000
rect 19510 -1100 19610 -1060
rect 19510 -1160 19530 -1100
rect 19590 -1160 19610 -1100
rect 19510 -1200 19610 -1160
rect 19510 -1260 19530 -1200
rect 19590 -1260 19610 -1200
rect 19510 -1300 19610 -1260
rect 19510 -1360 19530 -1300
rect 19590 -1360 19610 -1300
rect 19510 -1380 19610 -1360
rect 19680 -1000 19780 -980
rect 19680 -1060 19700 -1000
rect 19760 -1060 19780 -1000
rect 19680 -1100 19780 -1060
rect 19680 -1160 19700 -1100
rect 19760 -1160 19780 -1100
rect 19680 -1200 19780 -1160
rect 19680 -1260 19700 -1200
rect 19760 -1260 19780 -1200
rect 19680 -1300 19780 -1260
rect 19680 -1360 19700 -1300
rect 19760 -1360 19780 -1300
rect 19680 -1380 19780 -1360
rect 19850 -1000 19950 -980
rect 19850 -1060 19870 -1000
rect 19930 -1060 19950 -1000
rect 19850 -1100 19950 -1060
rect 19850 -1160 19870 -1100
rect 19930 -1160 19950 -1100
rect 19850 -1200 19950 -1160
rect 19850 -1260 19870 -1200
rect 19930 -1260 19950 -1200
rect 19850 -1300 19950 -1260
rect 19850 -1360 19870 -1300
rect 19930 -1360 19950 -1300
rect 19850 -1380 19950 -1360
rect 20020 -1000 20120 -980
rect 20020 -1060 20040 -1000
rect 20100 -1060 20120 -1000
rect 20020 -1100 20120 -1060
rect 20020 -1160 20040 -1100
rect 20100 -1160 20120 -1100
rect 20020 -1200 20120 -1160
rect 20020 -1260 20040 -1200
rect 20100 -1260 20120 -1200
rect 20020 -1300 20120 -1260
rect 20020 -1360 20040 -1300
rect 20100 -1360 20120 -1300
rect 20020 -1380 20120 -1360
rect 20190 -1000 20290 -980
rect 20190 -1060 20210 -1000
rect 20270 -1060 20290 -1000
rect 20190 -1100 20290 -1060
rect 20190 -1160 20210 -1100
rect 20270 -1160 20290 -1100
rect 20190 -1200 20290 -1160
rect 20190 -1260 20210 -1200
rect 20270 -1260 20290 -1200
rect 20190 -1300 20290 -1260
rect 20190 -1360 20210 -1300
rect 20270 -1360 20290 -1300
rect 20190 -1380 20290 -1360
rect 20360 -1000 20460 -980
rect 20360 -1060 20380 -1000
rect 20440 -1060 20460 -1000
rect 20360 -1100 20460 -1060
rect 20360 -1160 20380 -1100
rect 20440 -1160 20460 -1100
rect 20360 -1200 20460 -1160
rect 20360 -1260 20380 -1200
rect 20440 -1260 20460 -1200
rect 20360 -1300 20460 -1260
rect 20360 -1360 20380 -1300
rect 20440 -1360 20460 -1300
rect 20360 -1380 20460 -1360
rect 20530 -1000 20630 -980
rect 20530 -1060 20550 -1000
rect 20610 -1060 20630 -1000
rect 20530 -1100 20630 -1060
rect 20530 -1160 20550 -1100
rect 20610 -1160 20630 -1100
rect 20530 -1200 20630 -1160
rect 20530 -1260 20550 -1200
rect 20610 -1260 20630 -1200
rect 20530 -1300 20630 -1260
rect 20530 -1360 20550 -1300
rect 20610 -1360 20630 -1300
rect 20530 -1380 20630 -1360
rect 20700 -1000 20800 -980
rect 20700 -1060 20720 -1000
rect 20780 -1060 20800 -1000
rect 20700 -1100 20800 -1060
rect 20700 -1160 20720 -1100
rect 20780 -1160 20800 -1100
rect 20700 -1200 20800 -1160
rect 20700 -1260 20720 -1200
rect 20780 -1260 20800 -1200
rect 20700 -1300 20800 -1260
rect 20700 -1360 20720 -1300
rect 20780 -1360 20800 -1300
rect 20700 -1380 20800 -1360
rect 20870 -1000 20970 -980
rect 20870 -1060 20890 -1000
rect 20950 -1060 20970 -1000
rect 20870 -1100 20970 -1060
rect 20870 -1160 20890 -1100
rect 20950 -1160 20970 -1100
rect 20870 -1200 20970 -1160
rect 20870 -1260 20890 -1200
rect 20950 -1260 20970 -1200
rect 20870 -1300 20970 -1260
rect 20870 -1360 20890 -1300
rect 20950 -1360 20970 -1300
rect 20870 -1380 20970 -1360
rect 21040 -1000 21140 -980
rect 21040 -1060 21060 -1000
rect 21120 -1060 21140 -1000
rect 21040 -1100 21140 -1060
rect 21040 -1160 21060 -1100
rect 21120 -1160 21140 -1100
rect 21040 -1200 21140 -1160
rect 21040 -1260 21060 -1200
rect 21120 -1260 21140 -1200
rect 21040 -1300 21140 -1260
rect 21040 -1360 21060 -1300
rect 21120 -1360 21140 -1300
rect 21040 -1380 21140 -1360
rect 21210 -1000 21310 -980
rect 21210 -1060 21230 -1000
rect 21290 -1060 21310 -1000
rect 21210 -1100 21310 -1060
rect 21210 -1160 21230 -1100
rect 21290 -1160 21310 -1100
rect 21210 -1200 21310 -1160
rect 21210 -1260 21230 -1200
rect 21290 -1260 21310 -1200
rect 21210 -1300 21310 -1260
rect 21210 -1360 21230 -1300
rect 21290 -1360 21310 -1300
rect 21210 -1380 21310 -1360
rect 21380 -1000 21480 -980
rect 21380 -1060 21400 -1000
rect 21460 -1060 21480 -1000
rect 21380 -1100 21480 -1060
rect 21380 -1160 21400 -1100
rect 21460 -1160 21480 -1100
rect 21380 -1200 21480 -1160
rect 21380 -1260 21400 -1200
rect 21460 -1260 21480 -1200
rect 21380 -1300 21480 -1260
rect 21380 -1360 21400 -1300
rect 21460 -1360 21480 -1300
rect 21380 -1380 21480 -1360
rect 21550 -1000 21650 -980
rect 21550 -1060 21570 -1000
rect 21630 -1060 21650 -1000
rect 21550 -1100 21650 -1060
rect 21550 -1160 21570 -1100
rect 21630 -1160 21650 -1100
rect 21550 -1200 21650 -1160
rect 21550 -1260 21570 -1200
rect 21630 -1260 21650 -1200
rect 21550 -1300 21650 -1260
rect 21550 -1360 21570 -1300
rect 21630 -1360 21650 -1300
rect 21550 -1380 21650 -1360
rect 21720 -1000 21820 -980
rect 21720 -1060 21740 -1000
rect 21800 -1060 21820 -1000
rect 21720 -1100 21820 -1060
rect 21720 -1160 21740 -1100
rect 21800 -1160 21820 -1100
rect 21720 -1200 21820 -1160
rect 21720 -1260 21740 -1200
rect 21800 -1260 21820 -1200
rect 21720 -1300 21820 -1260
rect 21720 -1360 21740 -1300
rect 21800 -1360 21820 -1300
rect 21720 -1380 21820 -1360
rect 21890 -1000 21990 -980
rect 21890 -1060 21910 -1000
rect 21970 -1060 21990 -1000
rect 21890 -1100 21990 -1060
rect 21890 -1160 21910 -1100
rect 21970 -1160 21990 -1100
rect 21890 -1200 21990 -1160
rect 21890 -1260 21910 -1200
rect 21970 -1260 21990 -1200
rect 21890 -1300 21990 -1260
rect 21890 -1360 21910 -1300
rect 21970 -1360 21990 -1300
rect 21890 -1380 21990 -1360
rect 22060 -1000 22160 -980
rect 22060 -1060 22080 -1000
rect 22140 -1060 22160 -1000
rect 22060 -1100 22160 -1060
rect 22060 -1160 22080 -1100
rect 22140 -1160 22160 -1100
rect 22060 -1200 22160 -1160
rect 22060 -1260 22080 -1200
rect 22140 -1260 22160 -1200
rect 22060 -1300 22160 -1260
rect 22060 -1360 22080 -1300
rect 22140 -1360 22160 -1300
rect 22060 -1380 22160 -1360
rect 22230 -1000 22330 -980
rect 22230 -1060 22250 -1000
rect 22310 -1060 22330 -1000
rect 22230 -1100 22330 -1060
rect 22230 -1160 22250 -1100
rect 22310 -1160 22330 -1100
rect 22230 -1200 22330 -1160
rect 22230 -1260 22250 -1200
rect 22310 -1260 22330 -1200
rect 22230 -1300 22330 -1260
rect 22230 -1360 22250 -1300
rect 22310 -1360 22330 -1300
rect 22230 -1380 22330 -1360
rect 22400 -1000 22500 -980
rect 22400 -1060 22420 -1000
rect 22480 -1060 22500 -1000
rect 22400 -1100 22500 -1060
rect 22400 -1160 22420 -1100
rect 22480 -1160 22500 -1100
rect 22400 -1200 22500 -1160
rect 22400 -1260 22420 -1200
rect 22480 -1260 22500 -1200
rect 22400 -1300 22500 -1260
rect 22400 -1360 22420 -1300
rect 22480 -1360 22500 -1300
rect 22400 -1380 22500 -1360
rect 22570 -1000 22670 -980
rect 22570 -1060 22590 -1000
rect 22650 -1060 22670 -1000
rect 22570 -1100 22670 -1060
rect 22570 -1160 22590 -1100
rect 22650 -1160 22670 -1100
rect 22570 -1200 22670 -1160
rect 22570 -1260 22590 -1200
rect 22650 -1260 22670 -1200
rect 22570 -1300 22670 -1260
rect 22570 -1360 22590 -1300
rect 22650 -1360 22670 -1300
rect 22570 -1380 22670 -1360
rect 22740 -1000 22840 -980
rect 22740 -1060 22760 -1000
rect 22820 -1060 22840 -1000
rect 22740 -1100 22840 -1060
rect 22740 -1160 22760 -1100
rect 22820 -1160 22840 -1100
rect 22740 -1200 22840 -1160
rect 22740 -1260 22760 -1200
rect 22820 -1260 22840 -1200
rect 22740 -1300 22840 -1260
rect 22740 -1360 22760 -1300
rect 22820 -1360 22840 -1300
rect 22740 -1380 22840 -1360
rect 22910 -1000 23010 -980
rect 22910 -1060 22930 -1000
rect 22990 -1060 23010 -1000
rect 22910 -1100 23010 -1060
rect 22910 -1160 22930 -1100
rect 22990 -1160 23010 -1100
rect 22910 -1200 23010 -1160
rect 22910 -1260 22930 -1200
rect 22990 -1260 23010 -1200
rect 22910 -1300 23010 -1260
rect 22910 -1360 22930 -1300
rect 22990 -1360 23010 -1300
rect 22910 -1380 23010 -1360
rect 23080 -1000 23180 -980
rect 23080 -1060 23100 -1000
rect 23160 -1060 23180 -1000
rect 23080 -1100 23180 -1060
rect 23080 -1160 23100 -1100
rect 23160 -1160 23180 -1100
rect 23080 -1200 23180 -1160
rect 23080 -1260 23100 -1200
rect 23160 -1260 23180 -1200
rect 23080 -1300 23180 -1260
rect 23080 -1360 23100 -1300
rect 23160 -1360 23180 -1300
rect 23080 -1380 23180 -1360
rect 23250 -1000 23350 -980
rect 23250 -1060 23270 -1000
rect 23330 -1060 23350 -1000
rect 23250 -1100 23350 -1060
rect 23250 -1160 23270 -1100
rect 23330 -1160 23350 -1100
rect 23250 -1200 23350 -1160
rect 23250 -1260 23270 -1200
rect 23330 -1260 23350 -1200
rect 23250 -1300 23350 -1260
rect 23250 -1360 23270 -1300
rect 23330 -1360 23350 -1300
rect 23250 -1380 23350 -1360
rect 23420 -1000 23520 -980
rect 23420 -1060 23440 -1000
rect 23500 -1060 23520 -1000
rect 23420 -1100 23520 -1060
rect 23420 -1160 23440 -1100
rect 23500 -1160 23520 -1100
rect 23420 -1200 23520 -1160
rect 23420 -1260 23440 -1200
rect 23500 -1260 23520 -1200
rect 23420 -1300 23520 -1260
rect 23420 -1360 23440 -1300
rect 23500 -1360 23520 -1300
rect 23420 -1380 23520 -1360
rect 23590 -1000 23690 -980
rect 23590 -1060 23610 -1000
rect 23670 -1060 23690 -1000
rect 23590 -1100 23690 -1060
rect 23590 -1160 23610 -1100
rect 23670 -1160 23690 -1100
rect 23590 -1200 23690 -1160
rect 23590 -1260 23610 -1200
rect 23670 -1260 23690 -1200
rect 23590 -1300 23690 -1260
rect 23590 -1360 23610 -1300
rect 23670 -1360 23690 -1300
rect 23590 -1380 23690 -1360
rect 23760 -1000 23860 -980
rect 23760 -1060 23780 -1000
rect 23840 -1060 23860 -1000
rect 23760 -1100 23860 -1060
rect 23760 -1160 23780 -1100
rect 23840 -1160 23860 -1100
rect 23760 -1200 23860 -1160
rect 23760 -1260 23780 -1200
rect 23840 -1260 23860 -1200
rect 23760 -1300 23860 -1260
rect 23760 -1360 23780 -1300
rect 23840 -1360 23860 -1300
rect 23760 -1380 23860 -1360
rect 23930 -1000 24030 -980
rect 23930 -1060 23950 -1000
rect 24010 -1060 24030 -1000
rect 23930 -1100 24030 -1060
rect 23930 -1160 23950 -1100
rect 24010 -1160 24030 -1100
rect 23930 -1200 24030 -1160
rect 23930 -1260 23950 -1200
rect 24010 -1260 24030 -1200
rect 23930 -1300 24030 -1260
rect 23930 -1360 23950 -1300
rect 24010 -1360 24030 -1300
rect 23930 -1380 24030 -1360
rect 24100 -1000 24200 -980
rect 24100 -1060 24120 -1000
rect 24180 -1060 24200 -1000
rect 24100 -1100 24200 -1060
rect 24100 -1160 24120 -1100
rect 24180 -1160 24200 -1100
rect 24100 -1200 24200 -1160
rect 24100 -1260 24120 -1200
rect 24180 -1260 24200 -1200
rect 24100 -1300 24200 -1260
rect 24100 -1360 24120 -1300
rect 24180 -1360 24200 -1300
rect 24100 -1380 24200 -1360
rect 24270 -1000 24370 -980
rect 24270 -1060 24290 -1000
rect 24350 -1060 24370 -1000
rect 24270 -1100 24370 -1060
rect 24270 -1160 24290 -1100
rect 24350 -1160 24370 -1100
rect 24270 -1200 24370 -1160
rect 24270 -1260 24290 -1200
rect 24350 -1260 24370 -1200
rect 24270 -1300 24370 -1260
rect 24270 -1360 24290 -1300
rect 24350 -1360 24370 -1300
rect 24270 -1380 24370 -1360
rect 24440 -1000 24540 -980
rect 24440 -1060 24460 -1000
rect 24520 -1060 24540 -1000
rect 24440 -1100 24540 -1060
rect 24440 -1160 24460 -1100
rect 24520 -1160 24540 -1100
rect 24440 -1200 24540 -1160
rect 24440 -1260 24460 -1200
rect 24520 -1260 24540 -1200
rect 24440 -1300 24540 -1260
rect 24440 -1360 24460 -1300
rect 24520 -1360 24540 -1300
rect 24440 -1380 24540 -1360
rect 24610 -1000 24710 -980
rect 24610 -1060 24630 -1000
rect 24690 -1060 24710 -1000
rect 24610 -1100 24710 -1060
rect 24610 -1160 24630 -1100
rect 24690 -1160 24710 -1100
rect 24610 -1200 24710 -1160
rect 24610 -1260 24630 -1200
rect 24690 -1260 24710 -1200
rect 24610 -1300 24710 -1260
rect 24610 -1360 24630 -1300
rect 24690 -1360 24710 -1300
rect 24610 -1380 24710 -1360
rect 24780 -1000 24880 -980
rect 24780 -1060 24800 -1000
rect 24860 -1060 24880 -1000
rect 24780 -1100 24880 -1060
rect 24780 -1160 24800 -1100
rect 24860 -1160 24880 -1100
rect 24780 -1200 24880 -1160
rect 24780 -1260 24800 -1200
rect 24860 -1260 24880 -1200
rect 24780 -1300 24880 -1260
rect 24780 -1360 24800 -1300
rect 24860 -1360 24880 -1300
rect 24780 -1380 24880 -1360
rect 24950 -1000 25050 -980
rect 24950 -1060 24970 -1000
rect 25030 -1060 25050 -1000
rect 24950 -1100 25050 -1060
rect 24950 -1160 24970 -1100
rect 25030 -1160 25050 -1100
rect 24950 -1200 25050 -1160
rect 24950 -1260 24970 -1200
rect 25030 -1260 25050 -1200
rect 24950 -1300 25050 -1260
rect 24950 -1360 24970 -1300
rect 25030 -1360 25050 -1300
rect 24950 -1380 25050 -1360
rect 25120 -1000 25220 -980
rect 25120 -1060 25140 -1000
rect 25200 -1060 25220 -1000
rect 25120 -1100 25220 -1060
rect 25120 -1160 25140 -1100
rect 25200 -1160 25220 -1100
rect 25120 -1200 25220 -1160
rect 25120 -1260 25140 -1200
rect 25200 -1260 25220 -1200
rect 25120 -1300 25220 -1260
rect 25120 -1360 25140 -1300
rect 25200 -1360 25220 -1300
rect 25120 -1380 25220 -1360
rect 25290 -1000 25390 -980
rect 25290 -1060 25310 -1000
rect 25370 -1060 25390 -1000
rect 25290 -1100 25390 -1060
rect 25290 -1160 25310 -1100
rect 25370 -1160 25390 -1100
rect 25290 -1200 25390 -1160
rect 25290 -1260 25310 -1200
rect 25370 -1260 25390 -1200
rect 25290 -1300 25390 -1260
rect 25290 -1360 25310 -1300
rect 25370 -1360 25390 -1300
rect 25290 -1380 25390 -1360
rect 25460 -1000 25560 -980
rect 25460 -1060 25480 -1000
rect 25540 -1060 25560 -1000
rect 25460 -1100 25560 -1060
rect 25460 -1160 25480 -1100
rect 25540 -1160 25560 -1100
rect 25460 -1200 25560 -1160
rect 25460 -1260 25480 -1200
rect 25540 -1260 25560 -1200
rect 25460 -1300 25560 -1260
rect 25460 -1360 25480 -1300
rect 25540 -1360 25560 -1300
rect 25460 -1380 25560 -1360
rect 25630 -1000 25730 -980
rect 25630 -1060 25650 -1000
rect 25710 -1060 25730 -1000
rect 25630 -1100 25730 -1060
rect 25630 -1160 25650 -1100
rect 25710 -1160 25730 -1100
rect 25630 -1200 25730 -1160
rect 25630 -1260 25650 -1200
rect 25710 -1260 25730 -1200
rect 25630 -1300 25730 -1260
rect 25630 -1360 25650 -1300
rect 25710 -1360 25730 -1300
rect 25630 -1380 25730 -1360
rect 25800 -1000 25900 -980
rect 25800 -1060 25820 -1000
rect 25880 -1060 25900 -1000
rect 25800 -1100 25900 -1060
rect 25800 -1160 25820 -1100
rect 25880 -1160 25900 -1100
rect 25800 -1200 25900 -1160
rect 25800 -1260 25820 -1200
rect 25880 -1260 25900 -1200
rect 25800 -1300 25900 -1260
rect 25800 -1360 25820 -1300
rect 25880 -1360 25900 -1300
rect 25800 -1380 25900 -1360
rect 25970 -1000 26070 -980
rect 25970 -1060 25990 -1000
rect 26050 -1060 26070 -1000
rect 25970 -1100 26070 -1060
rect 25970 -1160 25990 -1100
rect 26050 -1160 26070 -1100
rect 25970 -1200 26070 -1160
rect 25970 -1260 25990 -1200
rect 26050 -1260 26070 -1200
rect 25970 -1300 26070 -1260
rect 25970 -1360 25990 -1300
rect 26050 -1360 26070 -1300
rect 25970 -1380 26070 -1360
rect 26140 -1000 26240 -980
rect 26140 -1060 26160 -1000
rect 26220 -1060 26240 -1000
rect 26140 -1100 26240 -1060
rect 26140 -1160 26160 -1100
rect 26220 -1160 26240 -1100
rect 26140 -1200 26240 -1160
rect 26140 -1260 26160 -1200
rect 26220 -1260 26240 -1200
rect 26140 -1300 26240 -1260
rect 26140 -1360 26160 -1300
rect 26220 -1360 26240 -1300
rect 26140 -1380 26240 -1360
rect 26310 -1000 26410 -980
rect 26310 -1060 26330 -1000
rect 26390 -1060 26410 -1000
rect 26310 -1100 26410 -1060
rect 26310 -1160 26330 -1100
rect 26390 -1160 26410 -1100
rect 26310 -1200 26410 -1160
rect 26310 -1260 26330 -1200
rect 26390 -1260 26410 -1200
rect 26310 -1300 26410 -1260
rect 26310 -1360 26330 -1300
rect 26390 -1360 26410 -1300
rect 26310 -1380 26410 -1360
rect 26480 -1000 26580 -980
rect 26480 -1060 26500 -1000
rect 26560 -1060 26580 -1000
rect 26480 -1100 26580 -1060
rect 26480 -1160 26500 -1100
rect 26560 -1160 26580 -1100
rect 26480 -1200 26580 -1160
rect 26480 -1260 26500 -1200
rect 26560 -1260 26580 -1200
rect 26480 -1300 26580 -1260
rect 26480 -1360 26500 -1300
rect 26560 -1360 26580 -1300
rect 26480 -1380 26580 -1360
rect 26650 -1000 26750 -980
rect 26650 -1060 26670 -1000
rect 26730 -1060 26750 -1000
rect 26650 -1100 26750 -1060
rect 26650 -1160 26670 -1100
rect 26730 -1160 26750 -1100
rect 26650 -1200 26750 -1160
rect 26650 -1260 26670 -1200
rect 26730 -1260 26750 -1200
rect 26650 -1300 26750 -1260
rect 26650 -1360 26670 -1300
rect 26730 -1360 26750 -1300
rect 26650 -1380 26750 -1360
rect 26820 -1000 26920 -980
rect 26820 -1060 26840 -1000
rect 26900 -1060 26920 -1000
rect 26820 -1100 26920 -1060
rect 26820 -1160 26840 -1100
rect 26900 -1160 26920 -1100
rect 26820 -1200 26920 -1160
rect 26820 -1260 26840 -1200
rect 26900 -1260 26920 -1200
rect 26820 -1300 26920 -1260
rect 26820 -1360 26840 -1300
rect 26900 -1360 26920 -1300
rect 26820 -1380 26920 -1360
rect 26990 -1000 27090 -980
rect 26990 -1060 27010 -1000
rect 27070 -1060 27090 -1000
rect 26990 -1100 27090 -1060
rect 26990 -1160 27010 -1100
rect 27070 -1160 27090 -1100
rect 26990 -1200 27090 -1160
rect 26990 -1260 27010 -1200
rect 27070 -1260 27090 -1200
rect 26990 -1300 27090 -1260
rect 26990 -1360 27010 -1300
rect 27070 -1360 27090 -1300
rect 26990 -1380 27090 -1360
rect 27160 -1000 27260 -980
rect 27160 -1060 27180 -1000
rect 27240 -1060 27260 -1000
rect 27160 -1100 27260 -1060
rect 27160 -1160 27180 -1100
rect 27240 -1160 27260 -1100
rect 27160 -1200 27260 -1160
rect 27160 -1260 27180 -1200
rect 27240 -1260 27260 -1200
rect 27160 -1300 27260 -1260
rect 27160 -1360 27180 -1300
rect 27240 -1360 27260 -1300
rect 27160 -1380 27260 -1360
rect 27330 -1000 27430 -980
rect 27330 -1060 27350 -1000
rect 27410 -1060 27430 -1000
rect 27330 -1100 27430 -1060
rect 27330 -1160 27350 -1100
rect 27410 -1160 27430 -1100
rect 27330 -1200 27430 -1160
rect 27330 -1260 27350 -1200
rect 27410 -1260 27430 -1200
rect 27330 -1300 27430 -1260
rect 27330 -1360 27350 -1300
rect 27410 -1360 27430 -1300
rect 27330 -1380 27430 -1360
rect 27500 -1000 27600 -980
rect 27500 -1060 27520 -1000
rect 27580 -1060 27600 -1000
rect 27500 -1100 27600 -1060
rect 27500 -1160 27520 -1100
rect 27580 -1160 27600 -1100
rect 27500 -1200 27600 -1160
rect 27500 -1260 27520 -1200
rect 27580 -1260 27600 -1200
rect 27500 -1300 27600 -1260
rect 27500 -1360 27520 -1300
rect 27580 -1360 27600 -1300
rect 27500 -1380 27600 -1360
rect 27670 -1000 27770 -980
rect 27670 -1060 27690 -1000
rect 27750 -1060 27770 -1000
rect 27670 -1100 27770 -1060
rect 27670 -1160 27690 -1100
rect 27750 -1160 27770 -1100
rect 27670 -1200 27770 -1160
rect 27670 -1260 27690 -1200
rect 27750 -1260 27770 -1200
rect 27670 -1300 27770 -1260
rect 27670 -1360 27690 -1300
rect 27750 -1360 27770 -1300
rect 27670 -1380 27770 -1360
rect 27840 -1000 27940 -980
rect 27840 -1060 27860 -1000
rect 27920 -1060 27940 -1000
rect 27840 -1100 27940 -1060
rect 27840 -1160 27860 -1100
rect 27920 -1160 27940 -1100
rect 27840 -1200 27940 -1160
rect 27840 -1260 27860 -1200
rect 27920 -1260 27940 -1200
rect 27840 -1300 27940 -1260
rect 27840 -1360 27860 -1300
rect 27920 -1360 27940 -1300
rect 27840 -1380 27940 -1360
rect 28010 -1000 28110 -980
rect 28010 -1060 28030 -1000
rect 28090 -1060 28110 -1000
rect 28010 -1100 28110 -1060
rect 28010 -1160 28030 -1100
rect 28090 -1160 28110 -1100
rect 28010 -1200 28110 -1160
rect 28010 -1260 28030 -1200
rect 28090 -1260 28110 -1200
rect 28010 -1300 28110 -1260
rect 28010 -1360 28030 -1300
rect 28090 -1360 28110 -1300
rect 28010 -1380 28110 -1360
rect 28180 -1000 28280 -980
rect 28180 -1060 28200 -1000
rect 28260 -1060 28280 -1000
rect 28180 -1100 28280 -1060
rect 28180 -1160 28200 -1100
rect 28260 -1160 28280 -1100
rect 28180 -1200 28280 -1160
rect 28180 -1260 28200 -1200
rect 28260 -1260 28280 -1200
rect 28180 -1300 28280 -1260
rect 28180 -1360 28200 -1300
rect 28260 -1360 28280 -1300
rect 28180 -1380 28280 -1360
rect 28350 -1000 28450 -980
rect 28350 -1060 28370 -1000
rect 28430 -1060 28450 -1000
rect 28350 -1100 28450 -1060
rect 28350 -1160 28370 -1100
rect 28430 -1160 28450 -1100
rect 28350 -1200 28450 -1160
rect 28350 -1260 28370 -1200
rect 28430 -1260 28450 -1200
rect 28350 -1300 28450 -1260
rect 28350 -1360 28370 -1300
rect 28430 -1360 28450 -1300
rect 28350 -1380 28450 -1360
rect 28520 -1000 28620 -980
rect 28520 -1060 28540 -1000
rect 28600 -1060 28620 -1000
rect 28520 -1100 28620 -1060
rect 28520 -1160 28540 -1100
rect 28600 -1160 28620 -1100
rect 28520 -1200 28620 -1160
rect 28520 -1260 28540 -1200
rect 28600 -1260 28620 -1200
rect 28520 -1300 28620 -1260
rect 28520 -1360 28540 -1300
rect 28600 -1360 28620 -1300
rect 28520 -1380 28620 -1360
rect 28690 -1000 28790 -980
rect 28690 -1060 28710 -1000
rect 28770 -1060 28790 -1000
rect 28690 -1100 28790 -1060
rect 28690 -1160 28710 -1100
rect 28770 -1160 28790 -1100
rect 28690 -1200 28790 -1160
rect 28690 -1260 28710 -1200
rect 28770 -1260 28790 -1200
rect 28690 -1300 28790 -1260
rect 28690 -1360 28710 -1300
rect 28770 -1360 28790 -1300
rect 28690 -1380 28790 -1360
rect 28860 -1000 28960 -980
rect 28860 -1060 28880 -1000
rect 28940 -1060 28960 -1000
rect 28860 -1100 28960 -1060
rect 28860 -1160 28880 -1100
rect 28940 -1160 28960 -1100
rect 28860 -1200 28960 -1160
rect 28860 -1260 28880 -1200
rect 28940 -1260 28960 -1200
rect 28860 -1300 28960 -1260
rect 28860 -1360 28880 -1300
rect 28940 -1360 28960 -1300
rect 28860 -1380 28960 -1360
rect 29030 -1000 29130 -980
rect 29030 -1060 29050 -1000
rect 29110 -1060 29130 -1000
rect 29030 -1100 29130 -1060
rect 29030 -1160 29050 -1100
rect 29110 -1160 29130 -1100
rect 29030 -1200 29130 -1160
rect 29030 -1260 29050 -1200
rect 29110 -1260 29130 -1200
rect 29030 -1300 29130 -1260
rect 29030 -1360 29050 -1300
rect 29110 -1360 29130 -1300
rect 29030 -1380 29130 -1360
rect 29200 -1000 29300 -980
rect 29200 -1060 29220 -1000
rect 29280 -1060 29300 -1000
rect 29200 -1100 29300 -1060
rect 29200 -1160 29220 -1100
rect 29280 -1160 29300 -1100
rect 29200 -1200 29300 -1160
rect 29200 -1260 29220 -1200
rect 29280 -1260 29300 -1200
rect 29200 -1300 29300 -1260
rect 29200 -1360 29220 -1300
rect 29280 -1360 29300 -1300
rect 29200 -1380 29300 -1360
rect 29370 -1000 29470 -980
rect 29370 -1060 29390 -1000
rect 29450 -1060 29470 -1000
rect 29370 -1100 29470 -1060
rect 29370 -1160 29390 -1100
rect 29450 -1160 29470 -1100
rect 29370 -1200 29470 -1160
rect 29370 -1260 29390 -1200
rect 29450 -1260 29470 -1200
rect 29370 -1300 29470 -1260
rect 29370 -1360 29390 -1300
rect 29450 -1360 29470 -1300
rect 29370 -1380 29470 -1360
rect 29540 -1000 29640 -980
rect 29540 -1060 29560 -1000
rect 29620 -1060 29640 -1000
rect 29540 -1100 29640 -1060
rect 29540 -1160 29560 -1100
rect 29620 -1160 29640 -1100
rect 29540 -1200 29640 -1160
rect 29540 -1260 29560 -1200
rect 29620 -1260 29640 -1200
rect 29540 -1300 29640 -1260
rect 29540 -1360 29560 -1300
rect 29620 -1360 29640 -1300
rect 29540 -1380 29640 -1360
rect 29710 -1000 29810 -980
rect 29710 -1060 29730 -1000
rect 29790 -1060 29810 -1000
rect 29710 -1100 29810 -1060
rect 29710 -1160 29730 -1100
rect 29790 -1160 29810 -1100
rect 29710 -1200 29810 -1160
rect 29710 -1260 29730 -1200
rect 29790 -1260 29810 -1200
rect 29710 -1300 29810 -1260
rect 29710 -1360 29730 -1300
rect 29790 -1360 29810 -1300
rect 29710 -1380 29810 -1360
rect 29880 -1000 29980 -980
rect 29880 -1060 29900 -1000
rect 29960 -1060 29980 -1000
rect 29880 -1100 29980 -1060
rect 29880 -1160 29900 -1100
rect 29960 -1160 29980 -1100
rect 29880 -1200 29980 -1160
rect 29880 -1260 29900 -1200
rect 29960 -1260 29980 -1200
rect 29880 -1300 29980 -1260
rect 29880 -1360 29900 -1300
rect 29960 -1360 29980 -1300
rect 29880 -1380 29980 -1360
rect 30050 -1000 30150 -980
rect 30050 -1060 30070 -1000
rect 30130 -1060 30150 -1000
rect 30050 -1100 30150 -1060
rect 30050 -1160 30070 -1100
rect 30130 -1160 30150 -1100
rect 30050 -1200 30150 -1160
rect 30050 -1260 30070 -1200
rect 30130 -1260 30150 -1200
rect 30050 -1300 30150 -1260
rect 30050 -1360 30070 -1300
rect 30130 -1360 30150 -1300
rect 30050 -1380 30150 -1360
rect 30220 -1000 30320 -980
rect 30220 -1060 30240 -1000
rect 30300 -1060 30320 -1000
rect 30220 -1100 30320 -1060
rect 30220 -1160 30240 -1100
rect 30300 -1160 30320 -1100
rect 30220 -1200 30320 -1160
rect 30220 -1260 30240 -1200
rect 30300 -1260 30320 -1200
rect 30220 -1300 30320 -1260
rect 30220 -1360 30240 -1300
rect 30300 -1360 30320 -1300
rect 30220 -1380 30320 -1360
rect 30390 -1000 30490 -980
rect 30390 -1060 30410 -1000
rect 30470 -1060 30490 -1000
rect 30390 -1100 30490 -1060
rect 30390 -1160 30410 -1100
rect 30470 -1160 30490 -1100
rect 30390 -1200 30490 -1160
rect 30390 -1260 30410 -1200
rect 30470 -1260 30490 -1200
rect 30390 -1300 30490 -1260
rect 30390 -1360 30410 -1300
rect 30470 -1360 30490 -1300
rect 30390 -1380 30490 -1360
rect 30560 -1000 30660 -980
rect 30560 -1060 30580 -1000
rect 30640 -1060 30660 -1000
rect 30560 -1100 30660 -1060
rect 30560 -1160 30580 -1100
rect 30640 -1160 30660 -1100
rect 30560 -1200 30660 -1160
rect 30560 -1260 30580 -1200
rect 30640 -1260 30660 -1200
rect 30560 -1300 30660 -1260
rect 30560 -1360 30580 -1300
rect 30640 -1360 30660 -1300
rect 30560 -1380 30660 -1360
rect 30730 -1000 30830 -980
rect 30730 -1060 30750 -1000
rect 30810 -1060 30830 -1000
rect 30730 -1100 30830 -1060
rect 30730 -1160 30750 -1100
rect 30810 -1160 30830 -1100
rect 30730 -1200 30830 -1160
rect 30730 -1260 30750 -1200
rect 30810 -1260 30830 -1200
rect 30730 -1300 30830 -1260
rect 30730 -1360 30750 -1300
rect 30810 -1360 30830 -1300
rect 30730 -1380 30830 -1360
rect 30900 -1000 31000 -980
rect 30900 -1060 30920 -1000
rect 30980 -1060 31000 -1000
rect 30900 -1100 31000 -1060
rect 30900 -1160 30920 -1100
rect 30980 -1160 31000 -1100
rect 30900 -1200 31000 -1160
rect 30900 -1260 30920 -1200
rect 30980 -1260 31000 -1200
rect 30900 -1300 31000 -1260
rect 30900 -1360 30920 -1300
rect 30980 -1360 31000 -1300
rect 30900 -1380 31000 -1360
rect 31070 -1000 31170 -980
rect 31070 -1060 31090 -1000
rect 31150 -1060 31170 -1000
rect 31070 -1100 31170 -1060
rect 31070 -1160 31090 -1100
rect 31150 -1160 31170 -1100
rect 31070 -1200 31170 -1160
rect 31070 -1260 31090 -1200
rect 31150 -1260 31170 -1200
rect 31070 -1300 31170 -1260
rect 31070 -1360 31090 -1300
rect 31150 -1360 31170 -1300
rect 31070 -1380 31170 -1360
rect 31240 -1000 31340 -980
rect 31240 -1060 31260 -1000
rect 31320 -1060 31340 -1000
rect 31240 -1100 31340 -1060
rect 31240 -1160 31260 -1100
rect 31320 -1160 31340 -1100
rect 31240 -1200 31340 -1160
rect 31240 -1260 31260 -1200
rect 31320 -1260 31340 -1200
rect 31240 -1300 31340 -1260
rect 31240 -1360 31260 -1300
rect 31320 -1360 31340 -1300
rect 31240 -1380 31340 -1360
rect 31410 -1000 31510 -980
rect 31410 -1060 31430 -1000
rect 31490 -1060 31510 -1000
rect 31410 -1100 31510 -1060
rect 31410 -1160 31430 -1100
rect 31490 -1160 31510 -1100
rect 31410 -1200 31510 -1160
rect 31410 -1260 31430 -1200
rect 31490 -1260 31510 -1200
rect 31410 -1300 31510 -1260
rect 31410 -1360 31430 -1300
rect 31490 -1360 31510 -1300
rect 31410 -1380 31510 -1360
rect 31580 -1000 31680 -980
rect 31580 -1060 31600 -1000
rect 31660 -1060 31680 -1000
rect 31580 -1100 31680 -1060
rect 31580 -1160 31600 -1100
rect 31660 -1160 31680 -1100
rect 31580 -1200 31680 -1160
rect 31580 -1260 31600 -1200
rect 31660 -1260 31680 -1200
rect 31580 -1300 31680 -1260
rect 31580 -1360 31600 -1300
rect 31660 -1360 31680 -1300
rect 31580 -1380 31680 -1360
rect 31750 -1000 31850 -980
rect 31750 -1060 31770 -1000
rect 31830 -1060 31850 -1000
rect 31750 -1100 31850 -1060
rect 31750 -1160 31770 -1100
rect 31830 -1160 31850 -1100
rect 31750 -1200 31850 -1160
rect 31750 -1260 31770 -1200
rect 31830 -1260 31850 -1200
rect 31750 -1300 31850 -1260
rect 31750 -1360 31770 -1300
rect 31830 -1360 31850 -1300
rect 31750 -1380 31850 -1360
rect 31920 -1000 32020 -980
rect 31920 -1060 31940 -1000
rect 32000 -1060 32020 -1000
rect 31920 -1100 32020 -1060
rect 31920 -1160 31940 -1100
rect 32000 -1160 32020 -1100
rect 31920 -1200 32020 -1160
rect 31920 -1260 31940 -1200
rect 32000 -1260 32020 -1200
rect 31920 -1300 32020 -1260
rect 31920 -1360 31940 -1300
rect 32000 -1360 32020 -1300
rect 31920 -1380 32020 -1360
rect 32090 -1000 32190 -980
rect 32090 -1060 32110 -1000
rect 32170 -1060 32190 -1000
rect 32090 -1100 32190 -1060
rect 32090 -1160 32110 -1100
rect 32170 -1160 32190 -1100
rect 32090 -1200 32190 -1160
rect 32090 -1260 32110 -1200
rect 32170 -1260 32190 -1200
rect 32090 -1300 32190 -1260
rect 32090 -1360 32110 -1300
rect 32170 -1360 32190 -1300
rect 32090 -1380 32190 -1360
rect 32260 -1000 32360 -980
rect 32260 -1060 32280 -1000
rect 32340 -1060 32360 -1000
rect 32260 -1100 32360 -1060
rect 32260 -1160 32280 -1100
rect 32340 -1160 32360 -1100
rect 32260 -1200 32360 -1160
rect 32260 -1260 32280 -1200
rect 32340 -1260 32360 -1200
rect 32260 -1300 32360 -1260
rect 32260 -1360 32280 -1300
rect 32340 -1360 32360 -1300
rect 32260 -1380 32360 -1360
rect 32430 -1000 32530 -980
rect 32430 -1060 32450 -1000
rect 32510 -1060 32530 -1000
rect 32430 -1100 32530 -1060
rect 32430 -1160 32450 -1100
rect 32510 -1160 32530 -1100
rect 32430 -1200 32530 -1160
rect 32430 -1260 32450 -1200
rect 32510 -1260 32530 -1200
rect 32430 -1300 32530 -1260
rect 32430 -1360 32450 -1300
rect 32510 -1360 32530 -1300
rect 32430 -1380 32530 -1360
rect 32600 -1000 32700 -980
rect 32600 -1060 32620 -1000
rect 32680 -1060 32700 -1000
rect 32600 -1100 32700 -1060
rect 32600 -1160 32620 -1100
rect 32680 -1160 32700 -1100
rect 32600 -1200 32700 -1160
rect 32600 -1260 32620 -1200
rect 32680 -1260 32700 -1200
rect 32600 -1300 32700 -1260
rect 32600 -1360 32620 -1300
rect 32680 -1360 32700 -1300
rect 32600 -1380 32700 -1360
rect 32770 -1000 32870 -980
rect 32770 -1060 32790 -1000
rect 32850 -1060 32870 -1000
rect 32770 -1100 32870 -1060
rect 32770 -1160 32790 -1100
rect 32850 -1160 32870 -1100
rect 32770 -1200 32870 -1160
rect 32770 -1260 32790 -1200
rect 32850 -1260 32870 -1200
rect 32770 -1300 32870 -1260
rect 32770 -1360 32790 -1300
rect 32850 -1360 32870 -1300
rect 32770 -1380 32870 -1360
rect 32940 -1000 33040 -980
rect 32940 -1060 32960 -1000
rect 33020 -1060 33040 -1000
rect 32940 -1100 33040 -1060
rect 32940 -1160 32960 -1100
rect 33020 -1160 33040 -1100
rect 32940 -1200 33040 -1160
rect 32940 -1260 32960 -1200
rect 33020 -1260 33040 -1200
rect 32940 -1300 33040 -1260
rect 32940 -1360 32960 -1300
rect 33020 -1360 33040 -1300
rect 32940 -1380 33040 -1360
rect 33110 -1000 33210 -980
rect 33110 -1060 33130 -1000
rect 33190 -1060 33210 -1000
rect 33110 -1100 33210 -1060
rect 33110 -1160 33130 -1100
rect 33190 -1160 33210 -1100
rect 33110 -1200 33210 -1160
rect 33110 -1260 33130 -1200
rect 33190 -1260 33210 -1200
rect 33110 -1300 33210 -1260
rect 33110 -1360 33130 -1300
rect 33190 -1360 33210 -1300
rect 33110 -1380 33210 -1360
rect 33280 -1000 33380 -980
rect 33280 -1060 33300 -1000
rect 33360 -1060 33380 -1000
rect 33280 -1100 33380 -1060
rect 33280 -1160 33300 -1100
rect 33360 -1160 33380 -1100
rect 33280 -1200 33380 -1160
rect 33280 -1260 33300 -1200
rect 33360 -1260 33380 -1200
rect 33280 -1300 33380 -1260
rect 33280 -1360 33300 -1300
rect 33360 -1360 33380 -1300
rect 33280 -1380 33380 -1360
rect 33450 -1000 33550 -980
rect 33450 -1060 33470 -1000
rect 33530 -1060 33550 -1000
rect 33450 -1100 33550 -1060
rect 33450 -1160 33470 -1100
rect 33530 -1160 33550 -1100
rect 33450 -1200 33550 -1160
rect 33450 -1260 33470 -1200
rect 33530 -1260 33550 -1200
rect 33450 -1300 33550 -1260
rect 33450 -1360 33470 -1300
rect 33530 -1360 33550 -1300
rect 33450 -1380 33550 -1360
rect 33620 -1000 33720 -980
rect 33620 -1060 33640 -1000
rect 33700 -1060 33720 -1000
rect 33620 -1100 33720 -1060
rect 33620 -1160 33640 -1100
rect 33700 -1160 33720 -1100
rect 33620 -1200 33720 -1160
rect 33620 -1260 33640 -1200
rect 33700 -1260 33720 -1200
rect 33620 -1300 33720 -1260
rect 33620 -1360 33640 -1300
rect 33700 -1360 33720 -1300
rect 33620 -1380 33720 -1360
rect 33790 -1000 33890 -980
rect 33790 -1060 33810 -1000
rect 33870 -1060 33890 -1000
rect 33790 -1100 33890 -1060
rect 33790 -1160 33810 -1100
rect 33870 -1160 33890 -1100
rect 33790 -1200 33890 -1160
rect 33790 -1260 33810 -1200
rect 33870 -1260 33890 -1200
rect 33790 -1300 33890 -1260
rect 33790 -1360 33810 -1300
rect 33870 -1360 33890 -1300
rect 33790 -1380 33890 -1360
rect 33960 -1000 34060 -980
rect 33960 -1060 33980 -1000
rect 34040 -1060 34060 -1000
rect 33960 -1100 34060 -1060
rect 33960 -1160 33980 -1100
rect 34040 -1160 34060 -1100
rect 33960 -1200 34060 -1160
rect 33960 -1260 33980 -1200
rect 34040 -1260 34060 -1200
rect 33960 -1300 34060 -1260
rect 33960 -1360 33980 -1300
rect 34040 -1360 34060 -1300
rect 33960 -1380 34060 -1360
rect 34130 -1000 34230 -980
rect 34130 -1060 34150 -1000
rect 34210 -1060 34230 -1000
rect 34130 -1100 34230 -1060
rect 34130 -1160 34150 -1100
rect 34210 -1160 34230 -1100
rect 34130 -1200 34230 -1160
rect 34130 -1260 34150 -1200
rect 34210 -1260 34230 -1200
rect 34130 -1300 34230 -1260
rect 34130 -1360 34150 -1300
rect 34210 -1360 34230 -1300
rect 34130 -1380 34230 -1360
rect 34300 -1000 34400 -980
rect 34300 -1060 34320 -1000
rect 34380 -1060 34400 -1000
rect 34300 -1100 34400 -1060
rect 34300 -1160 34320 -1100
rect 34380 -1160 34400 -1100
rect 34300 -1200 34400 -1160
rect 34300 -1260 34320 -1200
rect 34380 -1260 34400 -1200
rect 34300 -1300 34400 -1260
rect 34300 -1360 34320 -1300
rect 34380 -1360 34400 -1300
rect 34300 -1380 34400 -1360
rect 34470 -1000 34570 -980
rect 34470 -1060 34490 -1000
rect 34550 -1060 34570 -1000
rect 34470 -1100 34570 -1060
rect 34470 -1160 34490 -1100
rect 34550 -1160 34570 -1100
rect 34470 -1200 34570 -1160
rect 34470 -1260 34490 -1200
rect 34550 -1260 34570 -1200
rect 34470 -1300 34570 -1260
rect 34470 -1360 34490 -1300
rect 34550 -1360 34570 -1300
rect 34470 -1380 34570 -1360
rect 34640 -1000 34740 -980
rect 34640 -1060 34660 -1000
rect 34720 -1060 34740 -1000
rect 34640 -1100 34740 -1060
rect 34640 -1160 34660 -1100
rect 34720 -1160 34740 -1100
rect 34640 -1200 34740 -1160
rect 34640 -1260 34660 -1200
rect 34720 -1260 34740 -1200
rect 34640 -1300 34740 -1260
rect 34640 -1360 34660 -1300
rect 34720 -1360 34740 -1300
rect 34640 -1380 34740 -1360
rect 34810 -1000 34910 -980
rect 34810 -1060 34830 -1000
rect 34890 -1060 34910 -1000
rect 34810 -1100 34910 -1060
rect 34810 -1160 34830 -1100
rect 34890 -1160 34910 -1100
rect 34810 -1200 34910 -1160
rect 34810 -1260 34830 -1200
rect 34890 -1260 34910 -1200
rect 34810 -1300 34910 -1260
rect 34810 -1360 34830 -1300
rect 34890 -1360 34910 -1300
rect 34810 -1380 34910 -1360
rect 34980 -1000 35080 -980
rect 34980 -1060 35000 -1000
rect 35060 -1060 35080 -1000
rect 34980 -1100 35080 -1060
rect 34980 -1160 35000 -1100
rect 35060 -1160 35080 -1100
rect 34980 -1200 35080 -1160
rect 34980 -1260 35000 -1200
rect 35060 -1260 35080 -1200
rect 34980 -1300 35080 -1260
rect 34980 -1360 35000 -1300
rect 35060 -1360 35080 -1300
rect 34980 -1380 35080 -1360
rect 35150 -1000 35250 -980
rect 35150 -1060 35170 -1000
rect 35230 -1060 35250 -1000
rect 35150 -1100 35250 -1060
rect 35150 -1160 35170 -1100
rect 35230 -1160 35250 -1100
rect 35150 -1200 35250 -1160
rect 35150 -1260 35170 -1200
rect 35230 -1260 35250 -1200
rect 35150 -1300 35250 -1260
rect 35150 -1360 35170 -1300
rect 35230 -1360 35250 -1300
rect 35150 -1380 35250 -1360
rect 35320 -1000 35420 -980
rect 35320 -1060 35340 -1000
rect 35400 -1060 35420 -1000
rect 35320 -1100 35420 -1060
rect 35320 -1160 35340 -1100
rect 35400 -1160 35420 -1100
rect 35320 -1200 35420 -1160
rect 35320 -1260 35340 -1200
rect 35400 -1260 35420 -1200
rect 35320 -1300 35420 -1260
rect 35320 -1360 35340 -1300
rect 35400 -1360 35420 -1300
rect 35320 -1380 35420 -1360
rect 35490 -1000 35590 -980
rect 35490 -1060 35510 -1000
rect 35570 -1060 35590 -1000
rect 35490 -1100 35590 -1060
rect 35490 -1160 35510 -1100
rect 35570 -1160 35590 -1100
rect 35490 -1200 35590 -1160
rect 35490 -1260 35510 -1200
rect 35570 -1260 35590 -1200
rect 35490 -1300 35590 -1260
rect 35490 -1360 35510 -1300
rect 35570 -1360 35590 -1300
rect 35490 -1380 35590 -1360
rect 35660 -1000 35760 -980
rect 35660 -1060 35680 -1000
rect 35740 -1060 35760 -1000
rect 35660 -1100 35760 -1060
rect 35660 -1160 35680 -1100
rect 35740 -1160 35760 -1100
rect 35660 -1200 35760 -1160
rect 35660 -1260 35680 -1200
rect 35740 -1260 35760 -1200
rect 35660 -1300 35760 -1260
rect 35660 -1360 35680 -1300
rect 35740 -1360 35760 -1300
rect 35660 -1380 35760 -1360
rect 35830 -1000 35930 -980
rect 35830 -1060 35850 -1000
rect 35910 -1060 35930 -1000
rect 35830 -1100 35930 -1060
rect 35830 -1160 35850 -1100
rect 35910 -1160 35930 -1100
rect 35830 -1200 35930 -1160
rect 35830 -1260 35850 -1200
rect 35910 -1260 35930 -1200
rect 35830 -1300 35930 -1260
rect 35830 -1360 35850 -1300
rect 35910 -1360 35930 -1300
rect 35830 -1380 35930 -1360
rect 36000 -1000 36100 -980
rect 36000 -1060 36020 -1000
rect 36080 -1060 36100 -1000
rect 36000 -1100 36100 -1060
rect 36000 -1160 36020 -1100
rect 36080 -1160 36100 -1100
rect 36000 -1200 36100 -1160
rect 36000 -1260 36020 -1200
rect 36080 -1260 36100 -1200
rect 36000 -1300 36100 -1260
rect 36000 -1360 36020 -1300
rect 36080 -1360 36100 -1300
rect 36000 -1380 36100 -1360
rect 36170 -1000 36270 -980
rect 36170 -1060 36190 -1000
rect 36250 -1060 36270 -1000
rect 36170 -1100 36270 -1060
rect 36170 -1160 36190 -1100
rect 36250 -1160 36270 -1100
rect 36170 -1200 36270 -1160
rect 36170 -1260 36190 -1200
rect 36250 -1260 36270 -1200
rect 36170 -1300 36270 -1260
rect 36170 -1360 36190 -1300
rect 36250 -1360 36270 -1300
rect 36170 -1380 36270 -1360
rect 36340 -1000 36440 -980
rect 36340 -1060 36360 -1000
rect 36420 -1060 36440 -1000
rect 36340 -1100 36440 -1060
rect 36340 -1160 36360 -1100
rect 36420 -1160 36440 -1100
rect 36340 -1200 36440 -1160
rect 36340 -1260 36360 -1200
rect 36420 -1260 36440 -1200
rect 36340 -1300 36440 -1260
rect 36340 -1360 36360 -1300
rect 36420 -1360 36440 -1300
rect 36340 -1380 36440 -1360
rect 36510 -1000 36610 -980
rect 36510 -1060 36530 -1000
rect 36590 -1060 36610 -1000
rect 36510 -1100 36610 -1060
rect 36510 -1160 36530 -1100
rect 36590 -1160 36610 -1100
rect 36510 -1200 36610 -1160
rect 36510 -1260 36530 -1200
rect 36590 -1260 36610 -1200
rect 36510 -1300 36610 -1260
rect 36510 -1360 36530 -1300
rect 36590 -1360 36610 -1300
rect 36510 -1380 36610 -1360
rect 36680 -1000 36780 -980
rect 36680 -1060 36700 -1000
rect 36760 -1060 36780 -1000
rect 36680 -1100 36780 -1060
rect 36680 -1160 36700 -1100
rect 36760 -1160 36780 -1100
rect 36680 -1200 36780 -1160
rect 36680 -1260 36700 -1200
rect 36760 -1260 36780 -1200
rect 36680 -1300 36780 -1260
rect 36680 -1360 36700 -1300
rect 36760 -1360 36780 -1300
rect 36680 -1380 36780 -1360
rect 36850 -1000 36950 -980
rect 36850 -1060 36870 -1000
rect 36930 -1060 36950 -1000
rect 36850 -1100 36950 -1060
rect 36850 -1160 36870 -1100
rect 36930 -1160 36950 -1100
rect 36850 -1200 36950 -1160
rect 36850 -1260 36870 -1200
rect 36930 -1260 36950 -1200
rect 36850 -1300 36950 -1260
rect 36850 -1360 36870 -1300
rect 36930 -1360 36950 -1300
rect 36850 -1380 36950 -1360
rect 37020 -1000 37120 -980
rect 37020 -1060 37040 -1000
rect 37100 -1060 37120 -1000
rect 37020 -1100 37120 -1060
rect 37020 -1160 37040 -1100
rect 37100 -1160 37120 -1100
rect 37020 -1200 37120 -1160
rect 37020 -1260 37040 -1200
rect 37100 -1260 37120 -1200
rect 37020 -1300 37120 -1260
rect 37020 -1360 37040 -1300
rect 37100 -1360 37120 -1300
rect 37020 -1380 37120 -1360
rect 37190 -1000 37290 -980
rect 37190 -1060 37210 -1000
rect 37270 -1060 37290 -1000
rect 37190 -1100 37290 -1060
rect 37190 -1160 37210 -1100
rect 37270 -1160 37290 -1100
rect 37190 -1200 37290 -1160
rect 37190 -1260 37210 -1200
rect 37270 -1260 37290 -1200
rect 37190 -1300 37290 -1260
rect 37190 -1360 37210 -1300
rect 37270 -1360 37290 -1300
rect 37190 -1380 37290 -1360
rect 37360 -1000 37460 -980
rect 37360 -1060 37380 -1000
rect 37440 -1060 37460 -1000
rect 37360 -1100 37460 -1060
rect 37360 -1160 37380 -1100
rect 37440 -1160 37460 -1100
rect 37360 -1200 37460 -1160
rect 37360 -1260 37380 -1200
rect 37440 -1260 37460 -1200
rect 37360 -1300 37460 -1260
rect 37360 -1360 37380 -1300
rect 37440 -1360 37460 -1300
rect 37360 -1380 37460 -1360
rect 37530 -1000 37630 -980
rect 37530 -1060 37550 -1000
rect 37610 -1060 37630 -1000
rect 37530 -1100 37630 -1060
rect 37530 -1160 37550 -1100
rect 37610 -1160 37630 -1100
rect 37530 -1200 37630 -1160
rect 37530 -1260 37550 -1200
rect 37610 -1260 37630 -1200
rect 37530 -1300 37630 -1260
rect 37530 -1360 37550 -1300
rect 37610 -1360 37630 -1300
rect 37530 -1380 37630 -1360
rect 37700 -1000 37800 -980
rect 37700 -1060 37720 -1000
rect 37780 -1060 37800 -1000
rect 37700 -1100 37800 -1060
rect 37700 -1160 37720 -1100
rect 37780 -1160 37800 -1100
rect 37700 -1200 37800 -1160
rect 37700 -1260 37720 -1200
rect 37780 -1260 37800 -1200
rect 37700 -1300 37800 -1260
rect 37700 -1360 37720 -1300
rect 37780 -1360 37800 -1300
rect 37700 -1380 37800 -1360
rect 37870 -1000 37970 -980
rect 37870 -1060 37890 -1000
rect 37950 -1060 37970 -1000
rect 37870 -1100 37970 -1060
rect 37870 -1160 37890 -1100
rect 37950 -1160 37970 -1100
rect 37870 -1200 37970 -1160
rect 37870 -1260 37890 -1200
rect 37950 -1260 37970 -1200
rect 37870 -1300 37970 -1260
rect 37870 -1360 37890 -1300
rect 37950 -1360 37970 -1300
rect 37870 -1380 37970 -1360
rect 38040 -1000 38140 -980
rect 38040 -1060 38060 -1000
rect 38120 -1060 38140 -1000
rect 38040 -1100 38140 -1060
rect 38040 -1160 38060 -1100
rect 38120 -1160 38140 -1100
rect 38040 -1200 38140 -1160
rect 38040 -1260 38060 -1200
rect 38120 -1260 38140 -1200
rect 38040 -1300 38140 -1260
rect 38040 -1360 38060 -1300
rect 38120 -1360 38140 -1300
rect 38040 -1380 38140 -1360
rect 38210 -1000 38310 -980
rect 38210 -1060 38230 -1000
rect 38290 -1060 38310 -1000
rect 38210 -1100 38310 -1060
rect 38210 -1160 38230 -1100
rect 38290 -1160 38310 -1100
rect 38210 -1200 38310 -1160
rect 38210 -1260 38230 -1200
rect 38290 -1260 38310 -1200
rect 38210 -1300 38310 -1260
rect 38210 -1360 38230 -1300
rect 38290 -1360 38310 -1300
rect 38210 -1380 38310 -1360
rect 38380 -1000 38480 -980
rect 38380 -1060 38400 -1000
rect 38460 -1060 38480 -1000
rect 38380 -1100 38480 -1060
rect 38380 -1160 38400 -1100
rect 38460 -1160 38480 -1100
rect 38380 -1200 38480 -1160
rect 38380 -1260 38400 -1200
rect 38460 -1260 38480 -1200
rect 38380 -1300 38480 -1260
rect 38380 -1360 38400 -1300
rect 38460 -1360 38480 -1300
rect 38380 -1380 38480 -1360
rect 38550 -1000 38650 -980
rect 38550 -1060 38570 -1000
rect 38630 -1060 38650 -1000
rect 38550 -1100 38650 -1060
rect 38550 -1160 38570 -1100
rect 38630 -1160 38650 -1100
rect 38550 -1200 38650 -1160
rect 38550 -1260 38570 -1200
rect 38630 -1260 38650 -1200
rect 38550 -1300 38650 -1260
rect 38550 -1360 38570 -1300
rect 38630 -1360 38650 -1300
rect 38550 -1380 38650 -1360
rect 38720 -1000 38820 -980
rect 38720 -1060 38740 -1000
rect 38800 -1060 38820 -1000
rect 38720 -1100 38820 -1060
rect 38720 -1160 38740 -1100
rect 38800 -1160 38820 -1100
rect 38720 -1200 38820 -1160
rect 38720 -1260 38740 -1200
rect 38800 -1260 38820 -1200
rect 38720 -1300 38820 -1260
rect 38720 -1360 38740 -1300
rect 38800 -1360 38820 -1300
rect 38720 -1380 38820 -1360
rect 38890 -1000 38990 -980
rect 38890 -1060 38910 -1000
rect 38970 -1060 38990 -1000
rect 38890 -1100 38990 -1060
rect 38890 -1160 38910 -1100
rect 38970 -1160 38990 -1100
rect 38890 -1200 38990 -1160
rect 38890 -1260 38910 -1200
rect 38970 -1260 38990 -1200
rect 38890 -1300 38990 -1260
rect 38890 -1360 38910 -1300
rect 38970 -1360 38990 -1300
rect 38890 -1380 38990 -1360
rect 39060 -1000 39160 -980
rect 39060 -1060 39080 -1000
rect 39140 -1060 39160 -1000
rect 39060 -1100 39160 -1060
rect 39060 -1160 39080 -1100
rect 39140 -1160 39160 -1100
rect 39060 -1200 39160 -1160
rect 39060 -1260 39080 -1200
rect 39140 -1260 39160 -1200
rect 39060 -1300 39160 -1260
rect 39060 -1360 39080 -1300
rect 39140 -1360 39160 -1300
rect 39060 -1380 39160 -1360
rect 39230 -1000 39330 -980
rect 39230 -1060 39250 -1000
rect 39310 -1060 39330 -1000
rect 39230 -1100 39330 -1060
rect 39230 -1160 39250 -1100
rect 39310 -1160 39330 -1100
rect 39230 -1200 39330 -1160
rect 39230 -1260 39250 -1200
rect 39310 -1260 39330 -1200
rect 39230 -1300 39330 -1260
rect 39230 -1360 39250 -1300
rect 39310 -1360 39330 -1300
rect 39230 -1380 39330 -1360
rect 39400 -1000 39500 -980
rect 39400 -1060 39420 -1000
rect 39480 -1060 39500 -1000
rect 39400 -1100 39500 -1060
rect 39400 -1160 39420 -1100
rect 39480 -1160 39500 -1100
rect 39400 -1200 39500 -1160
rect 39400 -1260 39420 -1200
rect 39480 -1260 39500 -1200
rect 39400 -1300 39500 -1260
rect 39400 -1360 39420 -1300
rect 39480 -1360 39500 -1300
rect 39400 -1380 39500 -1360
rect 39570 -1000 39670 -980
rect 39570 -1060 39590 -1000
rect 39650 -1060 39670 -1000
rect 39570 -1100 39670 -1060
rect 39570 -1160 39590 -1100
rect 39650 -1160 39670 -1100
rect 39570 -1200 39670 -1160
rect 39570 -1260 39590 -1200
rect 39650 -1260 39670 -1200
rect 39570 -1300 39670 -1260
rect 39570 -1360 39590 -1300
rect 39650 -1360 39670 -1300
rect 39570 -1380 39670 -1360
rect 39740 -1000 39840 -980
rect 39740 -1060 39760 -1000
rect 39820 -1060 39840 -1000
rect 39740 -1100 39840 -1060
rect 39740 -1160 39760 -1100
rect 39820 -1160 39840 -1100
rect 39740 -1200 39840 -1160
rect 39740 -1260 39760 -1200
rect 39820 -1260 39840 -1200
rect 39740 -1300 39840 -1260
rect 39740 -1360 39760 -1300
rect 39820 -1360 39840 -1300
rect 39740 -1380 39840 -1360
rect 39910 -1000 40010 -980
rect 39910 -1060 39930 -1000
rect 39990 -1060 40010 -1000
rect 39910 -1100 40010 -1060
rect 39910 -1160 39930 -1100
rect 39990 -1160 40010 -1100
rect 39910 -1200 40010 -1160
rect 39910 -1260 39930 -1200
rect 39990 -1260 40010 -1200
rect 39910 -1300 40010 -1260
rect 39910 -1360 39930 -1300
rect 39990 -1360 40010 -1300
rect 39910 -1380 40010 -1360
rect 40080 -1000 40180 -980
rect 40080 -1060 40100 -1000
rect 40160 -1060 40180 -1000
rect 40080 -1100 40180 -1060
rect 40080 -1160 40100 -1100
rect 40160 -1160 40180 -1100
rect 40080 -1200 40180 -1160
rect 40080 -1260 40100 -1200
rect 40160 -1260 40180 -1200
rect 40080 -1300 40180 -1260
rect 40080 -1360 40100 -1300
rect 40160 -1360 40180 -1300
rect 40080 -1380 40180 -1360
rect 40250 -1000 40350 -980
rect 40250 -1060 40270 -1000
rect 40330 -1060 40350 -1000
rect 40250 -1100 40350 -1060
rect 40250 -1160 40270 -1100
rect 40330 -1160 40350 -1100
rect 40250 -1200 40350 -1160
rect 40250 -1260 40270 -1200
rect 40330 -1260 40350 -1200
rect 40250 -1300 40350 -1260
rect 40250 -1360 40270 -1300
rect 40330 -1360 40350 -1300
rect 40250 -1380 40350 -1360
rect 40420 -1000 40520 -980
rect 40420 -1060 40440 -1000
rect 40500 -1060 40520 -1000
rect 40420 -1100 40520 -1060
rect 40420 -1160 40440 -1100
rect 40500 -1160 40520 -1100
rect 40420 -1200 40520 -1160
rect 40420 -1260 40440 -1200
rect 40500 -1260 40520 -1200
rect 40420 -1300 40520 -1260
rect 40420 -1360 40440 -1300
rect 40500 -1360 40520 -1300
rect 40420 -1380 40520 -1360
rect 40590 -1000 40690 -980
rect 40590 -1060 40610 -1000
rect 40670 -1060 40690 -1000
rect 40590 -1100 40690 -1060
rect 40590 -1160 40610 -1100
rect 40670 -1160 40690 -1100
rect 40590 -1200 40690 -1160
rect 40590 -1260 40610 -1200
rect 40670 -1260 40690 -1200
rect 40590 -1300 40690 -1260
rect 40590 -1360 40610 -1300
rect 40670 -1360 40690 -1300
rect 40590 -1380 40690 -1360
rect 40760 -1000 40860 -980
rect 40760 -1060 40780 -1000
rect 40840 -1060 40860 -1000
rect 40760 -1100 40860 -1060
rect 40760 -1160 40780 -1100
rect 40840 -1160 40860 -1100
rect 40760 -1200 40860 -1160
rect 40760 -1260 40780 -1200
rect 40840 -1260 40860 -1200
rect 40760 -1300 40860 -1260
rect 40760 -1360 40780 -1300
rect 40840 -1360 40860 -1300
rect 40760 -1380 40860 -1360
rect 40930 -1000 41030 -980
rect 40930 -1060 40950 -1000
rect 41010 -1060 41030 -1000
rect 40930 -1100 41030 -1060
rect 40930 -1160 40950 -1100
rect 41010 -1160 41030 -1100
rect 40930 -1200 41030 -1160
rect 40930 -1260 40950 -1200
rect 41010 -1260 41030 -1200
rect 40930 -1300 41030 -1260
rect 40930 -1360 40950 -1300
rect 41010 -1360 41030 -1300
rect 40930 -1380 41030 -1360
rect 41100 -1000 41200 -980
rect 41100 -1060 41120 -1000
rect 41180 -1060 41200 -1000
rect 41100 -1100 41200 -1060
rect 41100 -1160 41120 -1100
rect 41180 -1160 41200 -1100
rect 41100 -1200 41200 -1160
rect 41100 -1260 41120 -1200
rect 41180 -1260 41200 -1200
rect 41100 -1300 41200 -1260
rect 41100 -1360 41120 -1300
rect 41180 -1360 41200 -1300
rect 41100 -1380 41200 -1360
rect 41270 -1000 41370 -980
rect 41270 -1060 41290 -1000
rect 41350 -1060 41370 -1000
rect 41270 -1100 41370 -1060
rect 41270 -1160 41290 -1100
rect 41350 -1160 41370 -1100
rect 41270 -1200 41370 -1160
rect 41270 -1260 41290 -1200
rect 41350 -1260 41370 -1200
rect 41270 -1300 41370 -1260
rect 41270 -1360 41290 -1300
rect 41350 -1360 41370 -1300
rect 41270 -1380 41370 -1360
rect 41440 -1000 41540 -980
rect 41440 -1060 41460 -1000
rect 41520 -1060 41540 -1000
rect 41440 -1100 41540 -1060
rect 41440 -1160 41460 -1100
rect 41520 -1160 41540 -1100
rect 41440 -1200 41540 -1160
rect 41440 -1260 41460 -1200
rect 41520 -1260 41540 -1200
rect 41440 -1300 41540 -1260
rect 41440 -1360 41460 -1300
rect 41520 -1360 41540 -1300
rect 41440 -1380 41540 -1360
rect 41610 -1000 41710 -980
rect 41610 -1060 41630 -1000
rect 41690 -1060 41710 -1000
rect 41610 -1100 41710 -1060
rect 41610 -1160 41630 -1100
rect 41690 -1160 41710 -1100
rect 41610 -1200 41710 -1160
rect 41610 -1260 41630 -1200
rect 41690 -1260 41710 -1200
rect 41610 -1300 41710 -1260
rect 41610 -1360 41630 -1300
rect 41690 -1360 41710 -1300
rect 41610 -1380 41710 -1360
rect 41780 -1000 41880 -980
rect 41780 -1060 41800 -1000
rect 41860 -1060 41880 -1000
rect 41780 -1100 41880 -1060
rect 41780 -1160 41800 -1100
rect 41860 -1160 41880 -1100
rect 41780 -1200 41880 -1160
rect 41780 -1260 41800 -1200
rect 41860 -1260 41880 -1200
rect 41780 -1300 41880 -1260
rect 41780 -1360 41800 -1300
rect 41860 -1360 41880 -1300
rect 41780 -1380 41880 -1360
rect 41950 -1000 42050 -980
rect 41950 -1060 41970 -1000
rect 42030 -1060 42050 -1000
rect 41950 -1100 42050 -1060
rect 41950 -1160 41970 -1100
rect 42030 -1160 42050 -1100
rect 41950 -1200 42050 -1160
rect 41950 -1260 41970 -1200
rect 42030 -1260 42050 -1200
rect 41950 -1300 42050 -1260
rect 41950 -1360 41970 -1300
rect 42030 -1360 42050 -1300
rect 41950 -1380 42050 -1360
rect 42120 -1000 42220 -980
rect 42120 -1060 42140 -1000
rect 42200 -1060 42220 -1000
rect 42120 -1100 42220 -1060
rect 42120 -1160 42140 -1100
rect 42200 -1160 42220 -1100
rect 42120 -1200 42220 -1160
rect 42120 -1260 42140 -1200
rect 42200 -1260 42220 -1200
rect 42120 -1300 42220 -1260
rect 42120 -1360 42140 -1300
rect 42200 -1360 42220 -1300
rect 42120 -1380 42220 -1360
rect 42290 -1000 42390 -980
rect 42290 -1060 42310 -1000
rect 42370 -1060 42390 -1000
rect 42290 -1100 42390 -1060
rect 42290 -1160 42310 -1100
rect 42370 -1160 42390 -1100
rect 42290 -1200 42390 -1160
rect 42290 -1260 42310 -1200
rect 42370 -1260 42390 -1200
rect 42290 -1300 42390 -1260
rect 42290 -1360 42310 -1300
rect 42370 -1360 42390 -1300
rect 42290 -1380 42390 -1360
rect 42460 -1000 42560 -980
rect 42460 -1060 42480 -1000
rect 42540 -1060 42560 -1000
rect 42460 -1100 42560 -1060
rect 42460 -1160 42480 -1100
rect 42540 -1160 42560 -1100
rect 42460 -1200 42560 -1160
rect 42460 -1260 42480 -1200
rect 42540 -1260 42560 -1200
rect 42460 -1300 42560 -1260
rect 42460 -1360 42480 -1300
rect 42540 -1360 42560 -1300
rect 42460 -1380 42560 -1360
rect 42630 -1000 42730 -980
rect 42630 -1060 42650 -1000
rect 42710 -1060 42730 -1000
rect 42630 -1100 42730 -1060
rect 42630 -1160 42650 -1100
rect 42710 -1160 42730 -1100
rect 42630 -1200 42730 -1160
rect 42630 -1260 42650 -1200
rect 42710 -1260 42730 -1200
rect 42630 -1300 42730 -1260
rect 42630 -1360 42650 -1300
rect 42710 -1360 42730 -1300
rect 42630 -1380 42730 -1360
rect 42800 -1000 42900 -980
rect 42800 -1060 42820 -1000
rect 42880 -1060 42900 -1000
rect 42800 -1100 42900 -1060
rect 42800 -1160 42820 -1100
rect 42880 -1160 42900 -1100
rect 42800 -1200 42900 -1160
rect 42800 -1260 42820 -1200
rect 42880 -1260 42900 -1200
rect 42800 -1300 42900 -1260
rect 42800 -1360 42820 -1300
rect 42880 -1360 42900 -1300
rect 42800 -1380 42900 -1360
rect 42970 -1000 43070 -980
rect 42970 -1060 42990 -1000
rect 43050 -1060 43070 -1000
rect 42970 -1100 43070 -1060
rect 42970 -1160 42990 -1100
rect 43050 -1160 43070 -1100
rect 42970 -1200 43070 -1160
rect 42970 -1260 42990 -1200
rect 43050 -1260 43070 -1200
rect 42970 -1300 43070 -1260
rect 42970 -1360 42990 -1300
rect 43050 -1360 43070 -1300
rect 42970 -1380 43070 -1360
rect 43140 -1000 43240 -980
rect 43140 -1060 43160 -1000
rect 43220 -1060 43240 -1000
rect 43140 -1100 43240 -1060
rect 43140 -1160 43160 -1100
rect 43220 -1160 43240 -1100
rect 43140 -1200 43240 -1160
rect 43140 -1260 43160 -1200
rect 43220 -1260 43240 -1200
rect 43140 -1300 43240 -1260
rect 43140 -1360 43160 -1300
rect 43220 -1360 43240 -1300
rect 43140 -1380 43240 -1360
rect 43310 -1000 43410 -980
rect 43310 -1060 43330 -1000
rect 43390 -1060 43410 -1000
rect 43310 -1100 43410 -1060
rect 43310 -1160 43330 -1100
rect 43390 -1160 43410 -1100
rect 43310 -1200 43410 -1160
rect 43310 -1260 43330 -1200
rect 43390 -1260 43410 -1200
rect 43310 -1300 43410 -1260
rect 43310 -1360 43330 -1300
rect 43390 -1360 43410 -1300
rect 43310 -1380 43410 -1360
rect 43480 -1000 43580 -980
rect 43480 -1060 43500 -1000
rect 43560 -1060 43580 -1000
rect 43480 -1100 43580 -1060
rect 43480 -1160 43500 -1100
rect 43560 -1160 43580 -1100
rect 43480 -1200 43580 -1160
rect 43480 -1260 43500 -1200
rect 43560 -1260 43580 -1200
rect 43480 -1300 43580 -1260
rect 43480 -1360 43500 -1300
rect 43560 -1360 43580 -1300
rect 43480 -1380 43580 -1360
rect 43650 -1000 43750 -980
rect 43650 -1060 43670 -1000
rect 43730 -1060 43750 -1000
rect 43650 -1100 43750 -1060
rect 43650 -1160 43670 -1100
rect 43730 -1160 43750 -1100
rect 43650 -1200 43750 -1160
rect 43650 -1260 43670 -1200
rect 43730 -1260 43750 -1200
rect 43650 -1300 43750 -1260
rect 43650 -1360 43670 -1300
rect 43730 -1360 43750 -1300
rect 43650 -1380 43750 -1360
rect 43820 -1000 43920 -980
rect 43820 -1060 43840 -1000
rect 43900 -1060 43920 -1000
rect 43820 -1100 43920 -1060
rect 43820 -1160 43840 -1100
rect 43900 -1160 43920 -1100
rect 43820 -1200 43920 -1160
rect 43820 -1260 43840 -1200
rect 43900 -1260 43920 -1200
rect 43820 -1300 43920 -1260
rect 43820 -1360 43840 -1300
rect 43900 -1360 43920 -1300
rect 43820 -1380 43920 -1360
rect 43990 -1000 44090 -980
rect 43990 -1060 44010 -1000
rect 44070 -1060 44090 -1000
rect 43990 -1100 44090 -1060
rect 43990 -1160 44010 -1100
rect 44070 -1160 44090 -1100
rect 43990 -1200 44090 -1160
rect 43990 -1260 44010 -1200
rect 44070 -1260 44090 -1200
rect 43990 -1300 44090 -1260
rect 43990 -1360 44010 -1300
rect 44070 -1360 44090 -1300
rect 43990 -1380 44090 -1360
rect 44160 -1000 44260 -980
rect 44160 -1060 44180 -1000
rect 44240 -1060 44260 -1000
rect 44160 -1100 44260 -1060
rect 44160 -1160 44180 -1100
rect 44240 -1160 44260 -1100
rect 44160 -1200 44260 -1160
rect 44160 -1260 44180 -1200
rect 44240 -1260 44260 -1200
rect 44160 -1300 44260 -1260
rect 44160 -1360 44180 -1300
rect 44240 -1360 44260 -1300
rect 44160 -1380 44260 -1360
rect 44330 -1000 44430 -980
rect 44330 -1060 44350 -1000
rect 44410 -1060 44430 -1000
rect 44330 -1100 44430 -1060
rect 44330 -1160 44350 -1100
rect 44410 -1160 44430 -1100
rect 44330 -1200 44430 -1160
rect 44330 -1260 44350 -1200
rect 44410 -1260 44430 -1200
rect 44330 -1300 44430 -1260
rect 44330 -1360 44350 -1300
rect 44410 -1360 44430 -1300
rect 44330 -1380 44430 -1360
rect 44500 -1000 44600 -980
rect 44500 -1060 44520 -1000
rect 44580 -1060 44600 -1000
rect 44500 -1100 44600 -1060
rect 44500 -1160 44520 -1100
rect 44580 -1160 44600 -1100
rect 44500 -1200 44600 -1160
rect 44500 -1260 44520 -1200
rect 44580 -1260 44600 -1200
rect 44500 -1300 44600 -1260
rect 44500 -1360 44520 -1300
rect 44580 -1360 44600 -1300
rect 44500 -1380 44600 -1360
rect 44670 -1000 44770 -980
rect 44670 -1060 44690 -1000
rect 44750 -1060 44770 -1000
rect 44670 -1100 44770 -1060
rect 44670 -1160 44690 -1100
rect 44750 -1160 44770 -1100
rect 44670 -1200 44770 -1160
rect 44670 -1260 44690 -1200
rect 44750 -1260 44770 -1200
rect 44670 -1300 44770 -1260
rect 44670 -1360 44690 -1300
rect 44750 -1360 44770 -1300
rect 44670 -1380 44770 -1360
rect 44840 -1000 44940 -980
rect 44840 -1060 44860 -1000
rect 44920 -1060 44940 -1000
rect 44840 -1100 44940 -1060
rect 44840 -1160 44860 -1100
rect 44920 -1160 44940 -1100
rect 44840 -1200 44940 -1160
rect 44840 -1260 44860 -1200
rect 44920 -1260 44940 -1200
rect 44840 -1300 44940 -1260
rect 44840 -1360 44860 -1300
rect 44920 -1360 44940 -1300
rect 44840 -1380 44940 -1360
rect 45010 -1000 45110 -980
rect 45010 -1060 45030 -1000
rect 45090 -1060 45110 -1000
rect 45010 -1100 45110 -1060
rect 45010 -1160 45030 -1100
rect 45090 -1160 45110 -1100
rect 45010 -1200 45110 -1160
rect 45010 -1260 45030 -1200
rect 45090 -1260 45110 -1200
rect 45010 -1300 45110 -1260
rect 45010 -1360 45030 -1300
rect 45090 -1360 45110 -1300
rect 45010 -1380 45110 -1360
rect 45180 -1000 45280 -980
rect 45180 -1060 45200 -1000
rect 45260 -1060 45280 -1000
rect 45180 -1100 45280 -1060
rect 45180 -1160 45200 -1100
rect 45260 -1160 45280 -1100
rect 45180 -1200 45280 -1160
rect 45180 -1260 45200 -1200
rect 45260 -1260 45280 -1200
rect 45180 -1300 45280 -1260
rect 45180 -1360 45200 -1300
rect 45260 -1360 45280 -1300
rect 45180 -1380 45280 -1360
rect 45350 -1000 45450 -980
rect 45350 -1060 45370 -1000
rect 45430 -1060 45450 -1000
rect 45350 -1100 45450 -1060
rect 45350 -1160 45370 -1100
rect 45430 -1160 45450 -1100
rect 45350 -1200 45450 -1160
rect 45350 -1260 45370 -1200
rect 45430 -1260 45450 -1200
rect 45350 -1300 45450 -1260
rect 45350 -1360 45370 -1300
rect 45430 -1360 45450 -1300
rect 45350 -1380 45450 -1360
rect 45520 -1000 45620 -980
rect 45520 -1060 45540 -1000
rect 45600 -1060 45620 -1000
rect 45520 -1100 45620 -1060
rect 45520 -1160 45540 -1100
rect 45600 -1160 45620 -1100
rect 45520 -1200 45620 -1160
rect 45520 -1260 45540 -1200
rect 45600 -1260 45620 -1200
rect 45520 -1300 45620 -1260
rect 45520 -1360 45540 -1300
rect 45600 -1360 45620 -1300
rect 45520 -1380 45620 -1360
rect 45690 -1000 45790 -980
rect 45690 -1060 45710 -1000
rect 45770 -1060 45790 -1000
rect 45690 -1100 45790 -1060
rect 45690 -1160 45710 -1100
rect 45770 -1160 45790 -1100
rect 45690 -1200 45790 -1160
rect 45690 -1260 45710 -1200
rect 45770 -1260 45790 -1200
rect 45690 -1300 45790 -1260
rect 45690 -1360 45710 -1300
rect 45770 -1360 45790 -1300
rect 45690 -1380 45790 -1360
rect 45860 -1000 45960 -980
rect 45860 -1060 45880 -1000
rect 45940 -1060 45960 -1000
rect 45860 -1100 45960 -1060
rect 45860 -1160 45880 -1100
rect 45940 -1160 45960 -1100
rect 45860 -1200 45960 -1160
rect 45860 -1260 45880 -1200
rect 45940 -1260 45960 -1200
rect 45860 -1300 45960 -1260
rect 45860 -1360 45880 -1300
rect 45940 -1360 45960 -1300
rect 45860 -1380 45960 -1360
rect 46030 -1000 46130 -980
rect 46030 -1060 46050 -1000
rect 46110 -1060 46130 -1000
rect 46030 -1100 46130 -1060
rect 46030 -1160 46050 -1100
rect 46110 -1160 46130 -1100
rect 46030 -1200 46130 -1160
rect 46030 -1260 46050 -1200
rect 46110 -1260 46130 -1200
rect 46030 -1300 46130 -1260
rect 46030 -1360 46050 -1300
rect 46110 -1360 46130 -1300
rect 46030 -1380 46130 -1360
rect 46200 -1000 46300 -980
rect 46200 -1060 46220 -1000
rect 46280 -1060 46300 -1000
rect 46200 -1100 46300 -1060
rect 46200 -1160 46220 -1100
rect 46280 -1160 46300 -1100
rect 46200 -1200 46300 -1160
rect 46200 -1260 46220 -1200
rect 46280 -1260 46300 -1200
rect 46200 -1300 46300 -1260
rect 46200 -1360 46220 -1300
rect 46280 -1360 46300 -1300
rect 46200 -1380 46300 -1360
rect 46370 -1000 46470 -980
rect 46370 -1060 46390 -1000
rect 46450 -1060 46470 -1000
rect 46370 -1100 46470 -1060
rect 46370 -1160 46390 -1100
rect 46450 -1160 46470 -1100
rect 46370 -1200 46470 -1160
rect 46370 -1260 46390 -1200
rect 46450 -1260 46470 -1200
rect 46370 -1300 46470 -1260
rect 46370 -1360 46390 -1300
rect 46450 -1360 46470 -1300
rect 46370 -1380 46470 -1360
rect 46540 -1000 46640 -980
rect 46540 -1060 46560 -1000
rect 46620 -1060 46640 -1000
rect 46540 -1100 46640 -1060
rect 46540 -1160 46560 -1100
rect 46620 -1160 46640 -1100
rect 46540 -1200 46640 -1160
rect 46540 -1260 46560 -1200
rect 46620 -1260 46640 -1200
rect 46540 -1300 46640 -1260
rect 46540 -1360 46560 -1300
rect 46620 -1360 46640 -1300
rect 46540 -1380 46640 -1360
rect 46710 -1000 46810 -980
rect 46710 -1060 46730 -1000
rect 46790 -1060 46810 -1000
rect 46710 -1100 46810 -1060
rect 46710 -1160 46730 -1100
rect 46790 -1160 46810 -1100
rect 46710 -1200 46810 -1160
rect 46710 -1260 46730 -1200
rect 46790 -1260 46810 -1200
rect 46710 -1300 46810 -1260
rect 46710 -1360 46730 -1300
rect 46790 -1360 46810 -1300
rect 46710 -1380 46810 -1360
rect 46880 -1000 46980 -980
rect 46880 -1060 46900 -1000
rect 46960 -1060 46980 -1000
rect 46880 -1100 46980 -1060
rect 46880 -1160 46900 -1100
rect 46960 -1160 46980 -1100
rect 46880 -1200 46980 -1160
rect 46880 -1260 46900 -1200
rect 46960 -1260 46980 -1200
rect 46880 -1300 46980 -1260
rect 46880 -1360 46900 -1300
rect 46960 -1360 46980 -1300
rect 46880 -1380 46980 -1360
rect 47050 -1000 47150 -980
rect 47050 -1060 47070 -1000
rect 47130 -1060 47150 -1000
rect 47050 -1100 47150 -1060
rect 47050 -1160 47070 -1100
rect 47130 -1160 47150 -1100
rect 47050 -1200 47150 -1160
rect 47050 -1260 47070 -1200
rect 47130 -1260 47150 -1200
rect 47050 -1300 47150 -1260
rect 47050 -1360 47070 -1300
rect 47130 -1360 47150 -1300
rect 47050 -1380 47150 -1360
rect 47220 -1000 47320 -980
rect 47220 -1060 47240 -1000
rect 47300 -1060 47320 -1000
rect 47220 -1100 47320 -1060
rect 47220 -1160 47240 -1100
rect 47300 -1160 47320 -1100
rect 47220 -1200 47320 -1160
rect 47220 -1260 47240 -1200
rect 47300 -1260 47320 -1200
rect 47220 -1300 47320 -1260
rect 47220 -1360 47240 -1300
rect 47300 -1360 47320 -1300
rect 47220 -1380 47320 -1360
rect 47390 -1000 47490 -980
rect 47390 -1060 47410 -1000
rect 47470 -1060 47490 -1000
rect 47390 -1100 47490 -1060
rect 47390 -1160 47410 -1100
rect 47470 -1160 47490 -1100
rect 47390 -1200 47490 -1160
rect 47390 -1260 47410 -1200
rect 47470 -1260 47490 -1200
rect 47390 -1300 47490 -1260
rect 47390 -1360 47410 -1300
rect 47470 -1360 47490 -1300
rect 47390 -1380 47490 -1360
rect 47560 -1000 47660 -980
rect 47560 -1060 47580 -1000
rect 47640 -1060 47660 -1000
rect 47560 -1100 47660 -1060
rect 47560 -1160 47580 -1100
rect 47640 -1160 47660 -1100
rect 47560 -1200 47660 -1160
rect 47560 -1260 47580 -1200
rect 47640 -1260 47660 -1200
rect 47560 -1300 47660 -1260
rect 47560 -1360 47580 -1300
rect 47640 -1360 47660 -1300
rect 47560 -1380 47660 -1360
rect 47730 -1000 47830 -980
rect 47730 -1060 47750 -1000
rect 47810 -1060 47830 -1000
rect 47730 -1100 47830 -1060
rect 47730 -1160 47750 -1100
rect 47810 -1160 47830 -1100
rect 47730 -1200 47830 -1160
rect 47730 -1260 47750 -1200
rect 47810 -1260 47830 -1200
rect 47730 -1300 47830 -1260
rect 47730 -1360 47750 -1300
rect 47810 -1360 47830 -1300
rect 47730 -1380 47830 -1360
rect 47900 -1000 48000 -980
rect 47900 -1060 47920 -1000
rect 47980 -1060 48000 -1000
rect 47900 -1100 48000 -1060
rect 47900 -1160 47920 -1100
rect 47980 -1160 48000 -1100
rect 47900 -1200 48000 -1160
rect 47900 -1260 47920 -1200
rect 47980 -1260 48000 -1200
rect 47900 -1300 48000 -1260
rect 47900 -1360 47920 -1300
rect 47980 -1360 48000 -1300
rect 47900 -1380 48000 -1360
rect 48070 -1000 48170 -980
rect 48070 -1060 48090 -1000
rect 48150 -1060 48170 -1000
rect 48070 -1100 48170 -1060
rect 48070 -1160 48090 -1100
rect 48150 -1160 48170 -1100
rect 48070 -1200 48170 -1160
rect 48070 -1260 48090 -1200
rect 48150 -1260 48170 -1200
rect 48070 -1300 48170 -1260
rect 48070 -1360 48090 -1300
rect 48150 -1360 48170 -1300
rect 48070 -1380 48170 -1360
rect 48240 -1000 48340 -980
rect 48240 -1060 48260 -1000
rect 48320 -1060 48340 -1000
rect 48240 -1100 48340 -1060
rect 48240 -1160 48260 -1100
rect 48320 -1160 48340 -1100
rect 48240 -1200 48340 -1160
rect 48240 -1260 48260 -1200
rect 48320 -1260 48340 -1200
rect 48240 -1300 48340 -1260
rect 48240 -1360 48260 -1300
rect 48320 -1360 48340 -1300
rect 48240 -1380 48340 -1360
rect 48410 -1000 48510 -980
rect 48410 -1060 48430 -1000
rect 48490 -1060 48510 -1000
rect 48410 -1100 48510 -1060
rect 48410 -1160 48430 -1100
rect 48490 -1160 48510 -1100
rect 48410 -1200 48510 -1160
rect 48410 -1260 48430 -1200
rect 48490 -1260 48510 -1200
rect 48410 -1300 48510 -1260
rect 48410 -1360 48430 -1300
rect 48490 -1360 48510 -1300
rect 48410 -1380 48510 -1360
rect 48580 -1000 48680 -980
rect 48580 -1060 48600 -1000
rect 48660 -1060 48680 -1000
rect 48580 -1100 48680 -1060
rect 48580 -1160 48600 -1100
rect 48660 -1160 48680 -1100
rect 48580 -1200 48680 -1160
rect 48580 -1260 48600 -1200
rect 48660 -1260 48680 -1200
rect 48580 -1300 48680 -1260
rect 48580 -1360 48600 -1300
rect 48660 -1360 48680 -1300
rect 48580 -1380 48680 -1360
rect 48750 -1000 48850 -980
rect 48750 -1060 48770 -1000
rect 48830 -1060 48850 -1000
rect 48750 -1100 48850 -1060
rect 48750 -1160 48770 -1100
rect 48830 -1160 48850 -1100
rect 48750 -1200 48850 -1160
rect 48750 -1260 48770 -1200
rect 48830 -1260 48850 -1200
rect 48750 -1300 48850 -1260
rect 48750 -1360 48770 -1300
rect 48830 -1360 48850 -1300
rect 48750 -1380 48850 -1360
rect 48920 -1000 49020 -980
rect 48920 -1060 48940 -1000
rect 49000 -1060 49020 -1000
rect 48920 -1100 49020 -1060
rect 48920 -1160 48940 -1100
rect 49000 -1160 49020 -1100
rect 48920 -1200 49020 -1160
rect 48920 -1260 48940 -1200
rect 49000 -1260 49020 -1200
rect 48920 -1300 49020 -1260
rect 48920 -1360 48940 -1300
rect 49000 -1360 49020 -1300
rect 48920 -1380 49020 -1360
rect 49090 -1000 49190 -980
rect 49090 -1060 49110 -1000
rect 49170 -1060 49190 -1000
rect 49090 -1100 49190 -1060
rect 49090 -1160 49110 -1100
rect 49170 -1160 49190 -1100
rect 49090 -1200 49190 -1160
rect 49090 -1260 49110 -1200
rect 49170 -1260 49190 -1200
rect 49090 -1300 49190 -1260
rect 49090 -1360 49110 -1300
rect 49170 -1360 49190 -1300
rect 49090 -1380 49190 -1360
rect 49260 -1000 49360 -980
rect 49260 -1060 49280 -1000
rect 49340 -1060 49360 -1000
rect 49260 -1100 49360 -1060
rect 49260 -1160 49280 -1100
rect 49340 -1160 49360 -1100
rect 49260 -1200 49360 -1160
rect 49260 -1260 49280 -1200
rect 49340 -1260 49360 -1200
rect 49260 -1300 49360 -1260
rect 49260 -1360 49280 -1300
rect 49340 -1360 49360 -1300
rect 49260 -1380 49360 -1360
rect 49430 -1000 49530 -980
rect 49430 -1060 49450 -1000
rect 49510 -1060 49530 -1000
rect 49430 -1100 49530 -1060
rect 49430 -1160 49450 -1100
rect 49510 -1160 49530 -1100
rect 49430 -1200 49530 -1160
rect 49430 -1260 49450 -1200
rect 49510 -1260 49530 -1200
rect 49430 -1300 49530 -1260
rect 49430 -1360 49450 -1300
rect 49510 -1360 49530 -1300
rect 49430 -1380 49530 -1360
rect 49600 -1000 49700 -980
rect 49600 -1060 49620 -1000
rect 49680 -1060 49700 -1000
rect 49600 -1100 49700 -1060
rect 49600 -1160 49620 -1100
rect 49680 -1160 49700 -1100
rect 49600 -1200 49700 -1160
rect 49600 -1260 49620 -1200
rect 49680 -1260 49700 -1200
rect 49600 -1300 49700 -1260
rect 49600 -1360 49620 -1300
rect 49680 -1360 49700 -1300
rect 49600 -1380 49700 -1360
rect 49770 -1000 49870 -980
rect 49770 -1060 49790 -1000
rect 49850 -1060 49870 -1000
rect 49770 -1100 49870 -1060
rect 49770 -1160 49790 -1100
rect 49850 -1160 49870 -1100
rect 49770 -1200 49870 -1160
rect 49770 -1260 49790 -1200
rect 49850 -1260 49870 -1200
rect 49770 -1300 49870 -1260
rect 49770 -1360 49790 -1300
rect 49850 -1360 49870 -1300
rect 49770 -1380 49870 -1360
rect 49940 -1000 50040 -980
rect 49940 -1060 49960 -1000
rect 50020 -1060 50040 -1000
rect 49940 -1100 50040 -1060
rect 49940 -1160 49960 -1100
rect 50020 -1160 50040 -1100
rect 49940 -1200 50040 -1160
rect 49940 -1260 49960 -1200
rect 50020 -1260 50040 -1200
rect 49940 -1300 50040 -1260
rect 49940 -1360 49960 -1300
rect 50020 -1360 50040 -1300
rect 49940 -1380 50040 -1360
rect 50110 -1000 50210 -980
rect 50110 -1060 50130 -1000
rect 50190 -1060 50210 -1000
rect 50110 -1100 50210 -1060
rect 50110 -1160 50130 -1100
rect 50190 -1160 50210 -1100
rect 50110 -1200 50210 -1160
rect 50110 -1260 50130 -1200
rect 50190 -1260 50210 -1200
rect 50110 -1300 50210 -1260
rect 50110 -1360 50130 -1300
rect 50190 -1360 50210 -1300
rect 50110 -1380 50210 -1360
rect 50280 -1000 50380 -980
rect 50280 -1060 50300 -1000
rect 50360 -1060 50380 -1000
rect 50280 -1100 50380 -1060
rect 50280 -1160 50300 -1100
rect 50360 -1160 50380 -1100
rect 50280 -1200 50380 -1160
rect 50280 -1260 50300 -1200
rect 50360 -1260 50380 -1200
rect 50280 -1300 50380 -1260
rect 50280 -1360 50300 -1300
rect 50360 -1360 50380 -1300
rect 50280 -1380 50380 -1360
rect 50450 -1000 50550 -980
rect 50450 -1060 50470 -1000
rect 50530 -1060 50550 -1000
rect 50450 -1100 50550 -1060
rect 50450 -1160 50470 -1100
rect 50530 -1160 50550 -1100
rect 50450 -1200 50550 -1160
rect 50450 -1260 50470 -1200
rect 50530 -1260 50550 -1200
rect 50450 -1300 50550 -1260
rect 50450 -1360 50470 -1300
rect 50530 -1360 50550 -1300
rect 50450 -1380 50550 -1360
rect 50620 -1000 50720 -980
rect 50620 -1060 50640 -1000
rect 50700 -1060 50720 -1000
rect 50620 -1100 50720 -1060
rect 50620 -1160 50640 -1100
rect 50700 -1160 50720 -1100
rect 50620 -1200 50720 -1160
rect 50620 -1260 50640 -1200
rect 50700 -1260 50720 -1200
rect 50620 -1300 50720 -1260
rect 50620 -1360 50640 -1300
rect 50700 -1360 50720 -1300
rect 50620 -1380 50720 -1360
rect 50790 -1000 50890 -980
rect 50790 -1060 50810 -1000
rect 50870 -1060 50890 -1000
rect 50790 -1100 50890 -1060
rect 50790 -1160 50810 -1100
rect 50870 -1160 50890 -1100
rect 50790 -1200 50890 -1160
rect 50790 -1260 50810 -1200
rect 50870 -1260 50890 -1200
rect 50790 -1300 50890 -1260
rect 50790 -1360 50810 -1300
rect 50870 -1360 50890 -1300
rect 50790 -1380 50890 -1360
rect 50960 -1000 51060 -980
rect 50960 -1060 50980 -1000
rect 51040 -1060 51060 -1000
rect 50960 -1100 51060 -1060
rect 50960 -1160 50980 -1100
rect 51040 -1160 51060 -1100
rect 50960 -1200 51060 -1160
rect 50960 -1260 50980 -1200
rect 51040 -1260 51060 -1200
rect 50960 -1300 51060 -1260
rect 50960 -1360 50980 -1300
rect 51040 -1360 51060 -1300
rect 50960 -1380 51060 -1360
rect 51130 -1000 51230 -980
rect 51130 -1060 51150 -1000
rect 51210 -1060 51230 -1000
rect 51130 -1100 51230 -1060
rect 51130 -1160 51150 -1100
rect 51210 -1160 51230 -1100
rect 51130 -1200 51230 -1160
rect 51130 -1260 51150 -1200
rect 51210 -1260 51230 -1200
rect 51130 -1300 51230 -1260
rect 51130 -1360 51150 -1300
rect 51210 -1360 51230 -1300
rect 51130 -1380 51230 -1360
rect 51300 -1000 51400 -980
rect 51300 -1060 51320 -1000
rect 51380 -1060 51400 -1000
rect 51300 -1100 51400 -1060
rect 51300 -1160 51320 -1100
rect 51380 -1160 51400 -1100
rect 51300 -1200 51400 -1160
rect 51300 -1260 51320 -1200
rect 51380 -1260 51400 -1200
rect 51300 -1300 51400 -1260
rect 51300 -1360 51320 -1300
rect 51380 -1360 51400 -1300
rect 51300 -1380 51400 -1360
rect 51470 -1000 51570 -980
rect 51470 -1060 51490 -1000
rect 51550 -1060 51570 -1000
rect 51470 -1100 51570 -1060
rect 51470 -1160 51490 -1100
rect 51550 -1160 51570 -1100
rect 51470 -1200 51570 -1160
rect 51470 -1260 51490 -1200
rect 51550 -1260 51570 -1200
rect 51470 -1300 51570 -1260
rect 51470 -1360 51490 -1300
rect 51550 -1360 51570 -1300
rect 51470 -1380 51570 -1360
rect 51640 -1000 51740 -980
rect 51640 -1060 51660 -1000
rect 51720 -1060 51740 -1000
rect 51640 -1100 51740 -1060
rect 51640 -1160 51660 -1100
rect 51720 -1160 51740 -1100
rect 51640 -1200 51740 -1160
rect 51640 -1260 51660 -1200
rect 51720 -1260 51740 -1200
rect 51640 -1300 51740 -1260
rect 51640 -1360 51660 -1300
rect 51720 -1360 51740 -1300
rect 51640 -1380 51740 -1360
rect 51810 -1000 51910 -980
rect 51810 -1060 51830 -1000
rect 51890 -1060 51910 -1000
rect 51810 -1100 51910 -1060
rect 51810 -1160 51830 -1100
rect 51890 -1160 51910 -1100
rect 51810 -1200 51910 -1160
rect 51810 -1260 51830 -1200
rect 51890 -1260 51910 -1200
rect 51810 -1300 51910 -1260
rect 51810 -1360 51830 -1300
rect 51890 -1360 51910 -1300
rect 51810 -1380 51910 -1360
rect 51980 -1000 52080 -980
rect 51980 -1060 52000 -1000
rect 52060 -1060 52080 -1000
rect 51980 -1100 52080 -1060
rect 51980 -1160 52000 -1100
rect 52060 -1160 52080 -1100
rect 51980 -1200 52080 -1160
rect 51980 -1260 52000 -1200
rect 52060 -1260 52080 -1200
rect 51980 -1300 52080 -1260
rect 51980 -1360 52000 -1300
rect 52060 -1360 52080 -1300
rect 51980 -1380 52080 -1360
rect 52150 -1000 52250 -980
rect 52150 -1060 52170 -1000
rect 52230 -1060 52250 -1000
rect 52150 -1100 52250 -1060
rect 52150 -1160 52170 -1100
rect 52230 -1160 52250 -1100
rect 52150 -1200 52250 -1160
rect 52150 -1260 52170 -1200
rect 52230 -1260 52250 -1200
rect 52150 -1300 52250 -1260
rect 52150 -1360 52170 -1300
rect 52230 -1360 52250 -1300
rect 52150 -1380 52250 -1360
rect 52320 -1000 52420 -980
rect 52320 -1060 52340 -1000
rect 52400 -1060 52420 -1000
rect 52320 -1100 52420 -1060
rect 52320 -1160 52340 -1100
rect 52400 -1160 52420 -1100
rect 52320 -1200 52420 -1160
rect 52320 -1260 52340 -1200
rect 52400 -1260 52420 -1200
rect 52320 -1300 52420 -1260
rect 52320 -1360 52340 -1300
rect 52400 -1360 52420 -1300
rect 52320 -1380 52420 -1360
rect 52490 -1000 52590 -980
rect 52490 -1060 52510 -1000
rect 52570 -1060 52590 -1000
rect 52490 -1100 52590 -1060
rect 52490 -1160 52510 -1100
rect 52570 -1160 52590 -1100
rect 52490 -1200 52590 -1160
rect 52490 -1260 52510 -1200
rect 52570 -1260 52590 -1200
rect 52490 -1300 52590 -1260
rect 52490 -1360 52510 -1300
rect 52570 -1360 52590 -1300
rect 52490 -1380 52590 -1360
rect 52660 -1000 52760 -980
rect 52660 -1060 52680 -1000
rect 52740 -1060 52760 -1000
rect 52660 -1100 52760 -1060
rect 52660 -1160 52680 -1100
rect 52740 -1160 52760 -1100
rect 52660 -1200 52760 -1160
rect 52660 -1260 52680 -1200
rect 52740 -1260 52760 -1200
rect 52660 -1300 52760 -1260
rect 52660 -1360 52680 -1300
rect 52740 -1360 52760 -1300
rect 52660 -1380 52760 -1360
rect 52830 -1000 52930 -980
rect 52830 -1060 52850 -1000
rect 52910 -1060 52930 -1000
rect 52830 -1100 52930 -1060
rect 52830 -1160 52850 -1100
rect 52910 -1160 52930 -1100
rect 52830 -1200 52930 -1160
rect 52830 -1260 52850 -1200
rect 52910 -1260 52930 -1200
rect 52830 -1300 52930 -1260
rect 52830 -1360 52850 -1300
rect 52910 -1360 52930 -1300
rect 52830 -1380 52930 -1360
rect 53000 -1000 53100 -980
rect 53000 -1060 53020 -1000
rect 53080 -1060 53100 -1000
rect 53000 -1100 53100 -1060
rect 53000 -1160 53020 -1100
rect 53080 -1160 53100 -1100
rect 53000 -1200 53100 -1160
rect 53000 -1260 53020 -1200
rect 53080 -1260 53100 -1200
rect 53000 -1300 53100 -1260
rect 53000 -1360 53020 -1300
rect 53080 -1360 53100 -1300
rect 53000 -1380 53100 -1360
rect 53170 -1000 53270 -980
rect 53170 -1060 53190 -1000
rect 53250 -1060 53270 -1000
rect 53170 -1100 53270 -1060
rect 53170 -1160 53190 -1100
rect 53250 -1160 53270 -1100
rect 53170 -1200 53270 -1160
rect 53170 -1260 53190 -1200
rect 53250 -1260 53270 -1200
rect 53170 -1300 53270 -1260
rect 53170 -1360 53190 -1300
rect 53250 -1360 53270 -1300
rect 53170 -1380 53270 -1360
rect 53340 -1000 53440 -980
rect 53340 -1060 53360 -1000
rect 53420 -1060 53440 -1000
rect 53340 -1100 53440 -1060
rect 53340 -1160 53360 -1100
rect 53420 -1160 53440 -1100
rect 53340 -1200 53440 -1160
rect 53340 -1260 53360 -1200
rect 53420 -1260 53440 -1200
rect 53340 -1300 53440 -1260
rect 53340 -1360 53360 -1300
rect 53420 -1360 53440 -1300
rect 53340 -1380 53440 -1360
rect 53510 -1000 53610 -980
rect 53510 -1060 53530 -1000
rect 53590 -1060 53610 -1000
rect 53510 -1100 53610 -1060
rect 53510 -1160 53530 -1100
rect 53590 -1160 53610 -1100
rect 53510 -1200 53610 -1160
rect 53510 -1260 53530 -1200
rect 53590 -1260 53610 -1200
rect 53510 -1300 53610 -1260
rect 53510 -1360 53530 -1300
rect 53590 -1360 53610 -1300
rect 53510 -1380 53610 -1360
rect 53680 -1000 53780 -980
rect 53680 -1060 53700 -1000
rect 53760 -1060 53780 -1000
rect 53680 -1100 53780 -1060
rect 53680 -1160 53700 -1100
rect 53760 -1160 53780 -1100
rect 53680 -1200 53780 -1160
rect 53680 -1260 53700 -1200
rect 53760 -1260 53780 -1200
rect 53680 -1300 53780 -1260
rect 53680 -1360 53700 -1300
rect 53760 -1360 53780 -1300
rect 53680 -1380 53780 -1360
rect 53850 -1000 53950 -980
rect 53850 -1060 53870 -1000
rect 53930 -1060 53950 -1000
rect 53850 -1100 53950 -1060
rect 53850 -1160 53870 -1100
rect 53930 -1160 53950 -1100
rect 53850 -1200 53950 -1160
rect 53850 -1260 53870 -1200
rect 53930 -1260 53950 -1200
rect 53850 -1300 53950 -1260
rect 53850 -1360 53870 -1300
rect 53930 -1360 53950 -1300
rect 53850 -1380 53950 -1360
rect 54020 -1000 54120 -980
rect 54020 -1060 54040 -1000
rect 54100 -1060 54120 -1000
rect 54020 -1100 54120 -1060
rect 54020 -1160 54040 -1100
rect 54100 -1160 54120 -1100
rect 54020 -1200 54120 -1160
rect 54020 -1260 54040 -1200
rect 54100 -1260 54120 -1200
rect 54020 -1300 54120 -1260
rect 54020 -1360 54040 -1300
rect 54100 -1360 54120 -1300
rect 54020 -1380 54120 -1360
rect 54190 -1000 54290 -980
rect 54190 -1060 54210 -1000
rect 54270 -1060 54290 -1000
rect 54190 -1100 54290 -1060
rect 54190 -1160 54210 -1100
rect 54270 -1160 54290 -1100
rect 54190 -1200 54290 -1160
rect 54190 -1260 54210 -1200
rect 54270 -1260 54290 -1200
rect 54190 -1300 54290 -1260
rect 54190 -1360 54210 -1300
rect 54270 -1360 54290 -1300
rect 54190 -1380 54290 -1360
rect 54360 -1000 54460 -980
rect 54360 -1060 54380 -1000
rect 54440 -1060 54460 -1000
rect 54360 -1100 54460 -1060
rect 54360 -1160 54380 -1100
rect 54440 -1160 54460 -1100
rect 54360 -1200 54460 -1160
rect 54360 -1260 54380 -1200
rect 54440 -1260 54460 -1200
rect 54360 -1300 54460 -1260
rect 54360 -1360 54380 -1300
rect 54440 -1360 54460 -1300
rect 54360 -1380 54460 -1360
rect 54530 -1000 54630 -980
rect 54530 -1060 54550 -1000
rect 54610 -1060 54630 -1000
rect 54530 -1100 54630 -1060
rect 54530 -1160 54550 -1100
rect 54610 -1160 54630 -1100
rect 54530 -1200 54630 -1160
rect 54530 -1260 54550 -1200
rect 54610 -1260 54630 -1200
rect 54530 -1300 54630 -1260
rect 54530 -1360 54550 -1300
rect 54610 -1360 54630 -1300
rect 54530 -1380 54630 -1360
rect 54700 -1000 54800 -980
rect 54700 -1060 54720 -1000
rect 54780 -1060 54800 -1000
rect 54700 -1100 54800 -1060
rect 54700 -1160 54720 -1100
rect 54780 -1160 54800 -1100
rect 54700 -1200 54800 -1160
rect 54700 -1260 54720 -1200
rect 54780 -1260 54800 -1200
rect 54700 -1300 54800 -1260
rect 54700 -1360 54720 -1300
rect 54780 -1360 54800 -1300
rect 54700 -1380 54800 -1360
rect 54870 -1000 54970 -980
rect 54870 -1060 54890 -1000
rect 54950 -1060 54970 -1000
rect 54870 -1100 54970 -1060
rect 54870 -1160 54890 -1100
rect 54950 -1160 54970 -1100
rect 54870 -1200 54970 -1160
rect 54870 -1260 54890 -1200
rect 54950 -1260 54970 -1200
rect 54870 -1300 54970 -1260
rect 54870 -1360 54890 -1300
rect 54950 -1360 54970 -1300
rect 54870 -1380 54970 -1360
rect 55040 -1000 55140 -980
rect 55040 -1060 55060 -1000
rect 55120 -1060 55140 -1000
rect 55040 -1100 55140 -1060
rect 55040 -1160 55060 -1100
rect 55120 -1160 55140 -1100
rect 55040 -1200 55140 -1160
rect 55040 -1260 55060 -1200
rect 55120 -1260 55140 -1200
rect 55040 -1300 55140 -1260
rect 55040 -1360 55060 -1300
rect 55120 -1360 55140 -1300
rect 55040 -1380 55140 -1360
rect 55210 -1000 55310 -980
rect 55210 -1060 55230 -1000
rect 55290 -1060 55310 -1000
rect 55210 -1100 55310 -1060
rect 55210 -1160 55230 -1100
rect 55290 -1160 55310 -1100
rect 55210 -1200 55310 -1160
rect 55210 -1260 55230 -1200
rect 55290 -1260 55310 -1200
rect 55210 -1300 55310 -1260
rect 55210 -1360 55230 -1300
rect 55290 -1360 55310 -1300
rect 55210 -1380 55310 -1360
rect 55380 -1000 55480 -980
rect 55380 -1060 55400 -1000
rect 55460 -1060 55480 -1000
rect 55380 -1100 55480 -1060
rect 55380 -1160 55400 -1100
rect 55460 -1160 55480 -1100
rect 55380 -1200 55480 -1160
rect 55380 -1260 55400 -1200
rect 55460 -1260 55480 -1200
rect 55380 -1300 55480 -1260
rect 55380 -1360 55400 -1300
rect 55460 -1360 55480 -1300
rect 55380 -1380 55480 -1360
rect 55550 -1000 55650 -980
rect 55550 -1060 55570 -1000
rect 55630 -1060 55650 -1000
rect 55550 -1100 55650 -1060
rect 55550 -1160 55570 -1100
rect 55630 -1160 55650 -1100
rect 55550 -1200 55650 -1160
rect 55550 -1260 55570 -1200
rect 55630 -1260 55650 -1200
rect 55550 -1300 55650 -1260
rect 55550 -1360 55570 -1300
rect 55630 -1360 55650 -1300
rect 55550 -1380 55650 -1360
rect 55720 -1000 55820 -980
rect 55720 -1060 55740 -1000
rect 55800 -1060 55820 -1000
rect 55720 -1100 55820 -1060
rect 55720 -1160 55740 -1100
rect 55800 -1160 55820 -1100
rect 55720 -1200 55820 -1160
rect 55720 -1260 55740 -1200
rect 55800 -1260 55820 -1200
rect 55720 -1300 55820 -1260
rect 55720 -1360 55740 -1300
rect 55800 -1360 55820 -1300
rect 55720 -1380 55820 -1360
rect 55890 -1000 55990 -980
rect 55890 -1060 55910 -1000
rect 55970 -1060 55990 -1000
rect 55890 -1100 55990 -1060
rect 55890 -1160 55910 -1100
rect 55970 -1160 55990 -1100
rect 55890 -1200 55990 -1160
rect 55890 -1260 55910 -1200
rect 55970 -1260 55990 -1200
rect 55890 -1300 55990 -1260
rect 55890 -1360 55910 -1300
rect 55970 -1360 55990 -1300
rect 55890 -1380 55990 -1360
rect 56060 -1000 56160 -980
rect 56060 -1060 56080 -1000
rect 56140 -1060 56160 -1000
rect 56060 -1100 56160 -1060
rect 56060 -1160 56080 -1100
rect 56140 -1160 56160 -1100
rect 56060 -1200 56160 -1160
rect 56060 -1260 56080 -1200
rect 56140 -1260 56160 -1200
rect 56060 -1300 56160 -1260
rect 56060 -1360 56080 -1300
rect 56140 -1360 56160 -1300
rect 56060 -1380 56160 -1360
rect 56230 -1000 56330 -980
rect 56230 -1060 56250 -1000
rect 56310 -1060 56330 -1000
rect 56230 -1100 56330 -1060
rect 56230 -1160 56250 -1100
rect 56310 -1160 56330 -1100
rect 56230 -1200 56330 -1160
rect 56230 -1260 56250 -1200
rect 56310 -1260 56330 -1200
rect 56230 -1300 56330 -1260
rect 56230 -1360 56250 -1300
rect 56310 -1360 56330 -1300
rect 56230 -1380 56330 -1360
rect 56400 -1000 56500 -980
rect 56400 -1060 56420 -1000
rect 56480 -1060 56500 -1000
rect 56400 -1100 56500 -1060
rect 56400 -1160 56420 -1100
rect 56480 -1160 56500 -1100
rect 56400 -1200 56500 -1160
rect 56400 -1260 56420 -1200
rect 56480 -1260 56500 -1200
rect 56400 -1300 56500 -1260
rect 56400 -1360 56420 -1300
rect 56480 -1360 56500 -1300
rect 56400 -1380 56500 -1360
rect 56570 -1000 56670 -980
rect 56570 -1060 56590 -1000
rect 56650 -1060 56670 -1000
rect 56570 -1100 56670 -1060
rect 56570 -1160 56590 -1100
rect 56650 -1160 56670 -1100
rect 56570 -1200 56670 -1160
rect 56570 -1260 56590 -1200
rect 56650 -1260 56670 -1200
rect 56570 -1300 56670 -1260
rect 56570 -1360 56590 -1300
rect 56650 -1360 56670 -1300
rect 56570 -1380 56670 -1360
rect 56740 -1000 56840 -980
rect 56740 -1060 56760 -1000
rect 56820 -1060 56840 -1000
rect 56740 -1100 56840 -1060
rect 56740 -1160 56760 -1100
rect 56820 -1160 56840 -1100
rect 56740 -1200 56840 -1160
rect 56740 -1260 56760 -1200
rect 56820 -1260 56840 -1200
rect 56740 -1300 56840 -1260
rect 56740 -1360 56760 -1300
rect 56820 -1360 56840 -1300
rect 56740 -1380 56840 -1360
rect 56910 -1000 57010 -980
rect 56910 -1060 56930 -1000
rect 56990 -1060 57010 -1000
rect 56910 -1100 57010 -1060
rect 56910 -1160 56930 -1100
rect 56990 -1160 57010 -1100
rect 56910 -1200 57010 -1160
rect 56910 -1260 56930 -1200
rect 56990 -1260 57010 -1200
rect 56910 -1300 57010 -1260
rect 56910 -1360 56930 -1300
rect 56990 -1360 57010 -1300
rect 56910 -1380 57010 -1360
rect 57080 -1000 57180 -980
rect 57080 -1060 57100 -1000
rect 57160 -1060 57180 -1000
rect 57080 -1100 57180 -1060
rect 57080 -1160 57100 -1100
rect 57160 -1160 57180 -1100
rect 57080 -1200 57180 -1160
rect 57080 -1260 57100 -1200
rect 57160 -1260 57180 -1200
rect 57080 -1300 57180 -1260
rect 57080 -1360 57100 -1300
rect 57160 -1360 57180 -1300
rect 57080 -1380 57180 -1360
rect 57250 -1000 57350 -980
rect 57250 -1060 57270 -1000
rect 57330 -1060 57350 -1000
rect 57250 -1100 57350 -1060
rect 57250 -1160 57270 -1100
rect 57330 -1160 57350 -1100
rect 57250 -1200 57350 -1160
rect 57250 -1260 57270 -1200
rect 57330 -1260 57350 -1200
rect 57250 -1300 57350 -1260
rect 57250 -1360 57270 -1300
rect 57330 -1360 57350 -1300
rect 57250 -1380 57350 -1360
rect 57420 -1000 57520 -980
rect 57420 -1060 57440 -1000
rect 57500 -1060 57520 -1000
rect 57420 -1100 57520 -1060
rect 57420 -1160 57440 -1100
rect 57500 -1160 57520 -1100
rect 57420 -1200 57520 -1160
rect 57420 -1260 57440 -1200
rect 57500 -1260 57520 -1200
rect 57420 -1300 57520 -1260
rect 57420 -1360 57440 -1300
rect 57500 -1360 57520 -1300
rect 57420 -1380 57520 -1360
rect 57590 -1000 57690 -980
rect 57590 -1060 57610 -1000
rect 57670 -1060 57690 -1000
rect 57590 -1100 57690 -1060
rect 57590 -1160 57610 -1100
rect 57670 -1160 57690 -1100
rect 57590 -1200 57690 -1160
rect 57590 -1260 57610 -1200
rect 57670 -1260 57690 -1200
rect 57590 -1300 57690 -1260
rect 57590 -1360 57610 -1300
rect 57670 -1360 57690 -1300
rect 57590 -1380 57690 -1360
rect 57760 -1000 57860 -980
rect 57760 -1060 57780 -1000
rect 57840 -1060 57860 -1000
rect 57760 -1100 57860 -1060
rect 57760 -1160 57780 -1100
rect 57840 -1160 57860 -1100
rect 57760 -1200 57860 -1160
rect 57760 -1260 57780 -1200
rect 57840 -1260 57860 -1200
rect 57760 -1300 57860 -1260
rect 57760 -1360 57780 -1300
rect 57840 -1360 57860 -1300
rect 57760 -1380 57860 -1360
rect 57930 -1000 58030 -980
rect 57930 -1060 57950 -1000
rect 58010 -1060 58030 -1000
rect 57930 -1100 58030 -1060
rect 57930 -1160 57950 -1100
rect 58010 -1160 58030 -1100
rect 57930 -1200 58030 -1160
rect 57930 -1260 57950 -1200
rect 58010 -1260 58030 -1200
rect 57930 -1300 58030 -1260
rect 57930 -1360 57950 -1300
rect 58010 -1360 58030 -1300
rect 57930 -1380 58030 -1360
rect 58100 -1000 58200 -980
rect 58100 -1060 58120 -1000
rect 58180 -1060 58200 -1000
rect 58100 -1100 58200 -1060
rect 58100 -1160 58120 -1100
rect 58180 -1160 58200 -1100
rect 58100 -1200 58200 -1160
rect 58100 -1260 58120 -1200
rect 58180 -1260 58200 -1200
rect 58100 -1300 58200 -1260
rect 58100 -1360 58120 -1300
rect 58180 -1360 58200 -1300
rect 58100 -1380 58200 -1360
rect 58270 -1000 58370 -980
rect 58270 -1060 58290 -1000
rect 58350 -1060 58370 -1000
rect 58270 -1100 58370 -1060
rect 58270 -1160 58290 -1100
rect 58350 -1160 58370 -1100
rect 58270 -1200 58370 -1160
rect 58270 -1260 58290 -1200
rect 58350 -1260 58370 -1200
rect 58270 -1300 58370 -1260
rect 58270 -1360 58290 -1300
rect 58350 -1360 58370 -1300
rect 58270 -1380 58370 -1360
rect 58440 -1000 58540 -980
rect 58440 -1060 58460 -1000
rect 58520 -1060 58540 -1000
rect 58440 -1100 58540 -1060
rect 58440 -1160 58460 -1100
rect 58520 -1160 58540 -1100
rect 58440 -1200 58540 -1160
rect 58440 -1260 58460 -1200
rect 58520 -1260 58540 -1200
rect 58440 -1300 58540 -1260
rect 58440 -1360 58460 -1300
rect 58520 -1360 58540 -1300
rect 58440 -1380 58540 -1360
rect 58610 -1000 58710 -980
rect 58610 -1060 58630 -1000
rect 58690 -1060 58710 -1000
rect 58610 -1100 58710 -1060
rect 58610 -1160 58630 -1100
rect 58690 -1160 58710 -1100
rect 58610 -1200 58710 -1160
rect 58610 -1260 58630 -1200
rect 58690 -1260 58710 -1200
rect 58610 -1300 58710 -1260
rect 58610 -1360 58630 -1300
rect 58690 -1360 58710 -1300
rect 58610 -1380 58710 -1360
rect 58780 -1000 58880 -980
rect 58780 -1060 58800 -1000
rect 58860 -1060 58880 -1000
rect 58780 -1100 58880 -1060
rect 58780 -1160 58800 -1100
rect 58860 -1160 58880 -1100
rect 58780 -1200 58880 -1160
rect 58780 -1260 58800 -1200
rect 58860 -1260 58880 -1200
rect 58780 -1300 58880 -1260
rect 58780 -1360 58800 -1300
rect 58860 -1360 58880 -1300
rect 58780 -1380 58880 -1360
rect 58950 -1000 59050 -980
rect 58950 -1060 58970 -1000
rect 59030 -1060 59050 -1000
rect 58950 -1100 59050 -1060
rect 58950 -1160 58970 -1100
rect 59030 -1160 59050 -1100
rect 58950 -1200 59050 -1160
rect 58950 -1260 58970 -1200
rect 59030 -1260 59050 -1200
rect 58950 -1300 59050 -1260
rect 58950 -1360 58970 -1300
rect 59030 -1360 59050 -1300
rect 58950 -1380 59050 -1360
rect 59120 -1000 59220 -980
rect 59120 -1060 59140 -1000
rect 59200 -1060 59220 -1000
rect 59120 -1100 59220 -1060
rect 59120 -1160 59140 -1100
rect 59200 -1160 59220 -1100
rect 59120 -1200 59220 -1160
rect 59120 -1260 59140 -1200
rect 59200 -1260 59220 -1200
rect 59120 -1300 59220 -1260
rect 59120 -1360 59140 -1300
rect 59200 -1360 59220 -1300
rect 59120 -1380 59220 -1360
rect 59290 -1000 59390 -980
rect 59290 -1060 59310 -1000
rect 59370 -1060 59390 -1000
rect 59290 -1100 59390 -1060
rect 59290 -1160 59310 -1100
rect 59370 -1160 59390 -1100
rect 59290 -1200 59390 -1160
rect 59290 -1260 59310 -1200
rect 59370 -1260 59390 -1200
rect 59290 -1300 59390 -1260
rect 59290 -1360 59310 -1300
rect 59370 -1360 59390 -1300
rect 59290 -1380 59390 -1360
rect 59460 -1000 59560 -980
rect 59460 -1060 59480 -1000
rect 59540 -1060 59560 -1000
rect 59460 -1100 59560 -1060
rect 59460 -1160 59480 -1100
rect 59540 -1160 59560 -1100
rect 59460 -1200 59560 -1160
rect 59460 -1260 59480 -1200
rect 59540 -1260 59560 -1200
rect 59460 -1300 59560 -1260
rect 59460 -1360 59480 -1300
rect 59540 -1360 59560 -1300
rect 59460 -1380 59560 -1360
rect 59630 -1000 59730 -980
rect 59630 -1060 59650 -1000
rect 59710 -1060 59730 -1000
rect 59630 -1100 59730 -1060
rect 59630 -1160 59650 -1100
rect 59710 -1160 59730 -1100
rect 59630 -1200 59730 -1160
rect 59630 -1260 59650 -1200
rect 59710 -1260 59730 -1200
rect 59630 -1300 59730 -1260
rect 59630 -1360 59650 -1300
rect 59710 -1360 59730 -1300
rect 59630 -1380 59730 -1360
rect 59800 -1000 59900 -980
rect 59800 -1060 59820 -1000
rect 59880 -1060 59900 -1000
rect 59800 -1100 59900 -1060
rect 59800 -1160 59820 -1100
rect 59880 -1160 59900 -1100
rect 59800 -1200 59900 -1160
rect 59800 -1260 59820 -1200
rect 59880 -1260 59900 -1200
rect 59800 -1300 59900 -1260
rect 59800 -1360 59820 -1300
rect 59880 -1360 59900 -1300
rect 59800 -1380 59900 -1360
rect 59970 -1000 60070 -980
rect 59970 -1060 59990 -1000
rect 60050 -1060 60070 -1000
rect 59970 -1100 60070 -1060
rect 59970 -1160 59990 -1100
rect 60050 -1160 60070 -1100
rect 59970 -1200 60070 -1160
rect 59970 -1260 59990 -1200
rect 60050 -1260 60070 -1200
rect 59970 -1300 60070 -1260
rect 59970 -1360 59990 -1300
rect 60050 -1360 60070 -1300
rect 59970 -1380 60070 -1360
rect 60140 -1000 60240 -980
rect 60140 -1060 60160 -1000
rect 60220 -1060 60240 -1000
rect 60140 -1100 60240 -1060
rect 60140 -1160 60160 -1100
rect 60220 -1160 60240 -1100
rect 60140 -1200 60240 -1160
rect 60140 -1260 60160 -1200
rect 60220 -1260 60240 -1200
rect 60140 -1300 60240 -1260
rect 60140 -1360 60160 -1300
rect 60220 -1360 60240 -1300
rect 60140 -1380 60240 -1360
rect 60310 -1000 60410 -980
rect 60310 -1060 60330 -1000
rect 60390 -1060 60410 -1000
rect 60310 -1100 60410 -1060
rect 60310 -1160 60330 -1100
rect 60390 -1160 60410 -1100
rect 60310 -1200 60410 -1160
rect 60310 -1260 60330 -1200
rect 60390 -1260 60410 -1200
rect 60310 -1300 60410 -1260
rect 60310 -1360 60330 -1300
rect 60390 -1360 60410 -1300
rect 60310 -1380 60410 -1360
rect 60480 -1000 60580 -980
rect 60480 -1060 60500 -1000
rect 60560 -1060 60580 -1000
rect 60480 -1100 60580 -1060
rect 60480 -1160 60500 -1100
rect 60560 -1160 60580 -1100
rect 60480 -1200 60580 -1160
rect 60480 -1260 60500 -1200
rect 60560 -1260 60580 -1200
rect 60480 -1300 60580 -1260
rect 60480 -1360 60500 -1300
rect 60560 -1360 60580 -1300
rect 60480 -1380 60580 -1360
rect 60650 -1000 60750 -980
rect 60650 -1060 60670 -1000
rect 60730 -1060 60750 -1000
rect 60650 -1100 60750 -1060
rect 60650 -1160 60670 -1100
rect 60730 -1160 60750 -1100
rect 60650 -1200 60750 -1160
rect 60650 -1260 60670 -1200
rect 60730 -1260 60750 -1200
rect 60650 -1300 60750 -1260
rect 60650 -1360 60670 -1300
rect 60730 -1360 60750 -1300
rect 60650 -1380 60750 -1360
rect 60820 -1000 60920 -980
rect 60820 -1060 60840 -1000
rect 60900 -1060 60920 -1000
rect 60820 -1100 60920 -1060
rect 60820 -1160 60840 -1100
rect 60900 -1160 60920 -1100
rect 60820 -1200 60920 -1160
rect 60820 -1260 60840 -1200
rect 60900 -1260 60920 -1200
rect 60820 -1300 60920 -1260
rect 60820 -1360 60840 -1300
rect 60900 -1360 60920 -1300
rect 60820 -1380 60920 -1360
rect 60990 -1000 61090 -980
rect 60990 -1060 61010 -1000
rect 61070 -1060 61090 -1000
rect 60990 -1100 61090 -1060
rect 60990 -1160 61010 -1100
rect 61070 -1160 61090 -1100
rect 60990 -1200 61090 -1160
rect 60990 -1260 61010 -1200
rect 61070 -1260 61090 -1200
rect 60990 -1300 61090 -1260
rect 60990 -1360 61010 -1300
rect 61070 -1360 61090 -1300
rect 60990 -1380 61090 -1360
rect 61160 -1000 61260 -980
rect 61160 -1060 61180 -1000
rect 61240 -1060 61260 -1000
rect 61160 -1100 61260 -1060
rect 61160 -1160 61180 -1100
rect 61240 -1160 61260 -1100
rect 61160 -1200 61260 -1160
rect 61160 -1260 61180 -1200
rect 61240 -1260 61260 -1200
rect 61160 -1300 61260 -1260
rect 61160 -1360 61180 -1300
rect 61240 -1360 61260 -1300
rect 61160 -1380 61260 -1360
rect 61330 -1000 61430 -980
rect 61330 -1060 61350 -1000
rect 61410 -1060 61430 -1000
rect 61330 -1100 61430 -1060
rect 61330 -1160 61350 -1100
rect 61410 -1160 61430 -1100
rect 61330 -1200 61430 -1160
rect 61330 -1260 61350 -1200
rect 61410 -1260 61430 -1200
rect 61330 -1300 61430 -1260
rect 61330 -1360 61350 -1300
rect 61410 -1360 61430 -1300
rect 61330 -1380 61430 -1360
rect 61500 -1000 61600 -980
rect 61500 -1060 61520 -1000
rect 61580 -1060 61600 -1000
rect 61500 -1100 61600 -1060
rect 61500 -1160 61520 -1100
rect 61580 -1160 61600 -1100
rect 61500 -1200 61600 -1160
rect 61500 -1260 61520 -1200
rect 61580 -1260 61600 -1200
rect 61500 -1300 61600 -1260
rect 61500 -1360 61520 -1300
rect 61580 -1360 61600 -1300
rect 61500 -1380 61600 -1360
rect 61670 -1000 61770 -980
rect 61670 -1060 61690 -1000
rect 61750 -1060 61770 -1000
rect 61670 -1100 61770 -1060
rect 61670 -1160 61690 -1100
rect 61750 -1160 61770 -1100
rect 61670 -1200 61770 -1160
rect 61670 -1260 61690 -1200
rect 61750 -1260 61770 -1200
rect 61670 -1300 61770 -1260
rect 61670 -1360 61690 -1300
rect 61750 -1360 61770 -1300
rect 61670 -1380 61770 -1360
rect 61840 -1000 61940 -980
rect 61840 -1060 61860 -1000
rect 61920 -1060 61940 -1000
rect 61840 -1100 61940 -1060
rect 61840 -1160 61860 -1100
rect 61920 -1160 61940 -1100
rect 61840 -1200 61940 -1160
rect 61840 -1260 61860 -1200
rect 61920 -1260 61940 -1200
rect 61840 -1300 61940 -1260
rect 61840 -1360 61860 -1300
rect 61920 -1360 61940 -1300
rect 61840 -1380 61940 -1360
rect 62010 -1000 62110 -980
rect 62010 -1060 62030 -1000
rect 62090 -1060 62110 -1000
rect 62010 -1100 62110 -1060
rect 62010 -1160 62030 -1100
rect 62090 -1160 62110 -1100
rect 62010 -1200 62110 -1160
rect 62010 -1260 62030 -1200
rect 62090 -1260 62110 -1200
rect 62010 -1300 62110 -1260
rect 62010 -1360 62030 -1300
rect 62090 -1360 62110 -1300
rect 62010 -1380 62110 -1360
rect 62180 -1000 62280 -980
rect 62180 -1060 62200 -1000
rect 62260 -1060 62280 -1000
rect 62180 -1100 62280 -1060
rect 62180 -1160 62200 -1100
rect 62260 -1160 62280 -1100
rect 62180 -1200 62280 -1160
rect 62180 -1260 62200 -1200
rect 62260 -1260 62280 -1200
rect 62180 -1300 62280 -1260
rect 62180 -1360 62200 -1300
rect 62260 -1360 62280 -1300
rect 62180 -1380 62280 -1360
rect 62350 -1000 62450 -980
rect 62350 -1060 62370 -1000
rect 62430 -1060 62450 -1000
rect 62350 -1100 62450 -1060
rect 62350 -1160 62370 -1100
rect 62430 -1160 62450 -1100
rect 62350 -1200 62450 -1160
rect 62350 -1260 62370 -1200
rect 62430 -1260 62450 -1200
rect 62350 -1300 62450 -1260
rect 62350 -1360 62370 -1300
rect 62430 -1360 62450 -1300
rect 62350 -1380 62450 -1360
rect 62520 -1000 62620 -980
rect 62520 -1060 62540 -1000
rect 62600 -1060 62620 -1000
rect 62520 -1100 62620 -1060
rect 62520 -1160 62540 -1100
rect 62600 -1160 62620 -1100
rect 62520 -1200 62620 -1160
rect 62520 -1260 62540 -1200
rect 62600 -1260 62620 -1200
rect 62520 -1300 62620 -1260
rect 62520 -1360 62540 -1300
rect 62600 -1360 62620 -1300
rect 62520 -1380 62620 -1360
rect 62690 -1000 62790 -980
rect 62690 -1060 62710 -1000
rect 62770 -1060 62790 -1000
rect 62690 -1100 62790 -1060
rect 62690 -1160 62710 -1100
rect 62770 -1160 62790 -1100
rect 62690 -1200 62790 -1160
rect 62690 -1260 62710 -1200
rect 62770 -1260 62790 -1200
rect 62690 -1300 62790 -1260
rect 62690 -1360 62710 -1300
rect 62770 -1360 62790 -1300
rect 62690 -1380 62790 -1360
rect 62860 -1000 62960 -980
rect 62860 -1060 62880 -1000
rect 62940 -1060 62960 -1000
rect 62860 -1100 62960 -1060
rect 62860 -1160 62880 -1100
rect 62940 -1160 62960 -1100
rect 62860 -1200 62960 -1160
rect 62860 -1260 62880 -1200
rect 62940 -1260 62960 -1200
rect 62860 -1300 62960 -1260
rect 62860 -1360 62880 -1300
rect 62940 -1360 62960 -1300
rect 62860 -1380 62960 -1360
rect 63030 -1000 63130 -980
rect 63030 -1060 63050 -1000
rect 63110 -1060 63130 -1000
rect 63030 -1100 63130 -1060
rect 63030 -1160 63050 -1100
rect 63110 -1160 63130 -1100
rect 63030 -1200 63130 -1160
rect 63030 -1260 63050 -1200
rect 63110 -1260 63130 -1200
rect 63030 -1300 63130 -1260
rect 63030 -1360 63050 -1300
rect 63110 -1360 63130 -1300
rect 63030 -1380 63130 -1360
rect 63200 -1000 63300 -980
rect 63200 -1060 63220 -1000
rect 63280 -1060 63300 -1000
rect 63200 -1100 63300 -1060
rect 63200 -1160 63220 -1100
rect 63280 -1160 63300 -1100
rect 63200 -1200 63300 -1160
rect 63200 -1260 63220 -1200
rect 63280 -1260 63300 -1200
rect 63200 -1300 63300 -1260
rect 63200 -1360 63220 -1300
rect 63280 -1360 63300 -1300
rect 63200 -1380 63300 -1360
rect 63370 -1000 63470 -980
rect 63370 -1060 63390 -1000
rect 63450 -1060 63470 -1000
rect 63370 -1100 63470 -1060
rect 63370 -1160 63390 -1100
rect 63450 -1160 63470 -1100
rect 63370 -1200 63470 -1160
rect 63370 -1260 63390 -1200
rect 63450 -1260 63470 -1200
rect 63370 -1300 63470 -1260
rect 63370 -1360 63390 -1300
rect 63450 -1360 63470 -1300
rect 63370 -1380 63470 -1360
rect 63540 -1000 63640 -980
rect 63540 -1060 63560 -1000
rect 63620 -1060 63640 -1000
rect 63540 -1100 63640 -1060
rect 63540 -1160 63560 -1100
rect 63620 -1160 63640 -1100
rect 63540 -1200 63640 -1160
rect 63540 -1260 63560 -1200
rect 63620 -1260 63640 -1200
rect 63540 -1300 63640 -1260
rect 63540 -1360 63560 -1300
rect 63620 -1360 63640 -1300
rect 63540 -1380 63640 -1360
rect 63710 -1000 63810 -980
rect 63710 -1060 63730 -1000
rect 63790 -1060 63810 -1000
rect 63710 -1100 63810 -1060
rect 63710 -1160 63730 -1100
rect 63790 -1160 63810 -1100
rect 63710 -1200 63810 -1160
rect 63710 -1260 63730 -1200
rect 63790 -1260 63810 -1200
rect 63710 -1300 63810 -1260
rect 63710 -1360 63730 -1300
rect 63790 -1360 63810 -1300
rect 63710 -1380 63810 -1360
rect 63880 -1000 63980 -980
rect 63880 -1060 63900 -1000
rect 63960 -1060 63980 -1000
rect 63880 -1100 63980 -1060
rect 63880 -1160 63900 -1100
rect 63960 -1160 63980 -1100
rect 63880 -1200 63980 -1160
rect 63880 -1260 63900 -1200
rect 63960 -1260 63980 -1200
rect 63880 -1300 63980 -1260
rect 63880 -1360 63900 -1300
rect 63960 -1360 63980 -1300
rect 63880 -1380 63980 -1360
rect 64050 -1000 64150 -980
rect 64050 -1060 64070 -1000
rect 64130 -1060 64150 -1000
rect 64050 -1100 64150 -1060
rect 64050 -1160 64070 -1100
rect 64130 -1160 64150 -1100
rect 64050 -1200 64150 -1160
rect 64050 -1260 64070 -1200
rect 64130 -1260 64150 -1200
rect 64050 -1300 64150 -1260
rect 64050 -1360 64070 -1300
rect 64130 -1360 64150 -1300
rect 64050 -1380 64150 -1360
rect 64220 -1000 64320 -980
rect 64220 -1060 64240 -1000
rect 64300 -1060 64320 -1000
rect 64220 -1100 64320 -1060
rect 64220 -1160 64240 -1100
rect 64300 -1160 64320 -1100
rect 64220 -1200 64320 -1160
rect 64220 -1260 64240 -1200
rect 64300 -1260 64320 -1200
rect 64220 -1300 64320 -1260
rect 64220 -1360 64240 -1300
rect 64300 -1360 64320 -1300
rect 64220 -1380 64320 -1360
rect 64390 -1000 64490 -980
rect 64390 -1060 64410 -1000
rect 64470 -1060 64490 -1000
rect 64390 -1100 64490 -1060
rect 64390 -1160 64410 -1100
rect 64470 -1160 64490 -1100
rect 64390 -1200 64490 -1160
rect 64390 -1260 64410 -1200
rect 64470 -1260 64490 -1200
rect 64390 -1300 64490 -1260
rect 64390 -1360 64410 -1300
rect 64470 -1360 64490 -1300
rect 64390 -1380 64490 -1360
rect 64560 -1000 64660 -980
rect 64560 -1060 64580 -1000
rect 64640 -1060 64660 -1000
rect 64560 -1100 64660 -1060
rect 64560 -1160 64580 -1100
rect 64640 -1160 64660 -1100
rect 64560 -1200 64660 -1160
rect 64560 -1260 64580 -1200
rect 64640 -1260 64660 -1200
rect 64560 -1300 64660 -1260
rect 64560 -1360 64580 -1300
rect 64640 -1360 64660 -1300
rect 64560 -1380 64660 -1360
rect 64730 -1000 64830 -980
rect 64730 -1060 64750 -1000
rect 64810 -1060 64830 -1000
rect 64730 -1100 64830 -1060
rect 64730 -1160 64750 -1100
rect 64810 -1160 64830 -1100
rect 64730 -1200 64830 -1160
rect 64730 -1260 64750 -1200
rect 64810 -1260 64830 -1200
rect 64730 -1300 64830 -1260
rect 64730 -1360 64750 -1300
rect 64810 -1360 64830 -1300
rect 64730 -1380 64830 -1360
rect 64900 -1000 65000 -980
rect 64900 -1060 64920 -1000
rect 64980 -1060 65000 -1000
rect 64900 -1100 65000 -1060
rect 64900 -1160 64920 -1100
rect 64980 -1160 65000 -1100
rect 64900 -1200 65000 -1160
rect 64900 -1260 64920 -1200
rect 64980 -1260 65000 -1200
rect 64900 -1300 65000 -1260
rect 64900 -1360 64920 -1300
rect 64980 -1360 65000 -1300
rect 64900 -1380 65000 -1360
rect 65070 -1000 65170 -980
rect 65070 -1060 65090 -1000
rect 65150 -1060 65170 -1000
rect 65070 -1100 65170 -1060
rect 65070 -1160 65090 -1100
rect 65150 -1160 65170 -1100
rect 65070 -1200 65170 -1160
rect 65070 -1260 65090 -1200
rect 65150 -1260 65170 -1200
rect 65070 -1300 65170 -1260
rect 65070 -1360 65090 -1300
rect 65150 -1360 65170 -1300
rect 65070 -1380 65170 -1360
rect 65240 -1000 65340 -980
rect 65240 -1060 65260 -1000
rect 65320 -1060 65340 -1000
rect 65240 -1100 65340 -1060
rect 65240 -1160 65260 -1100
rect 65320 -1160 65340 -1100
rect 65240 -1200 65340 -1160
rect 65240 -1260 65260 -1200
rect 65320 -1260 65340 -1200
rect 65240 -1300 65340 -1260
rect 65240 -1360 65260 -1300
rect 65320 -1360 65340 -1300
rect 65240 -1380 65340 -1360
rect 65410 -1000 65510 -980
rect 65410 -1060 65430 -1000
rect 65490 -1060 65510 -1000
rect 65410 -1100 65510 -1060
rect 65410 -1160 65430 -1100
rect 65490 -1160 65510 -1100
rect 65410 -1200 65510 -1160
rect 65410 -1260 65430 -1200
rect 65490 -1260 65510 -1200
rect 65410 -1300 65510 -1260
rect 65410 -1360 65430 -1300
rect 65490 -1360 65510 -1300
rect 65410 -1380 65510 -1360
rect 65580 -1000 65680 -980
rect 65580 -1060 65600 -1000
rect 65660 -1060 65680 -1000
rect 65580 -1100 65680 -1060
rect 65580 -1160 65600 -1100
rect 65660 -1160 65680 -1100
rect 65580 -1200 65680 -1160
rect 65580 -1260 65600 -1200
rect 65660 -1260 65680 -1200
rect 65580 -1300 65680 -1260
rect 65580 -1360 65600 -1300
rect 65660 -1360 65680 -1300
rect 65580 -1380 65680 -1360
rect 65750 -1000 65850 -980
rect 65750 -1060 65770 -1000
rect 65830 -1060 65850 -1000
rect 65750 -1100 65850 -1060
rect 65750 -1160 65770 -1100
rect 65830 -1160 65850 -1100
rect 65750 -1200 65850 -1160
rect 65750 -1260 65770 -1200
rect 65830 -1260 65850 -1200
rect 65750 -1300 65850 -1260
rect 65750 -1360 65770 -1300
rect 65830 -1360 65850 -1300
rect 65750 -1380 65850 -1360
rect 65920 -1000 66020 -980
rect 65920 -1060 65940 -1000
rect 66000 -1060 66020 -1000
rect 65920 -1100 66020 -1060
rect 65920 -1160 65940 -1100
rect 66000 -1160 66020 -1100
rect 65920 -1200 66020 -1160
rect 65920 -1260 65940 -1200
rect 66000 -1260 66020 -1200
rect 65920 -1300 66020 -1260
rect 65920 -1360 65940 -1300
rect 66000 -1360 66020 -1300
rect 65920 -1380 66020 -1360
rect 66090 -1000 66190 -980
rect 66090 -1060 66110 -1000
rect 66170 -1060 66190 -1000
rect 66090 -1100 66190 -1060
rect 66090 -1160 66110 -1100
rect 66170 -1160 66190 -1100
rect 66090 -1200 66190 -1160
rect 66090 -1260 66110 -1200
rect 66170 -1260 66190 -1200
rect 66090 -1300 66190 -1260
rect 66090 -1360 66110 -1300
rect 66170 -1360 66190 -1300
rect 66090 -1380 66190 -1360
rect 66260 -1000 66360 -980
rect 66260 -1060 66280 -1000
rect 66340 -1060 66360 -1000
rect 66260 -1100 66360 -1060
rect 66260 -1160 66280 -1100
rect 66340 -1160 66360 -1100
rect 66260 -1200 66360 -1160
rect 66260 -1260 66280 -1200
rect 66340 -1260 66360 -1200
rect 66260 -1300 66360 -1260
rect 66260 -1360 66280 -1300
rect 66340 -1360 66360 -1300
rect 66260 -1380 66360 -1360
rect 66430 -1000 66530 -980
rect 66430 -1060 66450 -1000
rect 66510 -1060 66530 -1000
rect 66430 -1100 66530 -1060
rect 66430 -1160 66450 -1100
rect 66510 -1160 66530 -1100
rect 66430 -1200 66530 -1160
rect 66430 -1260 66450 -1200
rect 66510 -1260 66530 -1200
rect 66430 -1300 66530 -1260
rect 66430 -1360 66450 -1300
rect 66510 -1360 66530 -1300
rect 66430 -1380 66530 -1360
rect 66600 -1000 66700 -980
rect 66600 -1060 66620 -1000
rect 66680 -1060 66700 -1000
rect 66600 -1100 66700 -1060
rect 66600 -1160 66620 -1100
rect 66680 -1160 66700 -1100
rect 66600 -1200 66700 -1160
rect 66600 -1260 66620 -1200
rect 66680 -1260 66700 -1200
rect 66600 -1300 66700 -1260
rect 66600 -1360 66620 -1300
rect 66680 -1360 66700 -1300
rect 66600 -1380 66700 -1360
rect 66770 -1000 66870 -980
rect 66770 -1060 66790 -1000
rect 66850 -1060 66870 -1000
rect 66770 -1100 66870 -1060
rect 66770 -1160 66790 -1100
rect 66850 -1160 66870 -1100
rect 66770 -1200 66870 -1160
rect 66770 -1260 66790 -1200
rect 66850 -1260 66870 -1200
rect 66770 -1300 66870 -1260
rect 66770 -1360 66790 -1300
rect 66850 -1360 66870 -1300
rect 66770 -1380 66870 -1360
rect 66940 -1000 67040 -980
rect 66940 -1060 66960 -1000
rect 67020 -1060 67040 -1000
rect 66940 -1100 67040 -1060
rect 66940 -1160 66960 -1100
rect 67020 -1160 67040 -1100
rect 66940 -1200 67040 -1160
rect 66940 -1260 66960 -1200
rect 67020 -1260 67040 -1200
rect 66940 -1300 67040 -1260
rect 66940 -1360 66960 -1300
rect 67020 -1360 67040 -1300
rect 66940 -1380 67040 -1360
rect 67110 -1000 67210 -980
rect 67110 -1060 67130 -1000
rect 67190 -1060 67210 -1000
rect 67110 -1100 67210 -1060
rect 67110 -1160 67130 -1100
rect 67190 -1160 67210 -1100
rect 67110 -1200 67210 -1160
rect 67110 -1260 67130 -1200
rect 67190 -1260 67210 -1200
rect 67110 -1300 67210 -1260
rect 67110 -1360 67130 -1300
rect 67190 -1360 67210 -1300
rect 67110 -1380 67210 -1360
rect 67280 -1000 67380 -980
rect 67280 -1060 67300 -1000
rect 67360 -1060 67380 -1000
rect 67280 -1100 67380 -1060
rect 67280 -1160 67300 -1100
rect 67360 -1160 67380 -1100
rect 67280 -1200 67380 -1160
rect 67280 -1260 67300 -1200
rect 67360 -1260 67380 -1200
rect 67280 -1300 67380 -1260
rect 67280 -1360 67300 -1300
rect 67360 -1360 67380 -1300
rect 67280 -1380 67380 -1360
rect 67450 -1000 67550 -980
rect 67450 -1060 67470 -1000
rect 67530 -1060 67550 -1000
rect 67450 -1100 67550 -1060
rect 67450 -1160 67470 -1100
rect 67530 -1160 67550 -1100
rect 67450 -1200 67550 -1160
rect 67450 -1260 67470 -1200
rect 67530 -1260 67550 -1200
rect 67450 -1300 67550 -1260
rect 67450 -1360 67470 -1300
rect 67530 -1360 67550 -1300
rect 67450 -1380 67550 -1360
rect 67620 -1000 67720 -980
rect 67620 -1060 67640 -1000
rect 67700 -1060 67720 -1000
rect 67620 -1100 67720 -1060
rect 67620 -1160 67640 -1100
rect 67700 -1160 67720 -1100
rect 67620 -1200 67720 -1160
rect 67620 -1260 67640 -1200
rect 67700 -1260 67720 -1200
rect 67620 -1300 67720 -1260
rect 67620 -1360 67640 -1300
rect 67700 -1360 67720 -1300
rect 67620 -1380 67720 -1360
rect 67790 -1000 67890 -980
rect 67790 -1060 67810 -1000
rect 67870 -1060 67890 -1000
rect 67790 -1100 67890 -1060
rect 67790 -1160 67810 -1100
rect 67870 -1160 67890 -1100
rect 67790 -1200 67890 -1160
rect 67790 -1260 67810 -1200
rect 67870 -1260 67890 -1200
rect 67790 -1300 67890 -1260
rect 67790 -1360 67810 -1300
rect 67870 -1360 67890 -1300
rect 67790 -1380 67890 -1360
rect 67960 -1000 68060 -980
rect 67960 -1060 67980 -1000
rect 68040 -1060 68060 -1000
rect 67960 -1100 68060 -1060
rect 67960 -1160 67980 -1100
rect 68040 -1160 68060 -1100
rect 67960 -1200 68060 -1160
rect 67960 -1260 67980 -1200
rect 68040 -1260 68060 -1200
rect 67960 -1300 68060 -1260
rect 67960 -1360 67980 -1300
rect 68040 -1360 68060 -1300
rect 67960 -1380 68060 -1360
rect 68130 -1000 68230 -980
rect 68130 -1060 68150 -1000
rect 68210 -1060 68230 -1000
rect 68130 -1100 68230 -1060
rect 68130 -1160 68150 -1100
rect 68210 -1160 68230 -1100
rect 68130 -1200 68230 -1160
rect 68130 -1260 68150 -1200
rect 68210 -1260 68230 -1200
rect 68130 -1300 68230 -1260
rect 68130 -1360 68150 -1300
rect 68210 -1360 68230 -1300
rect 68130 -1380 68230 -1360
rect 68300 -1000 68400 -980
rect 68300 -1060 68320 -1000
rect 68380 -1060 68400 -1000
rect 68300 -1100 68400 -1060
rect 68300 -1160 68320 -1100
rect 68380 -1160 68400 -1100
rect 68300 -1200 68400 -1160
rect 68300 -1260 68320 -1200
rect 68380 -1260 68400 -1200
rect 68300 -1300 68400 -1260
rect 68300 -1360 68320 -1300
rect 68380 -1360 68400 -1300
rect 68300 -1380 68400 -1360
rect 68470 -1000 68570 -980
rect 68470 -1060 68490 -1000
rect 68550 -1060 68570 -1000
rect 68470 -1100 68570 -1060
rect 68470 -1160 68490 -1100
rect 68550 -1160 68570 -1100
rect 68470 -1200 68570 -1160
rect 68470 -1260 68490 -1200
rect 68550 -1260 68570 -1200
rect 68470 -1300 68570 -1260
rect 68470 -1360 68490 -1300
rect 68550 -1360 68570 -1300
rect 68470 -1380 68570 -1360
rect 68640 -1000 68740 -980
rect 68640 -1060 68660 -1000
rect 68720 -1060 68740 -1000
rect 68640 -1100 68740 -1060
rect 68640 -1160 68660 -1100
rect 68720 -1160 68740 -1100
rect 68640 -1200 68740 -1160
rect 68640 -1260 68660 -1200
rect 68720 -1260 68740 -1200
rect 68640 -1300 68740 -1260
rect 68640 -1360 68660 -1300
rect 68720 -1360 68740 -1300
rect 68640 -1380 68740 -1360
rect 68810 -1000 68910 -980
rect 68810 -1060 68830 -1000
rect 68890 -1060 68910 -1000
rect 68810 -1100 68910 -1060
rect 68810 -1160 68830 -1100
rect 68890 -1160 68910 -1100
rect 68810 -1200 68910 -1160
rect 68810 -1260 68830 -1200
rect 68890 -1260 68910 -1200
rect 68810 -1300 68910 -1260
rect 68810 -1360 68830 -1300
rect 68890 -1360 68910 -1300
rect 68810 -1380 68910 -1360
rect 68980 -1000 69080 -980
rect 68980 -1060 69000 -1000
rect 69060 -1060 69080 -1000
rect 68980 -1100 69080 -1060
rect 68980 -1160 69000 -1100
rect 69060 -1160 69080 -1100
rect 68980 -1200 69080 -1160
rect 68980 -1260 69000 -1200
rect 69060 -1260 69080 -1200
rect 68980 -1300 69080 -1260
rect 68980 -1360 69000 -1300
rect 69060 -1360 69080 -1300
rect 68980 -1380 69080 -1360
rect 69150 -1000 69250 -980
rect 69150 -1060 69170 -1000
rect 69230 -1060 69250 -1000
rect 69150 -1100 69250 -1060
rect 69150 -1160 69170 -1100
rect 69230 -1160 69250 -1100
rect 69150 -1200 69250 -1160
rect 69150 -1260 69170 -1200
rect 69230 -1260 69250 -1200
rect 69150 -1300 69250 -1260
rect 69150 -1360 69170 -1300
rect 69230 -1360 69250 -1300
rect 69150 -1380 69250 -1360
rect 69320 -1000 69420 -980
rect 69320 -1060 69340 -1000
rect 69400 -1060 69420 -1000
rect 69320 -1100 69420 -1060
rect 69320 -1160 69340 -1100
rect 69400 -1160 69420 -1100
rect 69320 -1200 69420 -1160
rect 69320 -1260 69340 -1200
rect 69400 -1260 69420 -1200
rect 69320 -1300 69420 -1260
rect 69320 -1360 69340 -1300
rect 69400 -1360 69420 -1300
rect 69320 -1380 69420 -1360
rect 69490 -1000 69590 -980
rect 69490 -1060 69510 -1000
rect 69570 -1060 69590 -1000
rect 69490 -1100 69590 -1060
rect 69490 -1160 69510 -1100
rect 69570 -1160 69590 -1100
rect 69490 -1200 69590 -1160
rect 69490 -1260 69510 -1200
rect 69570 -1260 69590 -1200
rect 69490 -1300 69590 -1260
rect 69490 -1360 69510 -1300
rect 69570 -1360 69590 -1300
rect 69490 -1380 69590 -1360
rect 69660 -1000 69760 -980
rect 69660 -1060 69680 -1000
rect 69740 -1060 69760 -1000
rect 69660 -1100 69760 -1060
rect 69660 -1160 69680 -1100
rect 69740 -1160 69760 -1100
rect 69660 -1200 69760 -1160
rect 69660 -1260 69680 -1200
rect 69740 -1260 69760 -1200
rect 69660 -1300 69760 -1260
rect 69660 -1360 69680 -1300
rect 69740 -1360 69760 -1300
rect 69660 -1380 69760 -1360
rect 69830 -1000 69930 -980
rect 69830 -1060 69850 -1000
rect 69910 -1060 69930 -1000
rect 69830 -1100 69930 -1060
rect 69830 -1160 69850 -1100
rect 69910 -1160 69930 -1100
rect 69830 -1200 69930 -1160
rect 69830 -1260 69850 -1200
rect 69910 -1260 69930 -1200
rect 69830 -1300 69930 -1260
rect 69830 -1360 69850 -1300
rect 69910 -1360 69930 -1300
rect 69830 -1380 69930 -1360
rect 70000 -1000 70100 -980
rect 70000 -1060 70020 -1000
rect 70080 -1060 70100 -1000
rect 70000 -1100 70100 -1060
rect 70000 -1160 70020 -1100
rect 70080 -1160 70100 -1100
rect 70000 -1200 70100 -1160
rect 70000 -1260 70020 -1200
rect 70080 -1260 70100 -1200
rect 70000 -1300 70100 -1260
rect 70000 -1360 70020 -1300
rect 70080 -1360 70100 -1300
rect 70000 -1380 70100 -1360
rect 70170 -1000 70270 -980
rect 70170 -1060 70190 -1000
rect 70250 -1060 70270 -1000
rect 70170 -1100 70270 -1060
rect 70170 -1160 70190 -1100
rect 70250 -1160 70270 -1100
rect 70170 -1200 70270 -1160
rect 70170 -1260 70190 -1200
rect 70250 -1260 70270 -1200
rect 70170 -1300 70270 -1260
rect 70170 -1360 70190 -1300
rect 70250 -1360 70270 -1300
rect 70170 -1380 70270 -1360
rect 70340 -1000 70440 -980
rect 70340 -1060 70360 -1000
rect 70420 -1060 70440 -1000
rect 70340 -1100 70440 -1060
rect 70340 -1160 70360 -1100
rect 70420 -1160 70440 -1100
rect 70340 -1200 70440 -1160
rect 70340 -1260 70360 -1200
rect 70420 -1260 70440 -1200
rect 70340 -1300 70440 -1260
rect 70340 -1360 70360 -1300
rect 70420 -1360 70440 -1300
rect 70340 -1380 70440 -1360
rect 70510 -1000 70610 -980
rect 70510 -1060 70530 -1000
rect 70590 -1060 70610 -1000
rect 70510 -1100 70610 -1060
rect 70510 -1160 70530 -1100
rect 70590 -1160 70610 -1100
rect 70510 -1200 70610 -1160
rect 70510 -1260 70530 -1200
rect 70590 -1260 70610 -1200
rect 70510 -1300 70610 -1260
rect 70510 -1360 70530 -1300
rect 70590 -1360 70610 -1300
rect 70510 -1380 70610 -1360
rect 70680 -1000 70780 -980
rect 70680 -1060 70700 -1000
rect 70760 -1060 70780 -1000
rect 70680 -1100 70780 -1060
rect 70680 -1160 70700 -1100
rect 70760 -1160 70780 -1100
rect 70680 -1200 70780 -1160
rect 70680 -1260 70700 -1200
rect 70760 -1260 70780 -1200
rect 70680 -1300 70780 -1260
rect 70680 -1360 70700 -1300
rect 70760 -1360 70780 -1300
rect 70680 -1380 70780 -1360
rect 70850 -1000 70950 -980
rect 70850 -1060 70870 -1000
rect 70930 -1060 70950 -1000
rect 70850 -1100 70950 -1060
rect 70850 -1160 70870 -1100
rect 70930 -1160 70950 -1100
rect 70850 -1200 70950 -1160
rect 70850 -1260 70870 -1200
rect 70930 -1260 70950 -1200
rect 70850 -1300 70950 -1260
rect 70850 -1360 70870 -1300
rect 70930 -1360 70950 -1300
rect 70850 -1380 70950 -1360
rect 71020 -1000 71120 -980
rect 71020 -1060 71040 -1000
rect 71100 -1060 71120 -1000
rect 71020 -1100 71120 -1060
rect 71020 -1160 71040 -1100
rect 71100 -1160 71120 -1100
rect 71020 -1200 71120 -1160
rect 71020 -1260 71040 -1200
rect 71100 -1260 71120 -1200
rect 71020 -1300 71120 -1260
rect 71020 -1360 71040 -1300
rect 71100 -1360 71120 -1300
rect 71020 -1380 71120 -1360
rect 71190 -1000 71290 -980
rect 71190 -1060 71210 -1000
rect 71270 -1060 71290 -1000
rect 71190 -1100 71290 -1060
rect 71190 -1160 71210 -1100
rect 71270 -1160 71290 -1100
rect 71190 -1200 71290 -1160
rect 71190 -1260 71210 -1200
rect 71270 -1260 71290 -1200
rect 71190 -1300 71290 -1260
rect 71190 -1360 71210 -1300
rect 71270 -1360 71290 -1300
rect 71190 -1380 71290 -1360
rect 71360 -1000 71460 -980
rect 71360 -1060 71380 -1000
rect 71440 -1060 71460 -1000
rect 71360 -1100 71460 -1060
rect 71360 -1160 71380 -1100
rect 71440 -1160 71460 -1100
rect 71360 -1200 71460 -1160
rect 71360 -1260 71380 -1200
rect 71440 -1260 71460 -1200
rect 71360 -1300 71460 -1260
rect 71360 -1360 71380 -1300
rect 71440 -1360 71460 -1300
rect 71360 -1380 71460 -1360
rect 71530 -1000 71630 -980
rect 71530 -1060 71550 -1000
rect 71610 -1060 71630 -1000
rect 71530 -1100 71630 -1060
rect 71530 -1160 71550 -1100
rect 71610 -1160 71630 -1100
rect 71530 -1200 71630 -1160
rect 71530 -1260 71550 -1200
rect 71610 -1260 71630 -1200
rect 71530 -1300 71630 -1260
rect 71530 -1360 71550 -1300
rect 71610 -1360 71630 -1300
rect 71530 -1380 71630 -1360
rect 71700 -1000 71800 -980
rect 71700 -1060 71720 -1000
rect 71780 -1060 71800 -1000
rect 71700 -1100 71800 -1060
rect 71700 -1160 71720 -1100
rect 71780 -1160 71800 -1100
rect 71700 -1200 71800 -1160
rect 71700 -1260 71720 -1200
rect 71780 -1260 71800 -1200
rect 71700 -1300 71800 -1260
rect 71700 -1360 71720 -1300
rect 71780 -1360 71800 -1300
rect 71700 -1380 71800 -1360
rect 71870 -1000 71970 -980
rect 71870 -1060 71890 -1000
rect 71950 -1060 71970 -1000
rect 71870 -1100 71970 -1060
rect 71870 -1160 71890 -1100
rect 71950 -1160 71970 -1100
rect 71870 -1200 71970 -1160
rect 71870 -1260 71890 -1200
rect 71950 -1260 71970 -1200
rect 71870 -1300 71970 -1260
rect 71870 -1360 71890 -1300
rect 71950 -1360 71970 -1300
rect 71870 -1380 71970 -1360
rect 72040 -1000 72140 -980
rect 72040 -1060 72060 -1000
rect 72120 -1060 72140 -1000
rect 72040 -1100 72140 -1060
rect 72040 -1160 72060 -1100
rect 72120 -1160 72140 -1100
rect 72040 -1200 72140 -1160
rect 72040 -1260 72060 -1200
rect 72120 -1260 72140 -1200
rect 72040 -1300 72140 -1260
rect 72040 -1360 72060 -1300
rect 72120 -1360 72140 -1300
rect 72040 -1380 72140 -1360
rect 72210 -1000 72310 -980
rect 72210 -1060 72230 -1000
rect 72290 -1060 72310 -1000
rect 72210 -1100 72310 -1060
rect 72210 -1160 72230 -1100
rect 72290 -1160 72310 -1100
rect 72210 -1200 72310 -1160
rect 72210 -1260 72230 -1200
rect 72290 -1260 72310 -1200
rect 72210 -1300 72310 -1260
rect 72210 -1360 72230 -1300
rect 72290 -1360 72310 -1300
rect 72210 -1380 72310 -1360
rect 72380 -1000 72480 -980
rect 72380 -1060 72400 -1000
rect 72460 -1060 72480 -1000
rect 72380 -1100 72480 -1060
rect 72380 -1160 72400 -1100
rect 72460 -1160 72480 -1100
rect 72380 -1200 72480 -1160
rect 72380 -1260 72400 -1200
rect 72460 -1260 72480 -1200
rect 72380 -1300 72480 -1260
rect 72380 -1360 72400 -1300
rect 72460 -1360 72480 -1300
rect 72380 -1380 72480 -1360
rect 72550 -1000 72650 -980
rect 72550 -1060 72570 -1000
rect 72630 -1060 72650 -1000
rect 72550 -1100 72650 -1060
rect 72550 -1160 72570 -1100
rect 72630 -1160 72650 -1100
rect 72550 -1200 72650 -1160
rect 72550 -1260 72570 -1200
rect 72630 -1260 72650 -1200
rect 72550 -1300 72650 -1260
rect 72550 -1360 72570 -1300
rect 72630 -1360 72650 -1300
rect 72550 -1380 72650 -1360
rect 72720 -1000 72820 -980
rect 72720 -1060 72740 -1000
rect 72800 -1060 72820 -1000
rect 72720 -1100 72820 -1060
rect 72720 -1160 72740 -1100
rect 72800 -1160 72820 -1100
rect 72720 -1200 72820 -1160
rect 72720 -1260 72740 -1200
rect 72800 -1260 72820 -1200
rect 72720 -1300 72820 -1260
rect 72720 -1360 72740 -1300
rect 72800 -1360 72820 -1300
rect 72720 -1380 72820 -1360
rect 72890 -1000 72990 -980
rect 72890 -1060 72910 -1000
rect 72970 -1060 72990 -1000
rect 72890 -1100 72990 -1060
rect 72890 -1160 72910 -1100
rect 72970 -1160 72990 -1100
rect 72890 -1200 72990 -1160
rect 72890 -1260 72910 -1200
rect 72970 -1260 72990 -1200
rect 72890 -1300 72990 -1260
rect 72890 -1360 72910 -1300
rect 72970 -1360 72990 -1300
rect 72890 -1380 72990 -1360
rect 73060 -1000 73160 -980
rect 73060 -1060 73080 -1000
rect 73140 -1060 73160 -1000
rect 73060 -1100 73160 -1060
rect 73060 -1160 73080 -1100
rect 73140 -1160 73160 -1100
rect 73060 -1200 73160 -1160
rect 73060 -1260 73080 -1200
rect 73140 -1260 73160 -1200
rect 73060 -1300 73160 -1260
rect 73060 -1360 73080 -1300
rect 73140 -1360 73160 -1300
rect 73060 -1380 73160 -1360
rect 73230 -1000 73330 -980
rect 73230 -1060 73250 -1000
rect 73310 -1060 73330 -1000
rect 73230 -1100 73330 -1060
rect 73230 -1160 73250 -1100
rect 73310 -1160 73330 -1100
rect 73230 -1200 73330 -1160
rect 73230 -1260 73250 -1200
rect 73310 -1260 73330 -1200
rect 73230 -1300 73330 -1260
rect 73230 -1360 73250 -1300
rect 73310 -1360 73330 -1300
rect 73230 -1380 73330 -1360
rect 73400 -1000 73500 -980
rect 73400 -1060 73420 -1000
rect 73480 -1060 73500 -1000
rect 73400 -1100 73500 -1060
rect 73400 -1160 73420 -1100
rect 73480 -1160 73500 -1100
rect 73400 -1200 73500 -1160
rect 73400 -1260 73420 -1200
rect 73480 -1260 73500 -1200
rect 73400 -1300 73500 -1260
rect 73400 -1360 73420 -1300
rect 73480 -1360 73500 -1300
rect 73400 -1380 73500 -1360
rect 73570 -1000 73670 -980
rect 73570 -1060 73590 -1000
rect 73650 -1060 73670 -1000
rect 73570 -1100 73670 -1060
rect 73570 -1160 73590 -1100
rect 73650 -1160 73670 -1100
rect 73570 -1200 73670 -1160
rect 73570 -1260 73590 -1200
rect 73650 -1260 73670 -1200
rect 73570 -1300 73670 -1260
rect 73570 -1360 73590 -1300
rect 73650 -1360 73670 -1300
rect 73570 -1380 73670 -1360
rect 73740 -1000 73840 -980
rect 73740 -1060 73760 -1000
rect 73820 -1060 73840 -1000
rect 73740 -1100 73840 -1060
rect 73740 -1160 73760 -1100
rect 73820 -1160 73840 -1100
rect 73740 -1200 73840 -1160
rect 73740 -1260 73760 -1200
rect 73820 -1260 73840 -1200
rect 73740 -1300 73840 -1260
rect 73740 -1360 73760 -1300
rect 73820 -1360 73840 -1300
rect 73740 -1380 73840 -1360
rect 73910 -1000 74010 -980
rect 73910 -1060 73930 -1000
rect 73990 -1060 74010 -1000
rect 73910 -1100 74010 -1060
rect 73910 -1160 73930 -1100
rect 73990 -1160 74010 -1100
rect 73910 -1200 74010 -1160
rect 73910 -1260 73930 -1200
rect 73990 -1260 74010 -1200
rect 73910 -1300 74010 -1260
rect 73910 -1360 73930 -1300
rect 73990 -1360 74010 -1300
rect 73910 -1380 74010 -1360
rect 74080 -1000 74180 -980
rect 74080 -1060 74100 -1000
rect 74160 -1060 74180 -1000
rect 74080 -1100 74180 -1060
rect 74080 -1160 74100 -1100
rect 74160 -1160 74180 -1100
rect 74080 -1200 74180 -1160
rect 74080 -1260 74100 -1200
rect 74160 -1260 74180 -1200
rect 74080 -1300 74180 -1260
rect 74080 -1360 74100 -1300
rect 74160 -1360 74180 -1300
rect 74080 -1380 74180 -1360
rect 74250 -1000 74350 -980
rect 74250 -1060 74270 -1000
rect 74330 -1060 74350 -1000
rect 74250 -1100 74350 -1060
rect 74250 -1160 74270 -1100
rect 74330 -1160 74350 -1100
rect 74250 -1200 74350 -1160
rect 74250 -1260 74270 -1200
rect 74330 -1260 74350 -1200
rect 74250 -1300 74350 -1260
rect 74250 -1360 74270 -1300
rect 74330 -1360 74350 -1300
rect 74250 -1380 74350 -1360
rect 74420 -1000 74520 -980
rect 74420 -1060 74440 -1000
rect 74500 -1060 74520 -1000
rect 74420 -1100 74520 -1060
rect 74420 -1160 74440 -1100
rect 74500 -1160 74520 -1100
rect 74420 -1200 74520 -1160
rect 74420 -1260 74440 -1200
rect 74500 -1260 74520 -1200
rect 74420 -1300 74520 -1260
rect 74420 -1360 74440 -1300
rect 74500 -1360 74520 -1300
rect 74420 -1380 74520 -1360
rect 74590 -1000 74690 -980
rect 74590 -1060 74610 -1000
rect 74670 -1060 74690 -1000
rect 74590 -1100 74690 -1060
rect 74590 -1160 74610 -1100
rect 74670 -1160 74690 -1100
rect 74590 -1200 74690 -1160
rect 74590 -1260 74610 -1200
rect 74670 -1260 74690 -1200
rect 74590 -1300 74690 -1260
rect 74590 -1360 74610 -1300
rect 74670 -1360 74690 -1300
rect 74590 -1380 74690 -1360
rect 74760 -1000 74860 -980
rect 74760 -1060 74780 -1000
rect 74840 -1060 74860 -1000
rect 74760 -1100 74860 -1060
rect 74760 -1160 74780 -1100
rect 74840 -1160 74860 -1100
rect 74760 -1200 74860 -1160
rect 74760 -1260 74780 -1200
rect 74840 -1260 74860 -1200
rect 74760 -1300 74860 -1260
rect 74760 -1360 74780 -1300
rect 74840 -1360 74860 -1300
rect 74760 -1380 74860 -1360
rect 74930 -1000 75030 -980
rect 74930 -1060 74950 -1000
rect 75010 -1060 75030 -1000
rect 74930 -1100 75030 -1060
rect 74930 -1160 74950 -1100
rect 75010 -1160 75030 -1100
rect 74930 -1200 75030 -1160
rect 74930 -1260 74950 -1200
rect 75010 -1260 75030 -1200
rect 74930 -1300 75030 -1260
rect 74930 -1360 74950 -1300
rect 75010 -1360 75030 -1300
rect 74930 -1380 75030 -1360
rect 75100 -1000 75200 -980
rect 75100 -1060 75120 -1000
rect 75180 -1060 75200 -1000
rect 75100 -1100 75200 -1060
rect 75100 -1160 75120 -1100
rect 75180 -1160 75200 -1100
rect 75100 -1200 75200 -1160
rect 75100 -1260 75120 -1200
rect 75180 -1260 75200 -1200
rect 75100 -1300 75200 -1260
rect 75100 -1360 75120 -1300
rect 75180 -1360 75200 -1300
rect 75100 -1380 75200 -1360
rect 75270 -1000 75370 -980
rect 75270 -1060 75290 -1000
rect 75350 -1060 75370 -1000
rect 75270 -1100 75370 -1060
rect 75270 -1160 75290 -1100
rect 75350 -1160 75370 -1100
rect 75270 -1200 75370 -1160
rect 75270 -1260 75290 -1200
rect 75350 -1260 75370 -1200
rect 75270 -1300 75370 -1260
rect 75270 -1360 75290 -1300
rect 75350 -1360 75370 -1300
rect 75270 -1380 75370 -1360
rect 75440 -1000 75540 -980
rect 75440 -1060 75460 -1000
rect 75520 -1060 75540 -1000
rect 75440 -1100 75540 -1060
rect 75440 -1160 75460 -1100
rect 75520 -1160 75540 -1100
rect 75440 -1200 75540 -1160
rect 75440 -1260 75460 -1200
rect 75520 -1260 75540 -1200
rect 75440 -1300 75540 -1260
rect 75440 -1360 75460 -1300
rect 75520 -1360 75540 -1300
rect 75440 -1380 75540 -1360
rect 75610 -1000 75710 -980
rect 75610 -1060 75630 -1000
rect 75690 -1060 75710 -1000
rect 75610 -1100 75710 -1060
rect 75610 -1160 75630 -1100
rect 75690 -1160 75710 -1100
rect 75610 -1200 75710 -1160
rect 75610 -1260 75630 -1200
rect 75690 -1260 75710 -1200
rect 75610 -1300 75710 -1260
rect 75610 -1360 75630 -1300
rect 75690 -1360 75710 -1300
rect 75610 -1380 75710 -1360
rect 75780 -1000 75880 -980
rect 75780 -1060 75800 -1000
rect 75860 -1060 75880 -1000
rect 75780 -1100 75880 -1060
rect 75780 -1160 75800 -1100
rect 75860 -1160 75880 -1100
rect 75780 -1200 75880 -1160
rect 75780 -1260 75800 -1200
rect 75860 -1260 75880 -1200
rect 75780 -1300 75880 -1260
rect 75780 -1360 75800 -1300
rect 75860 -1360 75880 -1300
rect 75780 -1380 75880 -1360
rect 75950 -1000 76050 -980
rect 75950 -1060 75970 -1000
rect 76030 -1060 76050 -1000
rect 75950 -1100 76050 -1060
rect 75950 -1160 75970 -1100
rect 76030 -1160 76050 -1100
rect 75950 -1200 76050 -1160
rect 75950 -1260 75970 -1200
rect 76030 -1260 76050 -1200
rect 75950 -1300 76050 -1260
rect 75950 -1360 75970 -1300
rect 76030 -1360 76050 -1300
rect 75950 -1380 76050 -1360
rect 76120 -1000 76220 -980
rect 76120 -1060 76140 -1000
rect 76200 -1060 76220 -1000
rect 76120 -1100 76220 -1060
rect 76120 -1160 76140 -1100
rect 76200 -1160 76220 -1100
rect 76120 -1200 76220 -1160
rect 76120 -1260 76140 -1200
rect 76200 -1260 76220 -1200
rect 76120 -1300 76220 -1260
rect 76120 -1360 76140 -1300
rect 76200 -1360 76220 -1300
rect 76120 -1380 76220 -1360
rect 76290 -1000 76390 -980
rect 76290 -1060 76310 -1000
rect 76370 -1060 76390 -1000
rect 76290 -1100 76390 -1060
rect 76290 -1160 76310 -1100
rect 76370 -1160 76390 -1100
rect 76290 -1200 76390 -1160
rect 76290 -1260 76310 -1200
rect 76370 -1260 76390 -1200
rect 76290 -1300 76390 -1260
rect 76290 -1360 76310 -1300
rect 76370 -1360 76390 -1300
rect 76290 -1380 76390 -1360
rect 76460 -1000 76560 -980
rect 76460 -1060 76480 -1000
rect 76540 -1060 76560 -1000
rect 76460 -1100 76560 -1060
rect 76460 -1160 76480 -1100
rect 76540 -1160 76560 -1100
rect 76460 -1200 76560 -1160
rect 76460 -1260 76480 -1200
rect 76540 -1260 76560 -1200
rect 76460 -1300 76560 -1260
rect 76460 -1360 76480 -1300
rect 76540 -1360 76560 -1300
rect 76460 -1380 76560 -1360
rect 76630 -1000 76730 -980
rect 76630 -1060 76650 -1000
rect 76710 -1060 76730 -1000
rect 76630 -1100 76730 -1060
rect 76630 -1160 76650 -1100
rect 76710 -1160 76730 -1100
rect 76630 -1200 76730 -1160
rect 76630 -1260 76650 -1200
rect 76710 -1260 76730 -1200
rect 76630 -1300 76730 -1260
rect 76630 -1360 76650 -1300
rect 76710 -1360 76730 -1300
rect 76630 -1380 76730 -1360
rect 76800 -1000 76900 -980
rect 76800 -1060 76820 -1000
rect 76880 -1060 76900 -1000
rect 76800 -1100 76900 -1060
rect 76800 -1160 76820 -1100
rect 76880 -1160 76900 -1100
rect 76800 -1200 76900 -1160
rect 76800 -1260 76820 -1200
rect 76880 -1260 76900 -1200
rect 76800 -1300 76900 -1260
rect 76800 -1360 76820 -1300
rect 76880 -1360 76900 -1300
rect 76800 -1380 76900 -1360
rect 76970 -1000 77070 -980
rect 76970 -1060 76990 -1000
rect 77050 -1060 77070 -1000
rect 76970 -1100 77070 -1060
rect 76970 -1160 76990 -1100
rect 77050 -1160 77070 -1100
rect 76970 -1200 77070 -1160
rect 76970 -1260 76990 -1200
rect 77050 -1260 77070 -1200
rect 76970 -1300 77070 -1260
rect 76970 -1360 76990 -1300
rect 77050 -1360 77070 -1300
rect 76970 -1380 77070 -1360
rect 77140 -1000 77240 -980
rect 77140 -1060 77160 -1000
rect 77220 -1060 77240 -1000
rect 77140 -1100 77240 -1060
rect 77140 -1160 77160 -1100
rect 77220 -1160 77240 -1100
rect 77140 -1200 77240 -1160
rect 77140 -1260 77160 -1200
rect 77220 -1260 77240 -1200
rect 77140 -1300 77240 -1260
rect 77140 -1360 77160 -1300
rect 77220 -1360 77240 -1300
rect 77140 -1380 77240 -1360
rect 77310 -1000 77410 -980
rect 77310 -1060 77330 -1000
rect 77390 -1060 77410 -1000
rect 77310 -1100 77410 -1060
rect 77310 -1160 77330 -1100
rect 77390 -1160 77410 -1100
rect 77310 -1200 77410 -1160
rect 77310 -1260 77330 -1200
rect 77390 -1260 77410 -1200
rect 77310 -1300 77410 -1260
rect 77310 -1360 77330 -1300
rect 77390 -1360 77410 -1300
rect 77310 -1380 77410 -1360
rect 77480 -1000 77580 -980
rect 77480 -1060 77500 -1000
rect 77560 -1060 77580 -1000
rect 77480 -1100 77580 -1060
rect 77480 -1160 77500 -1100
rect 77560 -1160 77580 -1100
rect 77480 -1200 77580 -1160
rect 77480 -1260 77500 -1200
rect 77560 -1260 77580 -1200
rect 77480 -1300 77580 -1260
rect 77480 -1360 77500 -1300
rect 77560 -1360 77580 -1300
rect 77480 -1380 77580 -1360
rect 77650 -1000 77750 -980
rect 77650 -1060 77670 -1000
rect 77730 -1060 77750 -1000
rect 77650 -1100 77750 -1060
rect 77650 -1160 77670 -1100
rect 77730 -1160 77750 -1100
rect 77650 -1200 77750 -1160
rect 77650 -1260 77670 -1200
rect 77730 -1260 77750 -1200
rect 77650 -1300 77750 -1260
rect 77650 -1360 77670 -1300
rect 77730 -1360 77750 -1300
rect 77650 -1380 77750 -1360
rect 77820 -1000 77920 -980
rect 77820 -1060 77840 -1000
rect 77900 -1060 77920 -1000
rect 77820 -1100 77920 -1060
rect 77820 -1160 77840 -1100
rect 77900 -1160 77920 -1100
rect 77820 -1200 77920 -1160
rect 77820 -1260 77840 -1200
rect 77900 -1260 77920 -1200
rect 77820 -1300 77920 -1260
rect 77820 -1360 77840 -1300
rect 77900 -1360 77920 -1300
rect 77820 -1380 77920 -1360
rect 77990 -1000 78090 -980
rect 77990 -1060 78010 -1000
rect 78070 -1060 78090 -1000
rect 77990 -1100 78090 -1060
rect 77990 -1160 78010 -1100
rect 78070 -1160 78090 -1100
rect 77990 -1200 78090 -1160
rect 77990 -1260 78010 -1200
rect 78070 -1260 78090 -1200
rect 77990 -1300 78090 -1260
rect 77990 -1360 78010 -1300
rect 78070 -1360 78090 -1300
rect 77990 -1380 78090 -1360
rect 78160 -1000 78260 -980
rect 78160 -1060 78180 -1000
rect 78240 -1060 78260 -1000
rect 78160 -1100 78260 -1060
rect 78160 -1160 78180 -1100
rect 78240 -1160 78260 -1100
rect 78160 -1200 78260 -1160
rect 78160 -1260 78180 -1200
rect 78240 -1260 78260 -1200
rect 78160 -1300 78260 -1260
rect 78160 -1360 78180 -1300
rect 78240 -1360 78260 -1300
rect 78160 -1380 78260 -1360
rect 78330 -1000 78430 -980
rect 78330 -1060 78350 -1000
rect 78410 -1060 78430 -1000
rect 78330 -1100 78430 -1060
rect 78330 -1160 78350 -1100
rect 78410 -1160 78430 -1100
rect 78330 -1200 78430 -1160
rect 78330 -1260 78350 -1200
rect 78410 -1260 78430 -1200
rect 78330 -1300 78430 -1260
rect 78330 -1360 78350 -1300
rect 78410 -1360 78430 -1300
rect 78330 -1380 78430 -1360
rect 78500 -1000 78600 -980
rect 78500 -1060 78520 -1000
rect 78580 -1060 78600 -1000
rect 78500 -1100 78600 -1060
rect 78500 -1160 78520 -1100
rect 78580 -1160 78600 -1100
rect 78500 -1200 78600 -1160
rect 78500 -1260 78520 -1200
rect 78580 -1260 78600 -1200
rect 78500 -1300 78600 -1260
rect 78500 -1360 78520 -1300
rect 78580 -1360 78600 -1300
rect 78500 -1380 78600 -1360
rect 78670 -1000 78770 -980
rect 78670 -1060 78690 -1000
rect 78750 -1060 78770 -1000
rect 78670 -1100 78770 -1060
rect 78670 -1160 78690 -1100
rect 78750 -1160 78770 -1100
rect 78670 -1200 78770 -1160
rect 78670 -1260 78690 -1200
rect 78750 -1260 78770 -1200
rect 78670 -1300 78770 -1260
rect 78670 -1360 78690 -1300
rect 78750 -1360 78770 -1300
rect 78670 -1380 78770 -1360
rect 78840 -1000 78940 -980
rect 78840 -1060 78860 -1000
rect 78920 -1060 78940 -1000
rect 78840 -1100 78940 -1060
rect 78840 -1160 78860 -1100
rect 78920 -1160 78940 -1100
rect 78840 -1200 78940 -1160
rect 78840 -1260 78860 -1200
rect 78920 -1260 78940 -1200
rect 78840 -1300 78940 -1260
rect 78840 -1360 78860 -1300
rect 78920 -1360 78940 -1300
rect 78840 -1380 78940 -1360
rect 79010 -1000 79110 -980
rect 79010 -1060 79030 -1000
rect 79090 -1060 79110 -1000
rect 79010 -1100 79110 -1060
rect 79010 -1160 79030 -1100
rect 79090 -1160 79110 -1100
rect 79010 -1200 79110 -1160
rect 79010 -1260 79030 -1200
rect 79090 -1260 79110 -1200
rect 79010 -1300 79110 -1260
rect 79010 -1360 79030 -1300
rect 79090 -1360 79110 -1300
rect 79010 -1380 79110 -1360
rect 79180 -1000 79280 -980
rect 79180 -1060 79200 -1000
rect 79260 -1060 79280 -1000
rect 79180 -1100 79280 -1060
rect 79180 -1160 79200 -1100
rect 79260 -1160 79280 -1100
rect 79180 -1200 79280 -1160
rect 79180 -1260 79200 -1200
rect 79260 -1260 79280 -1200
rect 79180 -1300 79280 -1260
rect 79180 -1360 79200 -1300
rect 79260 -1360 79280 -1300
rect 79180 -1380 79280 -1360
rect 79350 -1000 79450 -980
rect 79350 -1060 79370 -1000
rect 79430 -1060 79450 -1000
rect 79350 -1100 79450 -1060
rect 79350 -1160 79370 -1100
rect 79430 -1160 79450 -1100
rect 79350 -1200 79450 -1160
rect 79350 -1260 79370 -1200
rect 79430 -1260 79450 -1200
rect 79350 -1300 79450 -1260
rect 79350 -1360 79370 -1300
rect 79430 -1360 79450 -1300
rect 79350 -1380 79450 -1360
rect 79520 -1000 79620 -980
rect 79520 -1060 79540 -1000
rect 79600 -1060 79620 -1000
rect 79520 -1100 79620 -1060
rect 79520 -1160 79540 -1100
rect 79600 -1160 79620 -1100
rect 79520 -1200 79620 -1160
rect 79520 -1260 79540 -1200
rect 79600 -1260 79620 -1200
rect 79520 -1300 79620 -1260
rect 79520 -1360 79540 -1300
rect 79600 -1360 79620 -1300
rect 79520 -1380 79620 -1360
rect 79690 -1000 79790 -980
rect 79690 -1060 79710 -1000
rect 79770 -1060 79790 -1000
rect 79690 -1100 79790 -1060
rect 79690 -1160 79710 -1100
rect 79770 -1160 79790 -1100
rect 79690 -1200 79790 -1160
rect 79690 -1260 79710 -1200
rect 79770 -1260 79790 -1200
rect 79690 -1300 79790 -1260
rect 79690 -1360 79710 -1300
rect 79770 -1360 79790 -1300
rect 79690 -1380 79790 -1360
rect 79860 -1000 79960 -980
rect 79860 -1060 79880 -1000
rect 79940 -1060 79960 -1000
rect 79860 -1100 79960 -1060
rect 79860 -1160 79880 -1100
rect 79940 -1160 79960 -1100
rect 79860 -1200 79960 -1160
rect 79860 -1260 79880 -1200
rect 79940 -1260 79960 -1200
rect 79860 -1300 79960 -1260
rect 79860 -1360 79880 -1300
rect 79940 -1360 79960 -1300
rect 79860 -1380 79960 -1360
rect 80030 -1000 80130 -980
rect 80030 -1060 80050 -1000
rect 80110 -1060 80130 -1000
rect 80030 -1100 80130 -1060
rect 80030 -1160 80050 -1100
rect 80110 -1160 80130 -1100
rect 80030 -1200 80130 -1160
rect 80030 -1260 80050 -1200
rect 80110 -1260 80130 -1200
rect 80030 -1300 80130 -1260
rect 80030 -1360 80050 -1300
rect 80110 -1360 80130 -1300
rect 80030 -1380 80130 -1360
rect 80200 -1000 80300 -980
rect 80200 -1060 80220 -1000
rect 80280 -1060 80300 -1000
rect 80200 -1100 80300 -1060
rect 80200 -1160 80220 -1100
rect 80280 -1160 80300 -1100
rect 80200 -1200 80300 -1160
rect 80200 -1260 80220 -1200
rect 80280 -1260 80300 -1200
rect 80200 -1300 80300 -1260
rect 80200 -1360 80220 -1300
rect 80280 -1360 80300 -1300
rect 80200 -1380 80300 -1360
rect 80370 -1000 80470 -980
rect 80370 -1060 80390 -1000
rect 80450 -1060 80470 -1000
rect 80370 -1100 80470 -1060
rect 80370 -1160 80390 -1100
rect 80450 -1160 80470 -1100
rect 80370 -1200 80470 -1160
rect 80370 -1260 80390 -1200
rect 80450 -1260 80470 -1200
rect 80370 -1300 80470 -1260
rect 80370 -1360 80390 -1300
rect 80450 -1360 80470 -1300
rect 80370 -1380 80470 -1360
rect 80540 -1000 80640 -980
rect 80540 -1060 80560 -1000
rect 80620 -1060 80640 -1000
rect 80540 -1100 80640 -1060
rect 80540 -1160 80560 -1100
rect 80620 -1160 80640 -1100
rect 80540 -1200 80640 -1160
rect 80540 -1260 80560 -1200
rect 80620 -1260 80640 -1200
rect 80540 -1300 80640 -1260
rect 80540 -1360 80560 -1300
rect 80620 -1360 80640 -1300
rect 80540 -1380 80640 -1360
rect 80710 -1000 80810 -980
rect 80710 -1060 80730 -1000
rect 80790 -1060 80810 -1000
rect 80710 -1100 80810 -1060
rect 80710 -1160 80730 -1100
rect 80790 -1160 80810 -1100
rect 80710 -1200 80810 -1160
rect 80710 -1260 80730 -1200
rect 80790 -1260 80810 -1200
rect 80710 -1300 80810 -1260
rect 80710 -1360 80730 -1300
rect 80790 -1360 80810 -1300
rect 80710 -1380 80810 -1360
rect 80880 -1000 80980 -980
rect 80880 -1060 80900 -1000
rect 80960 -1060 80980 -1000
rect 80880 -1100 80980 -1060
rect 80880 -1160 80900 -1100
rect 80960 -1160 80980 -1100
rect 80880 -1200 80980 -1160
rect 80880 -1260 80900 -1200
rect 80960 -1260 80980 -1200
rect 80880 -1300 80980 -1260
rect 80880 -1360 80900 -1300
rect 80960 -1360 80980 -1300
rect 80880 -1380 80980 -1360
rect 81050 -1000 81150 -980
rect 81050 -1060 81070 -1000
rect 81130 -1060 81150 -1000
rect 81050 -1100 81150 -1060
rect 81050 -1160 81070 -1100
rect 81130 -1160 81150 -1100
rect 81050 -1200 81150 -1160
rect 81050 -1260 81070 -1200
rect 81130 -1260 81150 -1200
rect 81050 -1300 81150 -1260
rect 81050 -1360 81070 -1300
rect 81130 -1360 81150 -1300
rect 81050 -1380 81150 -1360
rect 81220 -1000 81320 -980
rect 81220 -1060 81240 -1000
rect 81300 -1060 81320 -1000
rect 81220 -1100 81320 -1060
rect 81220 -1160 81240 -1100
rect 81300 -1160 81320 -1100
rect 81220 -1200 81320 -1160
rect 81220 -1260 81240 -1200
rect 81300 -1260 81320 -1200
rect 81220 -1300 81320 -1260
rect 81220 -1360 81240 -1300
rect 81300 -1360 81320 -1300
rect 81220 -1380 81320 -1360
rect 81390 -1000 81490 -980
rect 81390 -1060 81410 -1000
rect 81470 -1060 81490 -1000
rect 81390 -1100 81490 -1060
rect 81390 -1160 81410 -1100
rect 81470 -1160 81490 -1100
rect 81390 -1200 81490 -1160
rect 81390 -1260 81410 -1200
rect 81470 -1260 81490 -1200
rect 81390 -1300 81490 -1260
rect 81390 -1360 81410 -1300
rect 81470 -1360 81490 -1300
rect 81390 -1380 81490 -1360
rect 81560 -1000 81660 -980
rect 81560 -1060 81580 -1000
rect 81640 -1060 81660 -1000
rect 81560 -1100 81660 -1060
rect 81560 -1160 81580 -1100
rect 81640 -1160 81660 -1100
rect 81560 -1200 81660 -1160
rect 81560 -1260 81580 -1200
rect 81640 -1260 81660 -1200
rect 81560 -1300 81660 -1260
rect 81560 -1360 81580 -1300
rect 81640 -1360 81660 -1300
rect 81560 -1380 81660 -1360
rect 81730 -1000 81830 -980
rect 81730 -1060 81750 -1000
rect 81810 -1060 81830 -1000
rect 81730 -1100 81830 -1060
rect 81730 -1160 81750 -1100
rect 81810 -1160 81830 -1100
rect 81730 -1200 81830 -1160
rect 81730 -1260 81750 -1200
rect 81810 -1260 81830 -1200
rect 81730 -1300 81830 -1260
rect 81730 -1360 81750 -1300
rect 81810 -1360 81830 -1300
rect 81730 -1380 81830 -1360
rect 81900 -1000 82000 -980
rect 81900 -1060 81920 -1000
rect 81980 -1060 82000 -1000
rect 81900 -1100 82000 -1060
rect 81900 -1160 81920 -1100
rect 81980 -1160 82000 -1100
rect 81900 -1200 82000 -1160
rect 81900 -1260 81920 -1200
rect 81980 -1260 82000 -1200
rect 81900 -1300 82000 -1260
rect 81900 -1360 81920 -1300
rect 81980 -1360 82000 -1300
rect 81900 -1380 82000 -1360
rect 82070 -1000 82170 -980
rect 82070 -1060 82090 -1000
rect 82150 -1060 82170 -1000
rect 82070 -1100 82170 -1060
rect 82070 -1160 82090 -1100
rect 82150 -1160 82170 -1100
rect 82070 -1200 82170 -1160
rect 82070 -1260 82090 -1200
rect 82150 -1260 82170 -1200
rect 82070 -1300 82170 -1260
rect 82070 -1360 82090 -1300
rect 82150 -1360 82170 -1300
rect 82070 -1380 82170 -1360
rect 82240 -1000 82340 -980
rect 82240 -1060 82260 -1000
rect 82320 -1060 82340 -1000
rect 82240 -1100 82340 -1060
rect 82240 -1160 82260 -1100
rect 82320 -1160 82340 -1100
rect 82240 -1200 82340 -1160
rect 82240 -1260 82260 -1200
rect 82320 -1260 82340 -1200
rect 82240 -1300 82340 -1260
rect 82240 -1360 82260 -1300
rect 82320 -1360 82340 -1300
rect 82240 -1380 82340 -1360
rect 82410 -1000 82510 -980
rect 82410 -1060 82430 -1000
rect 82490 -1060 82510 -1000
rect 82410 -1100 82510 -1060
rect 82410 -1160 82430 -1100
rect 82490 -1160 82510 -1100
rect 82410 -1200 82510 -1160
rect 82410 -1260 82430 -1200
rect 82490 -1260 82510 -1200
rect 82410 -1300 82510 -1260
rect 82410 -1360 82430 -1300
rect 82490 -1360 82510 -1300
rect 82410 -1380 82510 -1360
rect 82580 -1000 82680 -980
rect 82580 -1060 82600 -1000
rect 82660 -1060 82680 -1000
rect 82580 -1100 82680 -1060
rect 82580 -1160 82600 -1100
rect 82660 -1160 82680 -1100
rect 82580 -1200 82680 -1160
rect 82580 -1260 82600 -1200
rect 82660 -1260 82680 -1200
rect 82580 -1300 82680 -1260
rect 82580 -1360 82600 -1300
rect 82660 -1360 82680 -1300
rect 82580 -1380 82680 -1360
rect 82750 -1000 82850 -980
rect 82750 -1060 82770 -1000
rect 82830 -1060 82850 -1000
rect 82750 -1100 82850 -1060
rect 82750 -1160 82770 -1100
rect 82830 -1160 82850 -1100
rect 82750 -1200 82850 -1160
rect 82750 -1260 82770 -1200
rect 82830 -1260 82850 -1200
rect 82750 -1300 82850 -1260
rect 82750 -1360 82770 -1300
rect 82830 -1360 82850 -1300
rect 82750 -1380 82850 -1360
rect 82920 -1000 83020 -980
rect 82920 -1060 82940 -1000
rect 83000 -1060 83020 -1000
rect 82920 -1100 83020 -1060
rect 82920 -1160 82940 -1100
rect 83000 -1160 83020 -1100
rect 82920 -1200 83020 -1160
rect 82920 -1260 82940 -1200
rect 83000 -1260 83020 -1200
rect 82920 -1300 83020 -1260
rect 82920 -1360 82940 -1300
rect 83000 -1360 83020 -1300
rect 82920 -1380 83020 -1360
rect 83090 -1000 83190 -980
rect 83090 -1060 83110 -1000
rect 83170 -1060 83190 -1000
rect 83090 -1100 83190 -1060
rect 83090 -1160 83110 -1100
rect 83170 -1160 83190 -1100
rect 83090 -1200 83190 -1160
rect 83090 -1260 83110 -1200
rect 83170 -1260 83190 -1200
rect 83090 -1300 83190 -1260
rect 83090 -1360 83110 -1300
rect 83170 -1360 83190 -1300
rect 83090 -1380 83190 -1360
rect 83260 -1000 83360 -980
rect 83260 -1060 83280 -1000
rect 83340 -1060 83360 -1000
rect 83260 -1100 83360 -1060
rect 83260 -1160 83280 -1100
rect 83340 -1160 83360 -1100
rect 83260 -1200 83360 -1160
rect 83260 -1260 83280 -1200
rect 83340 -1260 83360 -1200
rect 83260 -1300 83360 -1260
rect 83260 -1360 83280 -1300
rect 83340 -1360 83360 -1300
rect 83260 -1380 83360 -1360
rect 83430 -1000 83530 -980
rect 83430 -1060 83450 -1000
rect 83510 -1060 83530 -1000
rect 83430 -1100 83530 -1060
rect 83430 -1160 83450 -1100
rect 83510 -1160 83530 -1100
rect 83430 -1200 83530 -1160
rect 83430 -1260 83450 -1200
rect 83510 -1260 83530 -1200
rect 83430 -1300 83530 -1260
rect 83430 -1360 83450 -1300
rect 83510 -1360 83530 -1300
rect 83430 -1380 83530 -1360
rect 83600 -1000 83700 -980
rect 83600 -1060 83620 -1000
rect 83680 -1060 83700 -1000
rect 83600 -1100 83700 -1060
rect 83600 -1160 83620 -1100
rect 83680 -1160 83700 -1100
rect 83600 -1200 83700 -1160
rect 83600 -1260 83620 -1200
rect 83680 -1260 83700 -1200
rect 83600 -1300 83700 -1260
rect 83600 -1360 83620 -1300
rect 83680 -1360 83700 -1300
rect 83600 -1380 83700 -1360
rect 83770 -1000 83870 -980
rect 83770 -1060 83790 -1000
rect 83850 -1060 83870 -1000
rect 83770 -1100 83870 -1060
rect 83770 -1160 83790 -1100
rect 83850 -1160 83870 -1100
rect 83770 -1200 83870 -1160
rect 83770 -1260 83790 -1200
rect 83850 -1260 83870 -1200
rect 83770 -1300 83870 -1260
rect 83770 -1360 83790 -1300
rect 83850 -1360 83870 -1300
rect 83770 -1380 83870 -1360
rect 83940 -1000 84040 -980
rect 83940 -1060 83960 -1000
rect 84020 -1060 84040 -1000
rect 83940 -1100 84040 -1060
rect 83940 -1160 83960 -1100
rect 84020 -1160 84040 -1100
rect 83940 -1200 84040 -1160
rect 83940 -1260 83960 -1200
rect 84020 -1260 84040 -1200
rect 83940 -1300 84040 -1260
rect 83940 -1360 83960 -1300
rect 84020 -1360 84040 -1300
rect 83940 -1380 84040 -1360
rect 84110 -1000 84210 -980
rect 84110 -1060 84130 -1000
rect 84190 -1060 84210 -1000
rect 84110 -1100 84210 -1060
rect 84110 -1160 84130 -1100
rect 84190 -1160 84210 -1100
rect 84110 -1200 84210 -1160
rect 84110 -1260 84130 -1200
rect 84190 -1260 84210 -1200
rect 84110 -1300 84210 -1260
rect 84110 -1360 84130 -1300
rect 84190 -1360 84210 -1300
rect 84110 -1380 84210 -1360
rect 84280 -1000 84380 -980
rect 84280 -1060 84300 -1000
rect 84360 -1060 84380 -1000
rect 84280 -1100 84380 -1060
rect 84280 -1160 84300 -1100
rect 84360 -1160 84380 -1100
rect 84280 -1200 84380 -1160
rect 84280 -1260 84300 -1200
rect 84360 -1260 84380 -1200
rect 84280 -1300 84380 -1260
rect 84280 -1360 84300 -1300
rect 84360 -1360 84380 -1300
rect 84280 -1380 84380 -1360
rect 84450 -1000 84550 -980
rect 84450 -1060 84470 -1000
rect 84530 -1060 84550 -1000
rect 84450 -1100 84550 -1060
rect 84450 -1160 84470 -1100
rect 84530 -1160 84550 -1100
rect 84450 -1200 84550 -1160
rect 84450 -1260 84470 -1200
rect 84530 -1260 84550 -1200
rect 84450 -1300 84550 -1260
rect 84450 -1360 84470 -1300
rect 84530 -1360 84550 -1300
rect 84450 -1380 84550 -1360
rect 84620 -1000 84720 -980
rect 84620 -1060 84640 -1000
rect 84700 -1060 84720 -1000
rect 84620 -1100 84720 -1060
rect 84620 -1160 84640 -1100
rect 84700 -1160 84720 -1100
rect 84620 -1200 84720 -1160
rect 84620 -1260 84640 -1200
rect 84700 -1260 84720 -1200
rect 84620 -1300 84720 -1260
rect 84620 -1360 84640 -1300
rect 84700 -1360 84720 -1300
rect 84620 -1380 84720 -1360
rect 84790 -1000 84890 -980
rect 84790 -1060 84810 -1000
rect 84870 -1060 84890 -1000
rect 84790 -1100 84890 -1060
rect 84790 -1160 84810 -1100
rect 84870 -1160 84890 -1100
rect 84790 -1200 84890 -1160
rect 84790 -1260 84810 -1200
rect 84870 -1260 84890 -1200
rect 84790 -1300 84890 -1260
rect 84790 -1360 84810 -1300
rect 84870 -1360 84890 -1300
rect 84790 -1380 84890 -1360
rect 84960 -1000 85060 -980
rect 84960 -1060 84980 -1000
rect 85040 -1060 85060 -1000
rect 84960 -1100 85060 -1060
rect 84960 -1160 84980 -1100
rect 85040 -1160 85060 -1100
rect 84960 -1200 85060 -1160
rect 84960 -1260 84980 -1200
rect 85040 -1260 85060 -1200
rect 84960 -1300 85060 -1260
rect 84960 -1360 84980 -1300
rect 85040 -1360 85060 -1300
rect 84960 -1380 85060 -1360
rect 85130 -1000 85230 -980
rect 85130 -1060 85150 -1000
rect 85210 -1060 85230 -1000
rect 85130 -1100 85230 -1060
rect 85130 -1160 85150 -1100
rect 85210 -1160 85230 -1100
rect 85130 -1200 85230 -1160
rect 85130 -1260 85150 -1200
rect 85210 -1260 85230 -1200
rect 85130 -1300 85230 -1260
rect 85130 -1360 85150 -1300
rect 85210 -1360 85230 -1300
rect 85130 -1380 85230 -1360
rect 85300 -1000 85400 -980
rect 85300 -1060 85320 -1000
rect 85380 -1060 85400 -1000
rect 85300 -1100 85400 -1060
rect 85300 -1160 85320 -1100
rect 85380 -1160 85400 -1100
rect 85300 -1200 85400 -1160
rect 85300 -1260 85320 -1200
rect 85380 -1260 85400 -1200
rect 85300 -1300 85400 -1260
rect 85300 -1360 85320 -1300
rect 85380 -1360 85400 -1300
rect 85300 -1380 85400 -1360
rect 85470 -1000 85570 -980
rect 85470 -1060 85490 -1000
rect 85550 -1060 85570 -1000
rect 85470 -1100 85570 -1060
rect 85470 -1160 85490 -1100
rect 85550 -1160 85570 -1100
rect 85470 -1200 85570 -1160
rect 85470 -1260 85490 -1200
rect 85550 -1260 85570 -1200
rect 85470 -1300 85570 -1260
rect 85470 -1360 85490 -1300
rect 85550 -1360 85570 -1300
rect 85470 -1380 85570 -1360
rect 85640 -1000 85740 -980
rect 85640 -1060 85660 -1000
rect 85720 -1060 85740 -1000
rect 85640 -1100 85740 -1060
rect 85640 -1160 85660 -1100
rect 85720 -1160 85740 -1100
rect 85640 -1200 85740 -1160
rect 85640 -1260 85660 -1200
rect 85720 -1260 85740 -1200
rect 85640 -1300 85740 -1260
rect 85640 -1360 85660 -1300
rect 85720 -1360 85740 -1300
rect 85640 -1380 85740 -1360
rect 85810 -1000 85910 -980
rect 85810 -1060 85830 -1000
rect 85890 -1060 85910 -1000
rect 85810 -1100 85910 -1060
rect 85810 -1160 85830 -1100
rect 85890 -1160 85910 -1100
rect 85810 -1200 85910 -1160
rect 85810 -1260 85830 -1200
rect 85890 -1260 85910 -1200
rect 85810 -1300 85910 -1260
rect 85810 -1360 85830 -1300
rect 85890 -1360 85910 -1300
rect 85810 -1380 85910 -1360
rect 85980 -1000 86080 -980
rect 85980 -1060 86000 -1000
rect 86060 -1060 86080 -1000
rect 85980 -1100 86080 -1060
rect 85980 -1160 86000 -1100
rect 86060 -1160 86080 -1100
rect 85980 -1200 86080 -1160
rect 85980 -1260 86000 -1200
rect 86060 -1260 86080 -1200
rect 85980 -1300 86080 -1260
rect 85980 -1360 86000 -1300
rect 86060 -1360 86080 -1300
rect 85980 -1380 86080 -1360
rect 86150 -1000 86250 -980
rect 86150 -1060 86170 -1000
rect 86230 -1060 86250 -1000
rect 86150 -1100 86250 -1060
rect 86150 -1160 86170 -1100
rect 86230 -1160 86250 -1100
rect 86150 -1200 86250 -1160
rect 86150 -1260 86170 -1200
rect 86230 -1260 86250 -1200
rect 86150 -1300 86250 -1260
rect 86150 -1360 86170 -1300
rect 86230 -1360 86250 -1300
rect 86150 -1380 86250 -1360
rect 86320 -1000 86420 -980
rect 86320 -1060 86340 -1000
rect 86400 -1060 86420 -1000
rect 86320 -1100 86420 -1060
rect 86320 -1160 86340 -1100
rect 86400 -1160 86420 -1100
rect 86320 -1200 86420 -1160
rect 86320 -1260 86340 -1200
rect 86400 -1260 86420 -1200
rect 86320 -1300 86420 -1260
rect 86320 -1360 86340 -1300
rect 86400 -1360 86420 -1300
rect 86320 -1380 86420 -1360
rect 86490 -1000 86590 -980
rect 86490 -1060 86510 -1000
rect 86570 -1060 86590 -1000
rect 86490 -1100 86590 -1060
rect 86490 -1160 86510 -1100
rect 86570 -1160 86590 -1100
rect 86490 -1200 86590 -1160
rect 86490 -1260 86510 -1200
rect 86570 -1260 86590 -1200
rect 86490 -1300 86590 -1260
rect 86490 -1360 86510 -1300
rect 86570 -1360 86590 -1300
rect 86490 -1380 86590 -1360
rect 86660 -1000 86760 -980
rect 86660 -1060 86680 -1000
rect 86740 -1060 86760 -1000
rect 86660 -1100 86760 -1060
rect 86660 -1160 86680 -1100
rect 86740 -1160 86760 -1100
rect 86660 -1200 86760 -1160
rect 86660 -1260 86680 -1200
rect 86740 -1260 86760 -1200
rect 86660 -1300 86760 -1260
rect 86660 -1360 86680 -1300
rect 86740 -1360 86760 -1300
rect 86660 -1380 86760 -1360
rect 86830 -1000 86930 -980
rect 86830 -1060 86850 -1000
rect 86910 -1060 86930 -1000
rect 86830 -1100 86930 -1060
rect 86830 -1160 86850 -1100
rect 86910 -1160 86930 -1100
rect 86830 -1200 86930 -1160
rect 86830 -1260 86850 -1200
rect 86910 -1260 86930 -1200
rect 86830 -1300 86930 -1260
rect 86830 -1360 86850 -1300
rect 86910 -1360 86930 -1300
rect 86830 -1380 86930 -1360
rect 87000 -1000 87100 -980
rect 87000 -1060 87020 -1000
rect 87080 -1060 87100 -1000
rect 87000 -1100 87100 -1060
rect 87000 -1160 87020 -1100
rect 87080 -1160 87100 -1100
rect 87000 -1200 87100 -1160
rect 87000 -1260 87020 -1200
rect 87080 -1260 87100 -1200
rect 87000 -1300 87100 -1260
rect 87000 -1360 87020 -1300
rect 87080 -1360 87100 -1300
rect 87000 -1380 87100 -1360
rect 87170 -1000 87270 -980
rect 87170 -1060 87190 -1000
rect 87250 -1060 87270 -1000
rect 87170 -1100 87270 -1060
rect 87170 -1160 87190 -1100
rect 87250 -1160 87270 -1100
rect 87170 -1200 87270 -1160
rect 87170 -1260 87190 -1200
rect 87250 -1260 87270 -1200
rect 87170 -1300 87270 -1260
rect 87170 -1360 87190 -1300
rect 87250 -1360 87270 -1300
rect 87170 -1380 87270 -1360
rect 770 -1470 970 -1440
rect 770 -1540 830 -1470
rect 910 -1540 970 -1470
rect 770 -1570 970 -1540
rect 4940 -1470 5140 -1440
rect 4940 -1540 5000 -1470
rect 5080 -1540 5140 -1470
rect 4940 -1570 5140 -1540
rect 8970 -1470 9170 -1440
rect 8970 -1540 9030 -1470
rect 9110 -1540 9170 -1470
rect 8970 -1570 9170 -1540
rect 13000 -1470 13200 -1440
rect 13000 -1540 13060 -1470
rect 13140 -1540 13200 -1470
rect 13000 -1570 13200 -1540
rect 17040 -1470 17240 -1440
rect 17040 -1540 17100 -1470
rect 17180 -1540 17240 -1470
rect 17040 -1570 17240 -1540
rect 21140 -1470 21340 -1440
rect 21140 -1540 21200 -1470
rect 21280 -1540 21340 -1470
rect 21140 -1570 21340 -1540
rect 25250 -1470 25450 -1440
rect 25250 -1540 25310 -1470
rect 25390 -1540 25450 -1470
rect 25250 -1570 25450 -1540
rect 29350 -1470 29550 -1440
rect 29350 -1540 29410 -1470
rect 29490 -1540 29550 -1470
rect 29350 -1570 29550 -1540
rect 33380 -1470 33580 -1440
rect 33380 -1540 33440 -1470
rect 33520 -1540 33580 -1470
rect 33380 -1570 33580 -1540
rect 37490 -1470 37690 -1440
rect 37490 -1540 37550 -1470
rect 37630 -1540 37690 -1470
rect 37490 -1570 37690 -1540
rect 41590 -1470 41790 -1440
rect 41590 -1540 41650 -1470
rect 41730 -1540 41790 -1470
rect 41590 -1570 41790 -1540
rect 47040 -1470 47240 -1440
rect 47040 -1540 47100 -1470
rect 47180 -1540 47240 -1470
rect 47040 -1570 47240 -1540
rect 51120 -1470 51320 -1440
rect 51120 -1540 51180 -1470
rect 51260 -1540 51320 -1470
rect 51120 -1570 51320 -1540
rect 55230 -1470 55430 -1440
rect 55230 -1540 55290 -1470
rect 55370 -1540 55430 -1470
rect 55230 -1570 55430 -1540
rect 59260 -1470 59460 -1440
rect 59260 -1540 59320 -1470
rect 59400 -1540 59460 -1470
rect 59260 -1570 59460 -1540
rect 63360 -1470 63560 -1440
rect 63360 -1540 63420 -1470
rect 63500 -1540 63560 -1470
rect 63360 -1570 63560 -1540
rect 67470 -1470 67670 -1440
rect 67470 -1540 67530 -1470
rect 67610 -1540 67670 -1470
rect 67470 -1570 67670 -1540
rect 71500 -1470 71700 -1440
rect 71500 -1540 71560 -1470
rect 71640 -1540 71700 -1470
rect 71500 -1570 71700 -1540
rect 75750 -1470 75950 -1440
rect 75750 -1540 75810 -1470
rect 75890 -1540 75950 -1470
rect 75750 -1570 75950 -1540
rect 79710 -1470 79910 -1440
rect 79710 -1540 79770 -1470
rect 79850 -1540 79910 -1470
rect 79710 -1570 79910 -1540
rect 83890 -1470 84090 -1440
rect 83890 -1540 83950 -1470
rect 84030 -1540 84090 -1470
rect 83890 -1570 84090 -1540
rect 86450 -1474 86648 -1444
rect 86450 -1544 86508 -1474
rect 86588 -1544 86648 -1474
rect 86450 -1572 86648 -1544
<< viali >>
rect 543 935 577 995
rect 577 935 617 995
rect 1271 935 1311 995
rect 1311 935 1345 995
rect 5663 913 5697 973
rect 5697 913 5737 973
rect 6391 913 6431 973
rect 6431 913 6465 973
rect 520 630 610 690
rect 5630 630 5720 690
rect 790 520 870 590
rect 2170 520 2250 590
rect 3550 520 3630 590
rect 5210 520 5290 590
rect 8040 520 8120 590
rect 10800 520 10880 590
rect 13430 520 13510 590
rect 16470 520 16550 590
rect 20540 520 20620 590
rect 24680 520 24760 590
rect 28760 520 28840 590
rect 32910 520 32990 590
rect 36780 520 36860 590
rect 40920 520 41000 590
rect 44910 520 44990 590
rect 48990 520 49070 590
rect 53080 520 53160 590
rect 57240 520 57320 590
rect 30 350 90 410
rect 200 350 260 410
rect 200 250 260 310
rect 450 350 510 410
rect 620 250 680 310
rect 790 350 850 410
rect 960 250 1020 310
rect 1130 350 1190 410
rect 1520 350 1580 410
rect 1690 250 1750 310
rect 1860 350 1920 410
rect 2030 250 2090 310
rect 2200 350 2260 410
rect 2370 250 2430 310
rect 2540 350 2600 410
rect 2710 250 2770 310
rect 2880 350 2940 410
rect 3050 250 3110 310
rect 3220 350 3280 410
rect 3390 250 3450 310
rect 3560 350 3620 410
rect 3730 250 3790 310
rect 3900 350 3960 410
rect 4070 250 4130 310
rect 4240 350 4300 410
rect 4540 350 4600 410
rect 4710 250 4770 310
rect 4880 350 4940 410
rect 5050 250 5110 310
rect 5220 350 5280 410
rect 5390 250 5450 310
rect 5560 350 5620 410
rect 5730 250 5790 310
rect 5900 350 5960 410
rect 6070 250 6130 310
rect 6240 350 6300 410
rect 6410 250 6470 310
rect 6580 350 6640 410
rect 6750 250 6810 310
rect 6920 350 6980 410
rect 7090 250 7150 310
rect 7260 350 7320 410
rect 7430 250 7490 310
rect 7600 350 7660 410
rect 7770 250 7830 310
rect 7940 350 8000 410
rect 8110 250 8170 310
rect 8280 350 8340 410
rect 8450 250 8510 310
rect 8620 350 8680 410
rect 8790 250 8850 310
rect 8960 350 9020 410
rect 9130 250 9190 310
rect 9300 350 9360 410
rect 9470 250 9530 310
rect 9640 350 9700 410
rect 9810 250 9870 310
rect 9980 350 10040 410
rect 10150 250 10210 310
rect 10320 350 10380 410
rect 10490 250 10550 310
rect 10660 350 10720 410
rect 10830 250 10890 310
rect 11000 350 11060 410
rect 11170 250 11230 310
rect 11340 350 11400 410
rect 11510 250 11570 310
rect 11680 350 11740 410
rect 11850 250 11910 310
rect 12020 350 12080 410
rect 12190 250 12250 310
rect 12360 350 12420 410
rect 12530 250 12590 310
rect 12700 350 12760 410
rect 12870 250 12930 310
rect 13040 350 13100 410
rect 13210 250 13270 310
rect 13380 350 13440 410
rect 13550 250 13610 310
rect 13720 350 13780 410
rect 13890 250 13950 310
rect 14060 350 14120 410
rect 14230 250 14290 310
rect 14400 350 14460 410
rect 14570 250 14630 310
rect 14740 350 14800 410
rect 14910 250 14970 310
rect 15080 350 15140 410
rect 15250 250 15310 310
rect 15420 350 15480 410
rect 15720 350 15780 410
rect 15890 250 15950 310
rect 16060 350 16120 410
rect 16230 250 16290 310
rect 16400 350 16460 410
rect 16570 250 16630 310
rect 16740 350 16800 410
rect 16910 250 16970 310
rect 17080 350 17140 410
rect 17250 250 17310 310
rect 17420 350 17480 410
rect 17590 250 17650 310
rect 17760 350 17820 410
rect 17930 250 17990 310
rect 18100 350 18160 410
rect 18270 250 18330 310
rect 18440 350 18500 410
rect 18610 250 18670 310
rect 18780 350 18840 410
rect 18950 250 19010 310
rect 19120 350 19180 410
rect 19290 250 19350 310
rect 19460 350 19520 410
rect 19630 250 19690 310
rect 19800 350 19860 410
rect 19970 250 20030 310
rect 20140 350 20200 410
rect 20310 250 20370 310
rect 20480 350 20540 410
rect 20650 250 20710 310
rect 20820 350 20880 410
rect 20990 250 21050 310
rect 21160 350 21220 410
rect 21330 250 21390 310
rect 21500 350 21560 410
rect 21670 250 21730 310
rect 21840 350 21900 410
rect 22010 250 22070 310
rect 22180 350 22240 410
rect 22350 250 22410 310
rect 22520 350 22580 410
rect 22690 250 22750 310
rect 22860 350 22920 410
rect 23030 250 23090 310
rect 23200 350 23260 410
rect 23370 250 23430 310
rect 23540 350 23600 410
rect 23710 250 23770 310
rect 23880 350 23940 410
rect 24050 250 24110 310
rect 24220 350 24280 410
rect 24390 250 24450 310
rect 24560 350 24620 410
rect 24730 250 24790 310
rect 24900 350 24960 410
rect 25070 250 25130 310
rect 25240 350 25300 410
rect 25410 250 25470 310
rect 25580 350 25640 410
rect 25750 250 25810 310
rect 25920 350 25980 410
rect 26090 250 26150 310
rect 26260 350 26320 410
rect 26430 250 26490 310
rect 26600 350 26660 410
rect 26770 250 26830 310
rect 26940 350 27000 410
rect 27110 250 27170 310
rect 27280 350 27340 410
rect 27450 250 27510 310
rect 27620 350 27680 410
rect 27790 250 27850 310
rect 27960 350 28020 410
rect 28130 250 28190 310
rect 28300 350 28360 410
rect 28470 250 28530 310
rect 28640 350 28700 410
rect 28810 250 28870 310
rect 28980 350 29040 410
rect 29150 250 29210 310
rect 29320 350 29380 410
rect 29490 250 29550 310
rect 29660 350 29720 410
rect 29830 250 29890 310
rect 30000 350 30060 410
rect 30170 250 30230 310
rect 30340 350 30400 410
rect 30510 250 30570 310
rect 30680 350 30740 410
rect 30850 250 30910 310
rect 31020 350 31080 410
rect 31190 250 31250 310
rect 31360 350 31420 410
rect 31530 250 31590 310
rect 31700 350 31760 410
rect 31870 250 31930 310
rect 32040 350 32100 410
rect 32210 250 32270 310
rect 32380 350 32440 410
rect 32550 250 32610 310
rect 32720 350 32780 410
rect 32890 250 32950 310
rect 33060 350 33120 410
rect 33230 250 33290 310
rect 33400 350 33460 410
rect 33570 250 33630 310
rect 33740 350 33800 410
rect 33910 250 33970 310
rect 34080 350 34140 410
rect 34250 250 34310 310
rect 34420 350 34480 410
rect 34590 250 34650 310
rect 34760 350 34820 410
rect 34930 250 34990 310
rect 35100 350 35160 410
rect 35270 250 35330 310
rect 35440 350 35500 410
rect 35610 250 35670 310
rect 35780 350 35840 410
rect 35950 250 36010 310
rect 36120 350 36180 410
rect 36290 250 36350 310
rect 36460 350 36520 410
rect 36630 250 36690 310
rect 36800 350 36860 410
rect 36970 250 37030 310
rect 37140 350 37200 410
rect 37310 250 37370 310
rect 37480 350 37540 410
rect 37650 250 37710 310
rect 37820 350 37880 410
rect 37990 250 38050 310
rect 38160 350 38220 410
rect 38330 250 38390 310
rect 38500 350 38560 410
rect 38670 250 38730 310
rect 38840 350 38900 410
rect 39010 250 39070 310
rect 39180 350 39240 410
rect 39350 250 39410 310
rect 39520 350 39580 410
rect 39690 250 39750 310
rect 39860 350 39920 410
rect 40030 250 40090 310
rect 40200 350 40260 410
rect 40370 250 40430 310
rect 40540 350 40600 410
rect 40710 250 40770 310
rect 40880 350 40940 410
rect 41050 250 41110 310
rect 41220 350 41280 410
rect 41390 250 41450 310
rect 41560 350 41620 410
rect 41730 250 41790 310
rect 41900 350 41960 410
rect 42070 250 42130 310
rect 42240 350 42300 410
rect 42410 250 42470 310
rect 42580 350 42640 410
rect 42750 250 42810 310
rect 42920 350 42980 410
rect 43090 250 43150 310
rect 43260 350 43320 410
rect 43430 250 43490 310
rect 43600 350 43660 410
rect 43770 250 43830 310
rect 43940 350 44000 410
rect 44110 250 44170 310
rect 44280 350 44340 410
rect 44450 250 44510 310
rect 44620 350 44680 410
rect 44790 250 44850 310
rect 44960 350 45020 410
rect 45130 250 45190 310
rect 45300 350 45360 410
rect 45470 250 45530 310
rect 45640 350 45700 410
rect 45810 250 45870 310
rect 45980 350 46040 410
rect 46150 250 46210 310
rect 46320 350 46380 410
rect 46490 250 46550 310
rect 46660 350 46720 410
rect 46830 250 46890 310
rect 47000 350 47060 410
rect 47170 250 47230 310
rect 47340 350 47400 410
rect 47510 250 47570 310
rect 47680 350 47740 410
rect 47850 250 47910 310
rect 48020 350 48080 410
rect 48190 250 48250 310
rect 48360 350 48420 410
rect 48530 250 48590 310
rect 48700 350 48760 410
rect 48870 250 48930 310
rect 49040 350 49100 410
rect 49210 250 49270 310
rect 49380 350 49440 410
rect 49550 250 49610 310
rect 49720 350 49780 410
rect 49890 250 49950 310
rect 50060 350 50120 410
rect 50230 250 50290 310
rect 50400 350 50460 410
rect 50570 250 50630 310
rect 50740 350 50800 410
rect 50910 250 50970 310
rect 51080 350 51140 410
rect 51250 250 51310 310
rect 51420 350 51480 410
rect 51590 250 51650 310
rect 51760 350 51820 410
rect 51930 250 51990 310
rect 52100 350 52160 410
rect 52270 250 52330 310
rect 52440 350 52500 410
rect 52610 250 52670 310
rect 52780 350 52840 410
rect 52950 250 53010 310
rect 53120 350 53180 410
rect 53290 250 53350 310
rect 53460 350 53520 410
rect 53630 250 53690 310
rect 53800 350 53860 410
rect 53970 250 54030 310
rect 54140 350 54200 410
rect 54310 250 54370 310
rect 54480 350 54540 410
rect 54650 250 54710 310
rect 54820 350 54880 410
rect 54990 250 55050 310
rect 55160 350 55220 410
rect 55330 250 55390 310
rect 55500 350 55560 410
rect 55670 250 55730 310
rect 55840 350 55900 410
rect 56010 250 56070 310
rect 56180 350 56240 410
rect 56350 250 56410 310
rect 56520 350 56580 410
rect 56690 250 56750 310
rect 56860 350 56920 410
rect 57030 250 57090 310
rect 57200 350 57260 410
rect 57370 250 57430 310
rect 57540 350 57600 410
rect 57710 250 57770 310
rect 57880 350 57940 410
rect 58050 250 58110 310
rect 58220 350 58280 410
rect 58390 250 58450 310
rect 58560 350 58620 410
rect 58730 250 58790 310
rect 58900 350 58960 410
rect 59070 250 59130 310
rect 59240 350 59300 410
rect 70 30 130 110
rect 450 20 510 80
rect 620 20 680 80
rect 790 20 850 80
rect 960 20 1020 80
rect 1130 20 1190 80
rect 1520 20 1580 80
rect 1690 20 1750 80
rect 1860 20 1920 80
rect 2030 20 2090 80
rect 2200 20 2260 80
rect 2370 20 2430 80
rect 2540 20 2600 80
rect 2710 20 2770 80
rect 2880 20 2940 80
rect 3050 20 3110 80
rect 3220 20 3280 80
rect 3390 20 3450 80
rect 3560 20 3620 80
rect 3730 20 3790 80
rect 3900 20 3960 80
rect 4070 20 4130 80
rect 4240 20 4300 80
rect 4540 20 4600 80
rect 4710 20 4770 80
rect 4880 20 4940 80
rect 5050 20 5110 80
rect 5220 20 5280 80
rect 5390 20 5450 80
rect 5560 20 5620 80
rect 5730 20 5790 80
rect 5900 20 5960 80
rect 6070 20 6130 80
rect 6240 20 6300 80
rect 6410 20 6470 80
rect 6580 20 6640 80
rect 6750 20 6810 80
rect 6920 20 6980 80
rect 7090 20 7150 80
rect 7260 20 7320 80
rect 7430 20 7490 80
rect 7600 20 7660 80
rect 7770 20 7830 80
rect 7940 20 8000 80
rect 8110 20 8170 80
rect 8280 20 8340 80
rect 8450 20 8510 80
rect 8620 20 8680 80
rect 8790 20 8850 80
rect 8960 20 9020 80
rect 9130 20 9190 80
rect 9300 20 9360 80
rect 9470 20 9530 80
rect 9640 20 9700 80
rect 9810 20 9870 80
rect 9980 20 10040 80
rect 10150 20 10210 80
rect 10320 20 10380 80
rect 10490 20 10550 80
rect 10660 20 10720 80
rect 10830 20 10890 80
rect 11000 20 11060 80
rect 11170 20 11230 80
rect 11340 20 11400 80
rect 11510 20 11570 80
rect 11680 20 11740 80
rect 11850 20 11910 80
rect 12020 20 12080 80
rect 12190 20 12250 80
rect 12360 20 12420 80
rect 12530 20 12590 80
rect 12700 20 12760 80
rect 12870 20 12930 80
rect 13040 20 13100 80
rect 13210 20 13270 80
rect 13380 20 13440 80
rect 13550 20 13610 80
rect 13720 20 13780 80
rect 13890 20 13950 80
rect 14060 20 14120 80
rect 14230 20 14290 80
rect 14400 20 14460 80
rect 14570 20 14630 80
rect 14740 20 14800 80
rect 14910 20 14970 80
rect 15080 20 15140 80
rect 15250 20 15310 80
rect 15420 20 15480 80
rect 15720 20 15780 80
rect 15890 20 15950 80
rect 16060 20 16120 80
rect 16230 20 16290 80
rect 16400 20 16460 80
rect 16570 20 16630 80
rect 16740 20 16800 80
rect 16910 20 16970 80
rect 17080 20 17140 80
rect 17250 20 17310 80
rect 17420 20 17480 80
rect 17590 20 17650 80
rect 17760 20 17820 80
rect 17930 20 17990 80
rect 18100 20 18160 80
rect 18270 20 18330 80
rect 18440 20 18500 80
rect 18610 20 18670 80
rect 18780 20 18840 80
rect 18950 20 19010 80
rect 19120 20 19180 80
rect 19290 20 19350 80
rect 19460 20 19520 80
rect 19630 20 19690 80
rect 19800 20 19860 80
rect 19970 20 20030 80
rect 20140 20 20200 80
rect 20310 20 20370 80
rect 20480 20 20540 80
rect 20650 20 20710 80
rect 20820 20 20880 80
rect 20990 20 21050 80
rect 21160 20 21220 80
rect 21330 20 21390 80
rect 21500 20 21560 80
rect 21670 20 21730 80
rect 21840 20 21900 80
rect 22010 20 22070 80
rect 22180 20 22240 80
rect 22350 20 22410 80
rect 22520 20 22580 80
rect 22690 20 22750 80
rect 22860 20 22920 80
rect 23030 20 23090 80
rect 23200 20 23260 80
rect 23370 20 23430 80
rect 23540 20 23600 80
rect 23710 20 23770 80
rect 23880 20 23940 80
rect 24050 20 24110 80
rect 24220 20 24280 80
rect 24390 20 24450 80
rect 24560 20 24620 80
rect 24730 20 24790 80
rect 24900 20 24960 80
rect 25070 20 25130 80
rect 25240 20 25300 80
rect 25410 20 25470 80
rect 25580 20 25640 80
rect 25750 20 25810 80
rect 25920 20 25980 80
rect 26090 20 26150 80
rect 26260 20 26320 80
rect 26430 20 26490 80
rect 26600 20 26660 80
rect 26770 20 26830 80
rect 26940 20 27000 80
rect 27110 20 27170 80
rect 27280 20 27340 80
rect 27450 20 27510 80
rect 27620 20 27680 80
rect 27790 20 27850 80
rect 27960 20 28020 80
rect 28130 20 28190 80
rect 28300 20 28360 80
rect 28470 20 28530 80
rect 28640 20 28700 80
rect 28810 20 28870 80
rect 28980 20 29040 80
rect 29150 20 29210 80
rect 29320 20 29380 80
rect 29490 20 29550 80
rect 29660 20 29720 80
rect 29830 20 29890 80
rect 30000 20 30060 80
rect 30170 20 30230 80
rect 30340 20 30400 80
rect 30510 20 30570 80
rect 30680 20 30740 80
rect 30850 20 30910 80
rect 31020 20 31080 80
rect 31190 20 31250 80
rect 31360 20 31420 80
rect 31530 20 31590 80
rect 31700 20 31760 80
rect 31870 20 31930 80
rect 32040 20 32100 80
rect 32210 20 32270 80
rect 32380 20 32440 80
rect 32550 20 32610 80
rect 32720 20 32780 80
rect 32890 20 32950 80
rect 33060 20 33120 80
rect 33230 20 33290 80
rect 33400 20 33460 80
rect 33570 20 33630 80
rect 33740 20 33800 80
rect 33910 20 33970 80
rect 34080 20 34140 80
rect 34250 20 34310 80
rect 34420 20 34480 80
rect 34590 20 34650 80
rect 34760 20 34820 80
rect 34930 20 34990 80
rect 35100 20 35160 80
rect 35270 20 35330 80
rect 35440 20 35500 80
rect 35610 20 35670 80
rect 35780 20 35840 80
rect 35950 20 36010 80
rect 36120 20 36180 80
rect 36290 20 36350 80
rect 36460 20 36520 80
rect 36630 20 36690 80
rect 36800 20 36860 80
rect 36970 20 37030 80
rect 37140 20 37200 80
rect 37310 20 37370 80
rect 37480 20 37540 80
rect 37650 20 37710 80
rect 37820 20 37880 80
rect 37990 20 38050 80
rect 38160 20 38220 80
rect 38330 20 38390 80
rect 38500 20 38560 80
rect 38670 20 38730 80
rect 38840 20 38900 80
rect 39010 20 39070 80
rect 39180 20 39240 80
rect 39350 20 39410 80
rect 39520 20 39580 80
rect 39690 20 39750 80
rect 39860 20 39920 80
rect 40030 20 40090 80
rect 40200 20 40260 80
rect 40370 20 40430 80
rect 40540 20 40600 80
rect 40710 20 40770 80
rect 40880 20 40940 80
rect 41050 20 41110 80
rect 41220 20 41280 80
rect 41390 20 41450 80
rect 41560 20 41620 80
rect 41730 20 41790 80
rect 41900 20 41960 80
rect 42070 20 42130 80
rect 42240 20 42300 80
rect 42410 20 42470 80
rect 42580 20 42640 80
rect 42750 20 42810 80
rect 42920 20 42980 80
rect 43090 20 43150 80
rect 43260 20 43320 80
rect 43430 20 43490 80
rect 43600 20 43660 80
rect 43770 20 43830 80
rect 43940 20 44000 80
rect 44110 20 44170 80
rect 44280 20 44340 80
rect 44450 20 44510 80
rect 44620 20 44680 80
rect 44790 20 44850 80
rect 44960 20 45020 80
rect 45130 20 45190 80
rect 45300 20 45360 80
rect 45470 20 45530 80
rect 45640 20 45700 80
rect 45810 20 45870 80
rect 45980 20 46040 80
rect 46150 20 46210 80
rect 46320 20 46380 80
rect 46490 20 46550 80
rect 46660 20 46720 80
rect 46830 20 46890 80
rect 47000 20 47060 80
rect 47170 20 47230 80
rect 47340 20 47400 80
rect 47510 20 47570 80
rect 47680 20 47740 80
rect 47850 20 47910 80
rect 48020 20 48080 80
rect 48190 20 48250 80
rect 48360 20 48420 80
rect 48530 20 48590 80
rect 48700 20 48760 80
rect 48870 20 48930 80
rect 49040 20 49100 80
rect 49210 20 49270 80
rect 49380 20 49440 80
rect 49550 20 49610 80
rect 49720 20 49780 80
rect 49890 20 49950 80
rect 50060 20 50120 80
rect 50230 20 50290 80
rect 50400 20 50460 80
rect 50570 20 50630 80
rect 50740 20 50800 80
rect 50910 20 50970 80
rect 51080 20 51140 80
rect 51250 20 51310 80
rect 51420 20 51480 80
rect 51590 20 51650 80
rect 51760 20 51820 80
rect 51930 20 51990 80
rect 52100 20 52160 80
rect 52270 20 52330 80
rect 52440 20 52500 80
rect 52610 20 52670 80
rect 52780 20 52840 80
rect 52950 20 53010 80
rect 53120 20 53180 80
rect 53290 20 53350 80
rect 53460 20 53520 80
rect 53630 20 53690 80
rect 53800 20 53860 80
rect 53970 20 54030 80
rect 54140 20 54200 80
rect 54310 20 54370 80
rect 54480 20 54540 80
rect 54650 20 54710 80
rect 54820 20 54880 80
rect 54990 20 55050 80
rect 55160 20 55220 80
rect 55330 20 55390 80
rect 55500 20 55560 80
rect 55670 20 55730 80
rect 55840 20 55900 80
rect 56010 20 56070 80
rect 56180 20 56240 80
rect 56350 20 56410 80
rect 56520 20 56580 80
rect 56690 20 56750 80
rect 56860 20 56920 80
rect 57030 20 57090 80
rect 57200 20 57260 80
rect 57370 20 57430 80
rect 57540 20 57600 80
rect 57710 20 57770 80
rect 57880 20 57940 80
rect 58050 20 58110 80
rect 58220 20 58280 80
rect 58390 20 58450 80
rect 58560 20 58620 80
rect 58730 20 58790 80
rect 58900 20 58960 80
rect 59070 20 59130 80
rect 59240 20 59300 80
rect 30 -120 90 -60
rect 200 -120 260 -60
rect 530 -120 600 -60
rect 700 -120 770 -60
rect 870 -120 940 -60
rect 1040 -120 1110 -60
rect 1600 -120 1670 -60
rect 1770 -120 1840 -60
rect 1940 -120 2010 -60
rect 2110 -120 2180 -60
rect 2280 -120 2350 -60
rect 2450 -120 2520 -60
rect 2620 -120 2690 -60
rect 2790 -120 2860 -60
rect 2960 -120 3030 -60
rect 3130 -120 3200 -60
rect 3300 -120 3370 -60
rect 3470 -120 3540 -60
rect 3640 -120 3710 -60
rect 3810 -120 3880 -60
rect 3980 -120 4050 -60
rect 4150 -120 4220 -60
rect 4620 -120 4690 -60
rect 4790 -120 4860 -60
rect 4960 -120 5030 -60
rect 5130 -120 5200 -60
rect 5300 -120 5370 -60
rect 5470 -120 5540 -60
rect 5640 -120 5710 -60
rect 5810 -120 5880 -60
rect 5980 -120 6050 -60
rect 6150 -120 6220 -60
rect 6320 -120 6390 -60
rect 6490 -120 6560 -60
rect 6660 -120 6730 -60
rect 6830 -120 6900 -60
rect 7000 -120 7070 -60
rect 7170 -120 7240 -60
rect 7340 -120 7410 -60
rect 7510 -120 7580 -60
rect 7680 -120 7750 -60
rect 7850 -120 7920 -60
rect 8020 -120 8090 -60
rect 8190 -120 8260 -60
rect 8360 -120 8430 -60
rect 8530 -120 8600 -60
rect 8700 -120 8770 -60
rect 8870 -120 8940 -60
rect 9040 -120 9110 -60
rect 9210 -120 9280 -60
rect 9380 -120 9450 -60
rect 9550 -120 9620 -60
rect 9720 -120 9790 -60
rect 9890 -120 9960 -60
rect 10060 -120 10130 -60
rect 10230 -120 10300 -60
rect 10400 -120 10470 -60
rect 10570 -120 10640 -60
rect 10740 -120 10810 -60
rect 10910 -120 10980 -60
rect 11080 -120 11150 -60
rect 11250 -120 11320 -60
rect 11420 -120 11490 -60
rect 11590 -120 11660 -60
rect 11760 -120 11830 -60
rect 11930 -120 12000 -60
rect 12100 -120 12170 -60
rect 12270 -120 12340 -60
rect 12440 -120 12510 -60
rect 12610 -120 12680 -60
rect 12780 -120 12850 -60
rect 12950 -120 13020 -60
rect 13120 -120 13190 -60
rect 13290 -120 13360 -60
rect 13460 -120 13530 -60
rect 13630 -120 13700 -60
rect 13800 -120 13870 -60
rect 13970 -120 14040 -60
rect 14140 -120 14210 -60
rect 14310 -120 14380 -60
rect 14480 -120 14550 -60
rect 14650 -120 14720 -60
rect 14820 -120 14890 -60
rect 14990 -120 15060 -60
rect 15160 -120 15230 -60
rect 15330 -120 15400 -60
rect 15800 -120 15870 -60
rect 15970 -120 16040 -60
rect 16140 -120 16210 -60
rect 16310 -120 16380 -60
rect 16480 -120 16550 -60
rect 16650 -120 16720 -60
rect 16820 -120 16890 -60
rect 16990 -120 17060 -60
rect 17160 -120 17230 -60
rect 17330 -120 17400 -60
rect 17500 -120 17570 -60
rect 17670 -120 17740 -60
rect 17840 -120 17910 -60
rect 18010 -120 18080 -60
rect 18180 -120 18250 -60
rect 18350 -120 18420 -60
rect 18520 -120 18590 -60
rect 18690 -120 18760 -60
rect 18860 -120 18930 -60
rect 19030 -120 19100 -60
rect 19200 -120 19270 -60
rect 19370 -120 19440 -60
rect 19540 -120 19610 -60
rect 19710 -120 19780 -60
rect 19880 -120 19950 -60
rect 20050 -120 20120 -60
rect 20220 -120 20290 -60
rect 20390 -120 20460 -60
rect 20560 -120 20630 -60
rect 20730 -120 20800 -60
rect 20900 -120 20970 -60
rect 21070 -120 21140 -60
rect 21240 -120 21310 -60
rect 21410 -120 21480 -60
rect 21580 -120 21650 -60
rect 21750 -120 21820 -60
rect 21920 -120 21990 -60
rect 22090 -120 22160 -60
rect 22260 -120 22330 -60
rect 22430 -120 22500 -60
rect 22600 -120 22670 -60
rect 22770 -120 22840 -60
rect 22940 -120 23010 -60
rect 23110 -120 23180 -60
rect 23280 -120 23350 -60
rect 23450 -120 23520 -60
rect 23620 -120 23690 -60
rect 23790 -120 23860 -60
rect 23960 -120 24030 -60
rect 24130 -120 24200 -60
rect 24300 -120 24370 -60
rect 24470 -120 24540 -60
rect 24640 -120 24710 -60
rect 24810 -120 24880 -60
rect 24980 -120 25050 -60
rect 25150 -120 25220 -60
rect 25320 -120 25390 -60
rect 25490 -120 25560 -60
rect 25660 -120 25730 -60
rect 25830 -120 25900 -60
rect 26000 -120 26070 -60
rect 26170 -120 26240 -60
rect 26340 -120 26410 -60
rect 26510 -120 26580 -60
rect 26680 -120 26750 -60
rect 26850 -120 26920 -60
rect 27020 -120 27090 -60
rect 27190 -120 27260 -60
rect 27360 -120 27430 -60
rect 27530 -120 27600 -60
rect 27700 -120 27770 -60
rect 27870 -120 27940 -60
rect 28040 -120 28110 -60
rect 28210 -120 28280 -60
rect 28380 -120 28450 -60
rect 28550 -120 28620 -60
rect 28720 -120 28790 -60
rect 28890 -120 28960 -60
rect 29060 -120 29130 -60
rect 29230 -120 29300 -60
rect 29400 -120 29470 -60
rect 29570 -120 29640 -60
rect 29740 -120 29810 -60
rect 29910 -120 29980 -60
rect 30080 -120 30150 -60
rect 30250 -120 30320 -60
rect 30420 -120 30490 -60
rect 30590 -120 30660 -60
rect 30760 -120 30830 -60
rect 30930 -120 31000 -60
rect 31100 -120 31170 -60
rect 31270 -120 31340 -60
rect 31440 -120 31510 -60
rect 31610 -120 31680 -60
rect 31780 -120 31850 -60
rect 31950 -120 32020 -60
rect 32120 -120 32190 -60
rect 32290 -120 32360 -60
rect 32460 -120 32530 -60
rect 32630 -120 32700 -60
rect 32800 -120 32870 -60
rect 32970 -120 33040 -60
rect 33140 -120 33210 -60
rect 33310 -120 33380 -60
rect 33480 -120 33550 -60
rect 33650 -120 33720 -60
rect 33820 -120 33890 -60
rect 33990 -120 34060 -60
rect 34160 -120 34230 -60
rect 34330 -120 34400 -60
rect 34500 -120 34570 -60
rect 34670 -120 34740 -60
rect 34840 -120 34910 -60
rect 35010 -120 35080 -60
rect 35180 -120 35250 -60
rect 35350 -120 35420 -60
rect 35520 -120 35590 -60
rect 35690 -120 35760 -60
rect 35860 -120 35930 -60
rect 36030 -120 36100 -60
rect 36200 -120 36270 -60
rect 36370 -120 36440 -60
rect 36540 -120 36610 -60
rect 36710 -120 36780 -60
rect 36880 -120 36950 -60
rect 37050 -120 37120 -60
rect 37220 -120 37290 -60
rect 37390 -120 37460 -60
rect 37560 -120 37630 -60
rect 37730 -120 37800 -60
rect 37900 -120 37970 -60
rect 38070 -120 38140 -60
rect 38240 -120 38310 -60
rect 38410 -120 38480 -60
rect 38580 -120 38650 -60
rect 38750 -120 38820 -60
rect 38920 -120 38990 -60
rect 39090 -120 39160 -60
rect 39260 -120 39330 -60
rect 39430 -120 39500 -60
rect 39600 -120 39670 -60
rect 39770 -120 39840 -60
rect 39940 -120 40010 -60
rect 40110 -120 40180 -60
rect 40280 -120 40350 -60
rect 40450 -120 40520 -60
rect 40620 -120 40690 -60
rect 40790 -120 40860 -60
rect 40960 -120 41030 -60
rect 41130 -120 41200 -60
rect 41300 -120 41370 -60
rect 41470 -120 41540 -60
rect 41640 -120 41710 -60
rect 41810 -120 41880 -60
rect 41980 -120 42050 -60
rect 42150 -120 42220 -60
rect 42320 -120 42390 -60
rect 42490 -120 42560 -60
rect 42660 -120 42730 -60
rect 42830 -120 42900 -60
rect 43000 -120 43070 -60
rect 43170 -120 43240 -60
rect 43340 -120 43410 -60
rect 43510 -120 43580 -60
rect 43680 -120 43750 -60
rect 43850 -120 43920 -60
rect 44020 -120 44090 -60
rect 44190 -120 44260 -60
rect 44360 -120 44430 -60
rect 44530 -120 44600 -60
rect 44700 -120 44770 -60
rect 44870 -120 44940 -60
rect 45040 -120 45110 -60
rect 45210 -120 45280 -60
rect 45380 -120 45450 -60
rect 45550 -120 45620 -60
rect 45720 -120 45790 -60
rect 45890 -120 45960 -60
rect 46060 -120 46130 -60
rect 46230 -120 46300 -60
rect 46400 -120 46470 -60
rect 46570 -120 46640 -60
rect 46740 -120 46810 -60
rect 46910 -120 46980 -60
rect 47080 -120 47150 -60
rect 47250 -120 47320 -60
rect 47420 -120 47490 -60
rect 47590 -120 47660 -60
rect 47760 -120 47830 -60
rect 47930 -120 48000 -60
rect 48100 -120 48170 -60
rect 48270 -120 48340 -60
rect 48440 -120 48510 -60
rect 48610 -120 48680 -60
rect 48780 -120 48850 -60
rect 48950 -120 49020 -60
rect 49120 -120 49190 -60
rect 49290 -120 49360 -60
rect 49460 -120 49530 -60
rect 49630 -120 49700 -60
rect 49800 -120 49870 -60
rect 49970 -120 50040 -60
rect 50140 -120 50210 -60
rect 50310 -120 50380 -60
rect 50480 -120 50550 -60
rect 50650 -120 50720 -60
rect 50820 -120 50890 -60
rect 50990 -120 51060 -60
rect 51160 -120 51230 -60
rect 51330 -120 51400 -60
rect 51500 -120 51570 -60
rect 51670 -120 51740 -60
rect 51840 -120 51910 -60
rect 52010 -120 52080 -60
rect 52180 -120 52250 -60
rect 52350 -120 52420 -60
rect 52520 -120 52590 -60
rect 52690 -120 52760 -60
rect 52860 -120 52930 -60
rect 53030 -120 53100 -60
rect 53200 -120 53270 -60
rect 53370 -120 53440 -60
rect 53540 -120 53610 -60
rect 53710 -120 53780 -60
rect 53880 -120 53950 -60
rect 54050 -120 54120 -60
rect 54220 -120 54290 -60
rect 54390 -120 54460 -60
rect 54560 -120 54630 -60
rect 54730 -120 54800 -60
rect 54900 -120 54970 -60
rect 55070 -120 55140 -60
rect 55240 -120 55310 -60
rect 55410 -120 55480 -60
rect 55580 -120 55650 -60
rect 55750 -120 55820 -60
rect 55920 -120 55990 -60
rect 56090 -120 56160 -60
rect 56260 -120 56330 -60
rect 56430 -120 56500 -60
rect 56600 -120 56670 -60
rect 56770 -120 56840 -60
rect 56940 -120 57010 -60
rect 57110 -120 57180 -60
rect 57280 -120 57350 -60
rect 57450 -120 57520 -60
rect 57620 -120 57690 -60
rect 57790 -120 57860 -60
rect 57960 -120 58030 -60
rect 58130 -120 58200 -60
rect 58300 -120 58370 -60
rect 58470 -120 58540 -60
rect 58640 -120 58710 -60
rect 58810 -120 58880 -60
rect 58980 -120 59050 -60
rect 59150 -120 59220 -60
rect 2120 -390 2350 -260
rect 5138 -398 5368 -268
rect 7624 -398 7854 -268
rect 9044 -398 9274 -268
rect 13668 -394 13898 -264
rect 16868 -394 17098 -264
rect 20424 -394 20654 -264
rect 25758 -394 25988 -264
rect 28602 -394 28832 -264
rect 32514 -394 32744 -264
rect 34670 -394 34900 -264
rect 37492 -394 37722 -264
rect 40692 -394 40922 -264
rect 45668 -394 45898 -264
rect 48868 -394 49098 -264
rect 51002 -394 51232 -264
rect 54558 -394 54788 -264
rect 57402 -394 57632 -264
rect 61314 -394 61544 -264
rect 64158 -394 64388 -264
rect 67714 -394 67944 -264
rect 70558 -394 70788 -264
rect 74468 -394 74698 -264
rect 78380 -394 78610 -264
rect 82292 -394 82522 -264
rect 86202 -394 86432 -264
rect 230 -590 300 -530
rect 400 -590 470 -530
rect 570 -590 640 -530
rect 740 -590 810 -530
rect 910 -590 980 -530
rect 1080 -590 1150 -530
rect 1250 -590 1320 -530
rect 1420 -590 1490 -530
rect 1590 -590 1660 -530
rect 1760 -590 1830 -530
rect 1930 -590 2000 -530
rect 2100 -590 2170 -530
rect 2270 -590 2340 -530
rect 2440 -590 2510 -530
rect 2610 -590 2680 -530
rect 2780 -590 2850 -530
rect 2950 -590 3020 -530
rect 3120 -590 3190 -530
rect 3290 -590 3360 -530
rect 3460 -590 3530 -530
rect 3630 -590 3700 -530
rect 3800 -590 3870 -530
rect 3970 -590 4040 -530
rect 4140 -590 4210 -530
rect 4310 -590 4380 -530
rect 4480 -590 4550 -530
rect 4650 -590 4720 -530
rect 4820 -590 4890 -530
rect 4990 -590 5060 -530
rect 5160 -590 5230 -530
rect 5330 -590 5400 -530
rect 5500 -590 5570 -530
rect 5670 -590 5740 -530
rect 5840 -590 5910 -530
rect 6010 -590 6080 -530
rect 6180 -590 6250 -530
rect 6350 -590 6420 -530
rect 6520 -590 6590 -530
rect 6690 -590 6760 -530
rect 6860 -590 6930 -530
rect 7030 -590 7100 -530
rect 7200 -590 7270 -530
rect 7370 -590 7440 -530
rect 7540 -590 7610 -530
rect 7710 -590 7780 -530
rect 7880 -590 7950 -530
rect 8050 -590 8120 -530
rect 8220 -590 8290 -530
rect 8390 -590 8460 -530
rect 8560 -590 8630 -530
rect 8730 -590 8800 -530
rect 8900 -590 8970 -530
rect 9070 -590 9140 -530
rect 9240 -590 9310 -530
rect 9410 -590 9480 -530
rect 9580 -590 9650 -530
rect 9750 -590 9820 -530
rect 9920 -590 9990 -530
rect 10090 -590 10160 -530
rect 10260 -590 10330 -530
rect 10430 -590 10500 -530
rect 10600 -590 10670 -530
rect 10770 -590 10840 -530
rect 10940 -590 11010 -530
rect 11110 -590 11180 -530
rect 11280 -590 11350 -530
rect 11450 -590 11520 -530
rect 11620 -590 11690 -530
rect 11790 -590 11860 -530
rect 11960 -590 12030 -530
rect 12130 -590 12200 -530
rect 12300 -590 12370 -530
rect 12470 -590 12540 -530
rect 12640 -590 12710 -530
rect 12810 -590 12880 -530
rect 12980 -590 13050 -530
rect 13150 -590 13220 -530
rect 13320 -590 13390 -530
rect 13490 -590 13560 -530
rect 13660 -590 13730 -530
rect 13830 -590 13900 -530
rect 14000 -590 14070 -530
rect 14170 -590 14240 -530
rect 14340 -590 14410 -530
rect 14510 -590 14580 -530
rect 14680 -590 14750 -530
rect 14850 -590 14920 -530
rect 15020 -590 15090 -530
rect 15190 -590 15260 -530
rect 15360 -590 15430 -530
rect 15530 -590 15600 -530
rect 15700 -590 15770 -530
rect 15870 -590 15940 -530
rect 16040 -590 16110 -530
rect 16210 -590 16280 -530
rect 16380 -590 16450 -530
rect 16550 -590 16620 -530
rect 16720 -590 16790 -530
rect 16890 -590 16960 -530
rect 17060 -590 17130 -530
rect 17230 -590 17300 -530
rect 17400 -590 17470 -530
rect 17570 -590 17640 -530
rect 17740 -590 17810 -530
rect 17910 -590 17980 -530
rect 18080 -590 18150 -530
rect 18250 -590 18320 -530
rect 18420 -590 18490 -530
rect 18590 -590 18660 -530
rect 18760 -590 18830 -530
rect 18930 -590 19000 -530
rect 19100 -590 19170 -530
rect 19270 -590 19340 -530
rect 19440 -590 19510 -530
rect 19610 -590 19680 -530
rect 19780 -590 19850 -530
rect 19950 -590 20020 -530
rect 20120 -590 20190 -530
rect 20290 -590 20360 -530
rect 20460 -590 20530 -530
rect 20630 -590 20700 -530
rect 20800 -590 20870 -530
rect 20970 -590 21040 -530
rect 21140 -590 21210 -530
rect 21310 -590 21380 -530
rect 21480 -590 21550 -530
rect 21650 -590 21720 -530
rect 21820 -590 21890 -530
rect 21990 -590 22060 -530
rect 22160 -590 22230 -530
rect 22330 -590 22400 -530
rect 22500 -590 22570 -530
rect 22670 -590 22740 -530
rect 22840 -590 22910 -530
rect 23010 -590 23080 -530
rect 23180 -590 23250 -530
rect 23350 -590 23420 -530
rect 23520 -590 23590 -530
rect 23690 -590 23760 -530
rect 23860 -590 23930 -530
rect 24030 -590 24100 -530
rect 24200 -590 24270 -530
rect 24370 -590 24440 -530
rect 24540 -590 24610 -530
rect 24710 -590 24780 -530
rect 24880 -590 24950 -530
rect 25050 -590 25120 -530
rect 25220 -590 25290 -530
rect 25390 -590 25460 -530
rect 25560 -590 25630 -530
rect 25730 -590 25800 -530
rect 25900 -590 25970 -530
rect 26070 -590 26140 -530
rect 26240 -590 26310 -530
rect 26410 -590 26480 -530
rect 26580 -590 26650 -530
rect 26750 -590 26820 -530
rect 26920 -590 26990 -530
rect 27090 -590 27160 -530
rect 27260 -590 27330 -530
rect 27430 -590 27500 -530
rect 27600 -590 27670 -530
rect 27770 -590 27840 -530
rect 27940 -590 28010 -530
rect 28110 -590 28180 -530
rect 28280 -590 28350 -530
rect 28450 -590 28520 -530
rect 28620 -590 28690 -530
rect 28790 -590 28860 -530
rect 28960 -590 29030 -530
rect 29130 -590 29200 -530
rect 29300 -590 29370 -530
rect 29470 -590 29540 -530
rect 29640 -590 29710 -530
rect 29810 -590 29880 -530
rect 29980 -590 30050 -530
rect 30150 -590 30220 -530
rect 30320 -590 30390 -530
rect 30490 -590 30560 -530
rect 30660 -590 30730 -530
rect 30830 -590 30900 -530
rect 31000 -590 31070 -530
rect 31170 -590 31240 -530
rect 31340 -590 31410 -530
rect 31510 -590 31580 -530
rect 31680 -590 31750 -530
rect 31850 -590 31920 -530
rect 32020 -590 32090 -530
rect 32190 -590 32260 -530
rect 32360 -590 32430 -530
rect 32530 -590 32600 -530
rect 32700 -590 32770 -530
rect 32870 -590 32940 -530
rect 33040 -590 33110 -530
rect 33210 -590 33280 -530
rect 33380 -590 33450 -530
rect 33550 -590 33620 -530
rect 33720 -590 33790 -530
rect 33890 -590 33960 -530
rect 34060 -590 34130 -530
rect 34230 -590 34300 -530
rect 34400 -590 34470 -530
rect 34570 -590 34640 -530
rect 34740 -590 34810 -530
rect 34910 -590 34980 -530
rect 35080 -590 35150 -530
rect 35250 -590 35320 -530
rect 35420 -590 35490 -530
rect 35590 -590 35660 -530
rect 35760 -590 35830 -530
rect 35930 -590 36000 -530
rect 36100 -590 36170 -530
rect 36270 -590 36340 -530
rect 36440 -590 36510 -530
rect 36610 -590 36680 -530
rect 36780 -590 36850 -530
rect 36950 -590 37020 -530
rect 37120 -590 37190 -530
rect 37290 -590 37360 -530
rect 37460 -590 37530 -530
rect 37630 -590 37700 -530
rect 37800 -590 37870 -530
rect 37970 -590 38040 -530
rect 38140 -590 38210 -530
rect 38310 -590 38380 -530
rect 38480 -590 38550 -530
rect 38650 -590 38720 -530
rect 38820 -590 38890 -530
rect 38990 -590 39060 -530
rect 39160 -590 39230 -530
rect 39330 -590 39400 -530
rect 39500 -590 39570 -530
rect 39670 -590 39740 -530
rect 39840 -590 39910 -530
rect 40010 -590 40080 -530
rect 40180 -590 40250 -530
rect 40350 -590 40420 -530
rect 40520 -590 40590 -530
rect 40690 -590 40760 -530
rect 40860 -590 40930 -530
rect 41030 -590 41100 -530
rect 41200 -590 41270 -530
rect 41370 -590 41440 -530
rect 41540 -590 41610 -530
rect 41710 -590 41780 -530
rect 41880 -590 41950 -530
rect 42050 -590 42120 -530
rect 42220 -590 42290 -530
rect 42390 -590 42460 -530
rect 42560 -590 42630 -530
rect 42730 -590 42800 -530
rect 42900 -590 42970 -530
rect 43070 -590 43140 -530
rect 43240 -590 43310 -530
rect 43410 -590 43480 -530
rect 43580 -590 43650 -530
rect 43750 -590 43820 -530
rect 43920 -590 43990 -530
rect 44090 -590 44160 -530
rect 44260 -590 44330 -530
rect 44430 -590 44500 -530
rect 44600 -590 44670 -530
rect 44770 -590 44840 -530
rect 44940 -590 45010 -530
rect 45110 -590 45180 -530
rect 45280 -590 45350 -530
rect 45450 -590 45520 -530
rect 45620 -590 45690 -530
rect 45790 -590 45860 -530
rect 45960 -590 46030 -530
rect 46130 -590 46200 -530
rect 46300 -590 46370 -530
rect 46470 -590 46540 -530
rect 46640 -590 46710 -530
rect 46810 -590 46880 -530
rect 46980 -590 47050 -530
rect 47150 -590 47220 -530
rect 47320 -590 47390 -530
rect 47490 -590 47560 -530
rect 47660 -590 47730 -530
rect 47830 -590 47900 -530
rect 48000 -590 48070 -530
rect 48170 -590 48240 -530
rect 48340 -590 48410 -530
rect 48510 -590 48580 -530
rect 48680 -590 48750 -530
rect 48850 -590 48920 -530
rect 49020 -590 49090 -530
rect 49190 -590 49260 -530
rect 49360 -590 49430 -530
rect 49530 -590 49600 -530
rect 49700 -590 49770 -530
rect 49870 -590 49940 -530
rect 50040 -590 50110 -530
rect 50210 -590 50280 -530
rect 50380 -590 50450 -530
rect 50550 -590 50620 -530
rect 50720 -590 50790 -530
rect 50890 -590 50960 -530
rect 51060 -590 51130 -530
rect 51230 -590 51300 -530
rect 51400 -590 51470 -530
rect 51570 -590 51640 -530
rect 51740 -590 51810 -530
rect 51910 -590 51980 -530
rect 52080 -590 52150 -530
rect 52250 -590 52320 -530
rect 52420 -590 52490 -530
rect 52590 -590 52660 -530
rect 52760 -590 52830 -530
rect 52930 -590 53000 -530
rect 53100 -590 53170 -530
rect 53270 -590 53340 -530
rect 53440 -590 53510 -530
rect 53610 -590 53680 -530
rect 53780 -590 53850 -530
rect 53950 -590 54020 -530
rect 54120 -590 54190 -530
rect 54290 -590 54360 -530
rect 54460 -590 54530 -530
rect 54630 -590 54700 -530
rect 54800 -590 54870 -530
rect 54970 -590 55040 -530
rect 55140 -590 55210 -530
rect 55310 -590 55380 -530
rect 55480 -590 55550 -530
rect 55650 -590 55720 -530
rect 55820 -590 55890 -530
rect 55990 -590 56060 -530
rect 56160 -590 56230 -530
rect 56330 -590 56400 -530
rect 56500 -590 56570 -530
rect 56670 -590 56740 -530
rect 56840 -590 56910 -530
rect 57010 -590 57080 -530
rect 57180 -590 57250 -530
rect 57350 -590 57420 -530
rect 57520 -590 57590 -530
rect 57690 -590 57760 -530
rect 57860 -590 57930 -530
rect 58030 -590 58100 -530
rect 58200 -590 58270 -530
rect 58370 -590 58440 -530
rect 58540 -590 58610 -530
rect 58710 -590 58780 -530
rect 58880 -590 58950 -530
rect 59050 -590 59120 -530
rect 59220 -590 59290 -530
rect 59390 -590 59460 -530
rect 59560 -590 59630 -530
rect 59730 -590 59800 -530
rect 59900 -590 59970 -530
rect 60070 -590 60140 -530
rect 60240 -590 60310 -530
rect 60410 -590 60480 -530
rect 60580 -590 60650 -530
rect 60750 -590 60820 -530
rect 60920 -590 60990 -530
rect 61090 -590 61160 -530
rect 61260 -590 61330 -530
rect 61430 -590 61500 -530
rect 61600 -590 61670 -530
rect 61770 -590 61840 -530
rect 61940 -590 62010 -530
rect 62110 -590 62180 -530
rect 62280 -590 62350 -530
rect 62450 -590 62520 -530
rect 62620 -590 62690 -530
rect 62790 -590 62860 -530
rect 62960 -590 63030 -530
rect 63130 -590 63200 -530
rect 63300 -590 63370 -530
rect 63470 -590 63540 -530
rect 63640 -590 63710 -530
rect 63810 -590 63880 -530
rect 63980 -590 64050 -530
rect 64150 -590 64220 -530
rect 64320 -590 64390 -530
rect 64490 -590 64560 -530
rect 64660 -590 64730 -530
rect 64830 -590 64900 -530
rect 65000 -590 65070 -530
rect 65170 -590 65240 -530
rect 65340 -590 65410 -530
rect 65510 -590 65580 -530
rect 65680 -590 65750 -530
rect 65850 -590 65920 -530
rect 66020 -590 66090 -530
rect 66190 -590 66260 -530
rect 66360 -590 66430 -530
rect 66530 -590 66600 -530
rect 66700 -590 66770 -530
rect 66870 -590 66940 -530
rect 67040 -590 67110 -530
rect 67210 -590 67280 -530
rect 67380 -590 67450 -530
rect 67550 -590 67620 -530
rect 67720 -590 67790 -530
rect 67890 -590 67960 -530
rect 68060 -590 68130 -530
rect 68230 -590 68300 -530
rect 68400 -590 68470 -530
rect 68570 -590 68640 -530
rect 68740 -590 68810 -530
rect 68910 -590 68980 -530
rect 69080 -590 69150 -530
rect 69250 -590 69320 -530
rect 69420 -590 69490 -530
rect 69590 -590 69660 -530
rect 69760 -590 69830 -530
rect 69930 -590 70000 -530
rect 70100 -590 70170 -530
rect 70270 -590 70340 -530
rect 70440 -590 70510 -530
rect 70610 -590 70680 -530
rect 70780 -590 70850 -530
rect 70950 -590 71020 -530
rect 71120 -590 71190 -530
rect 71290 -590 71360 -530
rect 71460 -590 71530 -530
rect 71630 -590 71700 -530
rect 71800 -590 71870 -530
rect 71970 -590 72040 -530
rect 72140 -590 72210 -530
rect 72310 -590 72380 -530
rect 72480 -590 72550 -530
rect 72650 -590 72720 -530
rect 72820 -590 72890 -530
rect 72990 -590 73060 -530
rect 73160 -590 73230 -530
rect 73330 -590 73400 -530
rect 73500 -590 73570 -530
rect 73670 -590 73740 -530
rect 73840 -590 73910 -530
rect 74010 -590 74080 -530
rect 74180 -590 74250 -530
rect 74350 -590 74420 -530
rect 74520 -590 74590 -530
rect 74690 -590 74760 -530
rect 74860 -590 74930 -530
rect 75030 -590 75100 -530
rect 75200 -590 75270 -530
rect 75370 -590 75440 -530
rect 75540 -590 75610 -530
rect 75710 -590 75780 -530
rect 75880 -590 75950 -530
rect 76050 -590 76120 -530
rect 76220 -590 76290 -530
rect 76390 -590 76460 -530
rect 76560 -590 76630 -530
rect 76730 -590 76800 -530
rect 76900 -590 76970 -530
rect 77070 -590 77140 -530
rect 77240 -590 77310 -530
rect 77410 -590 77480 -530
rect 77580 -590 77650 -530
rect 77750 -590 77820 -530
rect 77920 -590 77990 -530
rect 78090 -590 78160 -530
rect 78260 -590 78330 -530
rect 78430 -590 78500 -530
rect 78600 -590 78670 -530
rect 78770 -590 78840 -530
rect 78940 -590 79010 -530
rect 79110 -590 79180 -530
rect 79280 -590 79350 -530
rect 79450 -590 79520 -530
rect 79620 -590 79690 -530
rect 79790 -590 79860 -530
rect 79960 -590 80030 -530
rect 80130 -590 80200 -530
rect 80300 -590 80370 -530
rect 80470 -590 80540 -530
rect 80640 -590 80710 -530
rect 80810 -590 80880 -530
rect 80980 -590 81050 -530
rect 81150 -590 81220 -530
rect 81320 -590 81390 -530
rect 81490 -590 81560 -530
rect 81660 -590 81730 -530
rect 81830 -590 81900 -530
rect 82000 -590 82070 -530
rect 82170 -590 82240 -530
rect 82340 -590 82410 -530
rect 82510 -590 82580 -530
rect 82680 -590 82750 -530
rect 82850 -590 82920 -530
rect 83020 -590 83090 -530
rect 83190 -590 83260 -530
rect 83360 -590 83430 -530
rect 83530 -590 83600 -530
rect 83700 -590 83770 -530
rect 83870 -590 83940 -530
rect 84040 -590 84110 -530
rect 84210 -590 84280 -530
rect 84380 -590 84450 -530
rect 84550 -590 84620 -530
rect 84720 -590 84790 -530
rect 84890 -590 84960 -530
rect 85060 -590 85130 -530
rect 85230 -590 85300 -530
rect 85400 -590 85470 -530
rect 85570 -590 85640 -530
rect 85740 -590 85810 -530
rect 85910 -590 85980 -530
rect 86080 -590 86150 -530
rect 86250 -590 86320 -530
rect 86420 -590 86490 -530
rect 86590 -590 86660 -530
rect 86760 -590 86830 -530
rect 86930 -590 87000 -530
rect 87100 -590 87170 -530
rect 150 -730 210 -670
rect 320 -830 380 -770
rect 490 -730 550 -670
rect 660 -830 720 -770
rect 830 -730 890 -670
rect 1000 -830 1060 -770
rect 1170 -730 1230 -670
rect 1340 -830 1400 -770
rect 1510 -730 1570 -670
rect 1680 -830 1740 -770
rect 1850 -730 1910 -670
rect 2020 -830 2080 -770
rect 2190 -730 2250 -670
rect 2360 -830 2420 -770
rect 2530 -730 2590 -670
rect 2700 -830 2760 -770
rect 2870 -730 2930 -670
rect 3040 -830 3100 -770
rect 3210 -730 3270 -670
rect 3380 -830 3440 -770
rect 3550 -730 3610 -670
rect 3720 -830 3780 -770
rect 3890 -730 3950 -670
rect 4060 -830 4120 -770
rect 4230 -730 4290 -670
rect 4400 -830 4460 -770
rect 4570 -730 4630 -670
rect 4740 -830 4800 -770
rect 4910 -730 4970 -670
rect 5080 -830 5140 -770
rect 5250 -730 5310 -670
rect 5420 -830 5480 -770
rect 5590 -730 5650 -670
rect 5760 -830 5820 -770
rect 5930 -730 5990 -670
rect 6100 -830 6160 -770
rect 6270 -730 6330 -670
rect 6440 -830 6500 -770
rect 6610 -730 6670 -670
rect 6780 -830 6840 -770
rect 6950 -730 7010 -670
rect 7120 -830 7180 -770
rect 7290 -730 7350 -670
rect 7460 -830 7520 -770
rect 7630 -730 7690 -670
rect 7800 -830 7860 -770
rect 7970 -730 8030 -670
rect 8140 -830 8200 -770
rect 8310 -730 8370 -670
rect 8480 -830 8540 -770
rect 8650 -730 8710 -670
rect 8820 -830 8880 -770
rect 8990 -730 9050 -670
rect 9160 -830 9220 -770
rect 9330 -730 9390 -670
rect 9500 -830 9560 -770
rect 9670 -730 9730 -670
rect 9840 -830 9900 -770
rect 10010 -730 10070 -670
rect 10180 -830 10240 -770
rect 10350 -730 10410 -670
rect 10520 -830 10580 -770
rect 10690 -730 10750 -670
rect 10860 -830 10920 -770
rect 11030 -730 11090 -670
rect 11200 -830 11260 -770
rect 11370 -730 11430 -670
rect 11540 -830 11600 -770
rect 11710 -730 11770 -670
rect 11880 -830 11940 -770
rect 12050 -730 12110 -670
rect 12220 -830 12280 -770
rect 12390 -730 12450 -670
rect 12560 -830 12620 -770
rect 12730 -730 12790 -670
rect 12900 -830 12960 -770
rect 13070 -730 13130 -670
rect 13240 -830 13300 -770
rect 13410 -730 13470 -670
rect 13580 -830 13640 -770
rect 13750 -730 13810 -670
rect 13920 -830 13980 -770
rect 14090 -730 14150 -670
rect 14260 -830 14320 -770
rect 14430 -730 14490 -670
rect 14600 -830 14660 -770
rect 14770 -730 14830 -670
rect 14940 -830 15000 -770
rect 15110 -730 15170 -670
rect 15280 -830 15340 -770
rect 15450 -730 15510 -670
rect 15620 -830 15680 -770
rect 15790 -730 15850 -670
rect 15960 -830 16020 -770
rect 16130 -730 16190 -670
rect 16300 -830 16360 -770
rect 16470 -730 16530 -670
rect 16640 -830 16700 -770
rect 16810 -730 16870 -670
rect 16980 -830 17040 -770
rect 17150 -730 17210 -670
rect 17320 -830 17380 -770
rect 17490 -730 17550 -670
rect 17660 -830 17720 -770
rect 17830 -730 17890 -670
rect 18000 -830 18060 -770
rect 18170 -730 18230 -670
rect 18340 -830 18400 -770
rect 18510 -730 18570 -670
rect 18680 -830 18740 -770
rect 18850 -730 18910 -670
rect 19020 -830 19080 -770
rect 19190 -730 19250 -670
rect 19360 -830 19420 -770
rect 19530 -730 19590 -670
rect 19700 -830 19760 -770
rect 19870 -730 19930 -670
rect 20040 -830 20100 -770
rect 20210 -730 20270 -670
rect 20380 -830 20440 -770
rect 20550 -730 20610 -670
rect 20720 -830 20780 -770
rect 20890 -730 20950 -670
rect 21060 -830 21120 -770
rect 21230 -730 21290 -670
rect 21400 -830 21460 -770
rect 21570 -730 21630 -670
rect 21740 -830 21800 -770
rect 21910 -730 21970 -670
rect 22080 -830 22140 -770
rect 22250 -730 22310 -670
rect 22420 -830 22480 -770
rect 22590 -730 22650 -670
rect 22760 -830 22820 -770
rect 22930 -730 22990 -670
rect 23100 -830 23160 -770
rect 23270 -730 23330 -670
rect 23440 -830 23500 -770
rect 23610 -730 23670 -670
rect 23780 -830 23840 -770
rect 23950 -730 24010 -670
rect 24120 -830 24180 -770
rect 24290 -730 24350 -670
rect 24460 -830 24520 -770
rect 24630 -730 24690 -670
rect 24800 -830 24860 -770
rect 24970 -730 25030 -670
rect 25140 -830 25200 -770
rect 25310 -730 25370 -670
rect 25480 -830 25540 -770
rect 25650 -730 25710 -670
rect 25820 -830 25880 -770
rect 25990 -730 26050 -670
rect 26160 -830 26220 -770
rect 26330 -730 26390 -670
rect 26500 -830 26560 -770
rect 26670 -730 26730 -670
rect 26840 -830 26900 -770
rect 27010 -730 27070 -670
rect 27180 -830 27240 -770
rect 27350 -730 27410 -670
rect 27520 -830 27580 -770
rect 27690 -730 27750 -670
rect 27860 -830 27920 -770
rect 28030 -730 28090 -670
rect 28200 -830 28260 -770
rect 28370 -730 28430 -670
rect 28540 -830 28600 -770
rect 28710 -730 28770 -670
rect 28880 -830 28940 -770
rect 29050 -730 29110 -670
rect 29220 -830 29280 -770
rect 29390 -730 29450 -670
rect 29560 -830 29620 -770
rect 29730 -730 29790 -670
rect 29900 -830 29960 -770
rect 30070 -730 30130 -670
rect 30240 -830 30300 -770
rect 30410 -730 30470 -670
rect 30580 -830 30640 -770
rect 30750 -730 30810 -670
rect 30920 -830 30980 -770
rect 31090 -730 31150 -670
rect 31260 -830 31320 -770
rect 31430 -730 31490 -670
rect 31600 -830 31660 -770
rect 31770 -730 31830 -670
rect 31940 -830 32000 -770
rect 32110 -730 32170 -670
rect 32280 -830 32340 -770
rect 32450 -730 32510 -670
rect 32620 -830 32680 -770
rect 32790 -730 32850 -670
rect 32960 -830 33020 -770
rect 33130 -730 33190 -670
rect 33300 -830 33360 -770
rect 33470 -730 33530 -670
rect 33640 -830 33700 -770
rect 33810 -730 33870 -670
rect 33980 -830 34040 -770
rect 34150 -730 34210 -670
rect 34320 -830 34380 -770
rect 34490 -730 34550 -670
rect 34660 -830 34720 -770
rect 34830 -730 34890 -670
rect 35000 -830 35060 -770
rect 35170 -730 35230 -670
rect 35340 -830 35400 -770
rect 35510 -730 35570 -670
rect 35680 -830 35740 -770
rect 35850 -730 35910 -670
rect 36020 -830 36080 -770
rect 36190 -730 36250 -670
rect 36360 -830 36420 -770
rect 36530 -730 36590 -670
rect 36700 -830 36760 -770
rect 36870 -730 36930 -670
rect 37040 -830 37100 -770
rect 37210 -730 37270 -670
rect 37380 -830 37440 -770
rect 37550 -730 37610 -670
rect 37720 -830 37780 -770
rect 37890 -730 37950 -670
rect 38060 -830 38120 -770
rect 38230 -730 38290 -670
rect 38400 -830 38460 -770
rect 38570 -730 38630 -670
rect 38740 -830 38800 -770
rect 38910 -730 38970 -670
rect 39080 -830 39140 -770
rect 39250 -730 39310 -670
rect 39420 -830 39480 -770
rect 39590 -730 39650 -670
rect 39760 -830 39820 -770
rect 39930 -730 39990 -670
rect 40100 -830 40160 -770
rect 40270 -730 40330 -670
rect 40440 -830 40500 -770
rect 40610 -730 40670 -670
rect 40780 -830 40840 -770
rect 40950 -730 41010 -670
rect 41120 -830 41180 -770
rect 41290 -730 41350 -670
rect 41460 -830 41520 -770
rect 41630 -730 41690 -670
rect 41800 -830 41860 -770
rect 41970 -730 42030 -670
rect 42140 -830 42200 -770
rect 42310 -730 42370 -670
rect 42480 -830 42540 -770
rect 42650 -730 42710 -670
rect 42820 -830 42880 -770
rect 42990 -730 43050 -670
rect 43160 -830 43220 -770
rect 43330 -730 43390 -670
rect 43500 -830 43560 -770
rect 43670 -730 43730 -670
rect 43840 -830 43900 -770
rect 44010 -730 44070 -670
rect 44180 -830 44240 -770
rect 44350 -730 44410 -670
rect 44520 -830 44580 -770
rect 44690 -730 44750 -670
rect 44860 -830 44920 -770
rect 45030 -730 45090 -670
rect 45200 -830 45260 -770
rect 45370 -730 45430 -670
rect 45540 -830 45600 -770
rect 45710 -730 45770 -670
rect 45880 -830 45940 -770
rect 46050 -730 46110 -670
rect 46220 -830 46280 -770
rect 46390 -730 46450 -670
rect 46560 -830 46620 -770
rect 46730 -730 46790 -670
rect 46900 -830 46960 -770
rect 47070 -730 47130 -670
rect 47240 -830 47300 -770
rect 47410 -730 47470 -670
rect 47580 -830 47640 -770
rect 47750 -730 47810 -670
rect 47920 -830 47980 -770
rect 48090 -730 48150 -670
rect 48260 -830 48320 -770
rect 48430 -730 48490 -670
rect 48600 -830 48660 -770
rect 48770 -730 48830 -670
rect 48940 -830 49000 -770
rect 49110 -730 49170 -670
rect 49280 -830 49340 -770
rect 49450 -730 49510 -670
rect 49620 -830 49680 -770
rect 49790 -730 49850 -670
rect 49960 -830 50020 -770
rect 50130 -730 50190 -670
rect 50300 -830 50360 -770
rect 50470 -730 50530 -670
rect 50640 -830 50700 -770
rect 50810 -730 50870 -670
rect 50980 -830 51040 -770
rect 51150 -730 51210 -670
rect 51320 -830 51380 -770
rect 51490 -730 51550 -670
rect 51660 -830 51720 -770
rect 51830 -730 51890 -670
rect 52000 -830 52060 -770
rect 52170 -730 52230 -670
rect 52340 -830 52400 -770
rect 52510 -730 52570 -670
rect 52680 -830 52740 -770
rect 52850 -730 52910 -670
rect 53020 -830 53080 -770
rect 53190 -730 53250 -670
rect 53360 -830 53420 -770
rect 53530 -730 53590 -670
rect 53700 -830 53760 -770
rect 53870 -730 53930 -670
rect 54040 -830 54100 -770
rect 54210 -730 54270 -670
rect 54380 -830 54440 -770
rect 54550 -730 54610 -670
rect 54720 -830 54780 -770
rect 54890 -730 54950 -670
rect 55060 -830 55120 -770
rect 55230 -730 55290 -670
rect 55400 -830 55460 -770
rect 55570 -730 55630 -670
rect 55740 -830 55800 -770
rect 55910 -730 55970 -670
rect 56080 -830 56140 -770
rect 56250 -730 56310 -670
rect 56420 -830 56480 -770
rect 56590 -730 56650 -670
rect 56760 -830 56820 -770
rect 56930 -730 56990 -670
rect 57100 -830 57160 -770
rect 57270 -730 57330 -670
rect 57440 -830 57500 -770
rect 57610 -730 57670 -670
rect 57780 -830 57840 -770
rect 57950 -730 58010 -670
rect 58120 -830 58180 -770
rect 58290 -730 58350 -670
rect 58460 -830 58520 -770
rect 58630 -730 58690 -670
rect 58800 -830 58860 -770
rect 58970 -730 59030 -670
rect 59140 -830 59200 -770
rect 59310 -730 59370 -670
rect 59480 -830 59540 -770
rect 59650 -730 59710 -670
rect 59820 -830 59880 -770
rect 59990 -730 60050 -670
rect 60160 -830 60220 -770
rect 60330 -730 60390 -670
rect 60500 -830 60560 -770
rect 60670 -730 60730 -670
rect 60840 -830 60900 -770
rect 61010 -730 61070 -670
rect 61180 -830 61240 -770
rect 61350 -730 61410 -670
rect 61520 -830 61580 -770
rect 61690 -730 61750 -670
rect 61860 -830 61920 -770
rect 62030 -730 62090 -670
rect 62200 -830 62260 -770
rect 62370 -730 62430 -670
rect 62540 -830 62600 -770
rect 62710 -730 62770 -670
rect 62880 -830 62940 -770
rect 63050 -730 63110 -670
rect 63220 -830 63280 -770
rect 63390 -730 63450 -670
rect 63560 -830 63620 -770
rect 63730 -730 63790 -670
rect 63900 -830 63960 -770
rect 64070 -730 64130 -670
rect 64240 -830 64300 -770
rect 64410 -730 64470 -670
rect 64580 -830 64640 -770
rect 64750 -730 64810 -670
rect 64920 -830 64980 -770
rect 65090 -730 65150 -670
rect 65260 -830 65320 -770
rect 65430 -730 65490 -670
rect 65600 -830 65660 -770
rect 65770 -730 65830 -670
rect 65940 -830 66000 -770
rect 66110 -730 66170 -670
rect 66280 -830 66340 -770
rect 66450 -730 66510 -670
rect 66620 -830 66680 -770
rect 66790 -730 66850 -670
rect 66960 -830 67020 -770
rect 67130 -730 67190 -670
rect 67300 -830 67360 -770
rect 67470 -730 67530 -670
rect 67640 -830 67700 -770
rect 67810 -730 67870 -670
rect 67980 -830 68040 -770
rect 68150 -730 68210 -670
rect 68320 -830 68380 -770
rect 68490 -730 68550 -670
rect 68660 -830 68720 -770
rect 68830 -730 68890 -670
rect 69000 -830 69060 -770
rect 69170 -730 69230 -670
rect 69340 -830 69400 -770
rect 69510 -730 69570 -670
rect 69680 -830 69740 -770
rect 69850 -730 69910 -670
rect 70020 -830 70080 -770
rect 70190 -730 70250 -670
rect 70360 -830 70420 -770
rect 70530 -730 70590 -670
rect 70700 -830 70760 -770
rect 70870 -730 70930 -670
rect 71040 -830 71100 -770
rect 71210 -730 71270 -670
rect 71380 -830 71440 -770
rect 71550 -730 71610 -670
rect 71720 -830 71780 -770
rect 71890 -730 71950 -670
rect 72060 -830 72120 -770
rect 72230 -730 72290 -670
rect 72400 -830 72460 -770
rect 72570 -730 72630 -670
rect 72740 -830 72800 -770
rect 72910 -730 72970 -670
rect 73080 -830 73140 -770
rect 73250 -730 73310 -670
rect 73420 -830 73480 -770
rect 73590 -730 73650 -670
rect 73760 -830 73820 -770
rect 73930 -730 73990 -670
rect 74100 -830 74160 -770
rect 74270 -730 74330 -670
rect 74440 -830 74500 -770
rect 74610 -730 74670 -670
rect 74780 -830 74840 -770
rect 74950 -730 75010 -670
rect 75120 -830 75180 -770
rect 75290 -730 75350 -670
rect 75460 -830 75520 -770
rect 75630 -730 75690 -670
rect 75800 -830 75860 -770
rect 75970 -730 76030 -670
rect 76140 -830 76200 -770
rect 76310 -730 76370 -670
rect 76480 -830 76540 -770
rect 76650 -730 76710 -670
rect 76820 -830 76880 -770
rect 76990 -730 77050 -670
rect 77160 -830 77220 -770
rect 77330 -730 77390 -670
rect 77500 -830 77560 -770
rect 77670 -730 77730 -670
rect 77840 -830 77900 -770
rect 78010 -730 78070 -670
rect 78180 -830 78240 -770
rect 78350 -730 78410 -670
rect 78520 -830 78580 -770
rect 78690 -730 78750 -670
rect 78860 -830 78920 -770
rect 79030 -730 79090 -670
rect 79200 -830 79260 -770
rect 79370 -730 79430 -670
rect 79540 -830 79600 -770
rect 79710 -730 79770 -670
rect 79880 -830 79940 -770
rect 80050 -730 80110 -670
rect 80220 -830 80280 -770
rect 80390 -730 80450 -670
rect 80560 -830 80620 -770
rect 80730 -730 80790 -670
rect 80900 -830 80960 -770
rect 81070 -730 81130 -670
rect 81240 -830 81300 -770
rect 81410 -730 81470 -670
rect 81580 -830 81640 -770
rect 81750 -730 81810 -670
rect 81920 -830 81980 -770
rect 82090 -730 82150 -670
rect 82260 -830 82320 -770
rect 82430 -730 82490 -670
rect 82600 -830 82660 -770
rect 82770 -730 82830 -670
rect 82940 -830 83000 -770
rect 83110 -730 83170 -670
rect 83280 -830 83340 -770
rect 83450 -730 83510 -670
rect 83620 -830 83680 -770
rect 83790 -730 83850 -670
rect 83960 -830 84020 -770
rect 84130 -730 84190 -670
rect 84300 -830 84360 -770
rect 84470 -730 84530 -670
rect 84640 -830 84700 -770
rect 84810 -730 84870 -670
rect 84980 -830 85040 -770
rect 85150 -730 85210 -670
rect 85320 -830 85380 -770
rect 85490 -730 85550 -670
rect 85660 -830 85720 -770
rect 85830 -730 85890 -670
rect 86000 -830 86060 -770
rect 86170 -730 86230 -670
rect 86340 -830 86400 -770
rect 86510 -730 86570 -670
rect 86680 -830 86740 -770
rect 86850 -730 86910 -670
rect 87020 -830 87080 -770
rect 87190 -730 87250 -670
rect 150 -1160 210 -1100
rect 150 -1360 210 -1300
rect 320 -1060 380 -1000
rect 320 -1260 380 -1200
rect 490 -1160 550 -1100
rect 490 -1360 550 -1300
rect 660 -1060 720 -1000
rect 660 -1260 720 -1200
rect 830 -1160 890 -1100
rect 830 -1360 890 -1300
rect 1000 -1060 1060 -1000
rect 1000 -1260 1060 -1200
rect 1170 -1160 1230 -1100
rect 1170 -1360 1230 -1300
rect 1340 -1060 1400 -1000
rect 1340 -1260 1400 -1200
rect 1510 -1160 1570 -1100
rect 1510 -1360 1570 -1300
rect 1680 -1060 1740 -1000
rect 1680 -1260 1740 -1200
rect 1850 -1160 1910 -1100
rect 1850 -1360 1910 -1300
rect 2020 -1060 2080 -1000
rect 2020 -1260 2080 -1200
rect 2190 -1160 2250 -1100
rect 2190 -1360 2250 -1300
rect 2360 -1060 2420 -1000
rect 2360 -1260 2420 -1200
rect 2530 -1160 2590 -1100
rect 2530 -1360 2590 -1300
rect 2700 -1060 2760 -1000
rect 2700 -1260 2760 -1200
rect 2870 -1160 2930 -1100
rect 2870 -1360 2930 -1300
rect 3040 -1060 3100 -1000
rect 3040 -1260 3100 -1200
rect 3210 -1160 3270 -1100
rect 3210 -1360 3270 -1300
rect 3380 -1060 3440 -1000
rect 3380 -1260 3440 -1200
rect 3550 -1160 3610 -1100
rect 3550 -1360 3610 -1300
rect 3720 -1060 3780 -1000
rect 3720 -1260 3780 -1200
rect 3890 -1160 3950 -1100
rect 3890 -1360 3950 -1300
rect 4060 -1060 4120 -1000
rect 4060 -1260 4120 -1200
rect 4230 -1160 4290 -1100
rect 4230 -1360 4290 -1300
rect 4400 -1060 4460 -1000
rect 4400 -1260 4460 -1200
rect 4570 -1160 4630 -1100
rect 4570 -1360 4630 -1300
rect 4740 -1060 4800 -1000
rect 4740 -1260 4800 -1200
rect 4910 -1160 4970 -1100
rect 4910 -1360 4970 -1300
rect 5080 -1060 5140 -1000
rect 5080 -1260 5140 -1200
rect 5250 -1160 5310 -1100
rect 5250 -1360 5310 -1300
rect 5420 -1060 5480 -1000
rect 5420 -1260 5480 -1200
rect 5590 -1160 5650 -1100
rect 5590 -1360 5650 -1300
rect 5760 -1060 5820 -1000
rect 5760 -1260 5820 -1200
rect 5930 -1160 5990 -1100
rect 5930 -1360 5990 -1300
rect 6100 -1060 6160 -1000
rect 6100 -1260 6160 -1200
rect 6270 -1160 6330 -1100
rect 6270 -1360 6330 -1300
rect 6440 -1060 6500 -1000
rect 6440 -1260 6500 -1200
rect 6610 -1160 6670 -1100
rect 6610 -1360 6670 -1300
rect 6780 -1060 6840 -1000
rect 6780 -1260 6840 -1200
rect 6950 -1160 7010 -1100
rect 6950 -1360 7010 -1300
rect 7120 -1060 7180 -1000
rect 7120 -1260 7180 -1200
rect 7290 -1160 7350 -1100
rect 7290 -1360 7350 -1300
rect 7460 -1060 7520 -1000
rect 7460 -1260 7520 -1200
rect 7630 -1160 7690 -1100
rect 7630 -1360 7690 -1300
rect 7800 -1060 7860 -1000
rect 7800 -1260 7860 -1200
rect 7970 -1160 8030 -1100
rect 7970 -1360 8030 -1300
rect 8140 -1060 8200 -1000
rect 8140 -1260 8200 -1200
rect 8310 -1160 8370 -1100
rect 8310 -1360 8370 -1300
rect 8480 -1060 8540 -1000
rect 8480 -1260 8540 -1200
rect 8650 -1160 8710 -1100
rect 8650 -1360 8710 -1300
rect 8820 -1060 8880 -1000
rect 8820 -1260 8880 -1200
rect 8990 -1160 9050 -1100
rect 8990 -1360 9050 -1300
rect 9160 -1060 9220 -1000
rect 9160 -1260 9220 -1200
rect 9330 -1160 9390 -1100
rect 9330 -1360 9390 -1300
rect 9500 -1060 9560 -1000
rect 9500 -1260 9560 -1200
rect 9670 -1160 9730 -1100
rect 9670 -1360 9730 -1300
rect 9840 -1060 9900 -1000
rect 9840 -1260 9900 -1200
rect 10010 -1160 10070 -1100
rect 10010 -1360 10070 -1300
rect 10180 -1060 10240 -1000
rect 10180 -1260 10240 -1200
rect 10350 -1160 10410 -1100
rect 10350 -1360 10410 -1300
rect 10520 -1060 10580 -1000
rect 10520 -1260 10580 -1200
rect 10690 -1160 10750 -1100
rect 10690 -1360 10750 -1300
rect 10860 -1060 10920 -1000
rect 10860 -1260 10920 -1200
rect 11030 -1160 11090 -1100
rect 11030 -1360 11090 -1300
rect 11200 -1060 11260 -1000
rect 11200 -1260 11260 -1200
rect 11370 -1160 11430 -1100
rect 11370 -1360 11430 -1300
rect 11540 -1060 11600 -1000
rect 11540 -1260 11600 -1200
rect 11710 -1160 11770 -1100
rect 11710 -1360 11770 -1300
rect 11880 -1060 11940 -1000
rect 11880 -1260 11940 -1200
rect 12050 -1160 12110 -1100
rect 12050 -1360 12110 -1300
rect 12220 -1060 12280 -1000
rect 12220 -1260 12280 -1200
rect 12390 -1160 12450 -1100
rect 12390 -1360 12450 -1300
rect 12560 -1060 12620 -1000
rect 12560 -1260 12620 -1200
rect 12730 -1160 12790 -1100
rect 12730 -1360 12790 -1300
rect 12900 -1060 12960 -1000
rect 12900 -1260 12960 -1200
rect 13070 -1160 13130 -1100
rect 13070 -1360 13130 -1300
rect 13240 -1060 13300 -1000
rect 13240 -1260 13300 -1200
rect 13410 -1160 13470 -1100
rect 13410 -1360 13470 -1300
rect 13580 -1060 13640 -1000
rect 13580 -1260 13640 -1200
rect 13750 -1160 13810 -1100
rect 13750 -1360 13810 -1300
rect 13920 -1060 13980 -1000
rect 13920 -1260 13980 -1200
rect 14090 -1160 14150 -1100
rect 14090 -1360 14150 -1300
rect 14260 -1060 14320 -1000
rect 14260 -1260 14320 -1200
rect 14430 -1160 14490 -1100
rect 14430 -1360 14490 -1300
rect 14600 -1060 14660 -1000
rect 14600 -1260 14660 -1200
rect 14770 -1160 14830 -1100
rect 14770 -1360 14830 -1300
rect 14940 -1060 15000 -1000
rect 14940 -1260 15000 -1200
rect 15110 -1160 15170 -1100
rect 15110 -1360 15170 -1300
rect 15280 -1060 15340 -1000
rect 15280 -1260 15340 -1200
rect 15450 -1160 15510 -1100
rect 15450 -1360 15510 -1300
rect 15620 -1060 15680 -1000
rect 15620 -1260 15680 -1200
rect 15790 -1160 15850 -1100
rect 15790 -1360 15850 -1300
rect 15960 -1060 16020 -1000
rect 15960 -1260 16020 -1200
rect 16130 -1160 16190 -1100
rect 16130 -1360 16190 -1300
rect 16300 -1060 16360 -1000
rect 16300 -1260 16360 -1200
rect 16470 -1160 16530 -1100
rect 16470 -1360 16530 -1300
rect 16640 -1060 16700 -1000
rect 16640 -1260 16700 -1200
rect 16810 -1160 16870 -1100
rect 16810 -1360 16870 -1300
rect 16980 -1060 17040 -1000
rect 16980 -1260 17040 -1200
rect 17150 -1160 17210 -1100
rect 17150 -1360 17210 -1300
rect 17320 -1060 17380 -1000
rect 17320 -1260 17380 -1200
rect 17490 -1160 17550 -1100
rect 17490 -1360 17550 -1300
rect 17660 -1060 17720 -1000
rect 17660 -1260 17720 -1200
rect 17830 -1160 17890 -1100
rect 17830 -1360 17890 -1300
rect 18000 -1060 18060 -1000
rect 18000 -1260 18060 -1200
rect 18170 -1160 18230 -1100
rect 18170 -1360 18230 -1300
rect 18340 -1060 18400 -1000
rect 18340 -1260 18400 -1200
rect 18510 -1160 18570 -1100
rect 18510 -1360 18570 -1300
rect 18680 -1060 18740 -1000
rect 18680 -1260 18740 -1200
rect 18850 -1160 18910 -1100
rect 18850 -1360 18910 -1300
rect 19020 -1060 19080 -1000
rect 19020 -1260 19080 -1200
rect 19190 -1160 19250 -1100
rect 19190 -1360 19250 -1300
rect 19360 -1060 19420 -1000
rect 19360 -1260 19420 -1200
rect 19530 -1160 19590 -1100
rect 19530 -1360 19590 -1300
rect 19700 -1060 19760 -1000
rect 19700 -1260 19760 -1200
rect 19870 -1160 19930 -1100
rect 19870 -1360 19930 -1300
rect 20040 -1060 20100 -1000
rect 20040 -1260 20100 -1200
rect 20210 -1160 20270 -1100
rect 20210 -1360 20270 -1300
rect 20380 -1060 20440 -1000
rect 20380 -1260 20440 -1200
rect 20550 -1160 20610 -1100
rect 20550 -1360 20610 -1300
rect 20720 -1060 20780 -1000
rect 20720 -1260 20780 -1200
rect 20890 -1160 20950 -1100
rect 20890 -1360 20950 -1300
rect 21060 -1060 21120 -1000
rect 21060 -1260 21120 -1200
rect 21230 -1160 21290 -1100
rect 21230 -1360 21290 -1300
rect 21400 -1060 21460 -1000
rect 21400 -1260 21460 -1200
rect 21570 -1160 21630 -1100
rect 21570 -1360 21630 -1300
rect 21740 -1060 21800 -1000
rect 21740 -1260 21800 -1200
rect 21910 -1160 21970 -1100
rect 21910 -1360 21970 -1300
rect 22080 -1060 22140 -1000
rect 22080 -1260 22140 -1200
rect 22250 -1160 22310 -1100
rect 22250 -1360 22310 -1300
rect 22420 -1060 22480 -1000
rect 22420 -1260 22480 -1200
rect 22590 -1160 22650 -1100
rect 22590 -1360 22650 -1300
rect 22760 -1060 22820 -1000
rect 22760 -1260 22820 -1200
rect 22930 -1160 22990 -1100
rect 22930 -1360 22990 -1300
rect 23100 -1060 23160 -1000
rect 23100 -1260 23160 -1200
rect 23270 -1160 23330 -1100
rect 23270 -1360 23330 -1300
rect 23440 -1060 23500 -1000
rect 23440 -1260 23500 -1200
rect 23610 -1160 23670 -1100
rect 23610 -1360 23670 -1300
rect 23780 -1060 23840 -1000
rect 23780 -1260 23840 -1200
rect 23950 -1160 24010 -1100
rect 23950 -1360 24010 -1300
rect 24120 -1060 24180 -1000
rect 24120 -1260 24180 -1200
rect 24290 -1160 24350 -1100
rect 24290 -1360 24350 -1300
rect 24460 -1060 24520 -1000
rect 24460 -1260 24520 -1200
rect 24630 -1160 24690 -1100
rect 24630 -1360 24690 -1300
rect 24800 -1060 24860 -1000
rect 24800 -1260 24860 -1200
rect 24970 -1160 25030 -1100
rect 24970 -1360 25030 -1300
rect 25140 -1060 25200 -1000
rect 25140 -1260 25200 -1200
rect 25310 -1160 25370 -1100
rect 25310 -1360 25370 -1300
rect 25480 -1060 25540 -1000
rect 25480 -1260 25540 -1200
rect 25650 -1160 25710 -1100
rect 25650 -1360 25710 -1300
rect 25820 -1060 25880 -1000
rect 25820 -1260 25880 -1200
rect 25990 -1160 26050 -1100
rect 25990 -1360 26050 -1300
rect 26160 -1060 26220 -1000
rect 26160 -1260 26220 -1200
rect 26330 -1160 26390 -1100
rect 26330 -1360 26390 -1300
rect 26500 -1060 26560 -1000
rect 26500 -1260 26560 -1200
rect 26670 -1160 26730 -1100
rect 26670 -1360 26730 -1300
rect 26840 -1060 26900 -1000
rect 26840 -1260 26900 -1200
rect 27010 -1160 27070 -1100
rect 27010 -1360 27070 -1300
rect 27180 -1060 27240 -1000
rect 27180 -1260 27240 -1200
rect 27350 -1160 27410 -1100
rect 27350 -1360 27410 -1300
rect 27520 -1060 27580 -1000
rect 27520 -1260 27580 -1200
rect 27690 -1160 27750 -1100
rect 27690 -1360 27750 -1300
rect 27860 -1060 27920 -1000
rect 27860 -1260 27920 -1200
rect 28030 -1160 28090 -1100
rect 28030 -1360 28090 -1300
rect 28200 -1060 28260 -1000
rect 28200 -1260 28260 -1200
rect 28370 -1160 28430 -1100
rect 28370 -1360 28430 -1300
rect 28540 -1060 28600 -1000
rect 28540 -1260 28600 -1200
rect 28710 -1160 28770 -1100
rect 28710 -1360 28770 -1300
rect 28880 -1060 28940 -1000
rect 28880 -1260 28940 -1200
rect 29050 -1160 29110 -1100
rect 29050 -1360 29110 -1300
rect 29220 -1060 29280 -1000
rect 29220 -1260 29280 -1200
rect 29390 -1160 29450 -1100
rect 29390 -1360 29450 -1300
rect 29560 -1060 29620 -1000
rect 29560 -1260 29620 -1200
rect 29730 -1160 29790 -1100
rect 29730 -1360 29790 -1300
rect 29900 -1060 29960 -1000
rect 29900 -1260 29960 -1200
rect 30070 -1160 30130 -1100
rect 30070 -1360 30130 -1300
rect 30240 -1060 30300 -1000
rect 30240 -1260 30300 -1200
rect 30410 -1160 30470 -1100
rect 30410 -1360 30470 -1300
rect 30580 -1060 30640 -1000
rect 30580 -1260 30640 -1200
rect 30750 -1160 30810 -1100
rect 30750 -1360 30810 -1300
rect 30920 -1060 30980 -1000
rect 30920 -1260 30980 -1200
rect 31090 -1160 31150 -1100
rect 31090 -1360 31150 -1300
rect 31260 -1060 31320 -1000
rect 31260 -1260 31320 -1200
rect 31430 -1160 31490 -1100
rect 31430 -1360 31490 -1300
rect 31600 -1060 31660 -1000
rect 31600 -1260 31660 -1200
rect 31770 -1160 31830 -1100
rect 31770 -1360 31830 -1300
rect 31940 -1060 32000 -1000
rect 31940 -1260 32000 -1200
rect 32110 -1160 32170 -1100
rect 32110 -1360 32170 -1300
rect 32280 -1060 32340 -1000
rect 32280 -1260 32340 -1200
rect 32450 -1160 32510 -1100
rect 32450 -1360 32510 -1300
rect 32620 -1060 32680 -1000
rect 32620 -1260 32680 -1200
rect 32790 -1160 32850 -1100
rect 32790 -1360 32850 -1300
rect 32960 -1060 33020 -1000
rect 32960 -1260 33020 -1200
rect 33130 -1160 33190 -1100
rect 33130 -1360 33190 -1300
rect 33300 -1060 33360 -1000
rect 33300 -1260 33360 -1200
rect 33470 -1160 33530 -1100
rect 33470 -1360 33530 -1300
rect 33640 -1060 33700 -1000
rect 33640 -1260 33700 -1200
rect 33810 -1160 33870 -1100
rect 33810 -1360 33870 -1300
rect 33980 -1060 34040 -1000
rect 33980 -1260 34040 -1200
rect 34150 -1160 34210 -1100
rect 34150 -1360 34210 -1300
rect 34320 -1060 34380 -1000
rect 34320 -1260 34380 -1200
rect 34490 -1160 34550 -1100
rect 34490 -1360 34550 -1300
rect 34660 -1060 34720 -1000
rect 34660 -1260 34720 -1200
rect 34830 -1160 34890 -1100
rect 34830 -1360 34890 -1300
rect 35000 -1060 35060 -1000
rect 35000 -1260 35060 -1200
rect 35170 -1160 35230 -1100
rect 35170 -1360 35230 -1300
rect 35340 -1060 35400 -1000
rect 35340 -1260 35400 -1200
rect 35510 -1160 35570 -1100
rect 35510 -1360 35570 -1300
rect 35680 -1060 35740 -1000
rect 35680 -1260 35740 -1200
rect 35850 -1160 35910 -1100
rect 35850 -1360 35910 -1300
rect 36020 -1060 36080 -1000
rect 36020 -1260 36080 -1200
rect 36190 -1160 36250 -1100
rect 36190 -1360 36250 -1300
rect 36360 -1060 36420 -1000
rect 36360 -1260 36420 -1200
rect 36530 -1160 36590 -1100
rect 36530 -1360 36590 -1300
rect 36700 -1060 36760 -1000
rect 36700 -1260 36760 -1200
rect 36870 -1160 36930 -1100
rect 36870 -1360 36930 -1300
rect 37040 -1060 37100 -1000
rect 37040 -1260 37100 -1200
rect 37210 -1160 37270 -1100
rect 37210 -1360 37270 -1300
rect 37380 -1060 37440 -1000
rect 37380 -1260 37440 -1200
rect 37550 -1160 37610 -1100
rect 37550 -1360 37610 -1300
rect 37720 -1060 37780 -1000
rect 37720 -1260 37780 -1200
rect 37890 -1160 37950 -1100
rect 37890 -1360 37950 -1300
rect 38060 -1060 38120 -1000
rect 38060 -1260 38120 -1200
rect 38230 -1160 38290 -1100
rect 38230 -1360 38290 -1300
rect 38400 -1060 38460 -1000
rect 38400 -1260 38460 -1200
rect 38570 -1160 38630 -1100
rect 38570 -1360 38630 -1300
rect 38740 -1060 38800 -1000
rect 38740 -1260 38800 -1200
rect 38910 -1160 38970 -1100
rect 38910 -1360 38970 -1300
rect 39080 -1060 39140 -1000
rect 39080 -1260 39140 -1200
rect 39250 -1160 39310 -1100
rect 39250 -1360 39310 -1300
rect 39420 -1060 39480 -1000
rect 39420 -1260 39480 -1200
rect 39590 -1160 39650 -1100
rect 39590 -1360 39650 -1300
rect 39760 -1060 39820 -1000
rect 39760 -1260 39820 -1200
rect 39930 -1160 39990 -1100
rect 39930 -1360 39990 -1300
rect 40100 -1060 40160 -1000
rect 40100 -1260 40160 -1200
rect 40270 -1160 40330 -1100
rect 40270 -1360 40330 -1300
rect 40440 -1060 40500 -1000
rect 40440 -1260 40500 -1200
rect 40610 -1160 40670 -1100
rect 40610 -1360 40670 -1300
rect 40780 -1060 40840 -1000
rect 40780 -1260 40840 -1200
rect 40950 -1160 41010 -1100
rect 40950 -1360 41010 -1300
rect 41120 -1060 41180 -1000
rect 41120 -1260 41180 -1200
rect 41290 -1160 41350 -1100
rect 41290 -1360 41350 -1300
rect 41460 -1060 41520 -1000
rect 41460 -1260 41520 -1200
rect 41630 -1160 41690 -1100
rect 41630 -1360 41690 -1300
rect 41800 -1060 41860 -1000
rect 41800 -1260 41860 -1200
rect 41970 -1160 42030 -1100
rect 41970 -1360 42030 -1300
rect 42140 -1060 42200 -1000
rect 42140 -1260 42200 -1200
rect 42310 -1160 42370 -1100
rect 42310 -1360 42370 -1300
rect 42480 -1060 42540 -1000
rect 42480 -1260 42540 -1200
rect 42650 -1160 42710 -1100
rect 42650 -1360 42710 -1300
rect 42820 -1060 42880 -1000
rect 42820 -1260 42880 -1200
rect 42990 -1160 43050 -1100
rect 42990 -1360 43050 -1300
rect 43160 -1060 43220 -1000
rect 43160 -1260 43220 -1200
rect 43330 -1160 43390 -1100
rect 43330 -1360 43390 -1300
rect 43500 -1060 43560 -1000
rect 43500 -1260 43560 -1200
rect 43670 -1160 43730 -1100
rect 43670 -1360 43730 -1300
rect 43840 -1060 43900 -1000
rect 43840 -1260 43900 -1200
rect 44010 -1160 44070 -1100
rect 44010 -1360 44070 -1300
rect 44180 -1060 44240 -1000
rect 44180 -1260 44240 -1200
rect 44350 -1160 44410 -1100
rect 44350 -1360 44410 -1300
rect 44520 -1060 44580 -1000
rect 44520 -1260 44580 -1200
rect 44690 -1160 44750 -1100
rect 44690 -1360 44750 -1300
rect 44860 -1060 44920 -1000
rect 44860 -1260 44920 -1200
rect 45030 -1160 45090 -1100
rect 45030 -1360 45090 -1300
rect 45200 -1060 45260 -1000
rect 45200 -1260 45260 -1200
rect 45370 -1160 45430 -1100
rect 45370 -1360 45430 -1300
rect 45540 -1060 45600 -1000
rect 45540 -1260 45600 -1200
rect 45710 -1160 45770 -1100
rect 45710 -1360 45770 -1300
rect 45880 -1060 45940 -1000
rect 45880 -1260 45940 -1200
rect 46050 -1160 46110 -1100
rect 46050 -1360 46110 -1300
rect 46220 -1060 46280 -1000
rect 46220 -1260 46280 -1200
rect 46390 -1160 46450 -1100
rect 46390 -1360 46450 -1300
rect 46560 -1060 46620 -1000
rect 46560 -1260 46620 -1200
rect 46730 -1160 46790 -1100
rect 46730 -1360 46790 -1300
rect 46900 -1060 46960 -1000
rect 46900 -1260 46960 -1200
rect 47070 -1160 47130 -1100
rect 47070 -1360 47130 -1300
rect 47240 -1060 47300 -1000
rect 47240 -1260 47300 -1200
rect 47410 -1160 47470 -1100
rect 47410 -1360 47470 -1300
rect 47580 -1060 47640 -1000
rect 47580 -1260 47640 -1200
rect 47750 -1160 47810 -1100
rect 47750 -1360 47810 -1300
rect 47920 -1060 47980 -1000
rect 47920 -1260 47980 -1200
rect 48090 -1160 48150 -1100
rect 48090 -1360 48150 -1300
rect 48260 -1060 48320 -1000
rect 48260 -1260 48320 -1200
rect 48430 -1160 48490 -1100
rect 48430 -1360 48490 -1300
rect 48600 -1060 48660 -1000
rect 48600 -1260 48660 -1200
rect 48770 -1160 48830 -1100
rect 48770 -1360 48830 -1300
rect 48940 -1060 49000 -1000
rect 48940 -1260 49000 -1200
rect 49110 -1160 49170 -1100
rect 49110 -1360 49170 -1300
rect 49280 -1060 49340 -1000
rect 49280 -1260 49340 -1200
rect 49450 -1160 49510 -1100
rect 49450 -1360 49510 -1300
rect 49620 -1060 49680 -1000
rect 49620 -1260 49680 -1200
rect 49790 -1160 49850 -1100
rect 49790 -1360 49850 -1300
rect 49960 -1060 50020 -1000
rect 49960 -1260 50020 -1200
rect 50130 -1160 50190 -1100
rect 50130 -1360 50190 -1300
rect 50300 -1060 50360 -1000
rect 50300 -1260 50360 -1200
rect 50470 -1160 50530 -1100
rect 50470 -1360 50530 -1300
rect 50640 -1060 50700 -1000
rect 50640 -1260 50700 -1200
rect 50810 -1160 50870 -1100
rect 50810 -1360 50870 -1300
rect 50980 -1060 51040 -1000
rect 50980 -1260 51040 -1200
rect 51150 -1160 51210 -1100
rect 51150 -1360 51210 -1300
rect 51320 -1060 51380 -1000
rect 51320 -1260 51380 -1200
rect 51490 -1160 51550 -1100
rect 51490 -1360 51550 -1300
rect 51660 -1060 51720 -1000
rect 51660 -1260 51720 -1200
rect 51830 -1160 51890 -1100
rect 51830 -1360 51890 -1300
rect 52000 -1060 52060 -1000
rect 52000 -1260 52060 -1200
rect 52170 -1160 52230 -1100
rect 52170 -1360 52230 -1300
rect 52340 -1060 52400 -1000
rect 52340 -1260 52400 -1200
rect 52510 -1160 52570 -1100
rect 52510 -1360 52570 -1300
rect 52680 -1060 52740 -1000
rect 52680 -1260 52740 -1200
rect 52850 -1160 52910 -1100
rect 52850 -1360 52910 -1300
rect 53020 -1060 53080 -1000
rect 53020 -1260 53080 -1200
rect 53190 -1160 53250 -1100
rect 53190 -1360 53250 -1300
rect 53360 -1060 53420 -1000
rect 53360 -1260 53420 -1200
rect 53530 -1160 53590 -1100
rect 53530 -1360 53590 -1300
rect 53700 -1060 53760 -1000
rect 53700 -1260 53760 -1200
rect 53870 -1160 53930 -1100
rect 53870 -1360 53930 -1300
rect 54040 -1060 54100 -1000
rect 54040 -1260 54100 -1200
rect 54210 -1160 54270 -1100
rect 54210 -1360 54270 -1300
rect 54380 -1060 54440 -1000
rect 54380 -1260 54440 -1200
rect 54550 -1160 54610 -1100
rect 54550 -1360 54610 -1300
rect 54720 -1060 54780 -1000
rect 54720 -1260 54780 -1200
rect 54890 -1160 54950 -1100
rect 54890 -1360 54950 -1300
rect 55060 -1060 55120 -1000
rect 55060 -1260 55120 -1200
rect 55230 -1160 55290 -1100
rect 55230 -1360 55290 -1300
rect 55400 -1060 55460 -1000
rect 55400 -1260 55460 -1200
rect 55570 -1160 55630 -1100
rect 55570 -1360 55630 -1300
rect 55740 -1060 55800 -1000
rect 55740 -1260 55800 -1200
rect 55910 -1160 55970 -1100
rect 55910 -1360 55970 -1300
rect 56080 -1060 56140 -1000
rect 56080 -1260 56140 -1200
rect 56250 -1160 56310 -1100
rect 56250 -1360 56310 -1300
rect 56420 -1060 56480 -1000
rect 56420 -1260 56480 -1200
rect 56590 -1160 56650 -1100
rect 56590 -1360 56650 -1300
rect 56760 -1060 56820 -1000
rect 56760 -1260 56820 -1200
rect 56930 -1160 56990 -1100
rect 56930 -1360 56990 -1300
rect 57100 -1060 57160 -1000
rect 57100 -1260 57160 -1200
rect 57270 -1160 57330 -1100
rect 57270 -1360 57330 -1300
rect 57440 -1060 57500 -1000
rect 57440 -1260 57500 -1200
rect 57610 -1160 57670 -1100
rect 57610 -1360 57670 -1300
rect 57780 -1060 57840 -1000
rect 57780 -1260 57840 -1200
rect 57950 -1160 58010 -1100
rect 57950 -1360 58010 -1300
rect 58120 -1060 58180 -1000
rect 58120 -1260 58180 -1200
rect 58290 -1160 58350 -1100
rect 58290 -1360 58350 -1300
rect 58460 -1060 58520 -1000
rect 58460 -1260 58520 -1200
rect 58630 -1160 58690 -1100
rect 58630 -1360 58690 -1300
rect 58800 -1060 58860 -1000
rect 58800 -1260 58860 -1200
rect 58970 -1160 59030 -1100
rect 58970 -1360 59030 -1300
rect 59140 -1060 59200 -1000
rect 59140 -1260 59200 -1200
rect 59310 -1160 59370 -1100
rect 59310 -1360 59370 -1300
rect 59480 -1060 59540 -1000
rect 59480 -1260 59540 -1200
rect 59650 -1160 59710 -1100
rect 59650 -1360 59710 -1300
rect 59820 -1060 59880 -1000
rect 59820 -1260 59880 -1200
rect 59990 -1160 60050 -1100
rect 59990 -1360 60050 -1300
rect 60160 -1060 60220 -1000
rect 60160 -1260 60220 -1200
rect 60330 -1160 60390 -1100
rect 60330 -1360 60390 -1300
rect 60500 -1060 60560 -1000
rect 60500 -1260 60560 -1200
rect 60670 -1160 60730 -1100
rect 60670 -1360 60730 -1300
rect 60840 -1060 60900 -1000
rect 60840 -1260 60900 -1200
rect 61010 -1160 61070 -1100
rect 61010 -1360 61070 -1300
rect 61180 -1060 61240 -1000
rect 61180 -1260 61240 -1200
rect 61350 -1160 61410 -1100
rect 61350 -1360 61410 -1300
rect 61520 -1060 61580 -1000
rect 61520 -1260 61580 -1200
rect 61690 -1160 61750 -1100
rect 61690 -1360 61750 -1300
rect 61860 -1060 61920 -1000
rect 61860 -1260 61920 -1200
rect 62030 -1160 62090 -1100
rect 62030 -1360 62090 -1300
rect 62200 -1060 62260 -1000
rect 62200 -1260 62260 -1200
rect 62370 -1160 62430 -1100
rect 62370 -1360 62430 -1300
rect 62540 -1060 62600 -1000
rect 62540 -1260 62600 -1200
rect 62710 -1160 62770 -1100
rect 62710 -1360 62770 -1300
rect 62880 -1060 62940 -1000
rect 62880 -1260 62940 -1200
rect 63050 -1160 63110 -1100
rect 63050 -1360 63110 -1300
rect 63220 -1060 63280 -1000
rect 63220 -1260 63280 -1200
rect 63390 -1160 63450 -1100
rect 63390 -1360 63450 -1300
rect 63560 -1060 63620 -1000
rect 63560 -1260 63620 -1200
rect 63730 -1160 63790 -1100
rect 63730 -1360 63790 -1300
rect 63900 -1060 63960 -1000
rect 63900 -1260 63960 -1200
rect 64070 -1160 64130 -1100
rect 64070 -1360 64130 -1300
rect 64240 -1060 64300 -1000
rect 64240 -1260 64300 -1200
rect 64410 -1160 64470 -1100
rect 64410 -1360 64470 -1300
rect 64580 -1060 64640 -1000
rect 64580 -1260 64640 -1200
rect 64750 -1160 64810 -1100
rect 64750 -1360 64810 -1300
rect 64920 -1060 64980 -1000
rect 64920 -1260 64980 -1200
rect 65090 -1160 65150 -1100
rect 65090 -1360 65150 -1300
rect 65260 -1060 65320 -1000
rect 65260 -1260 65320 -1200
rect 65430 -1160 65490 -1100
rect 65430 -1360 65490 -1300
rect 65600 -1060 65660 -1000
rect 65600 -1260 65660 -1200
rect 65770 -1160 65830 -1100
rect 65770 -1360 65830 -1300
rect 65940 -1060 66000 -1000
rect 65940 -1260 66000 -1200
rect 66110 -1160 66170 -1100
rect 66110 -1360 66170 -1300
rect 66280 -1060 66340 -1000
rect 66280 -1260 66340 -1200
rect 66450 -1160 66510 -1100
rect 66450 -1360 66510 -1300
rect 66620 -1060 66680 -1000
rect 66620 -1260 66680 -1200
rect 66790 -1160 66850 -1100
rect 66790 -1360 66850 -1300
rect 66960 -1060 67020 -1000
rect 66960 -1260 67020 -1200
rect 67130 -1160 67190 -1100
rect 67130 -1360 67190 -1300
rect 67300 -1060 67360 -1000
rect 67300 -1260 67360 -1200
rect 67470 -1160 67530 -1100
rect 67470 -1360 67530 -1300
rect 67640 -1060 67700 -1000
rect 67640 -1260 67700 -1200
rect 67810 -1160 67870 -1100
rect 67810 -1360 67870 -1300
rect 67980 -1060 68040 -1000
rect 67980 -1260 68040 -1200
rect 68150 -1160 68210 -1100
rect 68150 -1360 68210 -1300
rect 68320 -1060 68380 -1000
rect 68320 -1260 68380 -1200
rect 68490 -1160 68550 -1100
rect 68490 -1360 68550 -1300
rect 68660 -1060 68720 -1000
rect 68660 -1260 68720 -1200
rect 68830 -1160 68890 -1100
rect 68830 -1360 68890 -1300
rect 69000 -1060 69060 -1000
rect 69000 -1260 69060 -1200
rect 69170 -1160 69230 -1100
rect 69170 -1360 69230 -1300
rect 69340 -1060 69400 -1000
rect 69340 -1260 69400 -1200
rect 69510 -1160 69570 -1100
rect 69510 -1360 69570 -1300
rect 69680 -1060 69740 -1000
rect 69680 -1260 69740 -1200
rect 69850 -1160 69910 -1100
rect 69850 -1360 69910 -1300
rect 70020 -1060 70080 -1000
rect 70020 -1260 70080 -1200
rect 70190 -1160 70250 -1100
rect 70190 -1360 70250 -1300
rect 70360 -1060 70420 -1000
rect 70360 -1260 70420 -1200
rect 70530 -1160 70590 -1100
rect 70530 -1360 70590 -1300
rect 70700 -1060 70760 -1000
rect 70700 -1260 70760 -1200
rect 70870 -1160 70930 -1100
rect 70870 -1360 70930 -1300
rect 71040 -1060 71100 -1000
rect 71040 -1260 71100 -1200
rect 71210 -1160 71270 -1100
rect 71210 -1360 71270 -1300
rect 71380 -1060 71440 -1000
rect 71380 -1260 71440 -1200
rect 71550 -1160 71610 -1100
rect 71550 -1360 71610 -1300
rect 71720 -1060 71780 -1000
rect 71720 -1260 71780 -1200
rect 71890 -1160 71950 -1100
rect 71890 -1360 71950 -1300
rect 72060 -1060 72120 -1000
rect 72060 -1260 72120 -1200
rect 72230 -1160 72290 -1100
rect 72230 -1360 72290 -1300
rect 72400 -1060 72460 -1000
rect 72400 -1260 72460 -1200
rect 72570 -1160 72630 -1100
rect 72570 -1360 72630 -1300
rect 72740 -1060 72800 -1000
rect 72740 -1260 72800 -1200
rect 72910 -1160 72970 -1100
rect 72910 -1360 72970 -1300
rect 73080 -1060 73140 -1000
rect 73080 -1260 73140 -1200
rect 73250 -1160 73310 -1100
rect 73250 -1360 73310 -1300
rect 73420 -1060 73480 -1000
rect 73420 -1260 73480 -1200
rect 73590 -1160 73650 -1100
rect 73590 -1360 73650 -1300
rect 73760 -1060 73820 -1000
rect 73760 -1260 73820 -1200
rect 73930 -1160 73990 -1100
rect 73930 -1360 73990 -1300
rect 74100 -1060 74160 -1000
rect 74100 -1260 74160 -1200
rect 74270 -1160 74330 -1100
rect 74270 -1360 74330 -1300
rect 74440 -1060 74500 -1000
rect 74440 -1260 74500 -1200
rect 74610 -1160 74670 -1100
rect 74610 -1360 74670 -1300
rect 74780 -1060 74840 -1000
rect 74780 -1260 74840 -1200
rect 74950 -1160 75010 -1100
rect 74950 -1360 75010 -1300
rect 75120 -1060 75180 -1000
rect 75120 -1260 75180 -1200
rect 75290 -1160 75350 -1100
rect 75290 -1360 75350 -1300
rect 75460 -1060 75520 -1000
rect 75460 -1260 75520 -1200
rect 75630 -1160 75690 -1100
rect 75630 -1360 75690 -1300
rect 75800 -1060 75860 -1000
rect 75800 -1260 75860 -1200
rect 75970 -1160 76030 -1100
rect 75970 -1360 76030 -1300
rect 76140 -1060 76200 -1000
rect 76140 -1260 76200 -1200
rect 76310 -1160 76370 -1100
rect 76310 -1360 76370 -1300
rect 76480 -1060 76540 -1000
rect 76480 -1260 76540 -1200
rect 76650 -1160 76710 -1100
rect 76650 -1360 76710 -1300
rect 76820 -1060 76880 -1000
rect 76820 -1260 76880 -1200
rect 76990 -1160 77050 -1100
rect 76990 -1360 77050 -1300
rect 77160 -1060 77220 -1000
rect 77160 -1260 77220 -1200
rect 77330 -1160 77390 -1100
rect 77330 -1360 77390 -1300
rect 77500 -1060 77560 -1000
rect 77500 -1260 77560 -1200
rect 77670 -1160 77730 -1100
rect 77670 -1360 77730 -1300
rect 77840 -1060 77900 -1000
rect 77840 -1260 77900 -1200
rect 78010 -1160 78070 -1100
rect 78010 -1360 78070 -1300
rect 78180 -1060 78240 -1000
rect 78180 -1260 78240 -1200
rect 78350 -1160 78410 -1100
rect 78350 -1360 78410 -1300
rect 78520 -1060 78580 -1000
rect 78520 -1260 78580 -1200
rect 78690 -1160 78750 -1100
rect 78690 -1360 78750 -1300
rect 78860 -1060 78920 -1000
rect 78860 -1260 78920 -1200
rect 79030 -1160 79090 -1100
rect 79030 -1360 79090 -1300
rect 79200 -1060 79260 -1000
rect 79200 -1260 79260 -1200
rect 79370 -1160 79430 -1100
rect 79370 -1360 79430 -1300
rect 79540 -1060 79600 -1000
rect 79540 -1260 79600 -1200
rect 79710 -1160 79770 -1100
rect 79710 -1360 79770 -1300
rect 79880 -1060 79940 -1000
rect 79880 -1260 79940 -1200
rect 80050 -1160 80110 -1100
rect 80050 -1360 80110 -1300
rect 80220 -1060 80280 -1000
rect 80220 -1260 80280 -1200
rect 80390 -1160 80450 -1100
rect 80390 -1360 80450 -1300
rect 80560 -1060 80620 -1000
rect 80560 -1260 80620 -1200
rect 80730 -1160 80790 -1100
rect 80730 -1360 80790 -1300
rect 80900 -1060 80960 -1000
rect 80900 -1260 80960 -1200
rect 81070 -1160 81130 -1100
rect 81070 -1360 81130 -1300
rect 81240 -1060 81300 -1000
rect 81240 -1260 81300 -1200
rect 81410 -1160 81470 -1100
rect 81410 -1360 81470 -1300
rect 81580 -1060 81640 -1000
rect 81580 -1260 81640 -1200
rect 81750 -1160 81810 -1100
rect 81750 -1360 81810 -1300
rect 81920 -1060 81980 -1000
rect 81920 -1260 81980 -1200
rect 82090 -1160 82150 -1100
rect 82090 -1360 82150 -1300
rect 82260 -1060 82320 -1000
rect 82260 -1260 82320 -1200
rect 82430 -1160 82490 -1100
rect 82430 -1360 82490 -1300
rect 82600 -1060 82660 -1000
rect 82600 -1260 82660 -1200
rect 82770 -1160 82830 -1100
rect 82770 -1360 82830 -1300
rect 82940 -1060 83000 -1000
rect 82940 -1260 83000 -1200
rect 83110 -1160 83170 -1100
rect 83110 -1360 83170 -1300
rect 83280 -1060 83340 -1000
rect 83280 -1260 83340 -1200
rect 83450 -1160 83510 -1100
rect 83450 -1360 83510 -1300
rect 83620 -1060 83680 -1000
rect 83620 -1260 83680 -1200
rect 83790 -1160 83850 -1100
rect 83790 -1360 83850 -1300
rect 83960 -1060 84020 -1000
rect 83960 -1260 84020 -1200
rect 84130 -1160 84190 -1100
rect 84130 -1360 84190 -1300
rect 84300 -1060 84360 -1000
rect 84300 -1260 84360 -1200
rect 84470 -1160 84530 -1100
rect 84470 -1360 84530 -1300
rect 84640 -1060 84700 -1000
rect 84640 -1260 84700 -1200
rect 84810 -1160 84870 -1100
rect 84810 -1360 84870 -1300
rect 84980 -1060 85040 -1000
rect 84980 -1260 85040 -1200
rect 85150 -1160 85210 -1100
rect 85150 -1360 85210 -1300
rect 85320 -1060 85380 -1000
rect 85320 -1260 85380 -1200
rect 85490 -1160 85550 -1100
rect 85490 -1360 85550 -1300
rect 85660 -1060 85720 -1000
rect 85660 -1260 85720 -1200
rect 85830 -1160 85890 -1100
rect 85830 -1360 85890 -1300
rect 86000 -1060 86060 -1000
rect 86000 -1260 86060 -1200
rect 86170 -1160 86230 -1100
rect 86170 -1360 86230 -1300
rect 86340 -1060 86400 -1000
rect 86340 -1260 86400 -1200
rect 86510 -1160 86570 -1100
rect 86510 -1360 86570 -1300
rect 86680 -1060 86740 -1000
rect 86680 -1260 86740 -1200
rect 86850 -1160 86910 -1100
rect 86850 -1360 86910 -1300
rect 87020 -1060 87080 -1000
rect 87020 -1260 87080 -1200
rect 87190 -1160 87250 -1100
rect 87190 -1360 87250 -1300
rect 830 -1540 910 -1470
rect 5000 -1540 5080 -1470
rect 9030 -1540 9110 -1470
rect 13060 -1540 13140 -1470
rect 17100 -1540 17180 -1470
rect 21200 -1540 21280 -1470
rect 25310 -1540 25390 -1470
rect 29410 -1540 29490 -1470
rect 33440 -1540 33520 -1470
rect 37550 -1540 37630 -1470
rect 41650 -1540 41730 -1470
rect 47100 -1540 47180 -1470
rect 51180 -1540 51260 -1470
rect 55290 -1540 55370 -1470
rect 59320 -1540 59400 -1470
rect 63420 -1540 63500 -1470
rect 67530 -1540 67610 -1470
rect 71560 -1540 71640 -1470
rect 75810 -1540 75890 -1470
rect 79770 -1540 79850 -1470
rect 83950 -1540 84030 -1470
rect 86508 -1544 86588 -1474
<< metal1 >>
rect 540 1001 580 1010
rect 1310 1001 1350 1010
rect 531 995 629 1001
rect 531 935 543 995
rect 617 935 629 995
rect 531 929 629 935
rect 1259 995 1357 1001
rect 1259 935 1271 995
rect 1345 935 1357 995
rect 5660 979 5700 990
rect 6430 979 6470 990
rect 1259 929 1357 935
rect 5651 973 5749 979
rect 540 710 580 929
rect 1310 730 1350 929
rect 5651 913 5663 973
rect 5737 913 5749 973
rect 5651 907 5749 913
rect 6379 973 6477 979
rect 6379 913 6391 973
rect 6465 913 6477 973
rect 6379 907 6477 913
rect 1280 710 1410 730
rect 5660 710 5700 907
rect 6430 710 6470 907
rect 500 690 630 710
rect 500 630 520 690
rect 610 630 630 690
rect 1280 650 1300 710
rect 1390 650 1410 710
rect 1280 630 1410 650
rect 5610 690 5740 710
rect 5610 630 5630 690
rect 5720 630 5740 690
rect 500 610 630 630
rect 730 590 930 620
rect 730 520 790 590
rect 870 520 930 590
rect 730 490 930 520
rect 2110 590 2310 620
rect 2110 520 2170 590
rect 2250 520 2310 590
rect 2110 490 2310 520
rect 3490 590 3690 620
rect 3490 520 3550 590
rect 3630 520 3690 590
rect 3490 490 3690 520
rect 5150 590 5350 620
rect 5610 610 5740 630
rect 6370 690 6510 710
rect 6370 630 6390 690
rect 6490 630 6510 690
rect 6370 610 6510 630
rect 5150 520 5210 590
rect 5290 520 5350 590
rect 5150 490 5350 520
rect 7980 590 8180 620
rect 7980 520 8040 590
rect 8120 520 8180 590
rect 7980 490 8180 520
rect 10740 590 10940 620
rect 10740 520 10800 590
rect 10880 520 10940 590
rect 10740 490 10940 520
rect 13370 590 13570 620
rect 13370 520 13430 590
rect 13510 520 13570 590
rect 13370 490 13570 520
rect 16410 590 16610 620
rect 16410 520 16470 590
rect 16550 520 16610 590
rect 16410 490 16610 520
rect 20480 590 20680 620
rect 20480 520 20540 590
rect 20620 520 20680 590
rect 20480 490 20680 520
rect 24620 590 24820 620
rect 24620 520 24680 590
rect 24760 520 24820 590
rect 24620 490 24820 520
rect 28700 590 28900 620
rect 28700 520 28760 590
rect 28840 520 28900 590
rect 28700 490 28900 520
rect 32850 590 33050 620
rect 32850 520 32910 590
rect 32990 520 33050 590
rect 32850 490 33050 520
rect 36720 590 36920 620
rect 36720 520 36780 590
rect 36860 520 36920 590
rect 36720 490 36920 520
rect 40860 590 41060 620
rect 40860 520 40920 590
rect 41000 520 41060 590
rect 40860 490 41060 520
rect 44850 590 45050 620
rect 44850 520 44910 590
rect 44990 520 45050 590
rect 44850 490 45050 520
rect 48930 590 49130 620
rect 48930 520 48990 590
rect 49070 520 49130 590
rect 48930 490 49130 520
rect 53020 590 53220 620
rect 53020 520 53080 590
rect 53160 520 53220 590
rect 53020 490 53220 520
rect 57180 590 57380 620
rect 57180 520 57240 590
rect 57320 520 57380 590
rect 57180 490 57380 520
rect 10 410 110 430
rect 10 350 30 410
rect 90 350 110 410
rect 10 330 110 350
rect 180 410 280 430
rect 180 350 200 410
rect 260 350 280 410
rect 180 310 280 350
rect 430 410 530 430
rect 430 350 450 410
rect 510 350 530 410
rect 430 330 530 350
rect 770 410 870 430
rect 770 350 790 410
rect 850 350 870 410
rect 770 330 870 350
rect 1110 410 1210 430
rect 1110 350 1130 410
rect 1190 350 1210 410
rect 1110 330 1210 350
rect 1500 410 1600 430
rect 1500 350 1520 410
rect 1580 350 1600 410
rect 1500 330 1600 350
rect 1840 410 1940 430
rect 1840 350 1860 410
rect 1920 350 1940 410
rect 1840 330 1940 350
rect 2180 410 2280 430
rect 2180 350 2200 410
rect 2260 350 2280 410
rect 2180 330 2280 350
rect 2520 410 2620 430
rect 2520 350 2540 410
rect 2600 350 2620 410
rect 2520 330 2620 350
rect 2860 410 2960 430
rect 2860 350 2880 410
rect 2940 350 2960 410
rect 2860 330 2960 350
rect 3200 410 3300 430
rect 3200 350 3220 410
rect 3280 350 3300 410
rect 3200 330 3300 350
rect 3540 410 3640 430
rect 3540 350 3560 410
rect 3620 350 3640 410
rect 3540 330 3640 350
rect 3880 410 3980 430
rect 3880 350 3900 410
rect 3960 350 3980 410
rect 3880 330 3980 350
rect 4220 410 4320 430
rect 4220 350 4240 410
rect 4300 350 4320 410
rect 4220 330 4320 350
rect 4520 410 4620 430
rect 4520 350 4540 410
rect 4600 350 4620 410
rect 4520 330 4620 350
rect 4860 410 4960 430
rect 4860 350 4880 410
rect 4940 350 4960 410
rect 4860 330 4960 350
rect 5200 410 5300 430
rect 5200 350 5220 410
rect 5280 350 5300 410
rect 5200 330 5300 350
rect 5540 410 5640 430
rect 5540 350 5560 410
rect 5620 350 5640 410
rect 5540 330 5640 350
rect 5880 410 5980 430
rect 5880 350 5900 410
rect 5960 350 5980 410
rect 5880 330 5980 350
rect 6220 410 6320 430
rect 6220 350 6240 410
rect 6300 350 6320 410
rect 6220 330 6320 350
rect 6560 410 6660 430
rect 6560 350 6580 410
rect 6640 350 6660 410
rect 6560 330 6660 350
rect 6900 410 7000 430
rect 6900 350 6920 410
rect 6980 350 7000 410
rect 6900 330 7000 350
rect 7240 410 7340 430
rect 7240 350 7260 410
rect 7320 350 7340 410
rect 7240 330 7340 350
rect 7580 410 7680 430
rect 7580 350 7600 410
rect 7660 350 7680 410
rect 7580 330 7680 350
rect 7920 410 8020 430
rect 7920 350 7940 410
rect 8000 350 8020 410
rect 7920 330 8020 350
rect 8260 410 8360 430
rect 8260 350 8280 410
rect 8340 350 8360 410
rect 8260 330 8360 350
rect 8600 410 8700 430
rect 8600 350 8620 410
rect 8680 350 8700 410
rect 8600 330 8700 350
rect 8940 410 9040 430
rect 8940 350 8960 410
rect 9020 350 9040 410
rect 8940 330 9040 350
rect 9280 410 9380 430
rect 9280 350 9300 410
rect 9360 350 9380 410
rect 9280 330 9380 350
rect 9620 410 9720 430
rect 9620 350 9640 410
rect 9700 350 9720 410
rect 9620 330 9720 350
rect 9960 410 10060 430
rect 9960 350 9980 410
rect 10040 350 10060 410
rect 9960 330 10060 350
rect 10300 410 10400 430
rect 10300 350 10320 410
rect 10380 350 10400 410
rect 10300 330 10400 350
rect 10640 410 10740 430
rect 10640 350 10660 410
rect 10720 350 10740 410
rect 10640 330 10740 350
rect 10980 410 11080 430
rect 10980 350 11000 410
rect 11060 350 11080 410
rect 10980 330 11080 350
rect 11320 410 11420 430
rect 11320 350 11340 410
rect 11400 350 11420 410
rect 11320 330 11420 350
rect 11660 410 11760 430
rect 11660 350 11680 410
rect 11740 350 11760 410
rect 11660 330 11760 350
rect 12000 410 12100 430
rect 12000 350 12020 410
rect 12080 350 12100 410
rect 12000 330 12100 350
rect 12340 410 12440 430
rect 12340 350 12360 410
rect 12420 350 12440 410
rect 12340 330 12440 350
rect 12680 410 12780 430
rect 12680 350 12700 410
rect 12760 350 12780 410
rect 12680 330 12780 350
rect 13020 410 13120 430
rect 13020 350 13040 410
rect 13100 350 13120 410
rect 13020 330 13120 350
rect 13360 410 13460 430
rect 13360 350 13380 410
rect 13440 350 13460 410
rect 13360 330 13460 350
rect 13700 410 13800 430
rect 13700 350 13720 410
rect 13780 350 13800 410
rect 13700 330 13800 350
rect 14040 410 14140 430
rect 14040 350 14060 410
rect 14120 350 14140 410
rect 14040 330 14140 350
rect 14380 410 14480 430
rect 14380 350 14400 410
rect 14460 350 14480 410
rect 14380 330 14480 350
rect 14720 410 14820 430
rect 14720 350 14740 410
rect 14800 350 14820 410
rect 14720 330 14820 350
rect 15060 410 15160 430
rect 15060 350 15080 410
rect 15140 350 15160 410
rect 15060 330 15160 350
rect 15400 410 15500 430
rect 15400 350 15420 410
rect 15480 350 15500 410
rect 15400 330 15500 350
rect 15700 410 15800 430
rect 15700 350 15720 410
rect 15780 350 15800 410
rect 15700 330 15800 350
rect 16040 410 16140 430
rect 16040 350 16060 410
rect 16120 350 16140 410
rect 16040 330 16140 350
rect 16380 410 16480 430
rect 16380 350 16400 410
rect 16460 350 16480 410
rect 16380 330 16480 350
rect 16720 410 16820 430
rect 16720 350 16740 410
rect 16800 350 16820 410
rect 16720 330 16820 350
rect 17060 410 17160 430
rect 17060 350 17080 410
rect 17140 350 17160 410
rect 17060 330 17160 350
rect 17400 410 17500 430
rect 17400 350 17420 410
rect 17480 350 17500 410
rect 17400 330 17500 350
rect 17740 410 17840 430
rect 17740 350 17760 410
rect 17820 350 17840 410
rect 17740 330 17840 350
rect 18080 410 18180 430
rect 18080 350 18100 410
rect 18160 350 18180 410
rect 18080 330 18180 350
rect 18420 410 18520 430
rect 18420 350 18440 410
rect 18500 350 18520 410
rect 18420 330 18520 350
rect 18760 410 18860 430
rect 18760 350 18780 410
rect 18840 350 18860 410
rect 18760 330 18860 350
rect 19100 410 19200 430
rect 19100 350 19120 410
rect 19180 350 19200 410
rect 19100 330 19200 350
rect 19440 410 19540 430
rect 19440 350 19460 410
rect 19520 350 19540 410
rect 19440 330 19540 350
rect 19780 410 19880 430
rect 19780 350 19800 410
rect 19860 350 19880 410
rect 19780 330 19880 350
rect 20120 410 20220 430
rect 20120 350 20140 410
rect 20200 350 20220 410
rect 20120 330 20220 350
rect 20460 410 20560 430
rect 20460 350 20480 410
rect 20540 350 20560 410
rect 20460 330 20560 350
rect 20800 410 20900 430
rect 20800 350 20820 410
rect 20880 350 20900 410
rect 20800 330 20900 350
rect 21140 410 21240 430
rect 21140 350 21160 410
rect 21220 350 21240 410
rect 21140 330 21240 350
rect 21480 410 21580 430
rect 21480 350 21500 410
rect 21560 350 21580 410
rect 21480 330 21580 350
rect 21820 410 21920 430
rect 21820 350 21840 410
rect 21900 350 21920 410
rect 21820 330 21920 350
rect 22160 410 22260 430
rect 22160 350 22180 410
rect 22240 350 22260 410
rect 22160 330 22260 350
rect 22500 410 22600 430
rect 22500 350 22520 410
rect 22580 350 22600 410
rect 22500 330 22600 350
rect 22840 410 22940 430
rect 22840 350 22860 410
rect 22920 350 22940 410
rect 22840 330 22940 350
rect 23180 410 23280 430
rect 23180 350 23200 410
rect 23260 350 23280 410
rect 23180 330 23280 350
rect 23520 410 23620 430
rect 23520 350 23540 410
rect 23600 350 23620 410
rect 23520 330 23620 350
rect 23860 410 23960 430
rect 23860 350 23880 410
rect 23940 350 23960 410
rect 23860 330 23960 350
rect 24200 410 24300 430
rect 24200 350 24220 410
rect 24280 350 24300 410
rect 24200 330 24300 350
rect 24540 410 24640 430
rect 24540 350 24560 410
rect 24620 350 24640 410
rect 24540 330 24640 350
rect 24880 410 24980 430
rect 24880 350 24900 410
rect 24960 350 24980 410
rect 24880 330 24980 350
rect 25220 410 25320 430
rect 25220 350 25240 410
rect 25300 350 25320 410
rect 25220 330 25320 350
rect 25560 410 25660 430
rect 25560 350 25580 410
rect 25640 350 25660 410
rect 25560 330 25660 350
rect 25900 410 26000 430
rect 25900 350 25920 410
rect 25980 350 26000 410
rect 25900 330 26000 350
rect 26240 410 26340 430
rect 26240 350 26260 410
rect 26320 350 26340 410
rect 26240 330 26340 350
rect 26580 410 26680 430
rect 26580 350 26600 410
rect 26660 350 26680 410
rect 26580 330 26680 350
rect 26920 410 27020 430
rect 26920 350 26940 410
rect 27000 350 27020 410
rect 26920 330 27020 350
rect 27260 410 27360 430
rect 27260 350 27280 410
rect 27340 350 27360 410
rect 27260 330 27360 350
rect 27600 410 27700 430
rect 27600 350 27620 410
rect 27680 350 27700 410
rect 27600 330 27700 350
rect 27940 410 28040 430
rect 27940 350 27960 410
rect 28020 350 28040 410
rect 27940 330 28040 350
rect 28280 410 28380 430
rect 28280 350 28300 410
rect 28360 350 28380 410
rect 28280 330 28380 350
rect 28620 410 28720 430
rect 28620 350 28640 410
rect 28700 350 28720 410
rect 28620 330 28720 350
rect 28960 410 29060 430
rect 28960 350 28980 410
rect 29040 350 29060 410
rect 28960 330 29060 350
rect 29300 410 29400 430
rect 29300 350 29320 410
rect 29380 350 29400 410
rect 29300 330 29400 350
rect 29640 410 29740 430
rect 29640 350 29660 410
rect 29720 350 29740 410
rect 29640 330 29740 350
rect 29980 410 30080 430
rect 29980 350 30000 410
rect 30060 350 30080 410
rect 29980 330 30080 350
rect 30320 410 30420 430
rect 30320 350 30340 410
rect 30400 350 30420 410
rect 30320 330 30420 350
rect 30660 410 30760 430
rect 30660 350 30680 410
rect 30740 350 30760 410
rect 30660 330 30760 350
rect 31000 410 31100 430
rect 31000 350 31020 410
rect 31080 350 31100 410
rect 31000 330 31100 350
rect 31340 410 31440 430
rect 31340 350 31360 410
rect 31420 350 31440 410
rect 31340 330 31440 350
rect 31680 410 31780 430
rect 31680 350 31700 410
rect 31760 350 31780 410
rect 31680 330 31780 350
rect 32020 410 32120 430
rect 32020 350 32040 410
rect 32100 350 32120 410
rect 32020 330 32120 350
rect 32360 410 32460 430
rect 32360 350 32380 410
rect 32440 350 32460 410
rect 32360 330 32460 350
rect 32700 410 32800 430
rect 32700 350 32720 410
rect 32780 350 32800 410
rect 32700 330 32800 350
rect 33040 410 33140 430
rect 33040 350 33060 410
rect 33120 350 33140 410
rect 33040 330 33140 350
rect 33380 410 33480 430
rect 33380 350 33400 410
rect 33460 350 33480 410
rect 33380 330 33480 350
rect 33720 410 33820 430
rect 33720 350 33740 410
rect 33800 350 33820 410
rect 33720 330 33820 350
rect 34060 410 34160 430
rect 34060 350 34080 410
rect 34140 350 34160 410
rect 34060 330 34160 350
rect 34400 410 34500 430
rect 34400 350 34420 410
rect 34480 350 34500 410
rect 34400 330 34500 350
rect 34740 410 34840 430
rect 34740 350 34760 410
rect 34820 350 34840 410
rect 34740 330 34840 350
rect 35080 410 35180 430
rect 35080 350 35100 410
rect 35160 350 35180 410
rect 35080 330 35180 350
rect 35420 410 35520 430
rect 35420 350 35440 410
rect 35500 350 35520 410
rect 35420 330 35520 350
rect 35760 410 35860 430
rect 35760 350 35780 410
rect 35840 350 35860 410
rect 35760 330 35860 350
rect 36100 410 36200 430
rect 36100 350 36120 410
rect 36180 350 36200 410
rect 36100 330 36200 350
rect 36440 410 36540 430
rect 36440 350 36460 410
rect 36520 350 36540 410
rect 36440 330 36540 350
rect 36780 410 36880 430
rect 36780 350 36800 410
rect 36860 350 36880 410
rect 36780 330 36880 350
rect 37120 410 37220 430
rect 37120 350 37140 410
rect 37200 350 37220 410
rect 37120 330 37220 350
rect 37460 410 37560 430
rect 37460 350 37480 410
rect 37540 350 37560 410
rect 37460 330 37560 350
rect 37800 410 37900 430
rect 37800 350 37820 410
rect 37880 350 37900 410
rect 37800 330 37900 350
rect 38140 410 38240 430
rect 38140 350 38160 410
rect 38220 350 38240 410
rect 38140 330 38240 350
rect 38480 410 38580 430
rect 38480 350 38500 410
rect 38560 350 38580 410
rect 38480 330 38580 350
rect 38820 410 38920 430
rect 38820 350 38840 410
rect 38900 350 38920 410
rect 38820 330 38920 350
rect 39160 410 39260 430
rect 39160 350 39180 410
rect 39240 350 39260 410
rect 39160 330 39260 350
rect 39500 410 39600 430
rect 39500 350 39520 410
rect 39580 350 39600 410
rect 39500 330 39600 350
rect 39840 410 39940 430
rect 39840 350 39860 410
rect 39920 350 39940 410
rect 39840 330 39940 350
rect 40180 410 40280 430
rect 40180 350 40200 410
rect 40260 350 40280 410
rect 40180 330 40280 350
rect 40520 410 40620 430
rect 40520 350 40540 410
rect 40600 350 40620 410
rect 40520 330 40620 350
rect 40860 410 40960 430
rect 40860 350 40880 410
rect 40940 350 40960 410
rect 40860 330 40960 350
rect 41200 410 41300 430
rect 41200 350 41220 410
rect 41280 350 41300 410
rect 41200 330 41300 350
rect 41540 410 41640 430
rect 41540 350 41560 410
rect 41620 350 41640 410
rect 41540 330 41640 350
rect 41880 410 41980 430
rect 41880 350 41900 410
rect 41960 350 41980 410
rect 41880 330 41980 350
rect 42220 410 42320 430
rect 42220 350 42240 410
rect 42300 350 42320 410
rect 42220 330 42320 350
rect 42560 410 42660 430
rect 42560 350 42580 410
rect 42640 350 42660 410
rect 42560 330 42660 350
rect 42900 410 43000 430
rect 42900 350 42920 410
rect 42980 350 43000 410
rect 42900 330 43000 350
rect 43240 410 43340 430
rect 43240 350 43260 410
rect 43320 350 43340 410
rect 43240 330 43340 350
rect 43580 410 43680 430
rect 43580 350 43600 410
rect 43660 350 43680 410
rect 43580 330 43680 350
rect 43920 410 44020 430
rect 43920 350 43940 410
rect 44000 350 44020 410
rect 43920 330 44020 350
rect 44260 410 44360 430
rect 44260 350 44280 410
rect 44340 350 44360 410
rect 44260 330 44360 350
rect 44600 410 44700 430
rect 44600 350 44620 410
rect 44680 350 44700 410
rect 44600 330 44700 350
rect 44940 410 45040 430
rect 44940 350 44960 410
rect 45020 350 45040 410
rect 44940 330 45040 350
rect 45280 410 45380 430
rect 45280 350 45300 410
rect 45360 350 45380 410
rect 45280 330 45380 350
rect 45620 410 45720 430
rect 45620 350 45640 410
rect 45700 350 45720 410
rect 45620 330 45720 350
rect 45960 410 46060 430
rect 45960 350 45980 410
rect 46040 350 46060 410
rect 45960 330 46060 350
rect 46300 410 46400 430
rect 46300 350 46320 410
rect 46380 350 46400 410
rect 46300 330 46400 350
rect 46640 410 46740 430
rect 46640 350 46660 410
rect 46720 350 46740 410
rect 46640 330 46740 350
rect 46980 410 47080 430
rect 46980 350 47000 410
rect 47060 350 47080 410
rect 46980 330 47080 350
rect 47320 410 47420 430
rect 47320 350 47340 410
rect 47400 350 47420 410
rect 47320 330 47420 350
rect 47660 410 47760 430
rect 47660 350 47680 410
rect 47740 350 47760 410
rect 47660 330 47760 350
rect 48000 410 48100 430
rect 48000 350 48020 410
rect 48080 350 48100 410
rect 48000 330 48100 350
rect 48340 410 48440 430
rect 48340 350 48360 410
rect 48420 350 48440 410
rect 48340 330 48440 350
rect 48680 410 48780 430
rect 48680 350 48700 410
rect 48760 350 48780 410
rect 48680 330 48780 350
rect 49020 410 49120 430
rect 49020 350 49040 410
rect 49100 350 49120 410
rect 49020 330 49120 350
rect 49360 410 49460 430
rect 49360 350 49380 410
rect 49440 350 49460 410
rect 49360 330 49460 350
rect 49700 410 49800 430
rect 49700 350 49720 410
rect 49780 350 49800 410
rect 49700 330 49800 350
rect 50040 410 50140 430
rect 50040 350 50060 410
rect 50120 350 50140 410
rect 50040 330 50140 350
rect 50380 410 50480 430
rect 50380 350 50400 410
rect 50460 350 50480 410
rect 50380 330 50480 350
rect 50720 410 50820 430
rect 50720 350 50740 410
rect 50800 350 50820 410
rect 50720 330 50820 350
rect 51060 410 51160 430
rect 51060 350 51080 410
rect 51140 350 51160 410
rect 51060 330 51160 350
rect 51400 410 51500 430
rect 51400 350 51420 410
rect 51480 350 51500 410
rect 51400 330 51500 350
rect 51740 410 51840 430
rect 51740 350 51760 410
rect 51820 350 51840 410
rect 51740 330 51840 350
rect 52080 410 52180 430
rect 52080 350 52100 410
rect 52160 350 52180 410
rect 52080 330 52180 350
rect 52420 410 52520 430
rect 52420 350 52440 410
rect 52500 350 52520 410
rect 52420 330 52520 350
rect 52760 410 52860 430
rect 52760 350 52780 410
rect 52840 350 52860 410
rect 52760 330 52860 350
rect 53100 410 53200 430
rect 53100 350 53120 410
rect 53180 350 53200 410
rect 53100 330 53200 350
rect 53440 410 53540 430
rect 53440 350 53460 410
rect 53520 350 53540 410
rect 53440 330 53540 350
rect 53780 410 53880 430
rect 53780 350 53800 410
rect 53860 350 53880 410
rect 53780 330 53880 350
rect 54120 410 54220 430
rect 54120 350 54140 410
rect 54200 350 54220 410
rect 54120 330 54220 350
rect 54460 410 54560 430
rect 54460 350 54480 410
rect 54540 350 54560 410
rect 54460 330 54560 350
rect 54800 410 54900 430
rect 54800 350 54820 410
rect 54880 350 54900 410
rect 54800 330 54900 350
rect 55140 410 55240 430
rect 55140 350 55160 410
rect 55220 350 55240 410
rect 55140 330 55240 350
rect 55480 410 55580 430
rect 55480 350 55500 410
rect 55560 350 55580 410
rect 55480 330 55580 350
rect 55820 410 55920 430
rect 55820 350 55840 410
rect 55900 350 55920 410
rect 55820 330 55920 350
rect 56160 410 56260 430
rect 56160 350 56180 410
rect 56240 350 56260 410
rect 56160 330 56260 350
rect 56500 410 56600 430
rect 56500 350 56520 410
rect 56580 350 56600 410
rect 56500 330 56600 350
rect 56840 410 56940 430
rect 56840 350 56860 410
rect 56920 350 56940 410
rect 56840 330 56940 350
rect 57180 410 57280 430
rect 57180 350 57200 410
rect 57260 350 57280 410
rect 57180 330 57280 350
rect 57520 410 57620 430
rect 57520 350 57540 410
rect 57600 350 57620 410
rect 57520 330 57620 350
rect 57860 410 57960 430
rect 57860 350 57880 410
rect 57940 350 57960 410
rect 57860 330 57960 350
rect 58200 410 58300 430
rect 58200 350 58220 410
rect 58280 350 58300 410
rect 58200 330 58300 350
rect 58540 410 58640 430
rect 58540 350 58560 410
rect 58620 350 58640 410
rect 58540 330 58640 350
rect 58880 410 58980 430
rect 58880 350 58900 410
rect 58960 350 58980 410
rect 58880 330 58980 350
rect 59220 410 59320 430
rect 59220 350 59240 410
rect 59300 350 59320 410
rect 59220 330 59320 350
rect 180 250 200 310
rect 260 250 280 310
rect 50 110 150 130
rect 50 30 70 110
rect 130 30 150 110
rect 50 10 150 30
rect 10 -60 110 -40
rect 10 -120 30 -60
rect 90 -120 110 -60
rect 10 -140 110 -120
rect 180 -60 280 250
rect 600 310 700 320
rect 600 250 620 310
rect 680 250 700 310
rect 600 200 700 250
rect 600 130 620 200
rect 680 130 700 200
rect 430 80 530 100
rect 430 20 450 80
rect 510 20 530 80
rect 430 0 530 20
rect 600 80 700 130
rect 940 310 1040 320
rect 940 250 960 310
rect 1020 250 1040 310
rect 940 200 1040 250
rect 940 130 960 200
rect 1020 130 1040 200
rect 600 20 620 80
rect 680 20 700 80
rect 600 0 700 20
rect 770 80 870 100
rect 770 20 790 80
rect 850 20 870 80
rect 770 0 870 20
rect 940 80 1040 130
rect 1670 310 1770 320
rect 1670 250 1690 310
rect 1750 250 1770 310
rect 1670 200 1770 250
rect 1670 130 1690 200
rect 1750 130 1770 200
rect 940 20 960 80
rect 1020 20 1040 80
rect 940 0 1040 20
rect 1110 80 1210 100
rect 1110 20 1130 80
rect 1190 20 1210 80
rect 1110 0 1210 20
rect 1500 80 1600 100
rect 1500 20 1520 80
rect 1580 20 1600 80
rect 1500 0 1600 20
rect 1670 80 1770 130
rect 2010 310 2110 320
rect 2010 250 2030 310
rect 2090 250 2110 310
rect 2010 200 2110 250
rect 2010 130 2030 200
rect 2090 130 2110 200
rect 1670 20 1690 80
rect 1750 20 1770 80
rect 1670 0 1770 20
rect 1840 80 1940 100
rect 1840 20 1860 80
rect 1920 20 1940 80
rect 1840 0 1940 20
rect 2010 80 2110 130
rect 2350 310 2450 320
rect 2350 250 2370 310
rect 2430 250 2450 310
rect 2350 200 2450 250
rect 2350 130 2370 200
rect 2430 130 2450 200
rect 2010 20 2030 80
rect 2090 20 2110 80
rect 2010 0 2110 20
rect 2180 80 2280 100
rect 2180 20 2200 80
rect 2260 20 2280 80
rect 2180 0 2280 20
rect 2350 80 2450 130
rect 2690 310 2790 320
rect 2690 250 2710 310
rect 2770 250 2790 310
rect 2690 200 2790 250
rect 2690 130 2710 200
rect 2770 130 2790 200
rect 2350 20 2370 80
rect 2430 20 2450 80
rect 2350 0 2450 20
rect 2520 80 2620 100
rect 2520 20 2540 80
rect 2600 20 2620 80
rect 2520 0 2620 20
rect 2690 80 2790 130
rect 3030 310 3130 320
rect 3030 250 3050 310
rect 3110 250 3130 310
rect 3030 200 3130 250
rect 3030 130 3050 200
rect 3110 130 3130 200
rect 2690 20 2710 80
rect 2770 20 2790 80
rect 2690 0 2790 20
rect 2860 80 2960 100
rect 2860 20 2880 80
rect 2940 20 2960 80
rect 2860 0 2960 20
rect 3030 80 3130 130
rect 3370 310 3470 320
rect 3370 250 3390 310
rect 3450 250 3470 310
rect 3370 200 3470 250
rect 3370 130 3390 200
rect 3450 130 3470 200
rect 3030 20 3050 80
rect 3110 20 3130 80
rect 3030 0 3130 20
rect 3200 80 3300 100
rect 3200 20 3220 80
rect 3280 20 3300 80
rect 3200 0 3300 20
rect 3370 80 3470 130
rect 3710 310 3810 320
rect 3710 250 3730 310
rect 3790 250 3810 310
rect 3710 200 3810 250
rect 3710 130 3730 200
rect 3790 130 3810 200
rect 3370 20 3390 80
rect 3450 20 3470 80
rect 3370 0 3470 20
rect 3540 80 3640 100
rect 3540 20 3560 80
rect 3620 20 3640 80
rect 3540 0 3640 20
rect 3710 80 3810 130
rect 4050 310 4150 320
rect 4050 250 4070 310
rect 4130 250 4150 310
rect 4050 200 4150 250
rect 4050 130 4070 200
rect 4130 130 4150 200
rect 3710 20 3730 80
rect 3790 20 3810 80
rect 3710 0 3810 20
rect 3880 80 3980 100
rect 3880 20 3900 80
rect 3960 20 3980 80
rect 3880 0 3980 20
rect 4050 80 4150 130
rect 4690 310 4790 320
rect 4690 250 4710 310
rect 4770 250 4790 310
rect 4690 200 4790 250
rect 4690 130 4710 200
rect 4770 130 4790 200
rect 4050 20 4070 80
rect 4130 20 4150 80
rect 4050 0 4150 20
rect 4220 80 4320 100
rect 4220 20 4240 80
rect 4300 20 4320 80
rect 4220 0 4320 20
rect 4520 80 4620 100
rect 4520 20 4540 80
rect 4600 20 4620 80
rect 4520 0 4620 20
rect 4690 80 4790 130
rect 5030 310 5130 320
rect 5030 250 5050 310
rect 5110 250 5130 310
rect 5030 200 5130 250
rect 5030 130 5050 200
rect 5110 130 5130 200
rect 4690 20 4710 80
rect 4770 20 4790 80
rect 4690 0 4790 20
rect 4860 80 4960 100
rect 4860 20 4880 80
rect 4940 20 4960 80
rect 4860 0 4960 20
rect 5030 80 5130 130
rect 5370 310 5470 320
rect 5370 250 5390 310
rect 5450 250 5470 310
rect 5370 200 5470 250
rect 5370 130 5390 200
rect 5450 130 5470 200
rect 5030 20 5050 80
rect 5110 20 5130 80
rect 5030 0 5130 20
rect 5200 80 5300 100
rect 5200 20 5220 80
rect 5280 20 5300 80
rect 5200 0 5300 20
rect 5370 80 5470 130
rect 5710 310 5810 320
rect 5710 250 5730 310
rect 5790 250 5810 310
rect 5710 200 5810 250
rect 5710 130 5730 200
rect 5790 130 5810 200
rect 5370 20 5390 80
rect 5450 20 5470 80
rect 5370 0 5470 20
rect 5540 80 5640 100
rect 5540 20 5560 80
rect 5620 20 5640 80
rect 5540 0 5640 20
rect 5710 80 5810 130
rect 6050 310 6150 320
rect 6050 250 6070 310
rect 6130 250 6150 310
rect 6050 200 6150 250
rect 6050 130 6070 200
rect 6130 130 6150 200
rect 5710 20 5730 80
rect 5790 20 5810 80
rect 5710 0 5810 20
rect 5880 80 5980 100
rect 5880 20 5900 80
rect 5960 20 5980 80
rect 5880 0 5980 20
rect 6050 80 6150 130
rect 6390 310 6490 320
rect 6390 250 6410 310
rect 6470 250 6490 310
rect 6390 200 6490 250
rect 6390 130 6410 200
rect 6470 130 6490 200
rect 6050 20 6070 80
rect 6130 20 6150 80
rect 6050 0 6150 20
rect 6220 80 6320 100
rect 6220 20 6240 80
rect 6300 20 6320 80
rect 6220 0 6320 20
rect 6390 80 6490 130
rect 6730 310 6830 320
rect 6730 250 6750 310
rect 6810 250 6830 310
rect 6730 200 6830 250
rect 6730 130 6750 200
rect 6810 130 6830 200
rect 6390 20 6410 80
rect 6470 20 6490 80
rect 6390 0 6490 20
rect 6560 80 6660 100
rect 6560 20 6580 80
rect 6640 20 6660 80
rect 6560 0 6660 20
rect 6730 80 6830 130
rect 7070 310 7170 320
rect 7070 250 7090 310
rect 7150 250 7170 310
rect 7070 200 7170 250
rect 7070 130 7090 200
rect 7150 130 7170 200
rect 6730 20 6750 80
rect 6810 20 6830 80
rect 6730 0 6830 20
rect 6900 80 7000 100
rect 6900 20 6920 80
rect 6980 20 7000 80
rect 6900 0 7000 20
rect 7070 80 7170 130
rect 7410 310 7510 320
rect 7410 250 7430 310
rect 7490 250 7510 310
rect 7410 200 7510 250
rect 7410 130 7430 200
rect 7490 130 7510 200
rect 7070 20 7090 80
rect 7150 20 7170 80
rect 7070 0 7170 20
rect 7240 80 7340 100
rect 7240 20 7260 80
rect 7320 20 7340 80
rect 7240 0 7340 20
rect 7410 80 7510 130
rect 7750 310 7850 320
rect 7750 250 7770 310
rect 7830 250 7850 310
rect 7750 200 7850 250
rect 7750 130 7770 200
rect 7830 130 7850 200
rect 7410 20 7430 80
rect 7490 20 7510 80
rect 7410 0 7510 20
rect 7580 80 7680 100
rect 7580 20 7600 80
rect 7660 20 7680 80
rect 7580 0 7680 20
rect 7750 80 7850 130
rect 8090 310 8190 320
rect 8090 250 8110 310
rect 8170 250 8190 310
rect 8090 200 8190 250
rect 8090 130 8110 200
rect 8170 130 8190 200
rect 7750 20 7770 80
rect 7830 20 7850 80
rect 7750 0 7850 20
rect 7920 80 8020 100
rect 7920 20 7940 80
rect 8000 20 8020 80
rect 7920 0 8020 20
rect 8090 80 8190 130
rect 8430 310 8530 320
rect 8430 250 8450 310
rect 8510 250 8530 310
rect 8430 200 8530 250
rect 8430 130 8450 200
rect 8510 130 8530 200
rect 8090 20 8110 80
rect 8170 20 8190 80
rect 8090 0 8190 20
rect 8260 80 8360 100
rect 8260 20 8280 80
rect 8340 20 8360 80
rect 8260 0 8360 20
rect 8430 80 8530 130
rect 8770 310 8870 320
rect 8770 250 8790 310
rect 8850 250 8870 310
rect 8770 200 8870 250
rect 8770 130 8790 200
rect 8850 130 8870 200
rect 8430 20 8450 80
rect 8510 20 8530 80
rect 8430 0 8530 20
rect 8600 80 8700 100
rect 8600 20 8620 80
rect 8680 20 8700 80
rect 8600 0 8700 20
rect 8770 80 8870 130
rect 9110 310 9210 320
rect 9110 250 9130 310
rect 9190 250 9210 310
rect 9110 200 9210 250
rect 9110 130 9130 200
rect 9190 130 9210 200
rect 8770 20 8790 80
rect 8850 20 8870 80
rect 8770 0 8870 20
rect 8940 80 9040 100
rect 8940 20 8960 80
rect 9020 20 9040 80
rect 8940 0 9040 20
rect 9110 80 9210 130
rect 9450 310 9550 320
rect 9450 250 9470 310
rect 9530 250 9550 310
rect 9450 200 9550 250
rect 9450 130 9470 200
rect 9530 130 9550 200
rect 9110 20 9130 80
rect 9190 20 9210 80
rect 9110 0 9210 20
rect 9280 80 9380 100
rect 9280 20 9300 80
rect 9360 20 9380 80
rect 9280 0 9380 20
rect 9450 80 9550 130
rect 9790 310 9890 320
rect 9790 250 9810 310
rect 9870 250 9890 310
rect 9790 200 9890 250
rect 9790 130 9810 200
rect 9870 130 9890 200
rect 9450 20 9470 80
rect 9530 20 9550 80
rect 9450 0 9550 20
rect 9620 80 9720 100
rect 9620 20 9640 80
rect 9700 20 9720 80
rect 9620 0 9720 20
rect 9790 80 9890 130
rect 10130 310 10230 320
rect 10130 250 10150 310
rect 10210 250 10230 310
rect 10130 200 10230 250
rect 10130 130 10150 200
rect 10210 130 10230 200
rect 9790 20 9810 80
rect 9870 20 9890 80
rect 9790 0 9890 20
rect 9960 80 10060 100
rect 9960 20 9980 80
rect 10040 20 10060 80
rect 9960 0 10060 20
rect 10130 80 10230 130
rect 10470 310 10570 320
rect 10470 250 10490 310
rect 10550 250 10570 310
rect 10470 200 10570 250
rect 10470 130 10490 200
rect 10550 130 10570 200
rect 10130 20 10150 80
rect 10210 20 10230 80
rect 10130 0 10230 20
rect 10300 80 10400 100
rect 10300 20 10320 80
rect 10380 20 10400 80
rect 10300 0 10400 20
rect 10470 80 10570 130
rect 10810 310 10910 320
rect 10810 250 10830 310
rect 10890 250 10910 310
rect 10810 200 10910 250
rect 10810 130 10830 200
rect 10890 130 10910 200
rect 10470 20 10490 80
rect 10550 20 10570 80
rect 10470 0 10570 20
rect 10640 80 10740 100
rect 10640 20 10660 80
rect 10720 20 10740 80
rect 10640 0 10740 20
rect 10810 80 10910 130
rect 11150 310 11250 320
rect 11150 250 11170 310
rect 11230 250 11250 310
rect 11150 200 11250 250
rect 11150 130 11170 200
rect 11230 130 11250 200
rect 10810 20 10830 80
rect 10890 20 10910 80
rect 10810 0 10910 20
rect 10980 80 11080 100
rect 10980 20 11000 80
rect 11060 20 11080 80
rect 10980 0 11080 20
rect 11150 80 11250 130
rect 11490 310 11590 320
rect 11490 250 11510 310
rect 11570 250 11590 310
rect 11490 200 11590 250
rect 11490 130 11510 200
rect 11570 130 11590 200
rect 11150 20 11170 80
rect 11230 20 11250 80
rect 11150 0 11250 20
rect 11320 80 11420 100
rect 11320 20 11340 80
rect 11400 20 11420 80
rect 11320 0 11420 20
rect 11490 80 11590 130
rect 11830 310 11930 320
rect 11830 250 11850 310
rect 11910 250 11930 310
rect 11830 200 11930 250
rect 11830 130 11850 200
rect 11910 130 11930 200
rect 11490 20 11510 80
rect 11570 20 11590 80
rect 11490 0 11590 20
rect 11660 80 11760 100
rect 11660 20 11680 80
rect 11740 20 11760 80
rect 11660 0 11760 20
rect 11830 80 11930 130
rect 12170 310 12270 320
rect 12170 250 12190 310
rect 12250 250 12270 310
rect 12170 200 12270 250
rect 12170 130 12190 200
rect 12250 130 12270 200
rect 11830 20 11850 80
rect 11910 20 11930 80
rect 11830 0 11930 20
rect 12000 80 12100 100
rect 12000 20 12020 80
rect 12080 20 12100 80
rect 12000 0 12100 20
rect 12170 80 12270 130
rect 12510 310 12610 320
rect 12510 250 12530 310
rect 12590 250 12610 310
rect 12510 200 12610 250
rect 12510 130 12530 200
rect 12590 130 12610 200
rect 12170 20 12190 80
rect 12250 20 12270 80
rect 12170 0 12270 20
rect 12340 80 12440 100
rect 12340 20 12360 80
rect 12420 20 12440 80
rect 12340 0 12440 20
rect 12510 80 12610 130
rect 12850 310 12950 320
rect 12850 250 12870 310
rect 12930 250 12950 310
rect 12850 200 12950 250
rect 12850 130 12870 200
rect 12930 130 12950 200
rect 12510 20 12530 80
rect 12590 20 12610 80
rect 12510 0 12610 20
rect 12680 80 12780 100
rect 12680 20 12700 80
rect 12760 20 12780 80
rect 12680 0 12780 20
rect 12850 80 12950 130
rect 13190 310 13290 320
rect 13190 250 13210 310
rect 13270 250 13290 310
rect 13190 200 13290 250
rect 13190 130 13210 200
rect 13270 130 13290 200
rect 12850 20 12870 80
rect 12930 20 12950 80
rect 12850 0 12950 20
rect 13020 80 13120 100
rect 13020 20 13040 80
rect 13100 20 13120 80
rect 13020 0 13120 20
rect 13190 80 13290 130
rect 13530 310 13630 320
rect 13530 250 13550 310
rect 13610 250 13630 310
rect 13530 200 13630 250
rect 13530 130 13550 200
rect 13610 130 13630 200
rect 13190 20 13210 80
rect 13270 20 13290 80
rect 13190 0 13290 20
rect 13360 80 13460 100
rect 13360 20 13380 80
rect 13440 20 13460 80
rect 13360 0 13460 20
rect 13530 80 13630 130
rect 13870 310 13970 320
rect 13870 250 13890 310
rect 13950 250 13970 310
rect 13870 200 13970 250
rect 13870 130 13890 200
rect 13950 130 13970 200
rect 13530 20 13550 80
rect 13610 20 13630 80
rect 13530 0 13630 20
rect 13700 80 13800 100
rect 13700 20 13720 80
rect 13780 20 13800 80
rect 13700 0 13800 20
rect 13870 80 13970 130
rect 14210 310 14310 320
rect 14210 250 14230 310
rect 14290 250 14310 310
rect 14210 200 14310 250
rect 14210 130 14230 200
rect 14290 130 14310 200
rect 13870 20 13890 80
rect 13950 20 13970 80
rect 13870 0 13970 20
rect 14040 80 14140 100
rect 14040 20 14060 80
rect 14120 20 14140 80
rect 14040 0 14140 20
rect 14210 80 14310 130
rect 14550 310 14650 320
rect 14550 250 14570 310
rect 14630 250 14650 310
rect 14550 200 14650 250
rect 14550 130 14570 200
rect 14630 130 14650 200
rect 14210 20 14230 80
rect 14290 20 14310 80
rect 14210 0 14310 20
rect 14380 80 14480 100
rect 14380 20 14400 80
rect 14460 20 14480 80
rect 14380 0 14480 20
rect 14550 80 14650 130
rect 14890 310 14990 320
rect 14890 250 14910 310
rect 14970 250 14990 310
rect 14890 200 14990 250
rect 14890 130 14910 200
rect 14970 130 14990 200
rect 14550 20 14570 80
rect 14630 20 14650 80
rect 14550 0 14650 20
rect 14720 80 14820 100
rect 14720 20 14740 80
rect 14800 20 14820 80
rect 14720 0 14820 20
rect 14890 80 14990 130
rect 15230 310 15330 320
rect 15230 250 15250 310
rect 15310 250 15330 310
rect 15230 200 15330 250
rect 15230 130 15250 200
rect 15310 130 15330 200
rect 14890 20 14910 80
rect 14970 20 14990 80
rect 14890 0 14990 20
rect 15060 80 15160 100
rect 15060 20 15080 80
rect 15140 20 15160 80
rect 15060 0 15160 20
rect 15230 80 15330 130
rect 15870 310 15970 320
rect 15870 250 15890 310
rect 15950 250 15970 310
rect 15870 200 15970 250
rect 15870 130 15890 200
rect 15950 130 15970 200
rect 15230 20 15250 80
rect 15310 20 15330 80
rect 15230 0 15330 20
rect 15400 80 15500 100
rect 15400 20 15420 80
rect 15480 20 15500 80
rect 15400 0 15500 20
rect 15700 80 15800 100
rect 15700 20 15720 80
rect 15780 20 15800 80
rect 15700 0 15800 20
rect 15870 80 15970 130
rect 16210 310 16310 320
rect 16210 250 16230 310
rect 16290 250 16310 310
rect 16210 200 16310 250
rect 16210 130 16230 200
rect 16290 130 16310 200
rect 15870 20 15890 80
rect 15950 20 15970 80
rect 15870 0 15970 20
rect 16040 80 16140 100
rect 16040 20 16060 80
rect 16120 20 16140 80
rect 16040 0 16140 20
rect 16210 80 16310 130
rect 16550 310 16650 320
rect 16550 250 16570 310
rect 16630 250 16650 310
rect 16550 200 16650 250
rect 16550 130 16570 200
rect 16630 130 16650 200
rect 16210 20 16230 80
rect 16290 20 16310 80
rect 16210 0 16310 20
rect 16380 80 16480 100
rect 16380 20 16400 80
rect 16460 20 16480 80
rect 16380 0 16480 20
rect 16550 80 16650 130
rect 16890 310 16990 320
rect 16890 250 16910 310
rect 16970 250 16990 310
rect 16890 200 16990 250
rect 16890 130 16910 200
rect 16970 130 16990 200
rect 16550 20 16570 80
rect 16630 20 16650 80
rect 16550 0 16650 20
rect 16720 80 16820 100
rect 16720 20 16740 80
rect 16800 20 16820 80
rect 16720 0 16820 20
rect 16890 80 16990 130
rect 17230 310 17330 320
rect 17230 250 17250 310
rect 17310 250 17330 310
rect 17230 200 17330 250
rect 17230 130 17250 200
rect 17310 130 17330 200
rect 16890 20 16910 80
rect 16970 20 16990 80
rect 16890 0 16990 20
rect 17060 80 17160 100
rect 17060 20 17080 80
rect 17140 20 17160 80
rect 17060 0 17160 20
rect 17230 80 17330 130
rect 17570 310 17670 320
rect 17570 250 17590 310
rect 17650 250 17670 310
rect 17570 200 17670 250
rect 17570 130 17590 200
rect 17650 130 17670 200
rect 17230 20 17250 80
rect 17310 20 17330 80
rect 17230 0 17330 20
rect 17400 80 17500 100
rect 17400 20 17420 80
rect 17480 20 17500 80
rect 17400 0 17500 20
rect 17570 80 17670 130
rect 17910 310 18010 320
rect 17910 250 17930 310
rect 17990 250 18010 310
rect 17910 200 18010 250
rect 17910 130 17930 200
rect 17990 130 18010 200
rect 17570 20 17590 80
rect 17650 20 17670 80
rect 17570 0 17670 20
rect 17740 80 17840 100
rect 17740 20 17760 80
rect 17820 20 17840 80
rect 17740 0 17840 20
rect 17910 80 18010 130
rect 18250 310 18350 320
rect 18250 250 18270 310
rect 18330 250 18350 310
rect 18250 200 18350 250
rect 18250 130 18270 200
rect 18330 130 18350 200
rect 17910 20 17930 80
rect 17990 20 18010 80
rect 17910 0 18010 20
rect 18080 80 18180 100
rect 18080 20 18100 80
rect 18160 20 18180 80
rect 18080 0 18180 20
rect 18250 80 18350 130
rect 18590 310 18690 320
rect 18590 250 18610 310
rect 18670 250 18690 310
rect 18590 200 18690 250
rect 18590 130 18610 200
rect 18670 130 18690 200
rect 18250 20 18270 80
rect 18330 20 18350 80
rect 18250 0 18350 20
rect 18420 80 18520 100
rect 18420 20 18440 80
rect 18500 20 18520 80
rect 18420 0 18520 20
rect 18590 80 18690 130
rect 18930 310 19030 320
rect 18930 250 18950 310
rect 19010 250 19030 310
rect 18930 200 19030 250
rect 18930 130 18950 200
rect 19010 130 19030 200
rect 18590 20 18610 80
rect 18670 20 18690 80
rect 18590 0 18690 20
rect 18760 80 18860 100
rect 18760 20 18780 80
rect 18840 20 18860 80
rect 18760 0 18860 20
rect 18930 80 19030 130
rect 19270 310 19370 320
rect 19270 250 19290 310
rect 19350 250 19370 310
rect 19270 200 19370 250
rect 19270 130 19290 200
rect 19350 130 19370 200
rect 18930 20 18950 80
rect 19010 20 19030 80
rect 18930 0 19030 20
rect 19100 80 19200 100
rect 19100 20 19120 80
rect 19180 20 19200 80
rect 19100 0 19200 20
rect 19270 80 19370 130
rect 19610 310 19710 320
rect 19610 250 19630 310
rect 19690 250 19710 310
rect 19610 200 19710 250
rect 19610 130 19630 200
rect 19690 130 19710 200
rect 19270 20 19290 80
rect 19350 20 19370 80
rect 19270 0 19370 20
rect 19440 80 19540 100
rect 19440 20 19460 80
rect 19520 20 19540 80
rect 19440 0 19540 20
rect 19610 80 19710 130
rect 19950 310 20050 320
rect 19950 250 19970 310
rect 20030 250 20050 310
rect 19950 200 20050 250
rect 19950 130 19970 200
rect 20030 130 20050 200
rect 19610 20 19630 80
rect 19690 20 19710 80
rect 19610 0 19710 20
rect 19780 80 19880 100
rect 19780 20 19800 80
rect 19860 20 19880 80
rect 19780 0 19880 20
rect 19950 80 20050 130
rect 20290 310 20390 320
rect 20290 250 20310 310
rect 20370 250 20390 310
rect 20290 200 20390 250
rect 20290 130 20310 200
rect 20370 130 20390 200
rect 19950 20 19970 80
rect 20030 20 20050 80
rect 19950 0 20050 20
rect 20120 80 20220 100
rect 20120 20 20140 80
rect 20200 20 20220 80
rect 20120 0 20220 20
rect 20290 80 20390 130
rect 20630 310 20730 320
rect 20630 250 20650 310
rect 20710 250 20730 310
rect 20630 200 20730 250
rect 20630 130 20650 200
rect 20710 130 20730 200
rect 20290 20 20310 80
rect 20370 20 20390 80
rect 20290 0 20390 20
rect 20460 80 20560 100
rect 20460 20 20480 80
rect 20540 20 20560 80
rect 20460 0 20560 20
rect 20630 80 20730 130
rect 20970 310 21070 320
rect 20970 250 20990 310
rect 21050 250 21070 310
rect 20970 200 21070 250
rect 20970 130 20990 200
rect 21050 130 21070 200
rect 20630 20 20650 80
rect 20710 20 20730 80
rect 20630 0 20730 20
rect 20800 80 20900 100
rect 20800 20 20820 80
rect 20880 20 20900 80
rect 20800 0 20900 20
rect 20970 80 21070 130
rect 21310 310 21410 320
rect 21310 250 21330 310
rect 21390 250 21410 310
rect 21310 200 21410 250
rect 21310 130 21330 200
rect 21390 130 21410 200
rect 20970 20 20990 80
rect 21050 20 21070 80
rect 20970 0 21070 20
rect 21140 80 21240 100
rect 21140 20 21160 80
rect 21220 20 21240 80
rect 21140 0 21240 20
rect 21310 80 21410 130
rect 21650 310 21750 320
rect 21650 250 21670 310
rect 21730 250 21750 310
rect 21650 200 21750 250
rect 21650 130 21670 200
rect 21730 130 21750 200
rect 21310 20 21330 80
rect 21390 20 21410 80
rect 21310 0 21410 20
rect 21480 80 21580 100
rect 21480 20 21500 80
rect 21560 20 21580 80
rect 21480 0 21580 20
rect 21650 80 21750 130
rect 21990 310 22090 320
rect 21990 250 22010 310
rect 22070 250 22090 310
rect 21990 200 22090 250
rect 21990 130 22010 200
rect 22070 130 22090 200
rect 21650 20 21670 80
rect 21730 20 21750 80
rect 21650 0 21750 20
rect 21820 80 21920 100
rect 21820 20 21840 80
rect 21900 20 21920 80
rect 21820 0 21920 20
rect 21990 80 22090 130
rect 22330 310 22430 320
rect 22330 250 22350 310
rect 22410 250 22430 310
rect 22330 200 22430 250
rect 22330 130 22350 200
rect 22410 130 22430 200
rect 21990 20 22010 80
rect 22070 20 22090 80
rect 21990 0 22090 20
rect 22160 80 22260 100
rect 22160 20 22180 80
rect 22240 20 22260 80
rect 22160 0 22260 20
rect 22330 80 22430 130
rect 22670 310 22770 320
rect 22670 250 22690 310
rect 22750 250 22770 310
rect 22670 200 22770 250
rect 22670 130 22690 200
rect 22750 130 22770 200
rect 22330 20 22350 80
rect 22410 20 22430 80
rect 22330 0 22430 20
rect 22500 80 22600 100
rect 22500 20 22520 80
rect 22580 20 22600 80
rect 22500 0 22600 20
rect 22670 80 22770 130
rect 23010 310 23110 320
rect 23010 250 23030 310
rect 23090 250 23110 310
rect 23010 200 23110 250
rect 23010 130 23030 200
rect 23090 130 23110 200
rect 22670 20 22690 80
rect 22750 20 22770 80
rect 22670 0 22770 20
rect 22840 80 22940 100
rect 22840 20 22860 80
rect 22920 20 22940 80
rect 22840 0 22940 20
rect 23010 80 23110 130
rect 23350 310 23450 320
rect 23350 250 23370 310
rect 23430 250 23450 310
rect 23350 200 23450 250
rect 23350 130 23370 200
rect 23430 130 23450 200
rect 23010 20 23030 80
rect 23090 20 23110 80
rect 23010 0 23110 20
rect 23180 80 23280 100
rect 23180 20 23200 80
rect 23260 20 23280 80
rect 23180 0 23280 20
rect 23350 80 23450 130
rect 23690 310 23790 320
rect 23690 250 23710 310
rect 23770 250 23790 310
rect 23690 200 23790 250
rect 23690 130 23710 200
rect 23770 130 23790 200
rect 23350 20 23370 80
rect 23430 20 23450 80
rect 23350 0 23450 20
rect 23520 80 23620 100
rect 23520 20 23540 80
rect 23600 20 23620 80
rect 23520 0 23620 20
rect 23690 80 23790 130
rect 24030 310 24130 320
rect 24030 250 24050 310
rect 24110 250 24130 310
rect 24030 200 24130 250
rect 24030 130 24050 200
rect 24110 130 24130 200
rect 23690 20 23710 80
rect 23770 20 23790 80
rect 23690 0 23790 20
rect 23860 80 23960 100
rect 23860 20 23880 80
rect 23940 20 23960 80
rect 23860 0 23960 20
rect 24030 80 24130 130
rect 24370 310 24470 320
rect 24370 250 24390 310
rect 24450 250 24470 310
rect 24370 200 24470 250
rect 24370 130 24390 200
rect 24450 130 24470 200
rect 24030 20 24050 80
rect 24110 20 24130 80
rect 24030 0 24130 20
rect 24200 80 24300 100
rect 24200 20 24220 80
rect 24280 20 24300 80
rect 24200 0 24300 20
rect 24370 80 24470 130
rect 24710 310 24810 320
rect 24710 250 24730 310
rect 24790 250 24810 310
rect 24710 200 24810 250
rect 24710 130 24730 200
rect 24790 130 24810 200
rect 24370 20 24390 80
rect 24450 20 24470 80
rect 24370 0 24470 20
rect 24540 80 24640 100
rect 24540 20 24560 80
rect 24620 20 24640 80
rect 24540 0 24640 20
rect 24710 80 24810 130
rect 25050 310 25150 320
rect 25050 250 25070 310
rect 25130 250 25150 310
rect 25050 200 25150 250
rect 25050 130 25070 200
rect 25130 130 25150 200
rect 24710 20 24730 80
rect 24790 20 24810 80
rect 24710 0 24810 20
rect 24880 80 24980 100
rect 24880 20 24900 80
rect 24960 20 24980 80
rect 24880 0 24980 20
rect 25050 80 25150 130
rect 25390 310 25490 320
rect 25390 250 25410 310
rect 25470 250 25490 310
rect 25390 200 25490 250
rect 25390 130 25410 200
rect 25470 130 25490 200
rect 25050 20 25070 80
rect 25130 20 25150 80
rect 25050 0 25150 20
rect 25220 80 25320 100
rect 25220 20 25240 80
rect 25300 20 25320 80
rect 25220 0 25320 20
rect 25390 80 25490 130
rect 25730 310 25830 320
rect 25730 250 25750 310
rect 25810 250 25830 310
rect 25730 200 25830 250
rect 25730 130 25750 200
rect 25810 130 25830 200
rect 25390 20 25410 80
rect 25470 20 25490 80
rect 25390 0 25490 20
rect 25560 80 25660 100
rect 25560 20 25580 80
rect 25640 20 25660 80
rect 25560 0 25660 20
rect 25730 80 25830 130
rect 26070 310 26170 320
rect 26070 250 26090 310
rect 26150 250 26170 310
rect 26070 200 26170 250
rect 26070 130 26090 200
rect 26150 130 26170 200
rect 25730 20 25750 80
rect 25810 20 25830 80
rect 25730 0 25830 20
rect 25900 80 26000 100
rect 25900 20 25920 80
rect 25980 20 26000 80
rect 25900 0 26000 20
rect 26070 80 26170 130
rect 26410 310 26510 320
rect 26410 250 26430 310
rect 26490 250 26510 310
rect 26410 200 26510 250
rect 26410 130 26430 200
rect 26490 130 26510 200
rect 26070 20 26090 80
rect 26150 20 26170 80
rect 26070 0 26170 20
rect 26240 80 26340 100
rect 26240 20 26260 80
rect 26320 20 26340 80
rect 26240 0 26340 20
rect 26410 80 26510 130
rect 26750 310 26850 320
rect 26750 250 26770 310
rect 26830 250 26850 310
rect 26750 200 26850 250
rect 26750 130 26770 200
rect 26830 130 26850 200
rect 26410 20 26430 80
rect 26490 20 26510 80
rect 26410 0 26510 20
rect 26580 80 26680 100
rect 26580 20 26600 80
rect 26660 20 26680 80
rect 26580 0 26680 20
rect 26750 80 26850 130
rect 27090 310 27190 320
rect 27090 250 27110 310
rect 27170 250 27190 310
rect 27090 200 27190 250
rect 27090 130 27110 200
rect 27170 130 27190 200
rect 26750 20 26770 80
rect 26830 20 26850 80
rect 26750 0 26850 20
rect 26920 80 27020 100
rect 26920 20 26940 80
rect 27000 20 27020 80
rect 26920 0 27020 20
rect 27090 80 27190 130
rect 27430 310 27530 320
rect 27430 250 27450 310
rect 27510 250 27530 310
rect 27430 200 27530 250
rect 27430 130 27450 200
rect 27510 130 27530 200
rect 27090 20 27110 80
rect 27170 20 27190 80
rect 27090 0 27190 20
rect 27260 80 27360 100
rect 27260 20 27280 80
rect 27340 20 27360 80
rect 27260 0 27360 20
rect 27430 80 27530 130
rect 27770 310 27870 320
rect 27770 250 27790 310
rect 27850 250 27870 310
rect 27770 200 27870 250
rect 27770 130 27790 200
rect 27850 130 27870 200
rect 27430 20 27450 80
rect 27510 20 27530 80
rect 27430 0 27530 20
rect 27600 80 27700 100
rect 27600 20 27620 80
rect 27680 20 27700 80
rect 27600 0 27700 20
rect 27770 80 27870 130
rect 28110 310 28210 320
rect 28110 250 28130 310
rect 28190 250 28210 310
rect 28110 200 28210 250
rect 28110 130 28130 200
rect 28190 130 28210 200
rect 27770 20 27790 80
rect 27850 20 27870 80
rect 27770 0 27870 20
rect 27940 80 28040 100
rect 27940 20 27960 80
rect 28020 20 28040 80
rect 27940 0 28040 20
rect 28110 80 28210 130
rect 28450 310 28550 320
rect 28450 250 28470 310
rect 28530 250 28550 310
rect 28450 200 28550 250
rect 28450 130 28470 200
rect 28530 130 28550 200
rect 28110 20 28130 80
rect 28190 20 28210 80
rect 28110 0 28210 20
rect 28280 80 28380 100
rect 28280 20 28300 80
rect 28360 20 28380 80
rect 28280 0 28380 20
rect 28450 80 28550 130
rect 28790 310 28890 320
rect 28790 250 28810 310
rect 28870 250 28890 310
rect 28790 200 28890 250
rect 28790 130 28810 200
rect 28870 130 28890 200
rect 28450 20 28470 80
rect 28530 20 28550 80
rect 28450 0 28550 20
rect 28620 80 28720 100
rect 28620 20 28640 80
rect 28700 20 28720 80
rect 28620 0 28720 20
rect 28790 80 28890 130
rect 29130 310 29230 320
rect 29130 250 29150 310
rect 29210 250 29230 310
rect 29130 200 29230 250
rect 29130 130 29150 200
rect 29210 130 29230 200
rect 28790 20 28810 80
rect 28870 20 28890 80
rect 28790 0 28890 20
rect 28960 80 29060 100
rect 28960 20 28980 80
rect 29040 20 29060 80
rect 28960 0 29060 20
rect 29130 80 29230 130
rect 29470 310 29570 320
rect 29470 250 29490 310
rect 29550 250 29570 310
rect 29470 200 29570 250
rect 29470 130 29490 200
rect 29550 130 29570 200
rect 29130 20 29150 80
rect 29210 20 29230 80
rect 29130 0 29230 20
rect 29300 80 29400 100
rect 29300 20 29320 80
rect 29380 20 29400 80
rect 29300 0 29400 20
rect 29470 80 29570 130
rect 29810 310 29910 320
rect 29810 250 29830 310
rect 29890 250 29910 310
rect 29810 200 29910 250
rect 29810 130 29830 200
rect 29890 130 29910 200
rect 29470 20 29490 80
rect 29550 20 29570 80
rect 29470 0 29570 20
rect 29640 80 29740 100
rect 29640 20 29660 80
rect 29720 20 29740 80
rect 29640 0 29740 20
rect 29810 80 29910 130
rect 30150 310 30250 320
rect 30150 250 30170 310
rect 30230 250 30250 310
rect 30150 200 30250 250
rect 30150 130 30170 200
rect 30230 130 30250 200
rect 29810 20 29830 80
rect 29890 20 29910 80
rect 29810 0 29910 20
rect 29980 80 30080 100
rect 29980 20 30000 80
rect 30060 20 30080 80
rect 29980 0 30080 20
rect 30150 80 30250 130
rect 30490 310 30590 320
rect 30490 250 30510 310
rect 30570 250 30590 310
rect 30490 200 30590 250
rect 30490 130 30510 200
rect 30570 130 30590 200
rect 30150 20 30170 80
rect 30230 20 30250 80
rect 30150 0 30250 20
rect 30320 80 30420 100
rect 30320 20 30340 80
rect 30400 20 30420 80
rect 30320 0 30420 20
rect 30490 80 30590 130
rect 30830 310 30930 320
rect 30830 250 30850 310
rect 30910 250 30930 310
rect 30830 200 30930 250
rect 30830 130 30850 200
rect 30910 130 30930 200
rect 30490 20 30510 80
rect 30570 20 30590 80
rect 30490 0 30590 20
rect 30660 80 30760 100
rect 30660 20 30680 80
rect 30740 20 30760 80
rect 30660 0 30760 20
rect 30830 80 30930 130
rect 31170 310 31270 320
rect 31170 250 31190 310
rect 31250 250 31270 310
rect 31170 200 31270 250
rect 31170 130 31190 200
rect 31250 130 31270 200
rect 30830 20 30850 80
rect 30910 20 30930 80
rect 30830 0 30930 20
rect 31000 80 31100 100
rect 31000 20 31020 80
rect 31080 20 31100 80
rect 31000 0 31100 20
rect 31170 80 31270 130
rect 31510 310 31610 320
rect 31510 250 31530 310
rect 31590 250 31610 310
rect 31510 200 31610 250
rect 31510 130 31530 200
rect 31590 130 31610 200
rect 31170 20 31190 80
rect 31250 20 31270 80
rect 31170 0 31270 20
rect 31340 80 31440 100
rect 31340 20 31360 80
rect 31420 20 31440 80
rect 31340 0 31440 20
rect 31510 80 31610 130
rect 31850 310 31950 320
rect 31850 250 31870 310
rect 31930 250 31950 310
rect 31850 200 31950 250
rect 31850 130 31870 200
rect 31930 130 31950 200
rect 31510 20 31530 80
rect 31590 20 31610 80
rect 31510 0 31610 20
rect 31680 80 31780 100
rect 31680 20 31700 80
rect 31760 20 31780 80
rect 31680 0 31780 20
rect 31850 80 31950 130
rect 32190 310 32290 320
rect 32190 250 32210 310
rect 32270 250 32290 310
rect 32190 200 32290 250
rect 32190 130 32210 200
rect 32270 130 32290 200
rect 31850 20 31870 80
rect 31930 20 31950 80
rect 31850 0 31950 20
rect 32020 80 32120 100
rect 32020 20 32040 80
rect 32100 20 32120 80
rect 32020 0 32120 20
rect 32190 80 32290 130
rect 32530 310 32630 320
rect 32530 250 32550 310
rect 32610 250 32630 310
rect 32530 200 32630 250
rect 32530 130 32550 200
rect 32610 130 32630 200
rect 32190 20 32210 80
rect 32270 20 32290 80
rect 32190 0 32290 20
rect 32360 80 32460 100
rect 32360 20 32380 80
rect 32440 20 32460 80
rect 32360 0 32460 20
rect 32530 80 32630 130
rect 32870 310 32970 320
rect 32870 250 32890 310
rect 32950 250 32970 310
rect 32870 200 32970 250
rect 32870 130 32890 200
rect 32950 130 32970 200
rect 32530 20 32550 80
rect 32610 20 32630 80
rect 32530 0 32630 20
rect 32700 80 32800 100
rect 32700 20 32720 80
rect 32780 20 32800 80
rect 32700 0 32800 20
rect 32870 80 32970 130
rect 33210 310 33310 320
rect 33210 250 33230 310
rect 33290 250 33310 310
rect 33210 200 33310 250
rect 33210 130 33230 200
rect 33290 130 33310 200
rect 32870 20 32890 80
rect 32950 20 32970 80
rect 32870 0 32970 20
rect 33040 80 33140 100
rect 33040 20 33060 80
rect 33120 20 33140 80
rect 33040 0 33140 20
rect 33210 80 33310 130
rect 33550 310 33650 320
rect 33550 250 33570 310
rect 33630 250 33650 310
rect 33550 200 33650 250
rect 33550 130 33570 200
rect 33630 130 33650 200
rect 33210 20 33230 80
rect 33290 20 33310 80
rect 33210 0 33310 20
rect 33380 80 33480 100
rect 33380 20 33400 80
rect 33460 20 33480 80
rect 33380 0 33480 20
rect 33550 80 33650 130
rect 33890 310 33990 320
rect 33890 250 33910 310
rect 33970 250 33990 310
rect 33890 200 33990 250
rect 33890 130 33910 200
rect 33970 130 33990 200
rect 33550 20 33570 80
rect 33630 20 33650 80
rect 33550 0 33650 20
rect 33720 80 33820 100
rect 33720 20 33740 80
rect 33800 20 33820 80
rect 33720 0 33820 20
rect 33890 80 33990 130
rect 34230 310 34330 320
rect 34230 250 34250 310
rect 34310 250 34330 310
rect 34230 200 34330 250
rect 34230 130 34250 200
rect 34310 130 34330 200
rect 33890 20 33910 80
rect 33970 20 33990 80
rect 33890 0 33990 20
rect 34060 80 34160 100
rect 34060 20 34080 80
rect 34140 20 34160 80
rect 34060 0 34160 20
rect 34230 80 34330 130
rect 34570 310 34670 320
rect 34570 250 34590 310
rect 34650 250 34670 310
rect 34570 200 34670 250
rect 34570 130 34590 200
rect 34650 130 34670 200
rect 34230 20 34250 80
rect 34310 20 34330 80
rect 34230 0 34330 20
rect 34400 80 34500 100
rect 34400 20 34420 80
rect 34480 20 34500 80
rect 34400 0 34500 20
rect 34570 80 34670 130
rect 34910 310 35010 320
rect 34910 250 34930 310
rect 34990 250 35010 310
rect 34910 200 35010 250
rect 34910 130 34930 200
rect 34990 130 35010 200
rect 34570 20 34590 80
rect 34650 20 34670 80
rect 34570 0 34670 20
rect 34740 80 34840 100
rect 34740 20 34760 80
rect 34820 20 34840 80
rect 34740 0 34840 20
rect 34910 80 35010 130
rect 35250 310 35350 320
rect 35250 250 35270 310
rect 35330 250 35350 310
rect 35250 200 35350 250
rect 35250 130 35270 200
rect 35330 130 35350 200
rect 34910 20 34930 80
rect 34990 20 35010 80
rect 34910 0 35010 20
rect 35080 80 35180 100
rect 35080 20 35100 80
rect 35160 20 35180 80
rect 35080 0 35180 20
rect 35250 80 35350 130
rect 35590 310 35690 320
rect 35590 250 35610 310
rect 35670 250 35690 310
rect 35590 200 35690 250
rect 35590 130 35610 200
rect 35670 130 35690 200
rect 35250 20 35270 80
rect 35330 20 35350 80
rect 35250 0 35350 20
rect 35420 80 35520 100
rect 35420 20 35440 80
rect 35500 20 35520 80
rect 35420 0 35520 20
rect 35590 80 35690 130
rect 35930 310 36030 320
rect 35930 250 35950 310
rect 36010 250 36030 310
rect 35930 200 36030 250
rect 35930 130 35950 200
rect 36010 130 36030 200
rect 35590 20 35610 80
rect 35670 20 35690 80
rect 35590 0 35690 20
rect 35760 80 35860 100
rect 35760 20 35780 80
rect 35840 20 35860 80
rect 35760 0 35860 20
rect 35930 80 36030 130
rect 36270 310 36370 320
rect 36270 250 36290 310
rect 36350 250 36370 310
rect 36270 200 36370 250
rect 36270 130 36290 200
rect 36350 130 36370 200
rect 35930 20 35950 80
rect 36010 20 36030 80
rect 35930 0 36030 20
rect 36100 80 36200 100
rect 36100 20 36120 80
rect 36180 20 36200 80
rect 36100 0 36200 20
rect 36270 80 36370 130
rect 36610 310 36710 320
rect 36610 250 36630 310
rect 36690 250 36710 310
rect 36610 200 36710 250
rect 36610 130 36630 200
rect 36690 130 36710 200
rect 36270 20 36290 80
rect 36350 20 36370 80
rect 36270 0 36370 20
rect 36440 80 36540 100
rect 36440 20 36460 80
rect 36520 20 36540 80
rect 36440 0 36540 20
rect 36610 80 36710 130
rect 36950 310 37050 320
rect 36950 250 36970 310
rect 37030 250 37050 310
rect 36950 200 37050 250
rect 36950 130 36970 200
rect 37030 130 37050 200
rect 36610 20 36630 80
rect 36690 20 36710 80
rect 36610 0 36710 20
rect 36780 80 36880 100
rect 36780 20 36800 80
rect 36860 20 36880 80
rect 36780 0 36880 20
rect 36950 80 37050 130
rect 37290 310 37390 320
rect 37290 250 37310 310
rect 37370 250 37390 310
rect 37290 200 37390 250
rect 37290 130 37310 200
rect 37370 130 37390 200
rect 36950 20 36970 80
rect 37030 20 37050 80
rect 36950 0 37050 20
rect 37120 80 37220 100
rect 37120 20 37140 80
rect 37200 20 37220 80
rect 37120 0 37220 20
rect 37290 80 37390 130
rect 37630 310 37730 320
rect 37630 250 37650 310
rect 37710 250 37730 310
rect 37630 200 37730 250
rect 37630 130 37650 200
rect 37710 130 37730 200
rect 37290 20 37310 80
rect 37370 20 37390 80
rect 37290 0 37390 20
rect 37460 80 37560 100
rect 37460 20 37480 80
rect 37540 20 37560 80
rect 37460 0 37560 20
rect 37630 80 37730 130
rect 37970 310 38070 320
rect 37970 250 37990 310
rect 38050 250 38070 310
rect 37970 200 38070 250
rect 37970 130 37990 200
rect 38050 130 38070 200
rect 37630 20 37650 80
rect 37710 20 37730 80
rect 37630 0 37730 20
rect 37800 80 37900 100
rect 37800 20 37820 80
rect 37880 20 37900 80
rect 37800 0 37900 20
rect 37970 80 38070 130
rect 38310 310 38410 320
rect 38310 250 38330 310
rect 38390 250 38410 310
rect 38310 200 38410 250
rect 38310 130 38330 200
rect 38390 130 38410 200
rect 37970 20 37990 80
rect 38050 20 38070 80
rect 37970 0 38070 20
rect 38140 80 38240 100
rect 38140 20 38160 80
rect 38220 20 38240 80
rect 38140 0 38240 20
rect 38310 80 38410 130
rect 38650 310 38750 320
rect 38650 250 38670 310
rect 38730 250 38750 310
rect 38650 200 38750 250
rect 38650 130 38670 200
rect 38730 130 38750 200
rect 38310 20 38330 80
rect 38390 20 38410 80
rect 38310 0 38410 20
rect 38480 80 38580 100
rect 38480 20 38500 80
rect 38560 20 38580 80
rect 38480 0 38580 20
rect 38650 80 38750 130
rect 38990 310 39090 320
rect 38990 250 39010 310
rect 39070 250 39090 310
rect 38990 200 39090 250
rect 38990 130 39010 200
rect 39070 130 39090 200
rect 38650 20 38670 80
rect 38730 20 38750 80
rect 38650 0 38750 20
rect 38820 80 38920 100
rect 38820 20 38840 80
rect 38900 20 38920 80
rect 38820 0 38920 20
rect 38990 80 39090 130
rect 39330 310 39430 320
rect 39330 250 39350 310
rect 39410 250 39430 310
rect 39330 200 39430 250
rect 39330 130 39350 200
rect 39410 130 39430 200
rect 38990 20 39010 80
rect 39070 20 39090 80
rect 38990 0 39090 20
rect 39160 80 39260 100
rect 39160 20 39180 80
rect 39240 20 39260 80
rect 39160 0 39260 20
rect 39330 80 39430 130
rect 39670 310 39770 320
rect 39670 250 39690 310
rect 39750 250 39770 310
rect 39670 200 39770 250
rect 39670 130 39690 200
rect 39750 130 39770 200
rect 39330 20 39350 80
rect 39410 20 39430 80
rect 39330 0 39430 20
rect 39500 80 39600 100
rect 39500 20 39520 80
rect 39580 20 39600 80
rect 39500 0 39600 20
rect 39670 80 39770 130
rect 40010 310 40110 320
rect 40010 250 40030 310
rect 40090 250 40110 310
rect 40010 200 40110 250
rect 40010 130 40030 200
rect 40090 130 40110 200
rect 39670 20 39690 80
rect 39750 20 39770 80
rect 39670 0 39770 20
rect 39840 80 39940 100
rect 39840 20 39860 80
rect 39920 20 39940 80
rect 39840 0 39940 20
rect 40010 80 40110 130
rect 40350 310 40450 320
rect 40350 250 40370 310
rect 40430 250 40450 310
rect 40350 200 40450 250
rect 40350 130 40370 200
rect 40430 130 40450 200
rect 40010 20 40030 80
rect 40090 20 40110 80
rect 40010 0 40110 20
rect 40180 80 40280 100
rect 40180 20 40200 80
rect 40260 20 40280 80
rect 40180 0 40280 20
rect 40350 80 40450 130
rect 40690 310 40790 320
rect 40690 250 40710 310
rect 40770 250 40790 310
rect 40690 200 40790 250
rect 40690 130 40710 200
rect 40770 130 40790 200
rect 40350 20 40370 80
rect 40430 20 40450 80
rect 40350 0 40450 20
rect 40520 80 40620 100
rect 40520 20 40540 80
rect 40600 20 40620 80
rect 40520 0 40620 20
rect 40690 80 40790 130
rect 41030 310 41130 320
rect 41030 250 41050 310
rect 41110 250 41130 310
rect 41030 200 41130 250
rect 41030 130 41050 200
rect 41110 130 41130 200
rect 40690 20 40710 80
rect 40770 20 40790 80
rect 40690 0 40790 20
rect 40860 80 40960 100
rect 40860 20 40880 80
rect 40940 20 40960 80
rect 40860 0 40960 20
rect 41030 80 41130 130
rect 41370 310 41470 320
rect 41370 250 41390 310
rect 41450 250 41470 310
rect 41370 200 41470 250
rect 41370 130 41390 200
rect 41450 130 41470 200
rect 41030 20 41050 80
rect 41110 20 41130 80
rect 41030 0 41130 20
rect 41200 80 41300 100
rect 41200 20 41220 80
rect 41280 20 41300 80
rect 41200 0 41300 20
rect 41370 80 41470 130
rect 41710 310 41810 320
rect 41710 250 41730 310
rect 41790 250 41810 310
rect 41710 200 41810 250
rect 41710 130 41730 200
rect 41790 130 41810 200
rect 41370 20 41390 80
rect 41450 20 41470 80
rect 41370 0 41470 20
rect 41540 80 41640 100
rect 41540 20 41560 80
rect 41620 20 41640 80
rect 41540 0 41640 20
rect 41710 80 41810 130
rect 42050 310 42150 320
rect 42050 250 42070 310
rect 42130 250 42150 310
rect 42050 200 42150 250
rect 42050 130 42070 200
rect 42130 130 42150 200
rect 41710 20 41730 80
rect 41790 20 41810 80
rect 41710 0 41810 20
rect 41880 80 41980 100
rect 41880 20 41900 80
rect 41960 20 41980 80
rect 41880 0 41980 20
rect 42050 80 42150 130
rect 42390 310 42490 320
rect 42390 250 42410 310
rect 42470 250 42490 310
rect 42390 200 42490 250
rect 42390 130 42410 200
rect 42470 130 42490 200
rect 42050 20 42070 80
rect 42130 20 42150 80
rect 42050 0 42150 20
rect 42220 80 42320 100
rect 42220 20 42240 80
rect 42300 20 42320 80
rect 42220 0 42320 20
rect 42390 80 42490 130
rect 42730 310 42830 320
rect 42730 250 42750 310
rect 42810 250 42830 310
rect 42730 200 42830 250
rect 42730 130 42750 200
rect 42810 130 42830 200
rect 42390 20 42410 80
rect 42470 20 42490 80
rect 42390 0 42490 20
rect 42560 80 42660 100
rect 42560 20 42580 80
rect 42640 20 42660 80
rect 42560 0 42660 20
rect 42730 80 42830 130
rect 43070 310 43170 320
rect 43070 250 43090 310
rect 43150 250 43170 310
rect 43070 200 43170 250
rect 43070 130 43090 200
rect 43150 130 43170 200
rect 42730 20 42750 80
rect 42810 20 42830 80
rect 42730 0 42830 20
rect 42900 80 43000 100
rect 42900 20 42920 80
rect 42980 20 43000 80
rect 42900 0 43000 20
rect 43070 80 43170 130
rect 43410 310 43510 320
rect 43410 250 43430 310
rect 43490 250 43510 310
rect 43410 200 43510 250
rect 43410 130 43430 200
rect 43490 130 43510 200
rect 43070 20 43090 80
rect 43150 20 43170 80
rect 43070 0 43170 20
rect 43240 80 43340 100
rect 43240 20 43260 80
rect 43320 20 43340 80
rect 43240 0 43340 20
rect 43410 80 43510 130
rect 43750 310 43850 320
rect 43750 250 43770 310
rect 43830 250 43850 310
rect 43750 200 43850 250
rect 43750 130 43770 200
rect 43830 130 43850 200
rect 43410 20 43430 80
rect 43490 20 43510 80
rect 43410 0 43510 20
rect 43580 80 43680 100
rect 43580 20 43600 80
rect 43660 20 43680 80
rect 43580 0 43680 20
rect 43750 80 43850 130
rect 44090 310 44190 320
rect 44090 250 44110 310
rect 44170 250 44190 310
rect 44090 200 44190 250
rect 44090 130 44110 200
rect 44170 130 44190 200
rect 43750 20 43770 80
rect 43830 20 43850 80
rect 43750 0 43850 20
rect 43920 80 44020 100
rect 43920 20 43940 80
rect 44000 20 44020 80
rect 43920 0 44020 20
rect 44090 80 44190 130
rect 44430 310 44530 320
rect 44430 250 44450 310
rect 44510 250 44530 310
rect 44430 200 44530 250
rect 44430 130 44450 200
rect 44510 130 44530 200
rect 44090 20 44110 80
rect 44170 20 44190 80
rect 44090 0 44190 20
rect 44260 80 44360 100
rect 44260 20 44280 80
rect 44340 20 44360 80
rect 44260 0 44360 20
rect 44430 80 44530 130
rect 44770 310 44870 320
rect 44770 250 44790 310
rect 44850 250 44870 310
rect 44770 200 44870 250
rect 44770 130 44790 200
rect 44850 130 44870 200
rect 44430 20 44450 80
rect 44510 20 44530 80
rect 44430 0 44530 20
rect 44600 80 44700 100
rect 44600 20 44620 80
rect 44680 20 44700 80
rect 44600 0 44700 20
rect 44770 80 44870 130
rect 45110 310 45210 320
rect 45110 250 45130 310
rect 45190 250 45210 310
rect 45110 200 45210 250
rect 45110 130 45130 200
rect 45190 130 45210 200
rect 44770 20 44790 80
rect 44850 20 44870 80
rect 44770 0 44870 20
rect 44940 80 45040 100
rect 44940 20 44960 80
rect 45020 20 45040 80
rect 44940 0 45040 20
rect 45110 80 45210 130
rect 45450 310 45550 320
rect 45450 250 45470 310
rect 45530 250 45550 310
rect 45450 200 45550 250
rect 45450 130 45470 200
rect 45530 130 45550 200
rect 45110 20 45130 80
rect 45190 20 45210 80
rect 45110 0 45210 20
rect 45280 80 45380 100
rect 45280 20 45300 80
rect 45360 20 45380 80
rect 45280 0 45380 20
rect 45450 80 45550 130
rect 45790 310 45890 320
rect 45790 250 45810 310
rect 45870 250 45890 310
rect 45790 200 45890 250
rect 45790 130 45810 200
rect 45870 130 45890 200
rect 45450 20 45470 80
rect 45530 20 45550 80
rect 45450 0 45550 20
rect 45620 80 45720 100
rect 45620 20 45640 80
rect 45700 20 45720 80
rect 45620 0 45720 20
rect 45790 80 45890 130
rect 46130 310 46230 320
rect 46130 250 46150 310
rect 46210 250 46230 310
rect 46130 200 46230 250
rect 46130 130 46150 200
rect 46210 130 46230 200
rect 45790 20 45810 80
rect 45870 20 45890 80
rect 45790 0 45890 20
rect 45960 80 46060 100
rect 45960 20 45980 80
rect 46040 20 46060 80
rect 45960 0 46060 20
rect 46130 80 46230 130
rect 46470 310 46570 320
rect 46470 250 46490 310
rect 46550 250 46570 310
rect 46470 200 46570 250
rect 46470 130 46490 200
rect 46550 130 46570 200
rect 46130 20 46150 80
rect 46210 20 46230 80
rect 46130 0 46230 20
rect 46300 80 46400 100
rect 46300 20 46320 80
rect 46380 20 46400 80
rect 46300 0 46400 20
rect 46470 80 46570 130
rect 46810 310 46910 320
rect 46810 250 46830 310
rect 46890 250 46910 310
rect 46810 200 46910 250
rect 46810 130 46830 200
rect 46890 130 46910 200
rect 46470 20 46490 80
rect 46550 20 46570 80
rect 46470 0 46570 20
rect 46640 80 46740 100
rect 46640 20 46660 80
rect 46720 20 46740 80
rect 46640 0 46740 20
rect 46810 80 46910 130
rect 47150 310 47250 320
rect 47150 250 47170 310
rect 47230 250 47250 310
rect 47150 200 47250 250
rect 47150 130 47170 200
rect 47230 130 47250 200
rect 46810 20 46830 80
rect 46890 20 46910 80
rect 46810 0 46910 20
rect 46980 80 47080 100
rect 46980 20 47000 80
rect 47060 20 47080 80
rect 46980 0 47080 20
rect 47150 80 47250 130
rect 47490 310 47590 320
rect 47490 250 47510 310
rect 47570 250 47590 310
rect 47490 200 47590 250
rect 47490 130 47510 200
rect 47570 130 47590 200
rect 47150 20 47170 80
rect 47230 20 47250 80
rect 47150 0 47250 20
rect 47320 80 47420 100
rect 47320 20 47340 80
rect 47400 20 47420 80
rect 47320 0 47420 20
rect 47490 80 47590 130
rect 47830 310 47930 320
rect 47830 250 47850 310
rect 47910 250 47930 310
rect 47830 200 47930 250
rect 47830 130 47850 200
rect 47910 130 47930 200
rect 47490 20 47510 80
rect 47570 20 47590 80
rect 47490 0 47590 20
rect 47660 80 47760 100
rect 47660 20 47680 80
rect 47740 20 47760 80
rect 47660 0 47760 20
rect 47830 80 47930 130
rect 48170 310 48270 320
rect 48170 250 48190 310
rect 48250 250 48270 310
rect 48170 200 48270 250
rect 48170 130 48190 200
rect 48250 130 48270 200
rect 47830 20 47850 80
rect 47910 20 47930 80
rect 47830 0 47930 20
rect 48000 80 48100 100
rect 48000 20 48020 80
rect 48080 20 48100 80
rect 48000 0 48100 20
rect 48170 80 48270 130
rect 48510 310 48610 320
rect 48510 250 48530 310
rect 48590 250 48610 310
rect 48510 200 48610 250
rect 48510 130 48530 200
rect 48590 130 48610 200
rect 48170 20 48190 80
rect 48250 20 48270 80
rect 48170 0 48270 20
rect 48340 80 48440 100
rect 48340 20 48360 80
rect 48420 20 48440 80
rect 48340 0 48440 20
rect 48510 80 48610 130
rect 48850 310 48950 320
rect 48850 250 48870 310
rect 48930 250 48950 310
rect 48850 200 48950 250
rect 48850 130 48870 200
rect 48930 130 48950 200
rect 48510 20 48530 80
rect 48590 20 48610 80
rect 48510 0 48610 20
rect 48680 80 48780 100
rect 48680 20 48700 80
rect 48760 20 48780 80
rect 48680 0 48780 20
rect 48850 80 48950 130
rect 49190 310 49290 320
rect 49190 250 49210 310
rect 49270 250 49290 310
rect 49190 200 49290 250
rect 49190 130 49210 200
rect 49270 130 49290 200
rect 48850 20 48870 80
rect 48930 20 48950 80
rect 48850 0 48950 20
rect 49020 80 49120 100
rect 49020 20 49040 80
rect 49100 20 49120 80
rect 49020 0 49120 20
rect 49190 80 49290 130
rect 49530 310 49630 320
rect 49530 250 49550 310
rect 49610 250 49630 310
rect 49530 200 49630 250
rect 49530 130 49550 200
rect 49610 130 49630 200
rect 49190 20 49210 80
rect 49270 20 49290 80
rect 49190 0 49290 20
rect 49360 80 49460 100
rect 49360 20 49380 80
rect 49440 20 49460 80
rect 49360 0 49460 20
rect 49530 80 49630 130
rect 49870 310 49970 320
rect 49870 250 49890 310
rect 49950 250 49970 310
rect 49870 200 49970 250
rect 49870 130 49890 200
rect 49950 130 49970 200
rect 49530 20 49550 80
rect 49610 20 49630 80
rect 49530 0 49630 20
rect 49700 80 49800 100
rect 49700 20 49720 80
rect 49780 20 49800 80
rect 49700 0 49800 20
rect 49870 80 49970 130
rect 50210 310 50310 320
rect 50210 250 50230 310
rect 50290 250 50310 310
rect 50210 200 50310 250
rect 50210 130 50230 200
rect 50290 130 50310 200
rect 49870 20 49890 80
rect 49950 20 49970 80
rect 49870 0 49970 20
rect 50040 80 50140 100
rect 50040 20 50060 80
rect 50120 20 50140 80
rect 50040 0 50140 20
rect 50210 80 50310 130
rect 50550 310 50650 320
rect 50550 250 50570 310
rect 50630 250 50650 310
rect 50550 200 50650 250
rect 50550 130 50570 200
rect 50630 130 50650 200
rect 50210 20 50230 80
rect 50290 20 50310 80
rect 50210 0 50310 20
rect 50380 80 50480 100
rect 50380 20 50400 80
rect 50460 20 50480 80
rect 50380 0 50480 20
rect 50550 80 50650 130
rect 50890 310 50990 320
rect 50890 250 50910 310
rect 50970 250 50990 310
rect 50890 200 50990 250
rect 50890 130 50910 200
rect 50970 130 50990 200
rect 50550 20 50570 80
rect 50630 20 50650 80
rect 50550 0 50650 20
rect 50720 80 50820 100
rect 50720 20 50740 80
rect 50800 20 50820 80
rect 50720 0 50820 20
rect 50890 80 50990 130
rect 51230 310 51330 320
rect 51230 250 51250 310
rect 51310 250 51330 310
rect 51230 200 51330 250
rect 51230 130 51250 200
rect 51310 130 51330 200
rect 50890 20 50910 80
rect 50970 20 50990 80
rect 50890 0 50990 20
rect 51060 80 51160 100
rect 51060 20 51080 80
rect 51140 20 51160 80
rect 51060 0 51160 20
rect 51230 80 51330 130
rect 51570 310 51670 320
rect 51570 250 51590 310
rect 51650 250 51670 310
rect 51570 200 51670 250
rect 51570 130 51590 200
rect 51650 130 51670 200
rect 51230 20 51250 80
rect 51310 20 51330 80
rect 51230 0 51330 20
rect 51400 80 51500 100
rect 51400 20 51420 80
rect 51480 20 51500 80
rect 51400 0 51500 20
rect 51570 80 51670 130
rect 51910 310 52010 320
rect 51910 250 51930 310
rect 51990 250 52010 310
rect 51910 200 52010 250
rect 51910 130 51930 200
rect 51990 130 52010 200
rect 51570 20 51590 80
rect 51650 20 51670 80
rect 51570 0 51670 20
rect 51740 80 51840 100
rect 51740 20 51760 80
rect 51820 20 51840 80
rect 51740 0 51840 20
rect 51910 80 52010 130
rect 52250 310 52350 320
rect 52250 250 52270 310
rect 52330 250 52350 310
rect 52250 200 52350 250
rect 52250 130 52270 200
rect 52330 130 52350 200
rect 51910 20 51930 80
rect 51990 20 52010 80
rect 51910 0 52010 20
rect 52080 80 52180 100
rect 52080 20 52100 80
rect 52160 20 52180 80
rect 52080 0 52180 20
rect 52250 80 52350 130
rect 52590 310 52690 320
rect 52590 250 52610 310
rect 52670 250 52690 310
rect 52590 200 52690 250
rect 52590 130 52610 200
rect 52670 130 52690 200
rect 52250 20 52270 80
rect 52330 20 52350 80
rect 52250 0 52350 20
rect 52420 80 52520 100
rect 52420 20 52440 80
rect 52500 20 52520 80
rect 52420 0 52520 20
rect 52590 80 52690 130
rect 52930 310 53030 320
rect 52930 250 52950 310
rect 53010 250 53030 310
rect 52930 200 53030 250
rect 52930 130 52950 200
rect 53010 130 53030 200
rect 52590 20 52610 80
rect 52670 20 52690 80
rect 52590 0 52690 20
rect 52760 80 52860 100
rect 52760 20 52780 80
rect 52840 20 52860 80
rect 52760 0 52860 20
rect 52930 80 53030 130
rect 53270 310 53370 320
rect 53270 250 53290 310
rect 53350 250 53370 310
rect 53270 200 53370 250
rect 53270 130 53290 200
rect 53350 130 53370 200
rect 52930 20 52950 80
rect 53010 20 53030 80
rect 52930 0 53030 20
rect 53100 80 53200 100
rect 53100 20 53120 80
rect 53180 20 53200 80
rect 53100 0 53200 20
rect 53270 80 53370 130
rect 53610 310 53710 320
rect 53610 250 53630 310
rect 53690 250 53710 310
rect 53610 200 53710 250
rect 53610 130 53630 200
rect 53690 130 53710 200
rect 53270 20 53290 80
rect 53350 20 53370 80
rect 53270 0 53370 20
rect 53440 80 53540 100
rect 53440 20 53460 80
rect 53520 20 53540 80
rect 53440 0 53540 20
rect 53610 80 53710 130
rect 53950 310 54050 320
rect 53950 250 53970 310
rect 54030 250 54050 310
rect 53950 200 54050 250
rect 53950 130 53970 200
rect 54030 130 54050 200
rect 53610 20 53630 80
rect 53690 20 53710 80
rect 53610 0 53710 20
rect 53780 80 53880 100
rect 53780 20 53800 80
rect 53860 20 53880 80
rect 53780 0 53880 20
rect 53950 80 54050 130
rect 54290 310 54390 320
rect 54290 250 54310 310
rect 54370 250 54390 310
rect 54290 200 54390 250
rect 54290 130 54310 200
rect 54370 130 54390 200
rect 53950 20 53970 80
rect 54030 20 54050 80
rect 53950 0 54050 20
rect 54120 80 54220 100
rect 54120 20 54140 80
rect 54200 20 54220 80
rect 54120 0 54220 20
rect 54290 80 54390 130
rect 54630 310 54730 320
rect 54630 250 54650 310
rect 54710 250 54730 310
rect 54630 200 54730 250
rect 54630 130 54650 200
rect 54710 130 54730 200
rect 54290 20 54310 80
rect 54370 20 54390 80
rect 54290 0 54390 20
rect 54460 80 54560 100
rect 54460 20 54480 80
rect 54540 20 54560 80
rect 54460 0 54560 20
rect 54630 80 54730 130
rect 54970 310 55070 320
rect 54970 250 54990 310
rect 55050 250 55070 310
rect 54970 200 55070 250
rect 54970 130 54990 200
rect 55050 130 55070 200
rect 54630 20 54650 80
rect 54710 20 54730 80
rect 54630 0 54730 20
rect 54800 80 54900 100
rect 54800 20 54820 80
rect 54880 20 54900 80
rect 54800 0 54900 20
rect 54970 80 55070 130
rect 55310 310 55410 320
rect 55310 250 55330 310
rect 55390 250 55410 310
rect 55310 200 55410 250
rect 55310 130 55330 200
rect 55390 130 55410 200
rect 54970 20 54990 80
rect 55050 20 55070 80
rect 54970 0 55070 20
rect 55140 80 55240 100
rect 55140 20 55160 80
rect 55220 20 55240 80
rect 55140 0 55240 20
rect 55310 80 55410 130
rect 55650 310 55750 320
rect 55650 250 55670 310
rect 55730 250 55750 310
rect 55650 200 55750 250
rect 55650 130 55670 200
rect 55730 130 55750 200
rect 55310 20 55330 80
rect 55390 20 55410 80
rect 55310 0 55410 20
rect 55480 80 55580 100
rect 55480 20 55500 80
rect 55560 20 55580 80
rect 55480 0 55580 20
rect 55650 80 55750 130
rect 55990 310 56090 320
rect 55990 250 56010 310
rect 56070 250 56090 310
rect 55990 200 56090 250
rect 55990 130 56010 200
rect 56070 130 56090 200
rect 55650 20 55670 80
rect 55730 20 55750 80
rect 55650 0 55750 20
rect 55820 80 55920 100
rect 55820 20 55840 80
rect 55900 20 55920 80
rect 55820 0 55920 20
rect 55990 80 56090 130
rect 56330 310 56430 320
rect 56330 250 56350 310
rect 56410 250 56430 310
rect 56330 200 56430 250
rect 56330 130 56350 200
rect 56410 130 56430 200
rect 55990 20 56010 80
rect 56070 20 56090 80
rect 55990 0 56090 20
rect 56160 80 56260 100
rect 56160 20 56180 80
rect 56240 20 56260 80
rect 56160 0 56260 20
rect 56330 80 56430 130
rect 56670 310 56770 320
rect 56670 250 56690 310
rect 56750 250 56770 310
rect 56670 200 56770 250
rect 56670 130 56690 200
rect 56750 130 56770 200
rect 56330 20 56350 80
rect 56410 20 56430 80
rect 56330 0 56430 20
rect 56500 80 56600 100
rect 56500 20 56520 80
rect 56580 20 56600 80
rect 56500 0 56600 20
rect 56670 80 56770 130
rect 57010 310 57110 320
rect 57010 250 57030 310
rect 57090 250 57110 310
rect 57010 200 57110 250
rect 57010 130 57030 200
rect 57090 130 57110 200
rect 56670 20 56690 80
rect 56750 20 56770 80
rect 56670 0 56770 20
rect 56840 80 56940 100
rect 56840 20 56860 80
rect 56920 20 56940 80
rect 56840 0 56940 20
rect 57010 80 57110 130
rect 57350 310 57450 320
rect 57350 250 57370 310
rect 57430 250 57450 310
rect 57350 200 57450 250
rect 57350 130 57370 200
rect 57430 130 57450 200
rect 57010 20 57030 80
rect 57090 20 57110 80
rect 57010 0 57110 20
rect 57180 80 57280 100
rect 57180 20 57200 80
rect 57260 20 57280 80
rect 57180 0 57280 20
rect 57350 80 57450 130
rect 57690 310 57790 320
rect 57690 250 57710 310
rect 57770 250 57790 310
rect 57690 200 57790 250
rect 57690 130 57710 200
rect 57770 130 57790 200
rect 57350 20 57370 80
rect 57430 20 57450 80
rect 57350 0 57450 20
rect 57520 80 57620 100
rect 57520 20 57540 80
rect 57600 20 57620 80
rect 57520 0 57620 20
rect 57690 80 57790 130
rect 58030 310 58130 320
rect 58030 250 58050 310
rect 58110 250 58130 310
rect 58030 200 58130 250
rect 58030 130 58050 200
rect 58110 130 58130 200
rect 57690 20 57710 80
rect 57770 20 57790 80
rect 57690 0 57790 20
rect 57860 80 57960 100
rect 57860 20 57880 80
rect 57940 20 57960 80
rect 57860 0 57960 20
rect 58030 80 58130 130
rect 58370 310 58470 320
rect 58370 250 58390 310
rect 58450 250 58470 310
rect 58370 200 58470 250
rect 58370 130 58390 200
rect 58450 130 58470 200
rect 58030 20 58050 80
rect 58110 20 58130 80
rect 58030 0 58130 20
rect 58200 80 58300 100
rect 58200 20 58220 80
rect 58280 20 58300 80
rect 58200 0 58300 20
rect 58370 80 58470 130
rect 58710 310 58810 320
rect 58710 250 58730 310
rect 58790 250 58810 310
rect 58710 200 58810 250
rect 58710 130 58730 200
rect 58790 130 58810 200
rect 58370 20 58390 80
rect 58450 20 58470 80
rect 58370 0 58470 20
rect 58540 80 58640 100
rect 58540 20 58560 80
rect 58620 20 58640 80
rect 58540 0 58640 20
rect 58710 80 58810 130
rect 59050 310 59150 320
rect 59050 250 59070 310
rect 59130 250 59150 310
rect 59050 200 59150 250
rect 59050 130 59070 200
rect 59130 130 59150 200
rect 58710 20 58730 80
rect 58790 20 58810 80
rect 58710 0 58810 20
rect 58880 80 58980 100
rect 58880 20 58900 80
rect 58960 20 58980 80
rect 58880 0 58980 20
rect 59050 80 59150 130
rect 59050 20 59070 80
rect 59130 20 59150 80
rect 59050 0 59150 20
rect 59220 80 59320 100
rect 59220 20 59240 80
rect 59300 20 59320 80
rect 59220 0 59320 20
rect 180 -120 200 -60
rect 260 -120 280 -60
rect 180 -180 280 -120
rect 510 -60 620 -40
rect 510 -120 530 -60
rect 600 -120 620 -60
rect 510 -140 620 -120
rect 680 -60 790 -40
rect 680 -120 700 -60
rect 770 -120 790 -60
rect 680 -140 790 -120
rect 850 -60 960 -40
rect 850 -120 870 -60
rect 940 -120 960 -60
rect 850 -140 960 -120
rect 1020 -60 1130 -40
rect 1020 -120 1040 -60
rect 1110 -120 1130 -60
rect 1020 -140 1130 -120
rect 1580 -60 1690 -40
rect 1580 -120 1600 -60
rect 1670 -120 1690 -60
rect 1580 -140 1690 -120
rect 1750 -60 1860 -40
rect 1750 -120 1770 -60
rect 1840 -120 1860 -60
rect 1750 -140 1860 -120
rect 1920 -60 2030 -40
rect 1920 -120 1940 -60
rect 2010 -120 2030 -60
rect 1920 -140 2030 -120
rect 2090 -60 2200 -40
rect 2090 -120 2110 -60
rect 2180 -120 2200 -60
rect 2090 -140 2200 -120
rect 2260 -60 2370 -40
rect 2260 -120 2280 -60
rect 2350 -120 2370 -60
rect 2260 -140 2370 -120
rect 2430 -60 2540 -40
rect 2430 -120 2450 -60
rect 2520 -120 2540 -60
rect 2430 -140 2540 -120
rect 2600 -60 2710 -40
rect 2600 -120 2620 -60
rect 2690 -120 2710 -60
rect 2600 -140 2710 -120
rect 2770 -60 2880 -40
rect 2770 -120 2790 -60
rect 2860 -120 2880 -60
rect 2770 -140 2880 -120
rect 2940 -60 3050 -40
rect 2940 -120 2960 -60
rect 3030 -120 3050 -60
rect 2940 -140 3050 -120
rect 3110 -60 3220 -40
rect 3110 -120 3130 -60
rect 3200 -120 3220 -60
rect 3110 -140 3220 -120
rect 3280 -60 3390 -40
rect 3280 -120 3300 -60
rect 3370 -120 3390 -60
rect 3280 -140 3390 -120
rect 3450 -60 3560 -40
rect 3450 -120 3470 -60
rect 3540 -120 3560 -60
rect 3450 -140 3560 -120
rect 3620 -60 3730 -40
rect 3620 -120 3640 -60
rect 3710 -120 3730 -60
rect 3620 -140 3730 -120
rect 3790 -60 3900 -40
rect 3790 -120 3810 -60
rect 3880 -120 3900 -60
rect 3790 -140 3900 -120
rect 3960 -60 4070 -40
rect 3960 -120 3980 -60
rect 4050 -120 4070 -60
rect 3960 -140 4070 -120
rect 4130 -60 4240 -40
rect 4130 -120 4150 -60
rect 4220 -120 4240 -60
rect 4130 -140 4240 -120
rect 4600 -60 4710 -40
rect 4600 -120 4620 -60
rect 4690 -120 4710 -60
rect 4600 -140 4710 -120
rect 4770 -60 4880 -40
rect 4770 -120 4790 -60
rect 4860 -120 4880 -60
rect 4770 -140 4880 -120
rect 4940 -60 5050 -40
rect 4940 -120 4960 -60
rect 5030 -120 5050 -60
rect 4940 -140 5050 -120
rect 5110 -60 5220 -40
rect 5110 -120 5130 -60
rect 5200 -120 5220 -60
rect 5110 -140 5220 -120
rect 5280 -60 5390 -40
rect 5280 -120 5300 -60
rect 5370 -120 5390 -60
rect 5280 -140 5390 -120
rect 5450 -60 5560 -40
rect 5450 -120 5470 -60
rect 5540 -120 5560 -60
rect 5450 -140 5560 -120
rect 5620 -60 5730 -40
rect 5620 -120 5640 -60
rect 5710 -120 5730 -60
rect 5620 -140 5730 -120
rect 5790 -60 5900 -40
rect 5790 -120 5810 -60
rect 5880 -120 5900 -60
rect 5790 -140 5900 -120
rect 5960 -60 6070 -40
rect 5960 -120 5980 -60
rect 6050 -120 6070 -60
rect 5960 -140 6070 -120
rect 6130 -60 6240 -40
rect 6130 -120 6150 -60
rect 6220 -120 6240 -60
rect 6130 -140 6240 -120
rect 6300 -60 6410 -40
rect 6300 -120 6320 -60
rect 6390 -120 6410 -60
rect 6300 -140 6410 -120
rect 6470 -60 6580 -40
rect 6470 -120 6490 -60
rect 6560 -120 6580 -60
rect 6470 -140 6580 -120
rect 6640 -60 6750 -40
rect 6640 -120 6660 -60
rect 6730 -120 6750 -60
rect 6640 -140 6750 -120
rect 6810 -60 6920 -40
rect 6810 -120 6830 -60
rect 6900 -120 6920 -60
rect 6810 -140 6920 -120
rect 6980 -60 7090 -40
rect 6980 -120 7000 -60
rect 7070 -120 7090 -60
rect 6980 -140 7090 -120
rect 7150 -60 7260 -40
rect 7150 -120 7170 -60
rect 7240 -120 7260 -60
rect 7150 -140 7260 -120
rect 7320 -60 7430 -40
rect 7320 -120 7340 -60
rect 7410 -120 7430 -60
rect 7320 -140 7430 -120
rect 7490 -60 7600 -40
rect 7490 -120 7510 -60
rect 7580 -120 7600 -60
rect 7490 -140 7600 -120
rect 7660 -60 7770 -40
rect 7660 -120 7680 -60
rect 7750 -120 7770 -60
rect 7660 -140 7770 -120
rect 7830 -60 7940 -40
rect 7830 -120 7850 -60
rect 7920 -120 7940 -60
rect 7830 -140 7940 -120
rect 8000 -60 8110 -40
rect 8000 -120 8020 -60
rect 8090 -120 8110 -60
rect 8000 -140 8110 -120
rect 8170 -60 8280 -40
rect 8170 -120 8190 -60
rect 8260 -120 8280 -60
rect 8170 -140 8280 -120
rect 8340 -60 8450 -40
rect 8340 -120 8360 -60
rect 8430 -120 8450 -60
rect 8340 -140 8450 -120
rect 8510 -60 8620 -40
rect 8510 -120 8530 -60
rect 8600 -120 8620 -60
rect 8510 -140 8620 -120
rect 8680 -60 8790 -40
rect 8680 -120 8700 -60
rect 8770 -120 8790 -60
rect 8680 -140 8790 -120
rect 8850 -60 8960 -40
rect 8850 -120 8870 -60
rect 8940 -120 8960 -60
rect 8850 -140 8960 -120
rect 9020 -60 9130 -40
rect 9020 -120 9040 -60
rect 9110 -120 9130 -60
rect 9020 -140 9130 -120
rect 9190 -60 9300 -40
rect 9190 -120 9210 -60
rect 9280 -120 9300 -60
rect 9190 -140 9300 -120
rect 9360 -60 9470 -40
rect 9360 -120 9380 -60
rect 9450 -120 9470 -60
rect 9360 -140 9470 -120
rect 9530 -60 9640 -40
rect 9530 -120 9550 -60
rect 9620 -120 9640 -60
rect 9530 -140 9640 -120
rect 9700 -60 9810 -40
rect 9700 -120 9720 -60
rect 9790 -120 9810 -60
rect 9700 -140 9810 -120
rect 9870 -60 9980 -40
rect 9870 -120 9890 -60
rect 9960 -120 9980 -60
rect 9870 -140 9980 -120
rect 10040 -60 10150 -40
rect 10040 -120 10060 -60
rect 10130 -120 10150 -60
rect 10040 -140 10150 -120
rect 10210 -60 10320 -40
rect 10210 -120 10230 -60
rect 10300 -120 10320 -60
rect 10210 -140 10320 -120
rect 10380 -60 10490 -40
rect 10380 -120 10400 -60
rect 10470 -120 10490 -60
rect 10380 -140 10490 -120
rect 10550 -60 10660 -40
rect 10550 -120 10570 -60
rect 10640 -120 10660 -60
rect 10550 -140 10660 -120
rect 10720 -60 10830 -40
rect 10720 -120 10740 -60
rect 10810 -120 10830 -60
rect 10720 -140 10830 -120
rect 10890 -60 11000 -40
rect 10890 -120 10910 -60
rect 10980 -120 11000 -60
rect 10890 -140 11000 -120
rect 11060 -60 11170 -40
rect 11060 -120 11080 -60
rect 11150 -120 11170 -60
rect 11060 -140 11170 -120
rect 11230 -60 11340 -40
rect 11230 -120 11250 -60
rect 11320 -120 11340 -60
rect 11230 -140 11340 -120
rect 11400 -60 11510 -40
rect 11400 -120 11420 -60
rect 11490 -120 11510 -60
rect 11400 -140 11510 -120
rect 11570 -60 11680 -40
rect 11570 -120 11590 -60
rect 11660 -120 11680 -60
rect 11570 -140 11680 -120
rect 11740 -60 11850 -40
rect 11740 -120 11760 -60
rect 11830 -120 11850 -60
rect 11740 -140 11850 -120
rect 11910 -60 12020 -40
rect 11910 -120 11930 -60
rect 12000 -120 12020 -60
rect 11910 -140 12020 -120
rect 12080 -60 12190 -40
rect 12080 -120 12100 -60
rect 12170 -120 12190 -60
rect 12080 -140 12190 -120
rect 12250 -60 12360 -40
rect 12250 -120 12270 -60
rect 12340 -120 12360 -60
rect 12250 -140 12360 -120
rect 12420 -60 12530 -40
rect 12420 -120 12440 -60
rect 12510 -120 12530 -60
rect 12420 -140 12530 -120
rect 12590 -60 12700 -40
rect 12590 -120 12610 -60
rect 12680 -120 12700 -60
rect 12590 -140 12700 -120
rect 12760 -60 12870 -40
rect 12760 -120 12780 -60
rect 12850 -120 12870 -60
rect 12760 -140 12870 -120
rect 12930 -60 13040 -40
rect 12930 -120 12950 -60
rect 13020 -120 13040 -60
rect 12930 -140 13040 -120
rect 13100 -60 13210 -40
rect 13100 -120 13120 -60
rect 13190 -120 13210 -60
rect 13100 -140 13210 -120
rect 13270 -60 13380 -40
rect 13270 -120 13290 -60
rect 13360 -120 13380 -60
rect 13270 -140 13380 -120
rect 13440 -60 13550 -40
rect 13440 -120 13460 -60
rect 13530 -120 13550 -60
rect 13440 -140 13550 -120
rect 13610 -60 13720 -40
rect 13610 -120 13630 -60
rect 13700 -120 13720 -60
rect 13610 -140 13720 -120
rect 13780 -60 13890 -40
rect 13780 -120 13800 -60
rect 13870 -120 13890 -60
rect 13780 -140 13890 -120
rect 13950 -60 14060 -40
rect 13950 -120 13970 -60
rect 14040 -120 14060 -60
rect 13950 -140 14060 -120
rect 14120 -60 14230 -40
rect 14120 -120 14140 -60
rect 14210 -120 14230 -60
rect 14120 -140 14230 -120
rect 14290 -60 14400 -40
rect 14290 -120 14310 -60
rect 14380 -120 14400 -60
rect 14290 -140 14400 -120
rect 14460 -60 14570 -40
rect 14460 -120 14480 -60
rect 14550 -120 14570 -60
rect 14460 -140 14570 -120
rect 14630 -60 14740 -40
rect 14630 -120 14650 -60
rect 14720 -120 14740 -60
rect 14630 -140 14740 -120
rect 14800 -60 14910 -40
rect 14800 -120 14820 -60
rect 14890 -120 14910 -60
rect 14800 -140 14910 -120
rect 14970 -60 15080 -40
rect 14970 -120 14990 -60
rect 15060 -120 15080 -60
rect 14970 -140 15080 -120
rect 15140 -60 15250 -40
rect 15140 -120 15160 -60
rect 15230 -120 15250 -60
rect 15140 -140 15250 -120
rect 15310 -60 15420 -40
rect 15310 -120 15330 -60
rect 15400 -120 15420 -60
rect 15310 -140 15420 -120
rect 15780 -60 15890 -40
rect 15780 -120 15800 -60
rect 15870 -120 15890 -60
rect 15780 -140 15890 -120
rect 15950 -60 16060 -40
rect 15950 -120 15970 -60
rect 16040 -120 16060 -60
rect 15950 -140 16060 -120
rect 16120 -60 16230 -40
rect 16120 -120 16140 -60
rect 16210 -120 16230 -60
rect 16120 -140 16230 -120
rect 16290 -60 16400 -40
rect 16290 -120 16310 -60
rect 16380 -120 16400 -60
rect 16290 -140 16400 -120
rect 16460 -60 16570 -40
rect 16460 -120 16480 -60
rect 16550 -120 16570 -60
rect 16460 -140 16570 -120
rect 16630 -60 16740 -40
rect 16630 -120 16650 -60
rect 16720 -120 16740 -60
rect 16630 -140 16740 -120
rect 16800 -60 16910 -40
rect 16800 -120 16820 -60
rect 16890 -120 16910 -60
rect 16800 -140 16910 -120
rect 16970 -60 17080 -40
rect 16970 -120 16990 -60
rect 17060 -120 17080 -60
rect 16970 -140 17080 -120
rect 17140 -60 17250 -40
rect 17140 -120 17160 -60
rect 17230 -120 17250 -60
rect 17140 -140 17250 -120
rect 17310 -60 17420 -40
rect 17310 -120 17330 -60
rect 17400 -120 17420 -60
rect 17310 -140 17420 -120
rect 17480 -60 17590 -40
rect 17480 -120 17500 -60
rect 17570 -120 17590 -60
rect 17480 -140 17590 -120
rect 17650 -60 17760 -40
rect 17650 -120 17670 -60
rect 17740 -120 17760 -60
rect 17650 -140 17760 -120
rect 17820 -60 17930 -40
rect 17820 -120 17840 -60
rect 17910 -120 17930 -60
rect 17820 -140 17930 -120
rect 17990 -60 18100 -40
rect 17990 -120 18010 -60
rect 18080 -120 18100 -60
rect 17990 -140 18100 -120
rect 18160 -60 18270 -40
rect 18160 -120 18180 -60
rect 18250 -120 18270 -60
rect 18160 -140 18270 -120
rect 18330 -60 18440 -40
rect 18330 -120 18350 -60
rect 18420 -120 18440 -60
rect 18330 -140 18440 -120
rect 18500 -60 18610 -40
rect 18500 -120 18520 -60
rect 18590 -120 18610 -60
rect 18500 -140 18610 -120
rect 18670 -60 18780 -40
rect 18670 -120 18690 -60
rect 18760 -120 18780 -60
rect 18670 -140 18780 -120
rect 18840 -60 18950 -40
rect 18840 -120 18860 -60
rect 18930 -120 18950 -60
rect 18840 -140 18950 -120
rect 19010 -60 19120 -40
rect 19010 -120 19030 -60
rect 19100 -120 19120 -60
rect 19010 -140 19120 -120
rect 19180 -60 19290 -40
rect 19180 -120 19200 -60
rect 19270 -120 19290 -60
rect 19180 -140 19290 -120
rect 19350 -60 19460 -40
rect 19350 -120 19370 -60
rect 19440 -120 19460 -60
rect 19350 -140 19460 -120
rect 19520 -60 19630 -40
rect 19520 -120 19540 -60
rect 19610 -120 19630 -60
rect 19520 -140 19630 -120
rect 19690 -60 19800 -40
rect 19690 -120 19710 -60
rect 19780 -120 19800 -60
rect 19690 -140 19800 -120
rect 19860 -60 19970 -40
rect 19860 -120 19880 -60
rect 19950 -120 19970 -60
rect 19860 -140 19970 -120
rect 20030 -60 20140 -40
rect 20030 -120 20050 -60
rect 20120 -120 20140 -60
rect 20030 -140 20140 -120
rect 20200 -60 20310 -40
rect 20200 -120 20220 -60
rect 20290 -120 20310 -60
rect 20200 -140 20310 -120
rect 20370 -60 20480 -40
rect 20370 -120 20390 -60
rect 20460 -120 20480 -60
rect 20370 -140 20480 -120
rect 20540 -60 20650 -40
rect 20540 -120 20560 -60
rect 20630 -120 20650 -60
rect 20540 -140 20650 -120
rect 20710 -60 20820 -40
rect 20710 -120 20730 -60
rect 20800 -120 20820 -60
rect 20710 -140 20820 -120
rect 20880 -60 20990 -40
rect 20880 -120 20900 -60
rect 20970 -120 20990 -60
rect 20880 -140 20990 -120
rect 21050 -60 21160 -40
rect 21050 -120 21070 -60
rect 21140 -120 21160 -60
rect 21050 -140 21160 -120
rect 21220 -60 21330 -40
rect 21220 -120 21240 -60
rect 21310 -120 21330 -60
rect 21220 -140 21330 -120
rect 21390 -60 21500 -40
rect 21390 -120 21410 -60
rect 21480 -120 21500 -60
rect 21390 -140 21500 -120
rect 21560 -60 21670 -40
rect 21560 -120 21580 -60
rect 21650 -120 21670 -60
rect 21560 -140 21670 -120
rect 21730 -60 21840 -40
rect 21730 -120 21750 -60
rect 21820 -120 21840 -60
rect 21730 -140 21840 -120
rect 21900 -60 22010 -40
rect 21900 -120 21920 -60
rect 21990 -120 22010 -60
rect 21900 -140 22010 -120
rect 22070 -60 22180 -40
rect 22070 -120 22090 -60
rect 22160 -120 22180 -60
rect 22070 -140 22180 -120
rect 22240 -60 22350 -40
rect 22240 -120 22260 -60
rect 22330 -120 22350 -60
rect 22240 -140 22350 -120
rect 22410 -60 22520 -40
rect 22410 -120 22430 -60
rect 22500 -120 22520 -60
rect 22410 -140 22520 -120
rect 22580 -60 22690 -40
rect 22580 -120 22600 -60
rect 22670 -120 22690 -60
rect 22580 -140 22690 -120
rect 22750 -60 22860 -40
rect 22750 -120 22770 -60
rect 22840 -120 22860 -60
rect 22750 -140 22860 -120
rect 22920 -60 23030 -40
rect 22920 -120 22940 -60
rect 23010 -120 23030 -60
rect 22920 -140 23030 -120
rect 23090 -60 23200 -40
rect 23090 -120 23110 -60
rect 23180 -120 23200 -60
rect 23090 -140 23200 -120
rect 23260 -60 23370 -40
rect 23260 -120 23280 -60
rect 23350 -120 23370 -60
rect 23260 -140 23370 -120
rect 23430 -60 23540 -40
rect 23430 -120 23450 -60
rect 23520 -120 23540 -60
rect 23430 -140 23540 -120
rect 23600 -60 23710 -40
rect 23600 -120 23620 -60
rect 23690 -120 23710 -60
rect 23600 -140 23710 -120
rect 23770 -60 23880 -40
rect 23770 -120 23790 -60
rect 23860 -120 23880 -60
rect 23770 -140 23880 -120
rect 23940 -60 24050 -40
rect 23940 -120 23960 -60
rect 24030 -120 24050 -60
rect 23940 -140 24050 -120
rect 24110 -60 24220 -40
rect 24110 -120 24130 -60
rect 24200 -120 24220 -60
rect 24110 -140 24220 -120
rect 24280 -60 24390 -40
rect 24280 -120 24300 -60
rect 24370 -120 24390 -60
rect 24280 -140 24390 -120
rect 24450 -60 24560 -40
rect 24450 -120 24470 -60
rect 24540 -120 24560 -60
rect 24450 -140 24560 -120
rect 24620 -60 24730 -40
rect 24620 -120 24640 -60
rect 24710 -120 24730 -60
rect 24620 -140 24730 -120
rect 24790 -60 24900 -40
rect 24790 -120 24810 -60
rect 24880 -120 24900 -60
rect 24790 -140 24900 -120
rect 24960 -60 25070 -40
rect 24960 -120 24980 -60
rect 25050 -120 25070 -60
rect 24960 -140 25070 -120
rect 25130 -60 25240 -40
rect 25130 -120 25150 -60
rect 25220 -120 25240 -60
rect 25130 -140 25240 -120
rect 25300 -60 25410 -40
rect 25300 -120 25320 -60
rect 25390 -120 25410 -60
rect 25300 -140 25410 -120
rect 25470 -60 25580 -40
rect 25470 -120 25490 -60
rect 25560 -120 25580 -60
rect 25470 -140 25580 -120
rect 25640 -60 25750 -40
rect 25640 -120 25660 -60
rect 25730 -120 25750 -60
rect 25640 -140 25750 -120
rect 25810 -60 25920 -40
rect 25810 -120 25830 -60
rect 25900 -120 25920 -60
rect 25810 -140 25920 -120
rect 25980 -60 26090 -40
rect 25980 -120 26000 -60
rect 26070 -120 26090 -60
rect 25980 -140 26090 -120
rect 26150 -60 26260 -40
rect 26150 -120 26170 -60
rect 26240 -120 26260 -60
rect 26150 -140 26260 -120
rect 26320 -60 26430 -40
rect 26320 -120 26340 -60
rect 26410 -120 26430 -60
rect 26320 -140 26430 -120
rect 26490 -60 26600 -40
rect 26490 -120 26510 -60
rect 26580 -120 26600 -60
rect 26490 -140 26600 -120
rect 26660 -60 26770 -40
rect 26660 -120 26680 -60
rect 26750 -120 26770 -60
rect 26660 -140 26770 -120
rect 26830 -60 26940 -40
rect 26830 -120 26850 -60
rect 26920 -120 26940 -60
rect 26830 -140 26940 -120
rect 27000 -60 27110 -40
rect 27000 -120 27020 -60
rect 27090 -120 27110 -60
rect 27000 -140 27110 -120
rect 27170 -60 27280 -40
rect 27170 -120 27190 -60
rect 27260 -120 27280 -60
rect 27170 -140 27280 -120
rect 27340 -60 27450 -40
rect 27340 -120 27360 -60
rect 27430 -120 27450 -60
rect 27340 -140 27450 -120
rect 27510 -60 27620 -40
rect 27510 -120 27530 -60
rect 27600 -120 27620 -60
rect 27510 -140 27620 -120
rect 27680 -60 27790 -40
rect 27680 -120 27700 -60
rect 27770 -120 27790 -60
rect 27680 -140 27790 -120
rect 27850 -60 27960 -40
rect 27850 -120 27870 -60
rect 27940 -120 27960 -60
rect 27850 -140 27960 -120
rect 28020 -60 28130 -40
rect 28020 -120 28040 -60
rect 28110 -120 28130 -60
rect 28020 -140 28130 -120
rect 28190 -60 28300 -40
rect 28190 -120 28210 -60
rect 28280 -120 28300 -60
rect 28190 -140 28300 -120
rect 28360 -60 28470 -40
rect 28360 -120 28380 -60
rect 28450 -120 28470 -60
rect 28360 -140 28470 -120
rect 28530 -60 28640 -40
rect 28530 -120 28550 -60
rect 28620 -120 28640 -60
rect 28530 -140 28640 -120
rect 28700 -60 28810 -40
rect 28700 -120 28720 -60
rect 28790 -120 28810 -60
rect 28700 -140 28810 -120
rect 28870 -60 28980 -40
rect 28870 -120 28890 -60
rect 28960 -120 28980 -60
rect 28870 -140 28980 -120
rect 29040 -60 29150 -40
rect 29040 -120 29060 -60
rect 29130 -120 29150 -60
rect 29040 -140 29150 -120
rect 29210 -60 29320 -40
rect 29210 -120 29230 -60
rect 29300 -120 29320 -60
rect 29210 -140 29320 -120
rect 29380 -60 29490 -40
rect 29380 -120 29400 -60
rect 29470 -120 29490 -60
rect 29380 -140 29490 -120
rect 29550 -60 29660 -40
rect 29550 -120 29570 -60
rect 29640 -120 29660 -60
rect 29550 -140 29660 -120
rect 29720 -60 29830 -40
rect 29720 -120 29740 -60
rect 29810 -120 29830 -60
rect 29720 -140 29830 -120
rect 29890 -60 30000 -40
rect 29890 -120 29910 -60
rect 29980 -120 30000 -60
rect 29890 -140 30000 -120
rect 30060 -60 30170 -40
rect 30060 -120 30080 -60
rect 30150 -120 30170 -60
rect 30060 -140 30170 -120
rect 30230 -60 30340 -40
rect 30230 -120 30250 -60
rect 30320 -120 30340 -60
rect 30230 -140 30340 -120
rect 30400 -60 30510 -40
rect 30400 -120 30420 -60
rect 30490 -120 30510 -60
rect 30400 -140 30510 -120
rect 30570 -60 30680 -40
rect 30570 -120 30590 -60
rect 30660 -120 30680 -60
rect 30570 -140 30680 -120
rect 30740 -60 30850 -40
rect 30740 -120 30760 -60
rect 30830 -120 30850 -60
rect 30740 -140 30850 -120
rect 30910 -60 31020 -40
rect 30910 -120 30930 -60
rect 31000 -120 31020 -60
rect 30910 -140 31020 -120
rect 31080 -60 31190 -40
rect 31080 -120 31100 -60
rect 31170 -120 31190 -60
rect 31080 -140 31190 -120
rect 31250 -60 31360 -40
rect 31250 -120 31270 -60
rect 31340 -120 31360 -60
rect 31250 -140 31360 -120
rect 31420 -60 31530 -40
rect 31420 -120 31440 -60
rect 31510 -120 31530 -60
rect 31420 -140 31530 -120
rect 31590 -60 31700 -40
rect 31590 -120 31610 -60
rect 31680 -120 31700 -60
rect 31590 -140 31700 -120
rect 31760 -60 31870 -40
rect 31760 -120 31780 -60
rect 31850 -120 31870 -60
rect 31760 -140 31870 -120
rect 31930 -60 32040 -40
rect 31930 -120 31950 -60
rect 32020 -120 32040 -60
rect 31930 -140 32040 -120
rect 32100 -60 32210 -40
rect 32100 -120 32120 -60
rect 32190 -120 32210 -60
rect 32100 -140 32210 -120
rect 32270 -60 32380 -40
rect 32270 -120 32290 -60
rect 32360 -120 32380 -60
rect 32270 -140 32380 -120
rect 32440 -60 32550 -40
rect 32440 -120 32460 -60
rect 32530 -120 32550 -60
rect 32440 -140 32550 -120
rect 32610 -60 32720 -40
rect 32610 -120 32630 -60
rect 32700 -120 32720 -60
rect 32610 -140 32720 -120
rect 32780 -60 32890 -40
rect 32780 -120 32800 -60
rect 32870 -120 32890 -60
rect 32780 -140 32890 -120
rect 32950 -60 33060 -40
rect 32950 -120 32970 -60
rect 33040 -120 33060 -60
rect 32950 -140 33060 -120
rect 33120 -60 33230 -40
rect 33120 -120 33140 -60
rect 33210 -120 33230 -60
rect 33120 -140 33230 -120
rect 33290 -60 33400 -40
rect 33290 -120 33310 -60
rect 33380 -120 33400 -60
rect 33290 -140 33400 -120
rect 33460 -60 33570 -40
rect 33460 -120 33480 -60
rect 33550 -120 33570 -60
rect 33460 -140 33570 -120
rect 33630 -60 33740 -40
rect 33630 -120 33650 -60
rect 33720 -120 33740 -60
rect 33630 -140 33740 -120
rect 33800 -60 33910 -40
rect 33800 -120 33820 -60
rect 33890 -120 33910 -60
rect 33800 -140 33910 -120
rect 33970 -60 34080 -40
rect 33970 -120 33990 -60
rect 34060 -120 34080 -60
rect 33970 -140 34080 -120
rect 34140 -60 34250 -40
rect 34140 -120 34160 -60
rect 34230 -120 34250 -60
rect 34140 -140 34250 -120
rect 34310 -60 34420 -40
rect 34310 -120 34330 -60
rect 34400 -120 34420 -60
rect 34310 -140 34420 -120
rect 34480 -60 34590 -40
rect 34480 -120 34500 -60
rect 34570 -120 34590 -60
rect 34480 -140 34590 -120
rect 34650 -60 34760 -40
rect 34650 -120 34670 -60
rect 34740 -120 34760 -60
rect 34650 -140 34760 -120
rect 34820 -60 34930 -40
rect 34820 -120 34840 -60
rect 34910 -120 34930 -60
rect 34820 -140 34930 -120
rect 34990 -60 35100 -40
rect 34990 -120 35010 -60
rect 35080 -120 35100 -60
rect 34990 -140 35100 -120
rect 35160 -60 35270 -40
rect 35160 -120 35180 -60
rect 35250 -120 35270 -60
rect 35160 -140 35270 -120
rect 35330 -60 35440 -40
rect 35330 -120 35350 -60
rect 35420 -120 35440 -60
rect 35330 -140 35440 -120
rect 35500 -60 35610 -40
rect 35500 -120 35520 -60
rect 35590 -120 35610 -60
rect 35500 -140 35610 -120
rect 35670 -60 35780 -40
rect 35670 -120 35690 -60
rect 35760 -120 35780 -60
rect 35670 -140 35780 -120
rect 35840 -60 35950 -40
rect 35840 -120 35860 -60
rect 35930 -120 35950 -60
rect 35840 -140 35950 -120
rect 36010 -60 36120 -40
rect 36010 -120 36030 -60
rect 36100 -120 36120 -60
rect 36010 -140 36120 -120
rect 36180 -60 36290 -40
rect 36180 -120 36200 -60
rect 36270 -120 36290 -60
rect 36180 -140 36290 -120
rect 36350 -60 36460 -40
rect 36350 -120 36370 -60
rect 36440 -120 36460 -60
rect 36350 -140 36460 -120
rect 36520 -60 36630 -40
rect 36520 -120 36540 -60
rect 36610 -120 36630 -60
rect 36520 -140 36630 -120
rect 36690 -60 36800 -40
rect 36690 -120 36710 -60
rect 36780 -120 36800 -60
rect 36690 -140 36800 -120
rect 36860 -60 36970 -40
rect 36860 -120 36880 -60
rect 36950 -120 36970 -60
rect 36860 -140 36970 -120
rect 37030 -60 37140 -40
rect 37030 -120 37050 -60
rect 37120 -120 37140 -60
rect 37030 -140 37140 -120
rect 37200 -60 37310 -40
rect 37200 -120 37220 -60
rect 37290 -120 37310 -60
rect 37200 -140 37310 -120
rect 37370 -60 37480 -40
rect 37370 -120 37390 -60
rect 37460 -120 37480 -60
rect 37370 -140 37480 -120
rect 37540 -60 37650 -40
rect 37540 -120 37560 -60
rect 37630 -120 37650 -60
rect 37540 -140 37650 -120
rect 37710 -60 37820 -40
rect 37710 -120 37730 -60
rect 37800 -120 37820 -60
rect 37710 -140 37820 -120
rect 37880 -60 37990 -40
rect 37880 -120 37900 -60
rect 37970 -120 37990 -60
rect 37880 -140 37990 -120
rect 38050 -60 38160 -40
rect 38050 -120 38070 -60
rect 38140 -120 38160 -60
rect 38050 -140 38160 -120
rect 38220 -60 38330 -40
rect 38220 -120 38240 -60
rect 38310 -120 38330 -60
rect 38220 -140 38330 -120
rect 38390 -60 38500 -40
rect 38390 -120 38410 -60
rect 38480 -120 38500 -60
rect 38390 -140 38500 -120
rect 38560 -60 38670 -40
rect 38560 -120 38580 -60
rect 38650 -120 38670 -60
rect 38560 -140 38670 -120
rect 38730 -60 38840 -40
rect 38730 -120 38750 -60
rect 38820 -120 38840 -60
rect 38730 -140 38840 -120
rect 38900 -60 39010 -40
rect 38900 -120 38920 -60
rect 38990 -120 39010 -60
rect 38900 -140 39010 -120
rect 39070 -60 39180 -40
rect 39070 -120 39090 -60
rect 39160 -120 39180 -60
rect 39070 -140 39180 -120
rect 39240 -60 39350 -40
rect 39240 -120 39260 -60
rect 39330 -120 39350 -60
rect 39240 -140 39350 -120
rect 39410 -60 39520 -40
rect 39410 -120 39430 -60
rect 39500 -120 39520 -60
rect 39410 -140 39520 -120
rect 39580 -60 39690 -40
rect 39580 -120 39600 -60
rect 39670 -120 39690 -60
rect 39580 -140 39690 -120
rect 39750 -60 39860 -40
rect 39750 -120 39770 -60
rect 39840 -120 39860 -60
rect 39750 -140 39860 -120
rect 39920 -60 40030 -40
rect 39920 -120 39940 -60
rect 40010 -120 40030 -60
rect 39920 -140 40030 -120
rect 40090 -60 40200 -40
rect 40090 -120 40110 -60
rect 40180 -120 40200 -60
rect 40090 -140 40200 -120
rect 40260 -60 40370 -40
rect 40260 -120 40280 -60
rect 40350 -120 40370 -60
rect 40260 -140 40370 -120
rect 40430 -60 40540 -40
rect 40430 -120 40450 -60
rect 40520 -120 40540 -60
rect 40430 -140 40540 -120
rect 40600 -60 40710 -40
rect 40600 -120 40620 -60
rect 40690 -120 40710 -60
rect 40600 -140 40710 -120
rect 40770 -60 40880 -40
rect 40770 -120 40790 -60
rect 40860 -120 40880 -60
rect 40770 -140 40880 -120
rect 40940 -60 41050 -40
rect 40940 -120 40960 -60
rect 41030 -120 41050 -60
rect 40940 -140 41050 -120
rect 41110 -60 41220 -40
rect 41110 -120 41130 -60
rect 41200 -120 41220 -60
rect 41110 -140 41220 -120
rect 41280 -60 41390 -40
rect 41280 -120 41300 -60
rect 41370 -120 41390 -60
rect 41280 -140 41390 -120
rect 41450 -60 41560 -40
rect 41450 -120 41470 -60
rect 41540 -120 41560 -60
rect 41450 -140 41560 -120
rect 41620 -60 41730 -40
rect 41620 -120 41640 -60
rect 41710 -120 41730 -60
rect 41620 -140 41730 -120
rect 41790 -60 41900 -40
rect 41790 -120 41810 -60
rect 41880 -120 41900 -60
rect 41790 -140 41900 -120
rect 41960 -60 42070 -40
rect 41960 -120 41980 -60
rect 42050 -120 42070 -60
rect 41960 -140 42070 -120
rect 42130 -60 42240 -40
rect 42130 -120 42150 -60
rect 42220 -120 42240 -60
rect 42130 -140 42240 -120
rect 42300 -60 42410 -40
rect 42300 -120 42320 -60
rect 42390 -120 42410 -60
rect 42300 -140 42410 -120
rect 42470 -60 42580 -40
rect 42470 -120 42490 -60
rect 42560 -120 42580 -60
rect 42470 -140 42580 -120
rect 42640 -60 42750 -40
rect 42640 -120 42660 -60
rect 42730 -120 42750 -60
rect 42640 -140 42750 -120
rect 42810 -60 42920 -40
rect 42810 -120 42830 -60
rect 42900 -120 42920 -60
rect 42810 -140 42920 -120
rect 42980 -60 43090 -40
rect 42980 -120 43000 -60
rect 43070 -120 43090 -60
rect 42980 -140 43090 -120
rect 43150 -60 43260 -40
rect 43150 -120 43170 -60
rect 43240 -120 43260 -60
rect 43150 -140 43260 -120
rect 43320 -60 43430 -40
rect 43320 -120 43340 -60
rect 43410 -120 43430 -60
rect 43320 -140 43430 -120
rect 43490 -60 43600 -40
rect 43490 -120 43510 -60
rect 43580 -120 43600 -60
rect 43490 -140 43600 -120
rect 43660 -60 43770 -40
rect 43660 -120 43680 -60
rect 43750 -120 43770 -60
rect 43660 -140 43770 -120
rect 43830 -60 43940 -40
rect 43830 -120 43850 -60
rect 43920 -120 43940 -60
rect 43830 -140 43940 -120
rect 44000 -60 44110 -40
rect 44000 -120 44020 -60
rect 44090 -120 44110 -60
rect 44000 -140 44110 -120
rect 44170 -60 44280 -40
rect 44170 -120 44190 -60
rect 44260 -120 44280 -60
rect 44170 -140 44280 -120
rect 44340 -60 44450 -40
rect 44340 -120 44360 -60
rect 44430 -120 44450 -60
rect 44340 -140 44450 -120
rect 44510 -60 44620 -40
rect 44510 -120 44530 -60
rect 44600 -120 44620 -60
rect 44510 -140 44620 -120
rect 44680 -60 44790 -40
rect 44680 -120 44700 -60
rect 44770 -120 44790 -60
rect 44680 -140 44790 -120
rect 44850 -60 44960 -40
rect 44850 -120 44870 -60
rect 44940 -120 44960 -60
rect 44850 -140 44960 -120
rect 45020 -60 45130 -40
rect 45020 -120 45040 -60
rect 45110 -120 45130 -60
rect 45020 -140 45130 -120
rect 45190 -60 45300 -40
rect 45190 -120 45210 -60
rect 45280 -120 45300 -60
rect 45190 -140 45300 -120
rect 45360 -60 45470 -40
rect 45360 -120 45380 -60
rect 45450 -120 45470 -60
rect 45360 -140 45470 -120
rect 45530 -60 45640 -40
rect 45530 -120 45550 -60
rect 45620 -120 45640 -60
rect 45530 -140 45640 -120
rect 45700 -60 45810 -40
rect 45700 -120 45720 -60
rect 45790 -120 45810 -60
rect 45700 -140 45810 -120
rect 45870 -60 45980 -40
rect 45870 -120 45890 -60
rect 45960 -120 45980 -60
rect 45870 -140 45980 -120
rect 46040 -60 46150 -40
rect 46040 -120 46060 -60
rect 46130 -120 46150 -60
rect 46040 -140 46150 -120
rect 46210 -60 46320 -40
rect 46210 -120 46230 -60
rect 46300 -120 46320 -60
rect 46210 -140 46320 -120
rect 46380 -60 46490 -40
rect 46380 -120 46400 -60
rect 46470 -120 46490 -60
rect 46380 -140 46490 -120
rect 46550 -60 46660 -40
rect 46550 -120 46570 -60
rect 46640 -120 46660 -60
rect 46550 -140 46660 -120
rect 46720 -60 46830 -40
rect 46720 -120 46740 -60
rect 46810 -120 46830 -60
rect 46720 -140 46830 -120
rect 46890 -60 47000 -40
rect 46890 -120 46910 -60
rect 46980 -120 47000 -60
rect 46890 -140 47000 -120
rect 47060 -60 47170 -40
rect 47060 -120 47080 -60
rect 47150 -120 47170 -60
rect 47060 -140 47170 -120
rect 47230 -60 47340 -40
rect 47230 -120 47250 -60
rect 47320 -120 47340 -60
rect 47230 -140 47340 -120
rect 47400 -60 47510 -40
rect 47400 -120 47420 -60
rect 47490 -120 47510 -60
rect 47400 -140 47510 -120
rect 47570 -60 47680 -40
rect 47570 -120 47590 -60
rect 47660 -120 47680 -60
rect 47570 -140 47680 -120
rect 47740 -60 47850 -40
rect 47740 -120 47760 -60
rect 47830 -120 47850 -60
rect 47740 -140 47850 -120
rect 47910 -60 48020 -40
rect 47910 -120 47930 -60
rect 48000 -120 48020 -60
rect 47910 -140 48020 -120
rect 48080 -60 48190 -40
rect 48080 -120 48100 -60
rect 48170 -120 48190 -60
rect 48080 -140 48190 -120
rect 48250 -60 48360 -40
rect 48250 -120 48270 -60
rect 48340 -120 48360 -60
rect 48250 -140 48360 -120
rect 48420 -60 48530 -40
rect 48420 -120 48440 -60
rect 48510 -120 48530 -60
rect 48420 -140 48530 -120
rect 48590 -60 48700 -40
rect 48590 -120 48610 -60
rect 48680 -120 48700 -60
rect 48590 -140 48700 -120
rect 48760 -60 48870 -40
rect 48760 -120 48780 -60
rect 48850 -120 48870 -60
rect 48760 -140 48870 -120
rect 48930 -60 49040 -40
rect 48930 -120 48950 -60
rect 49020 -120 49040 -60
rect 48930 -140 49040 -120
rect 49100 -60 49210 -40
rect 49100 -120 49120 -60
rect 49190 -120 49210 -60
rect 49100 -140 49210 -120
rect 49270 -60 49380 -40
rect 49270 -120 49290 -60
rect 49360 -120 49380 -60
rect 49270 -140 49380 -120
rect 49440 -60 49550 -40
rect 49440 -120 49460 -60
rect 49530 -120 49550 -60
rect 49440 -140 49550 -120
rect 49610 -60 49720 -40
rect 49610 -120 49630 -60
rect 49700 -120 49720 -60
rect 49610 -140 49720 -120
rect 49780 -60 49890 -40
rect 49780 -120 49800 -60
rect 49870 -120 49890 -60
rect 49780 -140 49890 -120
rect 49950 -60 50060 -40
rect 49950 -120 49970 -60
rect 50040 -120 50060 -60
rect 49950 -140 50060 -120
rect 50120 -60 50230 -40
rect 50120 -120 50140 -60
rect 50210 -120 50230 -60
rect 50120 -140 50230 -120
rect 50290 -60 50400 -40
rect 50290 -120 50310 -60
rect 50380 -120 50400 -60
rect 50290 -140 50400 -120
rect 50460 -60 50570 -40
rect 50460 -120 50480 -60
rect 50550 -120 50570 -60
rect 50460 -140 50570 -120
rect 50630 -60 50740 -40
rect 50630 -120 50650 -60
rect 50720 -120 50740 -60
rect 50630 -140 50740 -120
rect 50800 -60 50910 -40
rect 50800 -120 50820 -60
rect 50890 -120 50910 -60
rect 50800 -140 50910 -120
rect 50970 -60 51080 -40
rect 50970 -120 50990 -60
rect 51060 -120 51080 -60
rect 50970 -140 51080 -120
rect 51140 -60 51250 -40
rect 51140 -120 51160 -60
rect 51230 -120 51250 -60
rect 51140 -140 51250 -120
rect 51310 -60 51420 -40
rect 51310 -120 51330 -60
rect 51400 -120 51420 -60
rect 51310 -140 51420 -120
rect 51480 -60 51590 -40
rect 51480 -120 51500 -60
rect 51570 -120 51590 -60
rect 51480 -140 51590 -120
rect 51650 -60 51760 -40
rect 51650 -120 51670 -60
rect 51740 -120 51760 -60
rect 51650 -140 51760 -120
rect 51820 -60 51930 -40
rect 51820 -120 51840 -60
rect 51910 -120 51930 -60
rect 51820 -140 51930 -120
rect 51990 -60 52100 -40
rect 51990 -120 52010 -60
rect 52080 -120 52100 -60
rect 51990 -140 52100 -120
rect 52160 -60 52270 -40
rect 52160 -120 52180 -60
rect 52250 -120 52270 -60
rect 52160 -140 52270 -120
rect 52330 -60 52440 -40
rect 52330 -120 52350 -60
rect 52420 -120 52440 -60
rect 52330 -140 52440 -120
rect 52500 -60 52610 -40
rect 52500 -120 52520 -60
rect 52590 -120 52610 -60
rect 52500 -140 52610 -120
rect 52670 -60 52780 -40
rect 52670 -120 52690 -60
rect 52760 -120 52780 -60
rect 52670 -140 52780 -120
rect 52840 -60 52950 -40
rect 52840 -120 52860 -60
rect 52930 -120 52950 -60
rect 52840 -140 52950 -120
rect 53010 -60 53120 -40
rect 53010 -120 53030 -60
rect 53100 -120 53120 -60
rect 53010 -140 53120 -120
rect 53180 -60 53290 -40
rect 53180 -120 53200 -60
rect 53270 -120 53290 -60
rect 53180 -140 53290 -120
rect 53350 -60 53460 -40
rect 53350 -120 53370 -60
rect 53440 -120 53460 -60
rect 53350 -140 53460 -120
rect 53520 -60 53630 -40
rect 53520 -120 53540 -60
rect 53610 -120 53630 -60
rect 53520 -140 53630 -120
rect 53690 -60 53800 -40
rect 53690 -120 53710 -60
rect 53780 -120 53800 -60
rect 53690 -140 53800 -120
rect 53860 -60 53970 -40
rect 53860 -120 53880 -60
rect 53950 -120 53970 -60
rect 53860 -140 53970 -120
rect 54030 -60 54140 -40
rect 54030 -120 54050 -60
rect 54120 -120 54140 -60
rect 54030 -140 54140 -120
rect 54200 -60 54310 -40
rect 54200 -120 54220 -60
rect 54290 -120 54310 -60
rect 54200 -140 54310 -120
rect 54370 -60 54480 -40
rect 54370 -120 54390 -60
rect 54460 -120 54480 -60
rect 54370 -140 54480 -120
rect 54540 -60 54650 -40
rect 54540 -120 54560 -60
rect 54630 -120 54650 -60
rect 54540 -140 54650 -120
rect 54710 -60 54820 -40
rect 54710 -120 54730 -60
rect 54800 -120 54820 -60
rect 54710 -140 54820 -120
rect 54880 -60 54990 -40
rect 54880 -120 54900 -60
rect 54970 -120 54990 -60
rect 54880 -140 54990 -120
rect 55050 -60 55160 -40
rect 55050 -120 55070 -60
rect 55140 -120 55160 -60
rect 55050 -140 55160 -120
rect 55220 -60 55330 -40
rect 55220 -120 55240 -60
rect 55310 -120 55330 -60
rect 55220 -140 55330 -120
rect 55390 -60 55500 -40
rect 55390 -120 55410 -60
rect 55480 -120 55500 -60
rect 55390 -140 55500 -120
rect 55560 -60 55670 -40
rect 55560 -120 55580 -60
rect 55650 -120 55670 -60
rect 55560 -140 55670 -120
rect 55730 -60 55840 -40
rect 55730 -120 55750 -60
rect 55820 -120 55840 -60
rect 55730 -140 55840 -120
rect 55900 -60 56010 -40
rect 55900 -120 55920 -60
rect 55990 -120 56010 -60
rect 55900 -140 56010 -120
rect 56070 -60 56180 -40
rect 56070 -120 56090 -60
rect 56160 -120 56180 -60
rect 56070 -140 56180 -120
rect 56240 -60 56350 -40
rect 56240 -120 56260 -60
rect 56330 -120 56350 -60
rect 56240 -140 56350 -120
rect 56410 -60 56520 -40
rect 56410 -120 56430 -60
rect 56500 -120 56520 -60
rect 56410 -140 56520 -120
rect 56580 -60 56690 -40
rect 56580 -120 56600 -60
rect 56670 -120 56690 -60
rect 56580 -140 56690 -120
rect 56750 -60 56860 -40
rect 56750 -120 56770 -60
rect 56840 -120 56860 -60
rect 56750 -140 56860 -120
rect 56920 -60 57030 -40
rect 56920 -120 56940 -60
rect 57010 -120 57030 -60
rect 56920 -140 57030 -120
rect 57090 -60 57200 -40
rect 57090 -120 57110 -60
rect 57180 -120 57200 -60
rect 57090 -140 57200 -120
rect 57260 -60 57370 -40
rect 57260 -120 57280 -60
rect 57350 -120 57370 -60
rect 57260 -140 57370 -120
rect 57430 -60 57540 -40
rect 57430 -120 57450 -60
rect 57520 -120 57540 -60
rect 57430 -140 57540 -120
rect 57600 -60 57710 -40
rect 57600 -120 57620 -60
rect 57690 -120 57710 -60
rect 57600 -140 57710 -120
rect 57770 -60 57880 -40
rect 57770 -120 57790 -60
rect 57860 -120 57880 -60
rect 57770 -140 57880 -120
rect 57940 -60 58050 -40
rect 57940 -120 57960 -60
rect 58030 -120 58050 -60
rect 57940 -140 58050 -120
rect 58110 -60 58220 -40
rect 58110 -120 58130 -60
rect 58200 -120 58220 -60
rect 58110 -140 58220 -120
rect 58280 -60 58390 -40
rect 58280 -120 58300 -60
rect 58370 -120 58390 -60
rect 58280 -140 58390 -120
rect 58450 -60 58560 -40
rect 58450 -120 58470 -60
rect 58540 -120 58560 -60
rect 58450 -140 58560 -120
rect 58620 -60 58730 -40
rect 58620 -120 58640 -60
rect 58710 -120 58730 -60
rect 58620 -140 58730 -120
rect 58790 -60 58900 -40
rect 58790 -120 58810 -60
rect 58880 -120 58900 -60
rect 58790 -140 58900 -120
rect 58960 -60 59070 -40
rect 58960 -120 58980 -60
rect 59050 -120 59070 -60
rect 58960 -140 59070 -120
rect 59130 -60 59240 -40
rect 59130 -120 59150 -60
rect 59220 -120 59240 -60
rect 59130 -140 59240 -120
rect 2070 -260 2400 -240
rect 2070 -390 2120 -260
rect 2350 -390 2400 -260
rect 2070 -410 2400 -390
rect 5088 -268 5418 -248
rect 5088 -398 5138 -268
rect 5368 -398 5418 -268
rect 5088 -418 5418 -398
rect 7574 -268 7904 -248
rect 7574 -398 7624 -268
rect 7854 -398 7904 -268
rect 7574 -418 7904 -398
rect 8994 -268 9324 -248
rect 8994 -398 9044 -268
rect 9274 -398 9324 -268
rect 8994 -418 9324 -398
rect 13618 -264 13948 -244
rect 13618 -394 13668 -264
rect 13898 -394 13948 -264
rect 13618 -414 13948 -394
rect 16818 -264 17148 -244
rect 16818 -394 16868 -264
rect 17098 -394 17148 -264
rect 16818 -414 17148 -394
rect 20374 -264 20704 -244
rect 20374 -394 20424 -264
rect 20654 -394 20704 -264
rect 20374 -414 20704 -394
rect 25708 -264 26038 -244
rect 25708 -394 25758 -264
rect 25988 -394 26038 -264
rect 25708 -414 26038 -394
rect 28552 -264 28882 -244
rect 28552 -394 28602 -264
rect 28832 -394 28882 -264
rect 28552 -414 28882 -394
rect 32464 -264 32794 -244
rect 32464 -394 32514 -264
rect 32744 -394 32794 -264
rect 32464 -414 32794 -394
rect 34620 -264 34950 -244
rect 34620 -394 34670 -264
rect 34900 -394 34950 -264
rect 34620 -414 34950 -394
rect 37442 -264 37772 -244
rect 37442 -394 37492 -264
rect 37722 -394 37772 -264
rect 37442 -414 37772 -394
rect 40642 -264 40972 -244
rect 40642 -394 40692 -264
rect 40922 -394 40972 -264
rect 40642 -414 40972 -394
rect 45618 -264 45948 -244
rect 45618 -394 45668 -264
rect 45898 -394 45948 -264
rect 45618 -414 45948 -394
rect 48818 -264 49148 -244
rect 48818 -394 48868 -264
rect 49098 -394 49148 -264
rect 48818 -414 49148 -394
rect 50952 -264 51282 -244
rect 50952 -394 51002 -264
rect 51232 -394 51282 -264
rect 50952 -414 51282 -394
rect 54508 -264 54838 -244
rect 54508 -394 54558 -264
rect 54788 -394 54838 -264
rect 54508 -414 54838 -394
rect 57352 -264 57682 -244
rect 57352 -394 57402 -264
rect 57632 -394 57682 -264
rect 57352 -414 57682 -394
rect 61264 -264 61594 -244
rect 61264 -394 61314 -264
rect 61544 -394 61594 -264
rect 61264 -414 61594 -394
rect 64108 -264 64438 -244
rect 64108 -394 64158 -264
rect 64388 -394 64438 -264
rect 64108 -414 64438 -394
rect 67664 -264 67994 -244
rect 67664 -394 67714 -264
rect 67944 -394 67994 -264
rect 67664 -414 67994 -394
rect 70508 -264 70838 -244
rect 70508 -394 70558 -264
rect 70788 -394 70838 -264
rect 70508 -414 70838 -394
rect 74418 -264 74748 -244
rect 74418 -394 74468 -264
rect 74698 -394 74748 -264
rect 74418 -414 74748 -394
rect 78330 -264 78660 -244
rect 78330 -394 78380 -264
rect 78610 -394 78660 -264
rect 78330 -414 78660 -394
rect 82242 -264 82572 -244
rect 82242 -394 82292 -264
rect 82522 -394 82572 -264
rect 82242 -414 82572 -394
rect 86152 -264 86482 -244
rect 86152 -394 86202 -264
rect 86432 -394 86482 -264
rect 86152 -414 86482 -394
rect 210 -530 320 -510
rect 210 -590 230 -530
rect 300 -590 320 -530
rect 210 -610 320 -590
rect 380 -530 490 -510
rect 380 -590 400 -530
rect 470 -590 490 -530
rect 380 -610 490 -590
rect 550 -530 660 -510
rect 550 -590 570 -530
rect 640 -590 660 -530
rect 550 -610 660 -590
rect 720 -530 830 -510
rect 720 -590 740 -530
rect 810 -590 830 -530
rect 720 -610 830 -590
rect 890 -530 1000 -510
rect 890 -590 910 -530
rect 980 -590 1000 -530
rect 890 -610 1000 -590
rect 1060 -530 1170 -510
rect 1060 -590 1080 -530
rect 1150 -590 1170 -530
rect 1060 -610 1170 -590
rect 1230 -530 1340 -510
rect 1230 -590 1250 -530
rect 1320 -590 1340 -530
rect 1230 -610 1340 -590
rect 1400 -530 1510 -510
rect 1400 -590 1420 -530
rect 1490 -590 1510 -530
rect 1400 -610 1510 -590
rect 1570 -530 1680 -510
rect 1570 -590 1590 -530
rect 1660 -590 1680 -530
rect 1570 -610 1680 -590
rect 1740 -530 1850 -510
rect 1740 -590 1760 -530
rect 1830 -590 1850 -530
rect 1740 -610 1850 -590
rect 1910 -530 2020 -510
rect 1910 -590 1930 -530
rect 2000 -590 2020 -530
rect 1910 -610 2020 -590
rect 2080 -530 2190 -510
rect 2080 -590 2100 -530
rect 2170 -590 2190 -530
rect 2080 -610 2190 -590
rect 2250 -530 2360 -510
rect 2250 -590 2270 -530
rect 2340 -590 2360 -530
rect 2250 -610 2360 -590
rect 2420 -530 2530 -510
rect 2420 -590 2440 -530
rect 2510 -590 2530 -530
rect 2420 -610 2530 -590
rect 2590 -530 2700 -510
rect 2590 -590 2610 -530
rect 2680 -590 2700 -530
rect 2590 -610 2700 -590
rect 2760 -530 2870 -510
rect 2760 -590 2780 -530
rect 2850 -590 2870 -530
rect 2760 -610 2870 -590
rect 2930 -530 3040 -510
rect 2930 -590 2950 -530
rect 3020 -590 3040 -530
rect 2930 -610 3040 -590
rect 3100 -530 3210 -510
rect 3100 -590 3120 -530
rect 3190 -590 3210 -530
rect 3100 -610 3210 -590
rect 3270 -530 3380 -510
rect 3270 -590 3290 -530
rect 3360 -590 3380 -530
rect 3270 -610 3380 -590
rect 3440 -530 3550 -510
rect 3440 -590 3460 -530
rect 3530 -590 3550 -530
rect 3440 -610 3550 -590
rect 3610 -530 3720 -510
rect 3610 -590 3630 -530
rect 3700 -590 3720 -530
rect 3610 -610 3720 -590
rect 3780 -530 3890 -510
rect 3780 -590 3800 -530
rect 3870 -590 3890 -530
rect 3780 -610 3890 -590
rect 3950 -530 4060 -510
rect 3950 -590 3970 -530
rect 4040 -590 4060 -530
rect 3950 -610 4060 -590
rect 4120 -530 4230 -510
rect 4120 -590 4140 -530
rect 4210 -590 4230 -530
rect 4120 -610 4230 -590
rect 4290 -530 4400 -510
rect 4290 -590 4310 -530
rect 4380 -590 4400 -530
rect 4290 -610 4400 -590
rect 4460 -530 4570 -510
rect 4460 -590 4480 -530
rect 4550 -590 4570 -530
rect 4460 -610 4570 -590
rect 4630 -530 4740 -510
rect 4630 -590 4650 -530
rect 4720 -590 4740 -530
rect 4630 -610 4740 -590
rect 4800 -530 4910 -510
rect 4800 -590 4820 -530
rect 4890 -590 4910 -530
rect 4800 -610 4910 -590
rect 4970 -530 5080 -510
rect 4970 -590 4990 -530
rect 5060 -590 5080 -530
rect 4970 -610 5080 -590
rect 5140 -530 5250 -510
rect 5140 -590 5160 -530
rect 5230 -590 5250 -530
rect 5140 -610 5250 -590
rect 5310 -530 5420 -510
rect 5310 -590 5330 -530
rect 5400 -590 5420 -530
rect 5310 -610 5420 -590
rect 5480 -530 5590 -510
rect 5480 -590 5500 -530
rect 5570 -590 5590 -530
rect 5480 -610 5590 -590
rect 5650 -530 5760 -510
rect 5650 -590 5670 -530
rect 5740 -590 5760 -530
rect 5650 -610 5760 -590
rect 5820 -530 5930 -510
rect 5820 -590 5840 -530
rect 5910 -590 5930 -530
rect 5820 -610 5930 -590
rect 5990 -530 6100 -510
rect 5990 -590 6010 -530
rect 6080 -590 6100 -530
rect 5990 -610 6100 -590
rect 6160 -530 6270 -510
rect 6160 -590 6180 -530
rect 6250 -590 6270 -530
rect 6160 -610 6270 -590
rect 6330 -530 6440 -510
rect 6330 -590 6350 -530
rect 6420 -590 6440 -530
rect 6330 -610 6440 -590
rect 6500 -530 6610 -510
rect 6500 -590 6520 -530
rect 6590 -590 6610 -530
rect 6500 -610 6610 -590
rect 6670 -530 6780 -510
rect 6670 -590 6690 -530
rect 6760 -590 6780 -530
rect 6670 -610 6780 -590
rect 6840 -530 6950 -510
rect 6840 -590 6860 -530
rect 6930 -590 6950 -530
rect 6840 -610 6950 -590
rect 7010 -530 7120 -510
rect 7010 -590 7030 -530
rect 7100 -590 7120 -530
rect 7010 -610 7120 -590
rect 7180 -530 7290 -510
rect 7180 -590 7200 -530
rect 7270 -590 7290 -530
rect 7180 -610 7290 -590
rect 7350 -530 7460 -510
rect 7350 -590 7370 -530
rect 7440 -590 7460 -530
rect 7350 -610 7460 -590
rect 7520 -530 7630 -510
rect 7520 -590 7540 -530
rect 7610 -590 7630 -530
rect 7520 -610 7630 -590
rect 7690 -530 7800 -510
rect 7690 -590 7710 -530
rect 7780 -590 7800 -530
rect 7690 -610 7800 -590
rect 7860 -530 7970 -510
rect 7860 -590 7880 -530
rect 7950 -590 7970 -530
rect 7860 -610 7970 -590
rect 8030 -530 8140 -510
rect 8030 -590 8050 -530
rect 8120 -590 8140 -530
rect 8030 -610 8140 -590
rect 8200 -530 8310 -510
rect 8200 -590 8220 -530
rect 8290 -590 8310 -530
rect 8200 -610 8310 -590
rect 8370 -530 8480 -510
rect 8370 -590 8390 -530
rect 8460 -590 8480 -530
rect 8370 -610 8480 -590
rect 8540 -530 8650 -510
rect 8540 -590 8560 -530
rect 8630 -590 8650 -530
rect 8540 -610 8650 -590
rect 8710 -530 8820 -510
rect 8710 -590 8730 -530
rect 8800 -590 8820 -530
rect 8710 -610 8820 -590
rect 8880 -530 8990 -510
rect 8880 -590 8900 -530
rect 8970 -590 8990 -530
rect 8880 -610 8990 -590
rect 9050 -530 9160 -510
rect 9050 -590 9070 -530
rect 9140 -590 9160 -530
rect 9050 -610 9160 -590
rect 9220 -530 9330 -510
rect 9220 -590 9240 -530
rect 9310 -590 9330 -530
rect 9220 -610 9330 -590
rect 9390 -530 9500 -510
rect 9390 -590 9410 -530
rect 9480 -590 9500 -530
rect 9390 -610 9500 -590
rect 9560 -530 9670 -510
rect 9560 -590 9580 -530
rect 9650 -590 9670 -530
rect 9560 -610 9670 -590
rect 9730 -530 9840 -510
rect 9730 -590 9750 -530
rect 9820 -590 9840 -530
rect 9730 -610 9840 -590
rect 9900 -530 10010 -510
rect 9900 -590 9920 -530
rect 9990 -590 10010 -530
rect 9900 -610 10010 -590
rect 10070 -530 10180 -510
rect 10070 -590 10090 -530
rect 10160 -590 10180 -530
rect 10070 -610 10180 -590
rect 10240 -530 10350 -510
rect 10240 -590 10260 -530
rect 10330 -590 10350 -530
rect 10240 -610 10350 -590
rect 10410 -530 10520 -510
rect 10410 -590 10430 -530
rect 10500 -590 10520 -530
rect 10410 -610 10520 -590
rect 10580 -530 10690 -510
rect 10580 -590 10600 -530
rect 10670 -590 10690 -530
rect 10580 -610 10690 -590
rect 10750 -530 10860 -510
rect 10750 -590 10770 -530
rect 10840 -590 10860 -530
rect 10750 -610 10860 -590
rect 10920 -530 11030 -510
rect 10920 -590 10940 -530
rect 11010 -590 11030 -530
rect 10920 -610 11030 -590
rect 11090 -530 11200 -510
rect 11090 -590 11110 -530
rect 11180 -590 11200 -530
rect 11090 -610 11200 -590
rect 11260 -530 11370 -510
rect 11260 -590 11280 -530
rect 11350 -590 11370 -530
rect 11260 -610 11370 -590
rect 11430 -530 11540 -510
rect 11430 -590 11450 -530
rect 11520 -590 11540 -530
rect 11430 -610 11540 -590
rect 11600 -530 11710 -510
rect 11600 -590 11620 -530
rect 11690 -590 11710 -530
rect 11600 -610 11710 -590
rect 11770 -530 11880 -510
rect 11770 -590 11790 -530
rect 11860 -590 11880 -530
rect 11770 -610 11880 -590
rect 11940 -530 12050 -510
rect 11940 -590 11960 -530
rect 12030 -590 12050 -530
rect 11940 -610 12050 -590
rect 12110 -530 12220 -510
rect 12110 -590 12130 -530
rect 12200 -590 12220 -530
rect 12110 -610 12220 -590
rect 12280 -530 12390 -510
rect 12280 -590 12300 -530
rect 12370 -590 12390 -530
rect 12280 -610 12390 -590
rect 12450 -530 12560 -510
rect 12450 -590 12470 -530
rect 12540 -590 12560 -530
rect 12450 -610 12560 -590
rect 12620 -530 12730 -510
rect 12620 -590 12640 -530
rect 12710 -590 12730 -530
rect 12620 -610 12730 -590
rect 12790 -530 12900 -510
rect 12790 -590 12810 -530
rect 12880 -590 12900 -530
rect 12790 -610 12900 -590
rect 12960 -530 13070 -510
rect 12960 -590 12980 -530
rect 13050 -590 13070 -530
rect 12960 -610 13070 -590
rect 13130 -530 13240 -510
rect 13130 -590 13150 -530
rect 13220 -590 13240 -530
rect 13130 -610 13240 -590
rect 13300 -530 13410 -510
rect 13300 -590 13320 -530
rect 13390 -590 13410 -530
rect 13300 -610 13410 -590
rect 13470 -530 13580 -510
rect 13470 -590 13490 -530
rect 13560 -590 13580 -530
rect 13470 -610 13580 -590
rect 13640 -530 13750 -510
rect 13640 -590 13660 -530
rect 13730 -590 13750 -530
rect 13640 -610 13750 -590
rect 13810 -530 13920 -510
rect 13810 -590 13830 -530
rect 13900 -590 13920 -530
rect 13810 -610 13920 -590
rect 13980 -530 14090 -510
rect 13980 -590 14000 -530
rect 14070 -590 14090 -530
rect 13980 -610 14090 -590
rect 14150 -530 14260 -510
rect 14150 -590 14170 -530
rect 14240 -590 14260 -530
rect 14150 -610 14260 -590
rect 14320 -530 14430 -510
rect 14320 -590 14340 -530
rect 14410 -590 14430 -530
rect 14320 -610 14430 -590
rect 14490 -530 14600 -510
rect 14490 -590 14510 -530
rect 14580 -590 14600 -530
rect 14490 -610 14600 -590
rect 14660 -530 14770 -510
rect 14660 -590 14680 -530
rect 14750 -590 14770 -530
rect 14660 -610 14770 -590
rect 14830 -530 14940 -510
rect 14830 -590 14850 -530
rect 14920 -590 14940 -530
rect 14830 -610 14940 -590
rect 15000 -530 15110 -510
rect 15000 -590 15020 -530
rect 15090 -590 15110 -530
rect 15000 -610 15110 -590
rect 15170 -530 15280 -510
rect 15170 -590 15190 -530
rect 15260 -590 15280 -530
rect 15170 -610 15280 -590
rect 15340 -530 15450 -510
rect 15340 -590 15360 -530
rect 15430 -590 15450 -530
rect 15340 -610 15450 -590
rect 15510 -530 15620 -510
rect 15510 -590 15530 -530
rect 15600 -590 15620 -530
rect 15510 -610 15620 -590
rect 15680 -530 15790 -510
rect 15680 -590 15700 -530
rect 15770 -590 15790 -530
rect 15680 -610 15790 -590
rect 15850 -530 15960 -510
rect 15850 -590 15870 -530
rect 15940 -590 15960 -530
rect 15850 -610 15960 -590
rect 16020 -530 16130 -510
rect 16020 -590 16040 -530
rect 16110 -590 16130 -530
rect 16020 -610 16130 -590
rect 16190 -530 16300 -510
rect 16190 -590 16210 -530
rect 16280 -590 16300 -530
rect 16190 -610 16300 -590
rect 16360 -530 16470 -510
rect 16360 -590 16380 -530
rect 16450 -590 16470 -530
rect 16360 -610 16470 -590
rect 16530 -530 16640 -510
rect 16530 -590 16550 -530
rect 16620 -590 16640 -530
rect 16530 -610 16640 -590
rect 16700 -530 16810 -510
rect 16700 -590 16720 -530
rect 16790 -590 16810 -530
rect 16700 -610 16810 -590
rect 16870 -530 16980 -510
rect 16870 -590 16890 -530
rect 16960 -590 16980 -530
rect 16870 -610 16980 -590
rect 17040 -530 17150 -510
rect 17040 -590 17060 -530
rect 17130 -590 17150 -530
rect 17040 -610 17150 -590
rect 17210 -530 17320 -510
rect 17210 -590 17230 -530
rect 17300 -590 17320 -530
rect 17210 -610 17320 -590
rect 17380 -530 17490 -510
rect 17380 -590 17400 -530
rect 17470 -590 17490 -530
rect 17380 -610 17490 -590
rect 17550 -530 17660 -510
rect 17550 -590 17570 -530
rect 17640 -590 17660 -530
rect 17550 -610 17660 -590
rect 17720 -530 17830 -510
rect 17720 -590 17740 -530
rect 17810 -590 17830 -530
rect 17720 -610 17830 -590
rect 17890 -530 18000 -510
rect 17890 -590 17910 -530
rect 17980 -590 18000 -530
rect 17890 -610 18000 -590
rect 18060 -530 18170 -510
rect 18060 -590 18080 -530
rect 18150 -590 18170 -530
rect 18060 -610 18170 -590
rect 18230 -530 18340 -510
rect 18230 -590 18250 -530
rect 18320 -590 18340 -530
rect 18230 -610 18340 -590
rect 18400 -530 18510 -510
rect 18400 -590 18420 -530
rect 18490 -590 18510 -530
rect 18400 -610 18510 -590
rect 18570 -530 18680 -510
rect 18570 -590 18590 -530
rect 18660 -590 18680 -530
rect 18570 -610 18680 -590
rect 18740 -530 18850 -510
rect 18740 -590 18760 -530
rect 18830 -590 18850 -530
rect 18740 -610 18850 -590
rect 18910 -530 19020 -510
rect 18910 -590 18930 -530
rect 19000 -590 19020 -530
rect 18910 -610 19020 -590
rect 19080 -530 19190 -510
rect 19080 -590 19100 -530
rect 19170 -590 19190 -530
rect 19080 -610 19190 -590
rect 19250 -530 19360 -510
rect 19250 -590 19270 -530
rect 19340 -590 19360 -530
rect 19250 -610 19360 -590
rect 19420 -530 19530 -510
rect 19420 -590 19440 -530
rect 19510 -590 19530 -530
rect 19420 -610 19530 -590
rect 19590 -530 19700 -510
rect 19590 -590 19610 -530
rect 19680 -590 19700 -530
rect 19590 -610 19700 -590
rect 19760 -530 19870 -510
rect 19760 -590 19780 -530
rect 19850 -590 19870 -530
rect 19760 -610 19870 -590
rect 19930 -530 20040 -510
rect 19930 -590 19950 -530
rect 20020 -590 20040 -530
rect 19930 -610 20040 -590
rect 20100 -530 20210 -510
rect 20100 -590 20120 -530
rect 20190 -590 20210 -530
rect 20100 -610 20210 -590
rect 20270 -530 20380 -510
rect 20270 -590 20290 -530
rect 20360 -590 20380 -530
rect 20270 -610 20380 -590
rect 20440 -530 20550 -510
rect 20440 -590 20460 -530
rect 20530 -590 20550 -530
rect 20440 -610 20550 -590
rect 20610 -530 20720 -510
rect 20610 -590 20630 -530
rect 20700 -590 20720 -530
rect 20610 -610 20720 -590
rect 20780 -530 20890 -510
rect 20780 -590 20800 -530
rect 20870 -590 20890 -530
rect 20780 -610 20890 -590
rect 20950 -530 21060 -510
rect 20950 -590 20970 -530
rect 21040 -590 21060 -530
rect 20950 -610 21060 -590
rect 21120 -530 21230 -510
rect 21120 -590 21140 -530
rect 21210 -590 21230 -530
rect 21120 -610 21230 -590
rect 21290 -530 21400 -510
rect 21290 -590 21310 -530
rect 21380 -590 21400 -530
rect 21290 -610 21400 -590
rect 21460 -530 21570 -510
rect 21460 -590 21480 -530
rect 21550 -590 21570 -530
rect 21460 -610 21570 -590
rect 21630 -530 21740 -510
rect 21630 -590 21650 -530
rect 21720 -590 21740 -530
rect 21630 -610 21740 -590
rect 21800 -530 21910 -510
rect 21800 -590 21820 -530
rect 21890 -590 21910 -530
rect 21800 -610 21910 -590
rect 21970 -530 22080 -510
rect 21970 -590 21990 -530
rect 22060 -590 22080 -530
rect 21970 -610 22080 -590
rect 22140 -530 22250 -510
rect 22140 -590 22160 -530
rect 22230 -590 22250 -530
rect 22140 -610 22250 -590
rect 22310 -530 22420 -510
rect 22310 -590 22330 -530
rect 22400 -590 22420 -530
rect 22310 -610 22420 -590
rect 22480 -530 22590 -510
rect 22480 -590 22500 -530
rect 22570 -590 22590 -530
rect 22480 -610 22590 -590
rect 22650 -530 22760 -510
rect 22650 -590 22670 -530
rect 22740 -590 22760 -530
rect 22650 -610 22760 -590
rect 22820 -530 22930 -510
rect 22820 -590 22840 -530
rect 22910 -590 22930 -530
rect 22820 -610 22930 -590
rect 22990 -530 23100 -510
rect 22990 -590 23010 -530
rect 23080 -590 23100 -530
rect 22990 -610 23100 -590
rect 23160 -530 23270 -510
rect 23160 -590 23180 -530
rect 23250 -590 23270 -530
rect 23160 -610 23270 -590
rect 23330 -530 23440 -510
rect 23330 -590 23350 -530
rect 23420 -590 23440 -530
rect 23330 -610 23440 -590
rect 23500 -530 23610 -510
rect 23500 -590 23520 -530
rect 23590 -590 23610 -530
rect 23500 -610 23610 -590
rect 23670 -530 23780 -510
rect 23670 -590 23690 -530
rect 23760 -590 23780 -530
rect 23670 -610 23780 -590
rect 23840 -530 23950 -510
rect 23840 -590 23860 -530
rect 23930 -590 23950 -530
rect 23840 -610 23950 -590
rect 24010 -530 24120 -510
rect 24010 -590 24030 -530
rect 24100 -590 24120 -530
rect 24010 -610 24120 -590
rect 24180 -530 24290 -510
rect 24180 -590 24200 -530
rect 24270 -590 24290 -530
rect 24180 -610 24290 -590
rect 24350 -530 24460 -510
rect 24350 -590 24370 -530
rect 24440 -590 24460 -530
rect 24350 -610 24460 -590
rect 24520 -530 24630 -510
rect 24520 -590 24540 -530
rect 24610 -590 24630 -530
rect 24520 -610 24630 -590
rect 24690 -530 24800 -510
rect 24690 -590 24710 -530
rect 24780 -590 24800 -530
rect 24690 -610 24800 -590
rect 24860 -530 24970 -510
rect 24860 -590 24880 -530
rect 24950 -590 24970 -530
rect 24860 -610 24970 -590
rect 25030 -530 25140 -510
rect 25030 -590 25050 -530
rect 25120 -590 25140 -530
rect 25030 -610 25140 -590
rect 25200 -530 25310 -510
rect 25200 -590 25220 -530
rect 25290 -590 25310 -530
rect 25200 -610 25310 -590
rect 25370 -530 25480 -510
rect 25370 -590 25390 -530
rect 25460 -590 25480 -530
rect 25370 -610 25480 -590
rect 25540 -530 25650 -510
rect 25540 -590 25560 -530
rect 25630 -590 25650 -530
rect 25540 -610 25650 -590
rect 25710 -530 25820 -510
rect 25710 -590 25730 -530
rect 25800 -590 25820 -530
rect 25710 -610 25820 -590
rect 25880 -530 25990 -510
rect 25880 -590 25900 -530
rect 25970 -590 25990 -530
rect 25880 -610 25990 -590
rect 26050 -530 26160 -510
rect 26050 -590 26070 -530
rect 26140 -590 26160 -530
rect 26050 -610 26160 -590
rect 26220 -530 26330 -510
rect 26220 -590 26240 -530
rect 26310 -590 26330 -530
rect 26220 -610 26330 -590
rect 26390 -530 26500 -510
rect 26390 -590 26410 -530
rect 26480 -590 26500 -530
rect 26390 -610 26500 -590
rect 26560 -530 26670 -510
rect 26560 -590 26580 -530
rect 26650 -590 26670 -530
rect 26560 -610 26670 -590
rect 26730 -530 26840 -510
rect 26730 -590 26750 -530
rect 26820 -590 26840 -530
rect 26730 -610 26840 -590
rect 26900 -530 27010 -510
rect 26900 -590 26920 -530
rect 26990 -590 27010 -530
rect 26900 -610 27010 -590
rect 27070 -530 27180 -510
rect 27070 -590 27090 -530
rect 27160 -590 27180 -530
rect 27070 -610 27180 -590
rect 27240 -530 27350 -510
rect 27240 -590 27260 -530
rect 27330 -590 27350 -530
rect 27240 -610 27350 -590
rect 27410 -530 27520 -510
rect 27410 -590 27430 -530
rect 27500 -590 27520 -530
rect 27410 -610 27520 -590
rect 27580 -530 27690 -510
rect 27580 -590 27600 -530
rect 27670 -590 27690 -530
rect 27580 -610 27690 -590
rect 27750 -530 27860 -510
rect 27750 -590 27770 -530
rect 27840 -590 27860 -530
rect 27750 -610 27860 -590
rect 27920 -530 28030 -510
rect 27920 -590 27940 -530
rect 28010 -590 28030 -530
rect 27920 -610 28030 -590
rect 28090 -530 28200 -510
rect 28090 -590 28110 -530
rect 28180 -590 28200 -530
rect 28090 -610 28200 -590
rect 28260 -530 28370 -510
rect 28260 -590 28280 -530
rect 28350 -590 28370 -530
rect 28260 -610 28370 -590
rect 28430 -530 28540 -510
rect 28430 -590 28450 -530
rect 28520 -590 28540 -530
rect 28430 -610 28540 -590
rect 28600 -530 28710 -510
rect 28600 -590 28620 -530
rect 28690 -590 28710 -530
rect 28600 -610 28710 -590
rect 28770 -530 28880 -510
rect 28770 -590 28790 -530
rect 28860 -590 28880 -530
rect 28770 -610 28880 -590
rect 28940 -530 29050 -510
rect 28940 -590 28960 -530
rect 29030 -590 29050 -530
rect 28940 -610 29050 -590
rect 29110 -530 29220 -510
rect 29110 -590 29130 -530
rect 29200 -590 29220 -530
rect 29110 -610 29220 -590
rect 29280 -530 29390 -510
rect 29280 -590 29300 -530
rect 29370 -590 29390 -530
rect 29280 -610 29390 -590
rect 29450 -530 29560 -510
rect 29450 -590 29470 -530
rect 29540 -590 29560 -530
rect 29450 -610 29560 -590
rect 29620 -530 29730 -510
rect 29620 -590 29640 -530
rect 29710 -590 29730 -530
rect 29620 -610 29730 -590
rect 29790 -530 29900 -510
rect 29790 -590 29810 -530
rect 29880 -590 29900 -530
rect 29790 -610 29900 -590
rect 29960 -530 30070 -510
rect 29960 -590 29980 -530
rect 30050 -590 30070 -530
rect 29960 -610 30070 -590
rect 30130 -530 30240 -510
rect 30130 -590 30150 -530
rect 30220 -590 30240 -530
rect 30130 -610 30240 -590
rect 30300 -530 30410 -510
rect 30300 -590 30320 -530
rect 30390 -590 30410 -530
rect 30300 -610 30410 -590
rect 30470 -530 30580 -510
rect 30470 -590 30490 -530
rect 30560 -590 30580 -530
rect 30470 -610 30580 -590
rect 30640 -530 30750 -510
rect 30640 -590 30660 -530
rect 30730 -590 30750 -530
rect 30640 -610 30750 -590
rect 30810 -530 30920 -510
rect 30810 -590 30830 -530
rect 30900 -590 30920 -530
rect 30810 -610 30920 -590
rect 30980 -530 31090 -510
rect 30980 -590 31000 -530
rect 31070 -590 31090 -530
rect 30980 -610 31090 -590
rect 31150 -530 31260 -510
rect 31150 -590 31170 -530
rect 31240 -590 31260 -530
rect 31150 -610 31260 -590
rect 31320 -530 31430 -510
rect 31320 -590 31340 -530
rect 31410 -590 31430 -530
rect 31320 -610 31430 -590
rect 31490 -530 31600 -510
rect 31490 -590 31510 -530
rect 31580 -590 31600 -530
rect 31490 -610 31600 -590
rect 31660 -530 31770 -510
rect 31660 -590 31680 -530
rect 31750 -590 31770 -530
rect 31660 -610 31770 -590
rect 31830 -530 31940 -510
rect 31830 -590 31850 -530
rect 31920 -590 31940 -530
rect 31830 -610 31940 -590
rect 32000 -530 32110 -510
rect 32000 -590 32020 -530
rect 32090 -590 32110 -530
rect 32000 -610 32110 -590
rect 32170 -530 32280 -510
rect 32170 -590 32190 -530
rect 32260 -590 32280 -530
rect 32170 -610 32280 -590
rect 32340 -530 32450 -510
rect 32340 -590 32360 -530
rect 32430 -590 32450 -530
rect 32340 -610 32450 -590
rect 32510 -530 32620 -510
rect 32510 -590 32530 -530
rect 32600 -590 32620 -530
rect 32510 -610 32620 -590
rect 32680 -530 32790 -510
rect 32680 -590 32700 -530
rect 32770 -590 32790 -530
rect 32680 -610 32790 -590
rect 32850 -530 32960 -510
rect 32850 -590 32870 -530
rect 32940 -590 32960 -530
rect 32850 -610 32960 -590
rect 33020 -530 33130 -510
rect 33020 -590 33040 -530
rect 33110 -590 33130 -530
rect 33020 -610 33130 -590
rect 33190 -530 33300 -510
rect 33190 -590 33210 -530
rect 33280 -590 33300 -530
rect 33190 -610 33300 -590
rect 33360 -530 33470 -510
rect 33360 -590 33380 -530
rect 33450 -590 33470 -530
rect 33360 -610 33470 -590
rect 33530 -530 33640 -510
rect 33530 -590 33550 -530
rect 33620 -590 33640 -530
rect 33530 -610 33640 -590
rect 33700 -530 33810 -510
rect 33700 -590 33720 -530
rect 33790 -590 33810 -530
rect 33700 -610 33810 -590
rect 33870 -530 33980 -510
rect 33870 -590 33890 -530
rect 33960 -590 33980 -530
rect 33870 -610 33980 -590
rect 34040 -530 34150 -510
rect 34040 -590 34060 -530
rect 34130 -590 34150 -530
rect 34040 -610 34150 -590
rect 34210 -530 34320 -510
rect 34210 -590 34230 -530
rect 34300 -590 34320 -530
rect 34210 -610 34320 -590
rect 34380 -530 34490 -510
rect 34380 -590 34400 -530
rect 34470 -590 34490 -530
rect 34380 -610 34490 -590
rect 34550 -530 34660 -510
rect 34550 -590 34570 -530
rect 34640 -590 34660 -530
rect 34550 -610 34660 -590
rect 34720 -530 34830 -510
rect 34720 -590 34740 -530
rect 34810 -590 34830 -530
rect 34720 -610 34830 -590
rect 34890 -530 35000 -510
rect 34890 -590 34910 -530
rect 34980 -590 35000 -530
rect 34890 -610 35000 -590
rect 35060 -530 35170 -510
rect 35060 -590 35080 -530
rect 35150 -590 35170 -530
rect 35060 -610 35170 -590
rect 35230 -530 35340 -510
rect 35230 -590 35250 -530
rect 35320 -590 35340 -530
rect 35230 -610 35340 -590
rect 35400 -530 35510 -510
rect 35400 -590 35420 -530
rect 35490 -590 35510 -530
rect 35400 -610 35510 -590
rect 35570 -530 35680 -510
rect 35570 -590 35590 -530
rect 35660 -590 35680 -530
rect 35570 -610 35680 -590
rect 35740 -530 35850 -510
rect 35740 -590 35760 -530
rect 35830 -590 35850 -530
rect 35740 -610 35850 -590
rect 35910 -530 36020 -510
rect 35910 -590 35930 -530
rect 36000 -590 36020 -530
rect 35910 -610 36020 -590
rect 36080 -530 36190 -510
rect 36080 -590 36100 -530
rect 36170 -590 36190 -530
rect 36080 -610 36190 -590
rect 36250 -530 36360 -510
rect 36250 -590 36270 -530
rect 36340 -590 36360 -530
rect 36250 -610 36360 -590
rect 36420 -530 36530 -510
rect 36420 -590 36440 -530
rect 36510 -590 36530 -530
rect 36420 -610 36530 -590
rect 36590 -530 36700 -510
rect 36590 -590 36610 -530
rect 36680 -590 36700 -530
rect 36590 -610 36700 -590
rect 36760 -530 36870 -510
rect 36760 -590 36780 -530
rect 36850 -590 36870 -530
rect 36760 -610 36870 -590
rect 36930 -530 37040 -510
rect 36930 -590 36950 -530
rect 37020 -590 37040 -530
rect 36930 -610 37040 -590
rect 37100 -530 37210 -510
rect 37100 -590 37120 -530
rect 37190 -590 37210 -530
rect 37100 -610 37210 -590
rect 37270 -530 37380 -510
rect 37270 -590 37290 -530
rect 37360 -590 37380 -530
rect 37270 -610 37380 -590
rect 37440 -530 37550 -510
rect 37440 -590 37460 -530
rect 37530 -590 37550 -530
rect 37440 -610 37550 -590
rect 37610 -530 37720 -510
rect 37610 -590 37630 -530
rect 37700 -590 37720 -530
rect 37610 -610 37720 -590
rect 37780 -530 37890 -510
rect 37780 -590 37800 -530
rect 37870 -590 37890 -530
rect 37780 -610 37890 -590
rect 37950 -530 38060 -510
rect 37950 -590 37970 -530
rect 38040 -590 38060 -530
rect 37950 -610 38060 -590
rect 38120 -530 38230 -510
rect 38120 -590 38140 -530
rect 38210 -590 38230 -530
rect 38120 -610 38230 -590
rect 38290 -530 38400 -510
rect 38290 -590 38310 -530
rect 38380 -590 38400 -530
rect 38290 -610 38400 -590
rect 38460 -530 38570 -510
rect 38460 -590 38480 -530
rect 38550 -590 38570 -530
rect 38460 -610 38570 -590
rect 38630 -530 38740 -510
rect 38630 -590 38650 -530
rect 38720 -590 38740 -530
rect 38630 -610 38740 -590
rect 38800 -530 38910 -510
rect 38800 -590 38820 -530
rect 38890 -590 38910 -530
rect 38800 -610 38910 -590
rect 38970 -530 39080 -510
rect 38970 -590 38990 -530
rect 39060 -590 39080 -530
rect 38970 -610 39080 -590
rect 39140 -530 39250 -510
rect 39140 -590 39160 -530
rect 39230 -590 39250 -530
rect 39140 -610 39250 -590
rect 39310 -530 39420 -510
rect 39310 -590 39330 -530
rect 39400 -590 39420 -530
rect 39310 -610 39420 -590
rect 39480 -530 39590 -510
rect 39480 -590 39500 -530
rect 39570 -590 39590 -530
rect 39480 -610 39590 -590
rect 39650 -530 39760 -510
rect 39650 -590 39670 -530
rect 39740 -590 39760 -530
rect 39650 -610 39760 -590
rect 39820 -530 39930 -510
rect 39820 -590 39840 -530
rect 39910 -590 39930 -530
rect 39820 -610 39930 -590
rect 39990 -530 40100 -510
rect 39990 -590 40010 -530
rect 40080 -590 40100 -530
rect 39990 -610 40100 -590
rect 40160 -530 40270 -510
rect 40160 -590 40180 -530
rect 40250 -590 40270 -530
rect 40160 -610 40270 -590
rect 40330 -530 40440 -510
rect 40330 -590 40350 -530
rect 40420 -590 40440 -530
rect 40330 -610 40440 -590
rect 40500 -530 40610 -510
rect 40500 -590 40520 -530
rect 40590 -590 40610 -530
rect 40500 -610 40610 -590
rect 40670 -530 40780 -510
rect 40670 -590 40690 -530
rect 40760 -590 40780 -530
rect 40670 -610 40780 -590
rect 40840 -530 40950 -510
rect 40840 -590 40860 -530
rect 40930 -590 40950 -530
rect 40840 -610 40950 -590
rect 41010 -530 41120 -510
rect 41010 -590 41030 -530
rect 41100 -590 41120 -530
rect 41010 -610 41120 -590
rect 41180 -530 41290 -510
rect 41180 -590 41200 -530
rect 41270 -590 41290 -530
rect 41180 -610 41290 -590
rect 41350 -530 41460 -510
rect 41350 -590 41370 -530
rect 41440 -590 41460 -530
rect 41350 -610 41460 -590
rect 41520 -530 41630 -510
rect 41520 -590 41540 -530
rect 41610 -590 41630 -530
rect 41520 -610 41630 -590
rect 41690 -530 41800 -510
rect 41690 -590 41710 -530
rect 41780 -590 41800 -530
rect 41690 -610 41800 -590
rect 41860 -530 41970 -510
rect 41860 -590 41880 -530
rect 41950 -590 41970 -530
rect 41860 -610 41970 -590
rect 42030 -530 42140 -510
rect 42030 -590 42050 -530
rect 42120 -590 42140 -530
rect 42030 -610 42140 -590
rect 42200 -530 42310 -510
rect 42200 -590 42220 -530
rect 42290 -590 42310 -530
rect 42200 -610 42310 -590
rect 42370 -530 42480 -510
rect 42370 -590 42390 -530
rect 42460 -590 42480 -530
rect 42370 -610 42480 -590
rect 42540 -530 42650 -510
rect 42540 -590 42560 -530
rect 42630 -590 42650 -530
rect 42540 -610 42650 -590
rect 42710 -530 42820 -510
rect 42710 -590 42730 -530
rect 42800 -590 42820 -530
rect 42710 -610 42820 -590
rect 42880 -530 42990 -510
rect 42880 -590 42900 -530
rect 42970 -590 42990 -530
rect 42880 -610 42990 -590
rect 43050 -530 43160 -510
rect 43050 -590 43070 -530
rect 43140 -590 43160 -530
rect 43050 -610 43160 -590
rect 43220 -530 43330 -510
rect 43220 -590 43240 -530
rect 43310 -590 43330 -530
rect 43220 -610 43330 -590
rect 43390 -530 43500 -510
rect 43390 -590 43410 -530
rect 43480 -590 43500 -530
rect 43390 -610 43500 -590
rect 43560 -530 43670 -510
rect 43560 -590 43580 -530
rect 43650 -590 43670 -530
rect 43560 -610 43670 -590
rect 43730 -530 43840 -510
rect 43730 -590 43750 -530
rect 43820 -590 43840 -530
rect 43730 -610 43840 -590
rect 43900 -530 44010 -510
rect 43900 -590 43920 -530
rect 43990 -590 44010 -530
rect 43900 -610 44010 -590
rect 44070 -530 44180 -510
rect 44070 -590 44090 -530
rect 44160 -590 44180 -530
rect 44070 -610 44180 -590
rect 44240 -530 44350 -510
rect 44240 -590 44260 -530
rect 44330 -590 44350 -530
rect 44240 -610 44350 -590
rect 44410 -530 44520 -510
rect 44410 -590 44430 -530
rect 44500 -590 44520 -530
rect 44410 -610 44520 -590
rect 44580 -530 44690 -510
rect 44580 -590 44600 -530
rect 44670 -590 44690 -530
rect 44580 -610 44690 -590
rect 44750 -530 44860 -510
rect 44750 -590 44770 -530
rect 44840 -590 44860 -530
rect 44750 -610 44860 -590
rect 44920 -530 45030 -510
rect 44920 -590 44940 -530
rect 45010 -590 45030 -530
rect 44920 -610 45030 -590
rect 45090 -530 45200 -510
rect 45090 -590 45110 -530
rect 45180 -590 45200 -530
rect 45090 -610 45200 -590
rect 45260 -530 45370 -510
rect 45260 -590 45280 -530
rect 45350 -590 45370 -530
rect 45260 -610 45370 -590
rect 45430 -530 45540 -510
rect 45430 -590 45450 -530
rect 45520 -590 45540 -530
rect 45430 -610 45540 -590
rect 45600 -530 45710 -510
rect 45600 -590 45620 -530
rect 45690 -590 45710 -530
rect 45600 -610 45710 -590
rect 45770 -530 45880 -510
rect 45770 -590 45790 -530
rect 45860 -590 45880 -530
rect 45770 -610 45880 -590
rect 45940 -530 46050 -510
rect 45940 -590 45960 -530
rect 46030 -590 46050 -530
rect 45940 -610 46050 -590
rect 46110 -530 46220 -510
rect 46110 -590 46130 -530
rect 46200 -590 46220 -530
rect 46110 -610 46220 -590
rect 46280 -530 46390 -510
rect 46280 -590 46300 -530
rect 46370 -590 46390 -530
rect 46280 -610 46390 -590
rect 46450 -530 46560 -510
rect 46450 -590 46470 -530
rect 46540 -590 46560 -530
rect 46450 -610 46560 -590
rect 46620 -530 46730 -510
rect 46620 -590 46640 -530
rect 46710 -590 46730 -530
rect 46620 -610 46730 -590
rect 46790 -530 46900 -510
rect 46790 -590 46810 -530
rect 46880 -590 46900 -530
rect 46790 -610 46900 -590
rect 46960 -530 47070 -510
rect 46960 -590 46980 -530
rect 47050 -590 47070 -530
rect 46960 -610 47070 -590
rect 47130 -530 47240 -510
rect 47130 -590 47150 -530
rect 47220 -590 47240 -530
rect 47130 -610 47240 -590
rect 47300 -530 47410 -510
rect 47300 -590 47320 -530
rect 47390 -590 47410 -530
rect 47300 -610 47410 -590
rect 47470 -530 47580 -510
rect 47470 -590 47490 -530
rect 47560 -590 47580 -530
rect 47470 -610 47580 -590
rect 47640 -530 47750 -510
rect 47640 -590 47660 -530
rect 47730 -590 47750 -530
rect 47640 -610 47750 -590
rect 47810 -530 47920 -510
rect 47810 -590 47830 -530
rect 47900 -590 47920 -530
rect 47810 -610 47920 -590
rect 47980 -530 48090 -510
rect 47980 -590 48000 -530
rect 48070 -590 48090 -530
rect 47980 -610 48090 -590
rect 48150 -530 48260 -510
rect 48150 -590 48170 -530
rect 48240 -590 48260 -530
rect 48150 -610 48260 -590
rect 48320 -530 48430 -510
rect 48320 -590 48340 -530
rect 48410 -590 48430 -530
rect 48320 -610 48430 -590
rect 48490 -530 48600 -510
rect 48490 -590 48510 -530
rect 48580 -590 48600 -530
rect 48490 -610 48600 -590
rect 48660 -530 48770 -510
rect 48660 -590 48680 -530
rect 48750 -590 48770 -530
rect 48660 -610 48770 -590
rect 48830 -530 48940 -510
rect 48830 -590 48850 -530
rect 48920 -590 48940 -530
rect 48830 -610 48940 -590
rect 49000 -530 49110 -510
rect 49000 -590 49020 -530
rect 49090 -590 49110 -530
rect 49000 -610 49110 -590
rect 49170 -530 49280 -510
rect 49170 -590 49190 -530
rect 49260 -590 49280 -530
rect 49170 -610 49280 -590
rect 49340 -530 49450 -510
rect 49340 -590 49360 -530
rect 49430 -590 49450 -530
rect 49340 -610 49450 -590
rect 49510 -530 49620 -510
rect 49510 -590 49530 -530
rect 49600 -590 49620 -530
rect 49510 -610 49620 -590
rect 49680 -530 49790 -510
rect 49680 -590 49700 -530
rect 49770 -590 49790 -530
rect 49680 -610 49790 -590
rect 49850 -530 49960 -510
rect 49850 -590 49870 -530
rect 49940 -590 49960 -530
rect 49850 -610 49960 -590
rect 50020 -530 50130 -510
rect 50020 -590 50040 -530
rect 50110 -590 50130 -530
rect 50020 -610 50130 -590
rect 50190 -530 50300 -510
rect 50190 -590 50210 -530
rect 50280 -590 50300 -530
rect 50190 -610 50300 -590
rect 50360 -530 50470 -510
rect 50360 -590 50380 -530
rect 50450 -590 50470 -530
rect 50360 -610 50470 -590
rect 50530 -530 50640 -510
rect 50530 -590 50550 -530
rect 50620 -590 50640 -530
rect 50530 -610 50640 -590
rect 50700 -530 50810 -510
rect 50700 -590 50720 -530
rect 50790 -590 50810 -530
rect 50700 -610 50810 -590
rect 50870 -530 50980 -510
rect 50870 -590 50890 -530
rect 50960 -590 50980 -530
rect 50870 -610 50980 -590
rect 51040 -530 51150 -510
rect 51040 -590 51060 -530
rect 51130 -590 51150 -530
rect 51040 -610 51150 -590
rect 51210 -530 51320 -510
rect 51210 -590 51230 -530
rect 51300 -590 51320 -530
rect 51210 -610 51320 -590
rect 51380 -530 51490 -510
rect 51380 -590 51400 -530
rect 51470 -590 51490 -530
rect 51380 -610 51490 -590
rect 51550 -530 51660 -510
rect 51550 -590 51570 -530
rect 51640 -590 51660 -530
rect 51550 -610 51660 -590
rect 51720 -530 51830 -510
rect 51720 -590 51740 -530
rect 51810 -590 51830 -530
rect 51720 -610 51830 -590
rect 51890 -530 52000 -510
rect 51890 -590 51910 -530
rect 51980 -590 52000 -530
rect 51890 -610 52000 -590
rect 52060 -530 52170 -510
rect 52060 -590 52080 -530
rect 52150 -590 52170 -530
rect 52060 -610 52170 -590
rect 52230 -530 52340 -510
rect 52230 -590 52250 -530
rect 52320 -590 52340 -530
rect 52230 -610 52340 -590
rect 52400 -530 52510 -510
rect 52400 -590 52420 -530
rect 52490 -590 52510 -530
rect 52400 -610 52510 -590
rect 52570 -530 52680 -510
rect 52570 -590 52590 -530
rect 52660 -590 52680 -530
rect 52570 -610 52680 -590
rect 52740 -530 52850 -510
rect 52740 -590 52760 -530
rect 52830 -590 52850 -530
rect 52740 -610 52850 -590
rect 52910 -530 53020 -510
rect 52910 -590 52930 -530
rect 53000 -590 53020 -530
rect 52910 -610 53020 -590
rect 53080 -530 53190 -510
rect 53080 -590 53100 -530
rect 53170 -590 53190 -530
rect 53080 -610 53190 -590
rect 53250 -530 53360 -510
rect 53250 -590 53270 -530
rect 53340 -590 53360 -530
rect 53250 -610 53360 -590
rect 53420 -530 53530 -510
rect 53420 -590 53440 -530
rect 53510 -590 53530 -530
rect 53420 -610 53530 -590
rect 53590 -530 53700 -510
rect 53590 -590 53610 -530
rect 53680 -590 53700 -530
rect 53590 -610 53700 -590
rect 53760 -530 53870 -510
rect 53760 -590 53780 -530
rect 53850 -590 53870 -530
rect 53760 -610 53870 -590
rect 53930 -530 54040 -510
rect 53930 -590 53950 -530
rect 54020 -590 54040 -530
rect 53930 -610 54040 -590
rect 54100 -530 54210 -510
rect 54100 -590 54120 -530
rect 54190 -590 54210 -530
rect 54100 -610 54210 -590
rect 54270 -530 54380 -510
rect 54270 -590 54290 -530
rect 54360 -590 54380 -530
rect 54270 -610 54380 -590
rect 54440 -530 54550 -510
rect 54440 -590 54460 -530
rect 54530 -590 54550 -530
rect 54440 -610 54550 -590
rect 54610 -530 54720 -510
rect 54610 -590 54630 -530
rect 54700 -590 54720 -530
rect 54610 -610 54720 -590
rect 54780 -530 54890 -510
rect 54780 -590 54800 -530
rect 54870 -590 54890 -530
rect 54780 -610 54890 -590
rect 54950 -530 55060 -510
rect 54950 -590 54970 -530
rect 55040 -590 55060 -530
rect 54950 -610 55060 -590
rect 55120 -530 55230 -510
rect 55120 -590 55140 -530
rect 55210 -590 55230 -530
rect 55120 -610 55230 -590
rect 55290 -530 55400 -510
rect 55290 -590 55310 -530
rect 55380 -590 55400 -530
rect 55290 -610 55400 -590
rect 55460 -530 55570 -510
rect 55460 -590 55480 -530
rect 55550 -590 55570 -530
rect 55460 -610 55570 -590
rect 55630 -530 55740 -510
rect 55630 -590 55650 -530
rect 55720 -590 55740 -530
rect 55630 -610 55740 -590
rect 55800 -530 55910 -510
rect 55800 -590 55820 -530
rect 55890 -590 55910 -530
rect 55800 -610 55910 -590
rect 55970 -530 56080 -510
rect 55970 -590 55990 -530
rect 56060 -590 56080 -530
rect 55970 -610 56080 -590
rect 56140 -530 56250 -510
rect 56140 -590 56160 -530
rect 56230 -590 56250 -530
rect 56140 -610 56250 -590
rect 56310 -530 56420 -510
rect 56310 -590 56330 -530
rect 56400 -590 56420 -530
rect 56310 -610 56420 -590
rect 56480 -530 56590 -510
rect 56480 -590 56500 -530
rect 56570 -590 56590 -530
rect 56480 -610 56590 -590
rect 56650 -530 56760 -510
rect 56650 -590 56670 -530
rect 56740 -590 56760 -530
rect 56650 -610 56760 -590
rect 56820 -530 56930 -510
rect 56820 -590 56840 -530
rect 56910 -590 56930 -530
rect 56820 -610 56930 -590
rect 56990 -530 57100 -510
rect 56990 -590 57010 -530
rect 57080 -590 57100 -530
rect 56990 -610 57100 -590
rect 57160 -530 57270 -510
rect 57160 -590 57180 -530
rect 57250 -590 57270 -530
rect 57160 -610 57270 -590
rect 57330 -530 57440 -510
rect 57330 -590 57350 -530
rect 57420 -590 57440 -530
rect 57330 -610 57440 -590
rect 57500 -530 57610 -510
rect 57500 -590 57520 -530
rect 57590 -590 57610 -530
rect 57500 -610 57610 -590
rect 57670 -530 57780 -510
rect 57670 -590 57690 -530
rect 57760 -590 57780 -530
rect 57670 -610 57780 -590
rect 57840 -530 57950 -510
rect 57840 -590 57860 -530
rect 57930 -590 57950 -530
rect 57840 -610 57950 -590
rect 58010 -530 58120 -510
rect 58010 -590 58030 -530
rect 58100 -590 58120 -530
rect 58010 -610 58120 -590
rect 58180 -530 58290 -510
rect 58180 -590 58200 -530
rect 58270 -590 58290 -530
rect 58180 -610 58290 -590
rect 58350 -530 58460 -510
rect 58350 -590 58370 -530
rect 58440 -590 58460 -530
rect 58350 -610 58460 -590
rect 58520 -530 58630 -510
rect 58520 -590 58540 -530
rect 58610 -590 58630 -530
rect 58520 -610 58630 -590
rect 58690 -530 58800 -510
rect 58690 -590 58710 -530
rect 58780 -590 58800 -530
rect 58690 -610 58800 -590
rect 58860 -530 58970 -510
rect 58860 -590 58880 -530
rect 58950 -590 58970 -530
rect 58860 -610 58970 -590
rect 59030 -530 59140 -510
rect 59030 -590 59050 -530
rect 59120 -590 59140 -530
rect 59030 -610 59140 -590
rect 59200 -530 59310 -510
rect 59200 -590 59220 -530
rect 59290 -590 59310 -530
rect 59200 -610 59310 -590
rect 59370 -530 59480 -510
rect 59370 -590 59390 -530
rect 59460 -590 59480 -530
rect 59370 -610 59480 -590
rect 59540 -530 59650 -510
rect 59540 -590 59560 -530
rect 59630 -590 59650 -530
rect 59540 -610 59650 -590
rect 59710 -530 59820 -510
rect 59710 -590 59730 -530
rect 59800 -590 59820 -530
rect 59710 -610 59820 -590
rect 59880 -530 59990 -510
rect 59880 -590 59900 -530
rect 59970 -590 59990 -530
rect 59880 -610 59990 -590
rect 60050 -530 60160 -510
rect 60050 -590 60070 -530
rect 60140 -590 60160 -530
rect 60050 -610 60160 -590
rect 60220 -530 60330 -510
rect 60220 -590 60240 -530
rect 60310 -590 60330 -530
rect 60220 -610 60330 -590
rect 60390 -530 60500 -510
rect 60390 -590 60410 -530
rect 60480 -590 60500 -530
rect 60390 -610 60500 -590
rect 60560 -530 60670 -510
rect 60560 -590 60580 -530
rect 60650 -590 60670 -530
rect 60560 -610 60670 -590
rect 60730 -530 60840 -510
rect 60730 -590 60750 -530
rect 60820 -590 60840 -530
rect 60730 -610 60840 -590
rect 60900 -530 61010 -510
rect 60900 -590 60920 -530
rect 60990 -590 61010 -530
rect 60900 -610 61010 -590
rect 61070 -530 61180 -510
rect 61070 -590 61090 -530
rect 61160 -590 61180 -530
rect 61070 -610 61180 -590
rect 61240 -530 61350 -510
rect 61240 -590 61260 -530
rect 61330 -590 61350 -530
rect 61240 -610 61350 -590
rect 61410 -530 61520 -510
rect 61410 -590 61430 -530
rect 61500 -590 61520 -530
rect 61410 -610 61520 -590
rect 61580 -530 61690 -510
rect 61580 -590 61600 -530
rect 61670 -590 61690 -530
rect 61580 -610 61690 -590
rect 61750 -530 61860 -510
rect 61750 -590 61770 -530
rect 61840 -590 61860 -530
rect 61750 -610 61860 -590
rect 61920 -530 62030 -510
rect 61920 -590 61940 -530
rect 62010 -590 62030 -530
rect 61920 -610 62030 -590
rect 62090 -530 62200 -510
rect 62090 -590 62110 -530
rect 62180 -590 62200 -530
rect 62090 -610 62200 -590
rect 62260 -530 62370 -510
rect 62260 -590 62280 -530
rect 62350 -590 62370 -530
rect 62260 -610 62370 -590
rect 62430 -530 62540 -510
rect 62430 -590 62450 -530
rect 62520 -590 62540 -530
rect 62430 -610 62540 -590
rect 62600 -530 62710 -510
rect 62600 -590 62620 -530
rect 62690 -590 62710 -530
rect 62600 -610 62710 -590
rect 62770 -530 62880 -510
rect 62770 -590 62790 -530
rect 62860 -590 62880 -530
rect 62770 -610 62880 -590
rect 62940 -530 63050 -510
rect 62940 -590 62960 -530
rect 63030 -590 63050 -530
rect 62940 -610 63050 -590
rect 63110 -530 63220 -510
rect 63110 -590 63130 -530
rect 63200 -590 63220 -530
rect 63110 -610 63220 -590
rect 63280 -530 63390 -510
rect 63280 -590 63300 -530
rect 63370 -590 63390 -530
rect 63280 -610 63390 -590
rect 63450 -530 63560 -510
rect 63450 -590 63470 -530
rect 63540 -590 63560 -530
rect 63450 -610 63560 -590
rect 63620 -530 63730 -510
rect 63620 -590 63640 -530
rect 63710 -590 63730 -530
rect 63620 -610 63730 -590
rect 63790 -530 63900 -510
rect 63790 -590 63810 -530
rect 63880 -590 63900 -530
rect 63790 -610 63900 -590
rect 63960 -530 64070 -510
rect 63960 -590 63980 -530
rect 64050 -590 64070 -530
rect 63960 -610 64070 -590
rect 64130 -530 64240 -510
rect 64130 -590 64150 -530
rect 64220 -590 64240 -530
rect 64130 -610 64240 -590
rect 64300 -530 64410 -510
rect 64300 -590 64320 -530
rect 64390 -590 64410 -530
rect 64300 -610 64410 -590
rect 64470 -530 64580 -510
rect 64470 -590 64490 -530
rect 64560 -590 64580 -530
rect 64470 -610 64580 -590
rect 64640 -530 64750 -510
rect 64640 -590 64660 -530
rect 64730 -590 64750 -530
rect 64640 -610 64750 -590
rect 64810 -530 64920 -510
rect 64810 -590 64830 -530
rect 64900 -590 64920 -530
rect 64810 -610 64920 -590
rect 64980 -530 65090 -510
rect 64980 -590 65000 -530
rect 65070 -590 65090 -530
rect 64980 -610 65090 -590
rect 65150 -530 65260 -510
rect 65150 -590 65170 -530
rect 65240 -590 65260 -530
rect 65150 -610 65260 -590
rect 65320 -530 65430 -510
rect 65320 -590 65340 -530
rect 65410 -590 65430 -530
rect 65320 -610 65430 -590
rect 65490 -530 65600 -510
rect 65490 -590 65510 -530
rect 65580 -590 65600 -530
rect 65490 -610 65600 -590
rect 65660 -530 65770 -510
rect 65660 -590 65680 -530
rect 65750 -590 65770 -530
rect 65660 -610 65770 -590
rect 65830 -530 65940 -510
rect 65830 -590 65850 -530
rect 65920 -590 65940 -530
rect 65830 -610 65940 -590
rect 66000 -530 66110 -510
rect 66000 -590 66020 -530
rect 66090 -590 66110 -530
rect 66000 -610 66110 -590
rect 66170 -530 66280 -510
rect 66170 -590 66190 -530
rect 66260 -590 66280 -530
rect 66170 -610 66280 -590
rect 66340 -530 66450 -510
rect 66340 -590 66360 -530
rect 66430 -590 66450 -530
rect 66340 -610 66450 -590
rect 66510 -530 66620 -510
rect 66510 -590 66530 -530
rect 66600 -590 66620 -530
rect 66510 -610 66620 -590
rect 66680 -530 66790 -510
rect 66680 -590 66700 -530
rect 66770 -590 66790 -530
rect 66680 -610 66790 -590
rect 66850 -530 66960 -510
rect 66850 -590 66870 -530
rect 66940 -590 66960 -530
rect 66850 -610 66960 -590
rect 67020 -530 67130 -510
rect 67020 -590 67040 -530
rect 67110 -590 67130 -530
rect 67020 -610 67130 -590
rect 67190 -530 67300 -510
rect 67190 -590 67210 -530
rect 67280 -590 67300 -530
rect 67190 -610 67300 -590
rect 67360 -530 67470 -510
rect 67360 -590 67380 -530
rect 67450 -590 67470 -530
rect 67360 -610 67470 -590
rect 67530 -530 67640 -510
rect 67530 -590 67550 -530
rect 67620 -590 67640 -530
rect 67530 -610 67640 -590
rect 67700 -530 67810 -510
rect 67700 -590 67720 -530
rect 67790 -590 67810 -530
rect 67700 -610 67810 -590
rect 67870 -530 67980 -510
rect 67870 -590 67890 -530
rect 67960 -590 67980 -530
rect 67870 -610 67980 -590
rect 68040 -530 68150 -510
rect 68040 -590 68060 -530
rect 68130 -590 68150 -530
rect 68040 -610 68150 -590
rect 68210 -530 68320 -510
rect 68210 -590 68230 -530
rect 68300 -590 68320 -530
rect 68210 -610 68320 -590
rect 68380 -530 68490 -510
rect 68380 -590 68400 -530
rect 68470 -590 68490 -530
rect 68380 -610 68490 -590
rect 68550 -530 68660 -510
rect 68550 -590 68570 -530
rect 68640 -590 68660 -530
rect 68550 -610 68660 -590
rect 68720 -530 68830 -510
rect 68720 -590 68740 -530
rect 68810 -590 68830 -530
rect 68720 -610 68830 -590
rect 68890 -530 69000 -510
rect 68890 -590 68910 -530
rect 68980 -590 69000 -530
rect 68890 -610 69000 -590
rect 69060 -530 69170 -510
rect 69060 -590 69080 -530
rect 69150 -590 69170 -530
rect 69060 -610 69170 -590
rect 69230 -530 69340 -510
rect 69230 -590 69250 -530
rect 69320 -590 69340 -530
rect 69230 -610 69340 -590
rect 69400 -530 69510 -510
rect 69400 -590 69420 -530
rect 69490 -590 69510 -530
rect 69400 -610 69510 -590
rect 69570 -530 69680 -510
rect 69570 -590 69590 -530
rect 69660 -590 69680 -530
rect 69570 -610 69680 -590
rect 69740 -530 69850 -510
rect 69740 -590 69760 -530
rect 69830 -590 69850 -530
rect 69740 -610 69850 -590
rect 69910 -530 70020 -510
rect 69910 -590 69930 -530
rect 70000 -590 70020 -530
rect 69910 -610 70020 -590
rect 70080 -530 70190 -510
rect 70080 -590 70100 -530
rect 70170 -590 70190 -530
rect 70080 -610 70190 -590
rect 70250 -530 70360 -510
rect 70250 -590 70270 -530
rect 70340 -590 70360 -530
rect 70250 -610 70360 -590
rect 70420 -530 70530 -510
rect 70420 -590 70440 -530
rect 70510 -590 70530 -530
rect 70420 -610 70530 -590
rect 70590 -530 70700 -510
rect 70590 -590 70610 -530
rect 70680 -590 70700 -530
rect 70590 -610 70700 -590
rect 70760 -530 70870 -510
rect 70760 -590 70780 -530
rect 70850 -590 70870 -530
rect 70760 -610 70870 -590
rect 70930 -530 71040 -510
rect 70930 -590 70950 -530
rect 71020 -590 71040 -530
rect 70930 -610 71040 -590
rect 71100 -530 71210 -510
rect 71100 -590 71120 -530
rect 71190 -590 71210 -530
rect 71100 -610 71210 -590
rect 71270 -530 71380 -510
rect 71270 -590 71290 -530
rect 71360 -590 71380 -530
rect 71270 -610 71380 -590
rect 71440 -530 71550 -510
rect 71440 -590 71460 -530
rect 71530 -590 71550 -530
rect 71440 -610 71550 -590
rect 71610 -530 71720 -510
rect 71610 -590 71630 -530
rect 71700 -590 71720 -530
rect 71610 -610 71720 -590
rect 71780 -530 71890 -510
rect 71780 -590 71800 -530
rect 71870 -590 71890 -530
rect 71780 -610 71890 -590
rect 71950 -530 72060 -510
rect 71950 -590 71970 -530
rect 72040 -590 72060 -530
rect 71950 -610 72060 -590
rect 72120 -530 72230 -510
rect 72120 -590 72140 -530
rect 72210 -590 72230 -530
rect 72120 -610 72230 -590
rect 72290 -530 72400 -510
rect 72290 -590 72310 -530
rect 72380 -590 72400 -530
rect 72290 -610 72400 -590
rect 72460 -530 72570 -510
rect 72460 -590 72480 -530
rect 72550 -590 72570 -530
rect 72460 -610 72570 -590
rect 72630 -530 72740 -510
rect 72630 -590 72650 -530
rect 72720 -590 72740 -530
rect 72630 -610 72740 -590
rect 72800 -530 72910 -510
rect 72800 -590 72820 -530
rect 72890 -590 72910 -530
rect 72800 -610 72910 -590
rect 72970 -530 73080 -510
rect 72970 -590 72990 -530
rect 73060 -590 73080 -530
rect 72970 -610 73080 -590
rect 73140 -530 73250 -510
rect 73140 -590 73160 -530
rect 73230 -590 73250 -530
rect 73140 -610 73250 -590
rect 73310 -530 73420 -510
rect 73310 -590 73330 -530
rect 73400 -590 73420 -530
rect 73310 -610 73420 -590
rect 73480 -530 73590 -510
rect 73480 -590 73500 -530
rect 73570 -590 73590 -530
rect 73480 -610 73590 -590
rect 73650 -530 73760 -510
rect 73650 -590 73670 -530
rect 73740 -590 73760 -530
rect 73650 -610 73760 -590
rect 73820 -530 73930 -510
rect 73820 -590 73840 -530
rect 73910 -590 73930 -530
rect 73820 -610 73930 -590
rect 73990 -530 74100 -510
rect 73990 -590 74010 -530
rect 74080 -590 74100 -530
rect 73990 -610 74100 -590
rect 74160 -530 74270 -510
rect 74160 -590 74180 -530
rect 74250 -590 74270 -530
rect 74160 -610 74270 -590
rect 74330 -530 74440 -510
rect 74330 -590 74350 -530
rect 74420 -590 74440 -530
rect 74330 -610 74440 -590
rect 74500 -530 74610 -510
rect 74500 -590 74520 -530
rect 74590 -590 74610 -530
rect 74500 -610 74610 -590
rect 74670 -530 74780 -510
rect 74670 -590 74690 -530
rect 74760 -590 74780 -530
rect 74670 -610 74780 -590
rect 74840 -530 74950 -510
rect 74840 -590 74860 -530
rect 74930 -590 74950 -530
rect 74840 -610 74950 -590
rect 75010 -530 75120 -510
rect 75010 -590 75030 -530
rect 75100 -590 75120 -530
rect 75010 -610 75120 -590
rect 75180 -530 75290 -510
rect 75180 -590 75200 -530
rect 75270 -590 75290 -530
rect 75180 -610 75290 -590
rect 75350 -530 75460 -510
rect 75350 -590 75370 -530
rect 75440 -590 75460 -530
rect 75350 -610 75460 -590
rect 75520 -530 75630 -510
rect 75520 -590 75540 -530
rect 75610 -590 75630 -530
rect 75520 -610 75630 -590
rect 75690 -530 75800 -510
rect 75690 -590 75710 -530
rect 75780 -590 75800 -530
rect 75690 -610 75800 -590
rect 75860 -530 75970 -510
rect 75860 -590 75880 -530
rect 75950 -590 75970 -530
rect 75860 -610 75970 -590
rect 76030 -530 76140 -510
rect 76030 -590 76050 -530
rect 76120 -590 76140 -530
rect 76030 -610 76140 -590
rect 76200 -530 76310 -510
rect 76200 -590 76220 -530
rect 76290 -590 76310 -530
rect 76200 -610 76310 -590
rect 76370 -530 76480 -510
rect 76370 -590 76390 -530
rect 76460 -590 76480 -530
rect 76370 -610 76480 -590
rect 76540 -530 76650 -510
rect 76540 -590 76560 -530
rect 76630 -590 76650 -530
rect 76540 -610 76650 -590
rect 76710 -530 76820 -510
rect 76710 -590 76730 -530
rect 76800 -590 76820 -530
rect 76710 -610 76820 -590
rect 76880 -530 76990 -510
rect 76880 -590 76900 -530
rect 76970 -590 76990 -530
rect 76880 -610 76990 -590
rect 77050 -530 77160 -510
rect 77050 -590 77070 -530
rect 77140 -590 77160 -530
rect 77050 -610 77160 -590
rect 77220 -530 77330 -510
rect 77220 -590 77240 -530
rect 77310 -590 77330 -530
rect 77220 -610 77330 -590
rect 77390 -530 77500 -510
rect 77390 -590 77410 -530
rect 77480 -590 77500 -530
rect 77390 -610 77500 -590
rect 77560 -530 77670 -510
rect 77560 -590 77580 -530
rect 77650 -590 77670 -530
rect 77560 -610 77670 -590
rect 77730 -530 77840 -510
rect 77730 -590 77750 -530
rect 77820 -590 77840 -530
rect 77730 -610 77840 -590
rect 77900 -530 78010 -510
rect 77900 -590 77920 -530
rect 77990 -590 78010 -530
rect 77900 -610 78010 -590
rect 78070 -530 78180 -510
rect 78070 -590 78090 -530
rect 78160 -590 78180 -530
rect 78070 -610 78180 -590
rect 78240 -530 78350 -510
rect 78240 -590 78260 -530
rect 78330 -590 78350 -530
rect 78240 -610 78350 -590
rect 78410 -530 78520 -510
rect 78410 -590 78430 -530
rect 78500 -590 78520 -530
rect 78410 -610 78520 -590
rect 78580 -530 78690 -510
rect 78580 -590 78600 -530
rect 78670 -590 78690 -530
rect 78580 -610 78690 -590
rect 78750 -530 78860 -510
rect 78750 -590 78770 -530
rect 78840 -590 78860 -530
rect 78750 -610 78860 -590
rect 78920 -530 79030 -510
rect 78920 -590 78940 -530
rect 79010 -590 79030 -530
rect 78920 -610 79030 -590
rect 79090 -530 79200 -510
rect 79090 -590 79110 -530
rect 79180 -590 79200 -530
rect 79090 -610 79200 -590
rect 79260 -530 79370 -510
rect 79260 -590 79280 -530
rect 79350 -590 79370 -530
rect 79260 -610 79370 -590
rect 79430 -530 79540 -510
rect 79430 -590 79450 -530
rect 79520 -590 79540 -530
rect 79430 -610 79540 -590
rect 79600 -530 79710 -510
rect 79600 -590 79620 -530
rect 79690 -590 79710 -530
rect 79600 -610 79710 -590
rect 79770 -530 79880 -510
rect 79770 -590 79790 -530
rect 79860 -590 79880 -530
rect 79770 -610 79880 -590
rect 79940 -530 80050 -510
rect 79940 -590 79960 -530
rect 80030 -590 80050 -530
rect 79940 -610 80050 -590
rect 80110 -530 80220 -510
rect 80110 -590 80130 -530
rect 80200 -590 80220 -530
rect 80110 -610 80220 -590
rect 80280 -530 80390 -510
rect 80280 -590 80300 -530
rect 80370 -590 80390 -530
rect 80280 -610 80390 -590
rect 80450 -530 80560 -510
rect 80450 -590 80470 -530
rect 80540 -590 80560 -530
rect 80450 -610 80560 -590
rect 80620 -530 80730 -510
rect 80620 -590 80640 -530
rect 80710 -590 80730 -530
rect 80620 -610 80730 -590
rect 80790 -530 80900 -510
rect 80790 -590 80810 -530
rect 80880 -590 80900 -530
rect 80790 -610 80900 -590
rect 80960 -530 81070 -510
rect 80960 -590 80980 -530
rect 81050 -590 81070 -530
rect 80960 -610 81070 -590
rect 81130 -530 81240 -510
rect 81130 -590 81150 -530
rect 81220 -590 81240 -530
rect 81130 -610 81240 -590
rect 81300 -530 81410 -510
rect 81300 -590 81320 -530
rect 81390 -590 81410 -530
rect 81300 -610 81410 -590
rect 81470 -530 81580 -510
rect 81470 -590 81490 -530
rect 81560 -590 81580 -530
rect 81470 -610 81580 -590
rect 81640 -530 81750 -510
rect 81640 -590 81660 -530
rect 81730 -590 81750 -530
rect 81640 -610 81750 -590
rect 81810 -530 81920 -510
rect 81810 -590 81830 -530
rect 81900 -590 81920 -530
rect 81810 -610 81920 -590
rect 81980 -530 82090 -510
rect 81980 -590 82000 -530
rect 82070 -590 82090 -530
rect 81980 -610 82090 -590
rect 82150 -530 82260 -510
rect 82150 -590 82170 -530
rect 82240 -590 82260 -530
rect 82150 -610 82260 -590
rect 82320 -530 82430 -510
rect 82320 -590 82340 -530
rect 82410 -590 82430 -530
rect 82320 -610 82430 -590
rect 82490 -530 82600 -510
rect 82490 -590 82510 -530
rect 82580 -590 82600 -530
rect 82490 -610 82600 -590
rect 82660 -530 82770 -510
rect 82660 -590 82680 -530
rect 82750 -590 82770 -530
rect 82660 -610 82770 -590
rect 82830 -530 82940 -510
rect 82830 -590 82850 -530
rect 82920 -590 82940 -530
rect 82830 -610 82940 -590
rect 83000 -530 83110 -510
rect 83000 -590 83020 -530
rect 83090 -590 83110 -530
rect 83000 -610 83110 -590
rect 83170 -530 83280 -510
rect 83170 -590 83190 -530
rect 83260 -590 83280 -530
rect 83170 -610 83280 -590
rect 83340 -530 83450 -510
rect 83340 -590 83360 -530
rect 83430 -590 83450 -530
rect 83340 -610 83450 -590
rect 83510 -530 83620 -510
rect 83510 -590 83530 -530
rect 83600 -590 83620 -530
rect 83510 -610 83620 -590
rect 83680 -530 83790 -510
rect 83680 -590 83700 -530
rect 83770 -590 83790 -530
rect 83680 -610 83790 -590
rect 83850 -530 83960 -510
rect 83850 -590 83870 -530
rect 83940 -590 83960 -530
rect 83850 -610 83960 -590
rect 84020 -530 84130 -510
rect 84020 -590 84040 -530
rect 84110 -590 84130 -530
rect 84020 -610 84130 -590
rect 84190 -530 84300 -510
rect 84190 -590 84210 -530
rect 84280 -590 84300 -530
rect 84190 -610 84300 -590
rect 84360 -530 84470 -510
rect 84360 -590 84380 -530
rect 84450 -590 84470 -530
rect 84360 -610 84470 -590
rect 84530 -530 84640 -510
rect 84530 -590 84550 -530
rect 84620 -590 84640 -530
rect 84530 -610 84640 -590
rect 84700 -530 84810 -510
rect 84700 -590 84720 -530
rect 84790 -590 84810 -530
rect 84700 -610 84810 -590
rect 84870 -530 84980 -510
rect 84870 -590 84890 -530
rect 84960 -590 84980 -530
rect 84870 -610 84980 -590
rect 85040 -530 85150 -510
rect 85040 -590 85060 -530
rect 85130 -590 85150 -530
rect 85040 -610 85150 -590
rect 85210 -530 85320 -510
rect 85210 -590 85230 -530
rect 85300 -590 85320 -530
rect 85210 -610 85320 -590
rect 85380 -530 85490 -510
rect 85380 -590 85400 -530
rect 85470 -590 85490 -530
rect 85380 -610 85490 -590
rect 85550 -530 85660 -510
rect 85550 -590 85570 -530
rect 85640 -590 85660 -530
rect 85550 -610 85660 -590
rect 85720 -530 85830 -510
rect 85720 -590 85740 -530
rect 85810 -590 85830 -530
rect 85720 -610 85830 -590
rect 85890 -530 86000 -510
rect 85890 -590 85910 -530
rect 85980 -590 86000 -530
rect 85890 -610 86000 -590
rect 86060 -530 86170 -510
rect 86060 -590 86080 -530
rect 86150 -590 86170 -530
rect 86060 -610 86170 -590
rect 86230 -530 86340 -510
rect 86230 -590 86250 -530
rect 86320 -590 86340 -530
rect 86230 -610 86340 -590
rect 86400 -530 86510 -510
rect 86400 -590 86420 -530
rect 86490 -590 86510 -530
rect 86400 -610 86510 -590
rect 86570 -530 86680 -510
rect 86570 -590 86590 -530
rect 86660 -590 86680 -530
rect 86570 -610 86680 -590
rect 86740 -530 86850 -510
rect 86740 -590 86760 -530
rect 86830 -590 86850 -530
rect 86740 -610 86850 -590
rect 86910 -530 87020 -510
rect 86910 -590 86930 -530
rect 87000 -590 87020 -530
rect 86910 -610 87020 -590
rect 87080 -530 87190 -510
rect 87080 -590 87100 -530
rect 87170 -590 87190 -530
rect 87080 -610 87190 -590
rect 130 -670 230 -650
rect 130 -730 150 -670
rect 210 -730 230 -670
rect 130 -750 230 -730
rect 470 -670 570 -650
rect 470 -730 490 -670
rect 550 -730 570 -670
rect 470 -750 570 -730
rect 810 -670 910 -650
rect 810 -730 830 -670
rect 890 -730 910 -670
rect 810 -750 910 -730
rect 1150 -670 1250 -650
rect 1150 -730 1170 -670
rect 1230 -730 1250 -670
rect 1150 -750 1250 -730
rect 1490 -670 1590 -650
rect 1490 -730 1510 -670
rect 1570 -730 1590 -670
rect 1490 -750 1590 -730
rect 1830 -670 1930 -650
rect 1830 -730 1850 -670
rect 1910 -730 1930 -670
rect 1830 -750 1930 -730
rect 2170 -670 2270 -650
rect 2170 -730 2190 -670
rect 2250 -730 2270 -670
rect 2170 -750 2270 -730
rect 2510 -670 2610 -650
rect 2510 -730 2530 -670
rect 2590 -730 2610 -670
rect 2510 -750 2610 -730
rect 2850 -670 2950 -650
rect 2850 -730 2870 -670
rect 2930 -730 2950 -670
rect 2850 -750 2950 -730
rect 3190 -670 3290 -650
rect 3190 -730 3210 -670
rect 3270 -730 3290 -670
rect 3190 -750 3290 -730
rect 3530 -670 3630 -650
rect 3530 -730 3550 -670
rect 3610 -730 3630 -670
rect 3530 -750 3630 -730
rect 3870 -670 3970 -650
rect 3870 -730 3890 -670
rect 3950 -730 3970 -670
rect 3870 -750 3970 -730
rect 4210 -670 4310 -650
rect 4210 -730 4230 -670
rect 4290 -730 4310 -670
rect 4210 -750 4310 -730
rect 4550 -670 4650 -650
rect 4550 -730 4570 -670
rect 4630 -730 4650 -670
rect 4550 -750 4650 -730
rect 4890 -670 4990 -650
rect 4890 -730 4910 -670
rect 4970 -730 4990 -670
rect 4890 -750 4990 -730
rect 5230 -670 5330 -650
rect 5230 -730 5250 -670
rect 5310 -730 5330 -670
rect 5230 -750 5330 -730
rect 5570 -670 5670 -650
rect 5570 -730 5590 -670
rect 5650 -730 5670 -670
rect 5570 -750 5670 -730
rect 5910 -670 6010 -650
rect 5910 -730 5930 -670
rect 5990 -730 6010 -670
rect 5910 -750 6010 -730
rect 6250 -670 6350 -650
rect 6250 -730 6270 -670
rect 6330 -730 6350 -670
rect 6250 -750 6350 -730
rect 6590 -670 6690 -650
rect 6590 -730 6610 -670
rect 6670 -730 6690 -670
rect 6590 -750 6690 -730
rect 6930 -670 7030 -650
rect 6930 -730 6950 -670
rect 7010 -730 7030 -670
rect 6930 -750 7030 -730
rect 7270 -670 7370 -650
rect 7270 -730 7290 -670
rect 7350 -730 7370 -670
rect 7270 -750 7370 -730
rect 7610 -670 7710 -650
rect 7610 -730 7630 -670
rect 7690 -730 7710 -670
rect 7610 -750 7710 -730
rect 7950 -670 8050 -650
rect 7950 -730 7970 -670
rect 8030 -730 8050 -670
rect 7950 -750 8050 -730
rect 8290 -670 8390 -650
rect 8290 -730 8310 -670
rect 8370 -730 8390 -670
rect 8290 -750 8390 -730
rect 8630 -670 8730 -650
rect 8630 -730 8650 -670
rect 8710 -730 8730 -670
rect 8630 -750 8730 -730
rect 8970 -670 9070 -650
rect 8970 -730 8990 -670
rect 9050 -730 9070 -670
rect 8970 -750 9070 -730
rect 9310 -670 9410 -650
rect 9310 -730 9330 -670
rect 9390 -730 9410 -670
rect 9310 -750 9410 -730
rect 9650 -670 9750 -650
rect 9650 -730 9670 -670
rect 9730 -730 9750 -670
rect 9650 -750 9750 -730
rect 9990 -670 10090 -650
rect 9990 -730 10010 -670
rect 10070 -730 10090 -670
rect 9990 -750 10090 -730
rect 10330 -670 10430 -650
rect 10330 -730 10350 -670
rect 10410 -730 10430 -670
rect 10330 -750 10430 -730
rect 10670 -670 10770 -650
rect 10670 -730 10690 -670
rect 10750 -730 10770 -670
rect 10670 -750 10770 -730
rect 11010 -670 11110 -650
rect 11010 -730 11030 -670
rect 11090 -730 11110 -670
rect 11010 -750 11110 -730
rect 11350 -670 11450 -650
rect 11350 -730 11370 -670
rect 11430 -730 11450 -670
rect 11350 -750 11450 -730
rect 11690 -670 11790 -650
rect 11690 -730 11710 -670
rect 11770 -730 11790 -670
rect 11690 -750 11790 -730
rect 12030 -670 12130 -650
rect 12030 -730 12050 -670
rect 12110 -730 12130 -670
rect 12030 -750 12130 -730
rect 12370 -670 12470 -650
rect 12370 -730 12390 -670
rect 12450 -730 12470 -670
rect 12370 -750 12470 -730
rect 12710 -670 12810 -650
rect 12710 -730 12730 -670
rect 12790 -730 12810 -670
rect 12710 -750 12810 -730
rect 13050 -670 13150 -650
rect 13050 -730 13070 -670
rect 13130 -730 13150 -670
rect 13050 -750 13150 -730
rect 13390 -670 13490 -650
rect 13390 -730 13410 -670
rect 13470 -730 13490 -670
rect 13390 -750 13490 -730
rect 13730 -670 13830 -650
rect 13730 -730 13750 -670
rect 13810 -730 13830 -670
rect 13730 -750 13830 -730
rect 14070 -670 14170 -650
rect 14070 -730 14090 -670
rect 14150 -730 14170 -670
rect 14070 -750 14170 -730
rect 14410 -670 14510 -650
rect 14410 -730 14430 -670
rect 14490 -730 14510 -670
rect 14410 -750 14510 -730
rect 14750 -670 14850 -650
rect 14750 -730 14770 -670
rect 14830 -730 14850 -670
rect 14750 -750 14850 -730
rect 15090 -670 15190 -650
rect 15090 -730 15110 -670
rect 15170 -730 15190 -670
rect 15090 -750 15190 -730
rect 15430 -670 15530 -650
rect 15430 -730 15450 -670
rect 15510 -730 15530 -670
rect 15430 -750 15530 -730
rect 15770 -670 15870 -650
rect 15770 -730 15790 -670
rect 15850 -730 15870 -670
rect 15770 -750 15870 -730
rect 16110 -670 16210 -650
rect 16110 -730 16130 -670
rect 16190 -730 16210 -670
rect 16110 -750 16210 -730
rect 16450 -670 16550 -650
rect 16450 -730 16470 -670
rect 16530 -730 16550 -670
rect 16450 -750 16550 -730
rect 16790 -670 16890 -650
rect 16790 -730 16810 -670
rect 16870 -730 16890 -670
rect 16790 -750 16890 -730
rect 17130 -670 17230 -650
rect 17130 -730 17150 -670
rect 17210 -730 17230 -670
rect 17130 -750 17230 -730
rect 17470 -670 17570 -650
rect 17470 -730 17490 -670
rect 17550 -730 17570 -670
rect 17470 -750 17570 -730
rect 17810 -670 17910 -650
rect 17810 -730 17830 -670
rect 17890 -730 17910 -670
rect 17810 -750 17910 -730
rect 18150 -670 18250 -650
rect 18150 -730 18170 -670
rect 18230 -730 18250 -670
rect 18150 -750 18250 -730
rect 18490 -670 18590 -650
rect 18490 -730 18510 -670
rect 18570 -730 18590 -670
rect 18490 -750 18590 -730
rect 18830 -670 18930 -650
rect 18830 -730 18850 -670
rect 18910 -730 18930 -670
rect 18830 -750 18930 -730
rect 19170 -670 19270 -650
rect 19170 -730 19190 -670
rect 19250 -730 19270 -670
rect 19170 -750 19270 -730
rect 19510 -670 19610 -650
rect 19510 -730 19530 -670
rect 19590 -730 19610 -670
rect 19510 -750 19610 -730
rect 19850 -670 19950 -650
rect 19850 -730 19870 -670
rect 19930 -730 19950 -670
rect 19850 -750 19950 -730
rect 20190 -670 20290 -650
rect 20190 -730 20210 -670
rect 20270 -730 20290 -670
rect 20190 -750 20290 -730
rect 20530 -670 20630 -650
rect 20530 -730 20550 -670
rect 20610 -730 20630 -670
rect 20530 -750 20630 -730
rect 20870 -670 20970 -650
rect 20870 -730 20890 -670
rect 20950 -730 20970 -670
rect 20870 -750 20970 -730
rect 21210 -670 21310 -650
rect 21210 -730 21230 -670
rect 21290 -730 21310 -670
rect 21210 -750 21310 -730
rect 21550 -670 21650 -650
rect 21550 -730 21570 -670
rect 21630 -730 21650 -670
rect 21550 -750 21650 -730
rect 21890 -670 21990 -650
rect 21890 -730 21910 -670
rect 21970 -730 21990 -670
rect 21890 -750 21990 -730
rect 22230 -670 22330 -650
rect 22230 -730 22250 -670
rect 22310 -730 22330 -670
rect 22230 -750 22330 -730
rect 22570 -670 22670 -650
rect 22570 -730 22590 -670
rect 22650 -730 22670 -670
rect 22570 -750 22670 -730
rect 22910 -670 23010 -650
rect 22910 -730 22930 -670
rect 22990 -730 23010 -670
rect 22910 -750 23010 -730
rect 23250 -670 23350 -650
rect 23250 -730 23270 -670
rect 23330 -730 23350 -670
rect 23250 -750 23350 -730
rect 23590 -670 23690 -650
rect 23590 -730 23610 -670
rect 23670 -730 23690 -670
rect 23590 -750 23690 -730
rect 23930 -670 24030 -650
rect 23930 -730 23950 -670
rect 24010 -730 24030 -670
rect 23930 -750 24030 -730
rect 24270 -670 24370 -650
rect 24270 -730 24290 -670
rect 24350 -730 24370 -670
rect 24270 -750 24370 -730
rect 24610 -670 24710 -650
rect 24610 -730 24630 -670
rect 24690 -730 24710 -670
rect 24610 -750 24710 -730
rect 24950 -670 25050 -650
rect 24950 -730 24970 -670
rect 25030 -730 25050 -670
rect 24950 -750 25050 -730
rect 25290 -670 25390 -650
rect 25290 -730 25310 -670
rect 25370 -730 25390 -670
rect 25290 -750 25390 -730
rect 25630 -670 25730 -650
rect 25630 -730 25650 -670
rect 25710 -730 25730 -670
rect 25630 -750 25730 -730
rect 25970 -670 26070 -650
rect 25970 -730 25990 -670
rect 26050 -730 26070 -670
rect 25970 -750 26070 -730
rect 26310 -670 26410 -650
rect 26310 -730 26330 -670
rect 26390 -730 26410 -670
rect 26310 -750 26410 -730
rect 26650 -670 26750 -650
rect 26650 -730 26670 -670
rect 26730 -730 26750 -670
rect 26650 -750 26750 -730
rect 26990 -670 27090 -650
rect 26990 -730 27010 -670
rect 27070 -730 27090 -670
rect 26990 -750 27090 -730
rect 27330 -670 27430 -650
rect 27330 -730 27350 -670
rect 27410 -730 27430 -670
rect 27330 -750 27430 -730
rect 27670 -670 27770 -650
rect 27670 -730 27690 -670
rect 27750 -730 27770 -670
rect 27670 -750 27770 -730
rect 28010 -670 28110 -650
rect 28010 -730 28030 -670
rect 28090 -730 28110 -670
rect 28010 -750 28110 -730
rect 28350 -670 28450 -650
rect 28350 -730 28370 -670
rect 28430 -730 28450 -670
rect 28350 -750 28450 -730
rect 28690 -670 28790 -650
rect 28690 -730 28710 -670
rect 28770 -730 28790 -670
rect 28690 -750 28790 -730
rect 29030 -670 29130 -650
rect 29030 -730 29050 -670
rect 29110 -730 29130 -670
rect 29030 -750 29130 -730
rect 29370 -670 29470 -650
rect 29370 -730 29390 -670
rect 29450 -730 29470 -670
rect 29370 -750 29470 -730
rect 29710 -670 29810 -650
rect 29710 -730 29730 -670
rect 29790 -730 29810 -670
rect 29710 -750 29810 -730
rect 30050 -670 30150 -650
rect 30050 -730 30070 -670
rect 30130 -730 30150 -670
rect 30050 -750 30150 -730
rect 30390 -670 30490 -650
rect 30390 -730 30410 -670
rect 30470 -730 30490 -670
rect 30390 -750 30490 -730
rect 30730 -670 30830 -650
rect 30730 -730 30750 -670
rect 30810 -730 30830 -670
rect 30730 -750 30830 -730
rect 31070 -670 31170 -650
rect 31070 -730 31090 -670
rect 31150 -730 31170 -670
rect 31070 -750 31170 -730
rect 31410 -670 31510 -650
rect 31410 -730 31430 -670
rect 31490 -730 31510 -670
rect 31410 -750 31510 -730
rect 31750 -670 31850 -650
rect 31750 -730 31770 -670
rect 31830 -730 31850 -670
rect 31750 -750 31850 -730
rect 32090 -670 32190 -650
rect 32090 -730 32110 -670
rect 32170 -730 32190 -670
rect 32090 -750 32190 -730
rect 32430 -670 32530 -650
rect 32430 -730 32450 -670
rect 32510 -730 32530 -670
rect 32430 -750 32530 -730
rect 32770 -670 32870 -650
rect 32770 -730 32790 -670
rect 32850 -730 32870 -670
rect 32770 -750 32870 -730
rect 33110 -670 33210 -650
rect 33110 -730 33130 -670
rect 33190 -730 33210 -670
rect 33110 -750 33210 -730
rect 33450 -670 33550 -650
rect 33450 -730 33470 -670
rect 33530 -730 33550 -670
rect 33450 -750 33550 -730
rect 33790 -670 33890 -650
rect 33790 -730 33810 -670
rect 33870 -730 33890 -670
rect 33790 -750 33890 -730
rect 34130 -670 34230 -650
rect 34130 -730 34150 -670
rect 34210 -730 34230 -670
rect 34130 -750 34230 -730
rect 34470 -670 34570 -650
rect 34470 -730 34490 -670
rect 34550 -730 34570 -670
rect 34470 -750 34570 -730
rect 34810 -670 34910 -650
rect 34810 -730 34830 -670
rect 34890 -730 34910 -670
rect 34810 -750 34910 -730
rect 35150 -670 35250 -650
rect 35150 -730 35170 -670
rect 35230 -730 35250 -670
rect 35150 -750 35250 -730
rect 35490 -670 35590 -650
rect 35490 -730 35510 -670
rect 35570 -730 35590 -670
rect 35490 -750 35590 -730
rect 35830 -670 35930 -650
rect 35830 -730 35850 -670
rect 35910 -730 35930 -670
rect 35830 -750 35930 -730
rect 36170 -670 36270 -650
rect 36170 -730 36190 -670
rect 36250 -730 36270 -670
rect 36170 -750 36270 -730
rect 36510 -670 36610 -650
rect 36510 -730 36530 -670
rect 36590 -730 36610 -670
rect 36510 -750 36610 -730
rect 36850 -670 36950 -650
rect 36850 -730 36870 -670
rect 36930 -730 36950 -670
rect 36850 -750 36950 -730
rect 37190 -670 37290 -650
rect 37190 -730 37210 -670
rect 37270 -730 37290 -670
rect 37190 -750 37290 -730
rect 37530 -670 37630 -650
rect 37530 -730 37550 -670
rect 37610 -730 37630 -670
rect 37530 -750 37630 -730
rect 37870 -670 37970 -650
rect 37870 -730 37890 -670
rect 37950 -730 37970 -670
rect 37870 -750 37970 -730
rect 38210 -670 38310 -650
rect 38210 -730 38230 -670
rect 38290 -730 38310 -670
rect 38210 -750 38310 -730
rect 38550 -670 38650 -650
rect 38550 -730 38570 -670
rect 38630 -730 38650 -670
rect 38550 -750 38650 -730
rect 38890 -670 38990 -650
rect 38890 -730 38910 -670
rect 38970 -730 38990 -670
rect 38890 -750 38990 -730
rect 39230 -670 39330 -650
rect 39230 -730 39250 -670
rect 39310 -730 39330 -670
rect 39230 -750 39330 -730
rect 39570 -670 39670 -650
rect 39570 -730 39590 -670
rect 39650 -730 39670 -670
rect 39570 -750 39670 -730
rect 39910 -670 40010 -650
rect 39910 -730 39930 -670
rect 39990 -730 40010 -670
rect 39910 -750 40010 -730
rect 40250 -670 40350 -650
rect 40250 -730 40270 -670
rect 40330 -730 40350 -670
rect 40250 -750 40350 -730
rect 40590 -670 40690 -650
rect 40590 -730 40610 -670
rect 40670 -730 40690 -670
rect 40590 -750 40690 -730
rect 40930 -670 41030 -650
rect 40930 -730 40950 -670
rect 41010 -730 41030 -670
rect 40930 -750 41030 -730
rect 41270 -670 41370 -650
rect 41270 -730 41290 -670
rect 41350 -730 41370 -670
rect 41270 -750 41370 -730
rect 41610 -670 41710 -650
rect 41610 -730 41630 -670
rect 41690 -730 41710 -670
rect 41610 -750 41710 -730
rect 41950 -670 42050 -650
rect 41950 -730 41970 -670
rect 42030 -730 42050 -670
rect 41950 -750 42050 -730
rect 42290 -670 42390 -650
rect 42290 -730 42310 -670
rect 42370 -730 42390 -670
rect 42290 -750 42390 -730
rect 42630 -670 42730 -650
rect 42630 -730 42650 -670
rect 42710 -730 42730 -670
rect 42630 -750 42730 -730
rect 42970 -670 43070 -650
rect 42970 -730 42990 -670
rect 43050 -730 43070 -670
rect 42970 -750 43070 -730
rect 43310 -670 43410 -650
rect 43310 -730 43330 -670
rect 43390 -730 43410 -670
rect 43310 -750 43410 -730
rect 43650 -670 43750 -650
rect 43650 -730 43670 -670
rect 43730 -730 43750 -670
rect 43650 -750 43750 -730
rect 43990 -670 44090 -650
rect 43990 -730 44010 -670
rect 44070 -730 44090 -670
rect 43990 -750 44090 -730
rect 44330 -670 44430 -650
rect 44330 -730 44350 -670
rect 44410 -730 44430 -670
rect 44330 -750 44430 -730
rect 44670 -670 44770 -650
rect 44670 -730 44690 -670
rect 44750 -730 44770 -670
rect 44670 -750 44770 -730
rect 45010 -670 45110 -650
rect 45010 -730 45030 -670
rect 45090 -730 45110 -670
rect 45010 -750 45110 -730
rect 45350 -670 45450 -650
rect 45350 -730 45370 -670
rect 45430 -730 45450 -670
rect 45350 -750 45450 -730
rect 45690 -670 45790 -650
rect 45690 -730 45710 -670
rect 45770 -730 45790 -670
rect 45690 -750 45790 -730
rect 46030 -670 46130 -650
rect 46030 -730 46050 -670
rect 46110 -730 46130 -670
rect 46030 -750 46130 -730
rect 46370 -670 46470 -650
rect 46370 -730 46390 -670
rect 46450 -730 46470 -670
rect 46370 -750 46470 -730
rect 46710 -670 46810 -650
rect 46710 -730 46730 -670
rect 46790 -730 46810 -670
rect 46710 -750 46810 -730
rect 47050 -670 47150 -650
rect 47050 -730 47070 -670
rect 47130 -730 47150 -670
rect 47050 -750 47150 -730
rect 47390 -670 47490 -650
rect 47390 -730 47410 -670
rect 47470 -730 47490 -670
rect 47390 -750 47490 -730
rect 47730 -670 47830 -650
rect 47730 -730 47750 -670
rect 47810 -730 47830 -670
rect 47730 -750 47830 -730
rect 48070 -670 48170 -650
rect 48070 -730 48090 -670
rect 48150 -730 48170 -670
rect 48070 -750 48170 -730
rect 48410 -670 48510 -650
rect 48410 -730 48430 -670
rect 48490 -730 48510 -670
rect 48410 -750 48510 -730
rect 48750 -670 48850 -650
rect 48750 -730 48770 -670
rect 48830 -730 48850 -670
rect 48750 -750 48850 -730
rect 49090 -670 49190 -650
rect 49090 -730 49110 -670
rect 49170 -730 49190 -670
rect 49090 -750 49190 -730
rect 49430 -670 49530 -650
rect 49430 -730 49450 -670
rect 49510 -730 49530 -670
rect 49430 -750 49530 -730
rect 49770 -670 49870 -650
rect 49770 -730 49790 -670
rect 49850 -730 49870 -670
rect 49770 -750 49870 -730
rect 50110 -670 50210 -650
rect 50110 -730 50130 -670
rect 50190 -730 50210 -670
rect 50110 -750 50210 -730
rect 50450 -670 50550 -650
rect 50450 -730 50470 -670
rect 50530 -730 50550 -670
rect 50450 -750 50550 -730
rect 50790 -670 50890 -650
rect 50790 -730 50810 -670
rect 50870 -730 50890 -670
rect 50790 -750 50890 -730
rect 51130 -670 51230 -650
rect 51130 -730 51150 -670
rect 51210 -730 51230 -670
rect 51130 -750 51230 -730
rect 51470 -670 51570 -650
rect 51470 -730 51490 -670
rect 51550 -730 51570 -670
rect 51470 -750 51570 -730
rect 51810 -670 51910 -650
rect 51810 -730 51830 -670
rect 51890 -730 51910 -670
rect 51810 -750 51910 -730
rect 52150 -670 52250 -650
rect 52150 -730 52170 -670
rect 52230 -730 52250 -670
rect 52150 -750 52250 -730
rect 52490 -670 52590 -650
rect 52490 -730 52510 -670
rect 52570 -730 52590 -670
rect 52490 -750 52590 -730
rect 52830 -670 52930 -650
rect 52830 -730 52850 -670
rect 52910 -730 52930 -670
rect 52830 -750 52930 -730
rect 53170 -670 53270 -650
rect 53170 -730 53190 -670
rect 53250 -730 53270 -670
rect 53170 -750 53270 -730
rect 53510 -670 53610 -650
rect 53510 -730 53530 -670
rect 53590 -730 53610 -670
rect 53510 -750 53610 -730
rect 53850 -670 53950 -650
rect 53850 -730 53870 -670
rect 53930 -730 53950 -670
rect 53850 -750 53950 -730
rect 54190 -670 54290 -650
rect 54190 -730 54210 -670
rect 54270 -730 54290 -670
rect 54190 -750 54290 -730
rect 54530 -670 54630 -650
rect 54530 -730 54550 -670
rect 54610 -730 54630 -670
rect 54530 -750 54630 -730
rect 54870 -670 54970 -650
rect 54870 -730 54890 -670
rect 54950 -730 54970 -670
rect 54870 -750 54970 -730
rect 55210 -670 55310 -650
rect 55210 -730 55230 -670
rect 55290 -730 55310 -670
rect 55210 -750 55310 -730
rect 55550 -670 55650 -650
rect 55550 -730 55570 -670
rect 55630 -730 55650 -670
rect 55550 -750 55650 -730
rect 55890 -670 55990 -650
rect 55890 -730 55910 -670
rect 55970 -730 55990 -670
rect 55890 -750 55990 -730
rect 56230 -670 56330 -650
rect 56230 -730 56250 -670
rect 56310 -730 56330 -670
rect 56230 -750 56330 -730
rect 56570 -670 56670 -650
rect 56570 -730 56590 -670
rect 56650 -730 56670 -670
rect 56570 -750 56670 -730
rect 56910 -670 57010 -650
rect 56910 -730 56930 -670
rect 56990 -730 57010 -670
rect 56910 -750 57010 -730
rect 57250 -670 57350 -650
rect 57250 -730 57270 -670
rect 57330 -730 57350 -670
rect 57250 -750 57350 -730
rect 57590 -670 57690 -650
rect 57590 -730 57610 -670
rect 57670 -730 57690 -670
rect 57590 -750 57690 -730
rect 57930 -670 58030 -650
rect 57930 -730 57950 -670
rect 58010 -730 58030 -670
rect 57930 -750 58030 -730
rect 58270 -670 58370 -650
rect 58270 -730 58290 -670
rect 58350 -730 58370 -670
rect 58270 -750 58370 -730
rect 58610 -670 58710 -650
rect 58610 -730 58630 -670
rect 58690 -730 58710 -670
rect 58610 -750 58710 -730
rect 58950 -670 59050 -650
rect 58950 -730 58970 -670
rect 59030 -730 59050 -670
rect 58950 -750 59050 -730
rect 59290 -670 59390 -650
rect 59290 -730 59310 -670
rect 59370 -730 59390 -670
rect 59290 -750 59390 -730
rect 59630 -670 59730 -650
rect 59630 -730 59650 -670
rect 59710 -730 59730 -670
rect 59630 -750 59730 -730
rect 59970 -670 60070 -650
rect 59970 -730 59990 -670
rect 60050 -730 60070 -670
rect 59970 -750 60070 -730
rect 60310 -670 60410 -650
rect 60310 -730 60330 -670
rect 60390 -730 60410 -670
rect 60310 -750 60410 -730
rect 60650 -670 60750 -650
rect 60650 -730 60670 -670
rect 60730 -730 60750 -670
rect 60650 -750 60750 -730
rect 60990 -670 61090 -650
rect 60990 -730 61010 -670
rect 61070 -730 61090 -670
rect 60990 -750 61090 -730
rect 61330 -670 61430 -650
rect 61330 -730 61350 -670
rect 61410 -730 61430 -670
rect 61330 -750 61430 -730
rect 61670 -670 61770 -650
rect 61670 -730 61690 -670
rect 61750 -730 61770 -670
rect 61670 -750 61770 -730
rect 62010 -670 62110 -650
rect 62010 -730 62030 -670
rect 62090 -730 62110 -670
rect 62010 -750 62110 -730
rect 62350 -670 62450 -650
rect 62350 -730 62370 -670
rect 62430 -730 62450 -670
rect 62350 -750 62450 -730
rect 62690 -670 62790 -650
rect 62690 -730 62710 -670
rect 62770 -730 62790 -670
rect 62690 -750 62790 -730
rect 63030 -670 63130 -650
rect 63030 -730 63050 -670
rect 63110 -730 63130 -670
rect 63030 -750 63130 -730
rect 63370 -670 63470 -650
rect 63370 -730 63390 -670
rect 63450 -730 63470 -670
rect 63370 -750 63470 -730
rect 63710 -670 63810 -650
rect 63710 -730 63730 -670
rect 63790 -730 63810 -670
rect 63710 -750 63810 -730
rect 64050 -670 64150 -650
rect 64050 -730 64070 -670
rect 64130 -730 64150 -670
rect 64050 -750 64150 -730
rect 64390 -670 64490 -650
rect 64390 -730 64410 -670
rect 64470 -730 64490 -670
rect 64390 -750 64490 -730
rect 64730 -670 64830 -650
rect 64730 -730 64750 -670
rect 64810 -730 64830 -670
rect 64730 -750 64830 -730
rect 65070 -670 65170 -650
rect 65070 -730 65090 -670
rect 65150 -730 65170 -670
rect 65070 -750 65170 -730
rect 65410 -670 65510 -650
rect 65410 -730 65430 -670
rect 65490 -730 65510 -670
rect 65410 -750 65510 -730
rect 65750 -670 65850 -650
rect 65750 -730 65770 -670
rect 65830 -730 65850 -670
rect 65750 -750 65850 -730
rect 66090 -670 66190 -650
rect 66090 -730 66110 -670
rect 66170 -730 66190 -670
rect 66090 -750 66190 -730
rect 66430 -670 66530 -650
rect 66430 -730 66450 -670
rect 66510 -730 66530 -670
rect 66430 -750 66530 -730
rect 66770 -670 66870 -650
rect 66770 -730 66790 -670
rect 66850 -730 66870 -670
rect 66770 -750 66870 -730
rect 67110 -670 67210 -650
rect 67110 -730 67130 -670
rect 67190 -730 67210 -670
rect 67110 -750 67210 -730
rect 67450 -670 67550 -650
rect 67450 -730 67470 -670
rect 67530 -730 67550 -670
rect 67450 -750 67550 -730
rect 67790 -670 67890 -650
rect 67790 -730 67810 -670
rect 67870 -730 67890 -670
rect 67790 -750 67890 -730
rect 68130 -670 68230 -650
rect 68130 -730 68150 -670
rect 68210 -730 68230 -670
rect 68130 -750 68230 -730
rect 68470 -670 68570 -650
rect 68470 -730 68490 -670
rect 68550 -730 68570 -670
rect 68470 -750 68570 -730
rect 68810 -670 68910 -650
rect 68810 -730 68830 -670
rect 68890 -730 68910 -670
rect 68810 -750 68910 -730
rect 69150 -670 69250 -650
rect 69150 -730 69170 -670
rect 69230 -730 69250 -670
rect 69150 -750 69250 -730
rect 69490 -670 69590 -650
rect 69490 -730 69510 -670
rect 69570 -730 69590 -670
rect 69490 -750 69590 -730
rect 69830 -670 69930 -650
rect 69830 -730 69850 -670
rect 69910 -730 69930 -670
rect 69830 -750 69930 -730
rect 70170 -670 70270 -650
rect 70170 -730 70190 -670
rect 70250 -730 70270 -670
rect 70170 -750 70270 -730
rect 70510 -670 70610 -650
rect 70510 -730 70530 -670
rect 70590 -730 70610 -670
rect 70510 -750 70610 -730
rect 70850 -670 70950 -650
rect 70850 -730 70870 -670
rect 70930 -730 70950 -670
rect 70850 -750 70950 -730
rect 71190 -670 71290 -650
rect 71190 -730 71210 -670
rect 71270 -730 71290 -670
rect 71190 -750 71290 -730
rect 71530 -670 71630 -650
rect 71530 -730 71550 -670
rect 71610 -730 71630 -670
rect 71530 -750 71630 -730
rect 71870 -670 71970 -650
rect 71870 -730 71890 -670
rect 71950 -730 71970 -670
rect 71870 -750 71970 -730
rect 72210 -670 72310 -650
rect 72210 -730 72230 -670
rect 72290 -730 72310 -670
rect 72210 -750 72310 -730
rect 72550 -670 72650 -650
rect 72550 -730 72570 -670
rect 72630 -730 72650 -670
rect 72550 -750 72650 -730
rect 72890 -670 72990 -650
rect 72890 -730 72910 -670
rect 72970 -730 72990 -670
rect 72890 -750 72990 -730
rect 73230 -670 73330 -650
rect 73230 -730 73250 -670
rect 73310 -730 73330 -670
rect 73230 -750 73330 -730
rect 73570 -670 73670 -650
rect 73570 -730 73590 -670
rect 73650 -730 73670 -670
rect 73570 -750 73670 -730
rect 73910 -670 74010 -650
rect 73910 -730 73930 -670
rect 73990 -730 74010 -670
rect 73910 -750 74010 -730
rect 74250 -670 74350 -650
rect 74250 -730 74270 -670
rect 74330 -730 74350 -670
rect 74250 -750 74350 -730
rect 74590 -670 74690 -650
rect 74590 -730 74610 -670
rect 74670 -730 74690 -670
rect 74590 -750 74690 -730
rect 74930 -670 75030 -650
rect 74930 -730 74950 -670
rect 75010 -730 75030 -670
rect 74930 -750 75030 -730
rect 75270 -670 75370 -650
rect 75270 -730 75290 -670
rect 75350 -730 75370 -670
rect 75270 -750 75370 -730
rect 75610 -670 75710 -650
rect 75610 -730 75630 -670
rect 75690 -730 75710 -670
rect 75610 -750 75710 -730
rect 75950 -670 76050 -650
rect 75950 -730 75970 -670
rect 76030 -730 76050 -670
rect 75950 -750 76050 -730
rect 76290 -670 76390 -650
rect 76290 -730 76310 -670
rect 76370 -730 76390 -670
rect 76290 -750 76390 -730
rect 76630 -670 76730 -650
rect 76630 -730 76650 -670
rect 76710 -730 76730 -670
rect 76630 -750 76730 -730
rect 76970 -670 77070 -650
rect 76970 -730 76990 -670
rect 77050 -730 77070 -670
rect 76970 -750 77070 -730
rect 77310 -670 77410 -650
rect 77310 -730 77330 -670
rect 77390 -730 77410 -670
rect 77310 -750 77410 -730
rect 77650 -670 77750 -650
rect 77650 -730 77670 -670
rect 77730 -730 77750 -670
rect 77650 -750 77750 -730
rect 77990 -670 78090 -650
rect 77990 -730 78010 -670
rect 78070 -730 78090 -670
rect 77990 -750 78090 -730
rect 78330 -670 78430 -650
rect 78330 -730 78350 -670
rect 78410 -730 78430 -670
rect 78330 -750 78430 -730
rect 78670 -670 78770 -650
rect 78670 -730 78690 -670
rect 78750 -730 78770 -670
rect 78670 -750 78770 -730
rect 79010 -670 79110 -650
rect 79010 -730 79030 -670
rect 79090 -730 79110 -670
rect 79010 -750 79110 -730
rect 79350 -670 79450 -650
rect 79350 -730 79370 -670
rect 79430 -730 79450 -670
rect 79350 -750 79450 -730
rect 79690 -670 79790 -650
rect 79690 -730 79710 -670
rect 79770 -730 79790 -670
rect 79690 -750 79790 -730
rect 80030 -670 80130 -650
rect 80030 -730 80050 -670
rect 80110 -730 80130 -670
rect 80030 -750 80130 -730
rect 80370 -670 80470 -650
rect 80370 -730 80390 -670
rect 80450 -730 80470 -670
rect 80370 -750 80470 -730
rect 80710 -670 80810 -650
rect 80710 -730 80730 -670
rect 80790 -730 80810 -670
rect 80710 -750 80810 -730
rect 81050 -670 81150 -650
rect 81050 -730 81070 -670
rect 81130 -730 81150 -670
rect 81050 -750 81150 -730
rect 81390 -670 81490 -650
rect 81390 -730 81410 -670
rect 81470 -730 81490 -670
rect 81390 -750 81490 -730
rect 81730 -670 81830 -650
rect 81730 -730 81750 -670
rect 81810 -730 81830 -670
rect 81730 -750 81830 -730
rect 82070 -670 82170 -650
rect 82070 -730 82090 -670
rect 82150 -730 82170 -670
rect 82070 -750 82170 -730
rect 82410 -670 82510 -650
rect 82410 -730 82430 -670
rect 82490 -730 82510 -670
rect 82410 -750 82510 -730
rect 82750 -670 82850 -650
rect 82750 -730 82770 -670
rect 82830 -730 82850 -670
rect 82750 -750 82850 -730
rect 83090 -670 83190 -650
rect 83090 -730 83110 -670
rect 83170 -730 83190 -670
rect 83090 -750 83190 -730
rect 83430 -670 83530 -650
rect 83430 -730 83450 -670
rect 83510 -730 83530 -670
rect 83430 -750 83530 -730
rect 83770 -670 83870 -650
rect 83770 -730 83790 -670
rect 83850 -730 83870 -670
rect 83770 -750 83870 -730
rect 84110 -670 84210 -650
rect 84110 -730 84130 -670
rect 84190 -730 84210 -670
rect 84110 -750 84210 -730
rect 84450 -670 84550 -650
rect 84450 -730 84470 -670
rect 84530 -730 84550 -670
rect 84450 -750 84550 -730
rect 84790 -670 84890 -650
rect 84790 -730 84810 -670
rect 84870 -730 84890 -670
rect 84790 -750 84890 -730
rect 85130 -670 85230 -650
rect 85130 -730 85150 -670
rect 85210 -730 85230 -670
rect 85130 -750 85230 -730
rect 85470 -670 85570 -650
rect 85470 -730 85490 -670
rect 85550 -730 85570 -670
rect 85470 -750 85570 -730
rect 85810 -670 85910 -650
rect 85810 -730 85830 -670
rect 85890 -730 85910 -670
rect 85810 -750 85910 -730
rect 86150 -670 86250 -650
rect 86150 -730 86170 -670
rect 86230 -730 86250 -670
rect 86150 -750 86250 -730
rect 86490 -670 86590 -650
rect 86490 -730 86510 -670
rect 86570 -730 86590 -670
rect 86490 -750 86590 -730
rect 86830 -670 86930 -650
rect 86830 -730 86850 -670
rect 86910 -730 86930 -670
rect 86830 -750 86930 -730
rect 87170 -670 87270 -650
rect 87170 -730 87190 -670
rect 87250 -730 87270 -670
rect 87170 -750 87270 -730
rect 300 -770 400 -750
rect 300 -830 320 -770
rect 380 -830 400 -770
rect 300 -880 400 -830
rect 300 -950 320 -880
rect 380 -950 400 -880
rect 300 -1000 400 -950
rect 300 -1060 320 -1000
rect 380 -1060 400 -1000
rect 130 -1100 230 -1080
rect 130 -1160 150 -1100
rect 210 -1160 230 -1100
rect 130 -1180 230 -1160
rect 300 -1200 400 -1060
rect 640 -770 740 -750
rect 640 -830 660 -770
rect 720 -830 740 -770
rect 640 -880 740 -830
rect 640 -950 660 -880
rect 720 -950 740 -880
rect 640 -1000 740 -950
rect 640 -1060 660 -1000
rect 720 -1060 740 -1000
rect 470 -1100 570 -1080
rect 470 -1160 490 -1100
rect 550 -1160 570 -1100
rect 470 -1180 570 -1160
rect 300 -1260 320 -1200
rect 380 -1260 400 -1200
rect 300 -1270 400 -1260
rect 640 -1200 740 -1060
rect 980 -770 1080 -750
rect 980 -830 1000 -770
rect 1060 -830 1080 -770
rect 980 -880 1080 -830
rect 980 -950 1000 -880
rect 1060 -950 1080 -880
rect 980 -1000 1080 -950
rect 980 -1060 1000 -1000
rect 1060 -1060 1080 -1000
rect 810 -1100 910 -1080
rect 810 -1160 830 -1100
rect 890 -1160 910 -1100
rect 810 -1180 910 -1160
rect 640 -1260 660 -1200
rect 720 -1260 740 -1200
rect 640 -1270 740 -1260
rect 980 -1200 1080 -1060
rect 1320 -770 1420 -750
rect 1320 -830 1340 -770
rect 1400 -830 1420 -770
rect 1320 -880 1420 -830
rect 1320 -950 1340 -880
rect 1400 -950 1420 -880
rect 1320 -1000 1420 -950
rect 1320 -1060 1340 -1000
rect 1400 -1060 1420 -1000
rect 1150 -1100 1250 -1080
rect 1150 -1160 1170 -1100
rect 1230 -1160 1250 -1100
rect 1150 -1180 1250 -1160
rect 980 -1260 1000 -1200
rect 1060 -1260 1080 -1200
rect 980 -1270 1080 -1260
rect 1320 -1200 1420 -1060
rect 1660 -770 1760 -750
rect 1660 -830 1680 -770
rect 1740 -830 1760 -770
rect 1660 -880 1760 -830
rect 1660 -950 1680 -880
rect 1740 -950 1760 -880
rect 1660 -1000 1760 -950
rect 1660 -1060 1680 -1000
rect 1740 -1060 1760 -1000
rect 1490 -1100 1590 -1080
rect 1490 -1160 1510 -1100
rect 1570 -1160 1590 -1100
rect 1490 -1180 1590 -1160
rect 1320 -1260 1340 -1200
rect 1400 -1260 1420 -1200
rect 1320 -1270 1420 -1260
rect 1660 -1200 1760 -1060
rect 2000 -770 2100 -750
rect 2000 -830 2020 -770
rect 2080 -830 2100 -770
rect 2000 -880 2100 -830
rect 2000 -950 2020 -880
rect 2080 -950 2100 -880
rect 2000 -1000 2100 -950
rect 2000 -1060 2020 -1000
rect 2080 -1060 2100 -1000
rect 1830 -1100 1930 -1080
rect 1830 -1160 1850 -1100
rect 1910 -1160 1930 -1100
rect 1830 -1180 1930 -1160
rect 1660 -1260 1680 -1200
rect 1740 -1260 1760 -1200
rect 1660 -1270 1760 -1260
rect 2000 -1200 2100 -1060
rect 2340 -770 2440 -750
rect 2340 -830 2360 -770
rect 2420 -830 2440 -770
rect 2340 -880 2440 -830
rect 2340 -950 2360 -880
rect 2420 -950 2440 -880
rect 2340 -1000 2440 -950
rect 2340 -1060 2360 -1000
rect 2420 -1060 2440 -1000
rect 2170 -1100 2270 -1080
rect 2170 -1160 2190 -1100
rect 2250 -1160 2270 -1100
rect 2170 -1180 2270 -1160
rect 2000 -1260 2020 -1200
rect 2080 -1260 2100 -1200
rect 2000 -1270 2100 -1260
rect 2340 -1200 2440 -1060
rect 2680 -770 2780 -750
rect 2680 -830 2700 -770
rect 2760 -830 2780 -770
rect 2680 -880 2780 -830
rect 2680 -950 2700 -880
rect 2760 -950 2780 -880
rect 2680 -1000 2780 -950
rect 2680 -1060 2700 -1000
rect 2760 -1060 2780 -1000
rect 2510 -1100 2610 -1080
rect 2510 -1160 2530 -1100
rect 2590 -1160 2610 -1100
rect 2510 -1180 2610 -1160
rect 2340 -1260 2360 -1200
rect 2420 -1260 2440 -1200
rect 2340 -1270 2440 -1260
rect 2680 -1200 2780 -1060
rect 3020 -770 3120 -750
rect 3020 -830 3040 -770
rect 3100 -830 3120 -770
rect 3020 -880 3120 -830
rect 3020 -950 3040 -880
rect 3100 -950 3120 -880
rect 3020 -1000 3120 -950
rect 3020 -1060 3040 -1000
rect 3100 -1060 3120 -1000
rect 2850 -1100 2950 -1080
rect 2850 -1160 2870 -1100
rect 2930 -1160 2950 -1100
rect 2850 -1180 2950 -1160
rect 2680 -1260 2700 -1200
rect 2760 -1260 2780 -1200
rect 2680 -1270 2780 -1260
rect 3020 -1200 3120 -1060
rect 3360 -770 3460 -750
rect 3360 -830 3380 -770
rect 3440 -830 3460 -770
rect 3360 -880 3460 -830
rect 3360 -950 3380 -880
rect 3440 -950 3460 -880
rect 3360 -1000 3460 -950
rect 3360 -1060 3380 -1000
rect 3440 -1060 3460 -1000
rect 3190 -1100 3290 -1080
rect 3190 -1160 3210 -1100
rect 3270 -1160 3290 -1100
rect 3190 -1180 3290 -1160
rect 3020 -1260 3040 -1200
rect 3100 -1260 3120 -1200
rect 3020 -1270 3120 -1260
rect 3360 -1200 3460 -1060
rect 3700 -770 3800 -750
rect 3700 -830 3720 -770
rect 3780 -830 3800 -770
rect 3700 -880 3800 -830
rect 3700 -950 3720 -880
rect 3780 -950 3800 -880
rect 3700 -1000 3800 -950
rect 3700 -1060 3720 -1000
rect 3780 -1060 3800 -1000
rect 3530 -1100 3630 -1080
rect 3530 -1160 3550 -1100
rect 3610 -1160 3630 -1100
rect 3530 -1180 3630 -1160
rect 3360 -1260 3380 -1200
rect 3440 -1260 3460 -1200
rect 3360 -1270 3460 -1260
rect 3700 -1200 3800 -1060
rect 4040 -770 4140 -750
rect 4040 -830 4060 -770
rect 4120 -830 4140 -770
rect 4040 -880 4140 -830
rect 4040 -950 4060 -880
rect 4120 -950 4140 -880
rect 4040 -1000 4140 -950
rect 4040 -1060 4060 -1000
rect 4120 -1060 4140 -1000
rect 3870 -1100 3970 -1080
rect 3870 -1160 3890 -1100
rect 3950 -1160 3970 -1100
rect 3870 -1180 3970 -1160
rect 3700 -1260 3720 -1200
rect 3780 -1260 3800 -1200
rect 3700 -1270 3800 -1260
rect 4040 -1200 4140 -1060
rect 4380 -770 4480 -750
rect 4380 -830 4400 -770
rect 4460 -830 4480 -770
rect 4380 -880 4480 -830
rect 4380 -950 4400 -880
rect 4460 -950 4480 -880
rect 4380 -1000 4480 -950
rect 4380 -1060 4400 -1000
rect 4460 -1060 4480 -1000
rect 4210 -1100 4310 -1080
rect 4210 -1160 4230 -1100
rect 4290 -1160 4310 -1100
rect 4210 -1180 4310 -1160
rect 4040 -1260 4060 -1200
rect 4120 -1260 4140 -1200
rect 4040 -1270 4140 -1260
rect 4380 -1200 4480 -1060
rect 4720 -770 4820 -750
rect 4720 -830 4740 -770
rect 4800 -830 4820 -770
rect 4720 -880 4820 -830
rect 4720 -950 4740 -880
rect 4800 -950 4820 -880
rect 4720 -1000 4820 -950
rect 4720 -1060 4740 -1000
rect 4800 -1060 4820 -1000
rect 4550 -1100 4650 -1080
rect 4550 -1160 4570 -1100
rect 4630 -1160 4650 -1100
rect 4550 -1180 4650 -1160
rect 4380 -1260 4400 -1200
rect 4460 -1260 4480 -1200
rect 4380 -1270 4480 -1260
rect 4720 -1200 4820 -1060
rect 5060 -770 5160 -750
rect 5060 -830 5080 -770
rect 5140 -830 5160 -770
rect 5060 -880 5160 -830
rect 5060 -950 5080 -880
rect 5140 -950 5160 -880
rect 5060 -1000 5160 -950
rect 5060 -1060 5080 -1000
rect 5140 -1060 5160 -1000
rect 4890 -1100 4990 -1080
rect 4890 -1160 4910 -1100
rect 4970 -1160 4990 -1100
rect 4890 -1180 4990 -1160
rect 4720 -1260 4740 -1200
rect 4800 -1260 4820 -1200
rect 4720 -1270 4820 -1260
rect 5060 -1200 5160 -1060
rect 5400 -770 5500 -750
rect 5400 -830 5420 -770
rect 5480 -830 5500 -770
rect 5400 -880 5500 -830
rect 5400 -950 5420 -880
rect 5480 -950 5500 -880
rect 5400 -1000 5500 -950
rect 5400 -1060 5420 -1000
rect 5480 -1060 5500 -1000
rect 5230 -1100 5330 -1080
rect 5230 -1160 5250 -1100
rect 5310 -1160 5330 -1100
rect 5230 -1180 5330 -1160
rect 5060 -1260 5080 -1200
rect 5140 -1260 5160 -1200
rect 5060 -1270 5160 -1260
rect 5400 -1200 5500 -1060
rect 5740 -770 5840 -750
rect 5740 -830 5760 -770
rect 5820 -830 5840 -770
rect 5740 -880 5840 -830
rect 5740 -950 5760 -880
rect 5820 -950 5840 -880
rect 5740 -1000 5840 -950
rect 5740 -1060 5760 -1000
rect 5820 -1060 5840 -1000
rect 5570 -1100 5670 -1080
rect 5570 -1160 5590 -1100
rect 5650 -1160 5670 -1100
rect 5570 -1180 5670 -1160
rect 5400 -1260 5420 -1200
rect 5480 -1260 5500 -1200
rect 5400 -1270 5500 -1260
rect 5740 -1200 5840 -1060
rect 6080 -770 6180 -750
rect 6080 -830 6100 -770
rect 6160 -830 6180 -770
rect 6080 -880 6180 -830
rect 6080 -950 6100 -880
rect 6160 -950 6180 -880
rect 6080 -1000 6180 -950
rect 6080 -1060 6100 -1000
rect 6160 -1060 6180 -1000
rect 5910 -1100 6010 -1080
rect 5910 -1160 5930 -1100
rect 5990 -1160 6010 -1100
rect 5910 -1180 6010 -1160
rect 5740 -1260 5760 -1200
rect 5820 -1260 5840 -1200
rect 5740 -1270 5840 -1260
rect 6080 -1200 6180 -1060
rect 6420 -770 6520 -750
rect 6420 -830 6440 -770
rect 6500 -830 6520 -770
rect 6420 -880 6520 -830
rect 6420 -950 6440 -880
rect 6500 -950 6520 -880
rect 6420 -1000 6520 -950
rect 6420 -1060 6440 -1000
rect 6500 -1060 6520 -1000
rect 6250 -1100 6350 -1080
rect 6250 -1160 6270 -1100
rect 6330 -1160 6350 -1100
rect 6250 -1180 6350 -1160
rect 6080 -1260 6100 -1200
rect 6160 -1260 6180 -1200
rect 6080 -1270 6180 -1260
rect 6420 -1200 6520 -1060
rect 6760 -770 6860 -750
rect 6760 -830 6780 -770
rect 6840 -830 6860 -770
rect 6760 -880 6860 -830
rect 6760 -950 6780 -880
rect 6840 -950 6860 -880
rect 6760 -1000 6860 -950
rect 6760 -1060 6780 -1000
rect 6840 -1060 6860 -1000
rect 6590 -1100 6690 -1080
rect 6590 -1160 6610 -1100
rect 6670 -1160 6690 -1100
rect 6590 -1180 6690 -1160
rect 6420 -1260 6440 -1200
rect 6500 -1260 6520 -1200
rect 6420 -1270 6520 -1260
rect 6760 -1200 6860 -1060
rect 7100 -770 7200 -750
rect 7100 -830 7120 -770
rect 7180 -830 7200 -770
rect 7100 -880 7200 -830
rect 7100 -950 7120 -880
rect 7180 -950 7200 -880
rect 7100 -1000 7200 -950
rect 7100 -1060 7120 -1000
rect 7180 -1060 7200 -1000
rect 6930 -1100 7030 -1080
rect 6930 -1160 6950 -1100
rect 7010 -1160 7030 -1100
rect 6930 -1180 7030 -1160
rect 6760 -1260 6780 -1200
rect 6840 -1260 6860 -1200
rect 6760 -1270 6860 -1260
rect 7100 -1200 7200 -1060
rect 7440 -770 7540 -750
rect 7440 -830 7460 -770
rect 7520 -830 7540 -770
rect 7440 -880 7540 -830
rect 7440 -950 7460 -880
rect 7520 -950 7540 -880
rect 7440 -1000 7540 -950
rect 7440 -1060 7460 -1000
rect 7520 -1060 7540 -1000
rect 7270 -1100 7370 -1080
rect 7270 -1160 7290 -1100
rect 7350 -1160 7370 -1100
rect 7270 -1180 7370 -1160
rect 7100 -1260 7120 -1200
rect 7180 -1260 7200 -1200
rect 7100 -1270 7200 -1260
rect 7440 -1200 7540 -1060
rect 7780 -770 7880 -750
rect 7780 -830 7800 -770
rect 7860 -830 7880 -770
rect 7780 -880 7880 -830
rect 7780 -950 7800 -880
rect 7860 -950 7880 -880
rect 7780 -1000 7880 -950
rect 7780 -1060 7800 -1000
rect 7860 -1060 7880 -1000
rect 7610 -1100 7710 -1080
rect 7610 -1160 7630 -1100
rect 7690 -1160 7710 -1100
rect 7610 -1180 7710 -1160
rect 7440 -1260 7460 -1200
rect 7520 -1260 7540 -1200
rect 7440 -1270 7540 -1260
rect 7780 -1200 7880 -1060
rect 8120 -770 8220 -750
rect 8120 -830 8140 -770
rect 8200 -830 8220 -770
rect 8120 -880 8220 -830
rect 8120 -950 8140 -880
rect 8200 -950 8220 -880
rect 8120 -1000 8220 -950
rect 8120 -1060 8140 -1000
rect 8200 -1060 8220 -1000
rect 7950 -1100 8050 -1080
rect 7950 -1160 7970 -1100
rect 8030 -1160 8050 -1100
rect 7950 -1180 8050 -1160
rect 7780 -1260 7800 -1200
rect 7860 -1260 7880 -1200
rect 7780 -1270 7880 -1260
rect 8120 -1200 8220 -1060
rect 8460 -770 8560 -750
rect 8460 -830 8480 -770
rect 8540 -830 8560 -770
rect 8460 -880 8560 -830
rect 8460 -950 8480 -880
rect 8540 -950 8560 -880
rect 8460 -1000 8560 -950
rect 8460 -1060 8480 -1000
rect 8540 -1060 8560 -1000
rect 8290 -1100 8390 -1080
rect 8290 -1160 8310 -1100
rect 8370 -1160 8390 -1100
rect 8290 -1180 8390 -1160
rect 8120 -1260 8140 -1200
rect 8200 -1260 8220 -1200
rect 8120 -1270 8220 -1260
rect 8460 -1200 8560 -1060
rect 8800 -770 8900 -750
rect 8800 -830 8820 -770
rect 8880 -830 8900 -770
rect 8800 -880 8900 -830
rect 8800 -950 8820 -880
rect 8880 -950 8900 -880
rect 8800 -1000 8900 -950
rect 8800 -1060 8820 -1000
rect 8880 -1060 8900 -1000
rect 8630 -1100 8730 -1080
rect 8630 -1160 8650 -1100
rect 8710 -1160 8730 -1100
rect 8630 -1180 8730 -1160
rect 8460 -1260 8480 -1200
rect 8540 -1260 8560 -1200
rect 8460 -1270 8560 -1260
rect 8800 -1200 8900 -1060
rect 9140 -770 9240 -750
rect 9140 -830 9160 -770
rect 9220 -830 9240 -770
rect 9140 -880 9240 -830
rect 9140 -950 9160 -880
rect 9220 -950 9240 -880
rect 9140 -1000 9240 -950
rect 9140 -1060 9160 -1000
rect 9220 -1060 9240 -1000
rect 8970 -1100 9070 -1080
rect 8970 -1160 8990 -1100
rect 9050 -1160 9070 -1100
rect 8970 -1180 9070 -1160
rect 8800 -1260 8820 -1200
rect 8880 -1260 8900 -1200
rect 8800 -1270 8900 -1260
rect 9140 -1200 9240 -1060
rect 9480 -770 9580 -750
rect 9480 -830 9500 -770
rect 9560 -830 9580 -770
rect 9480 -880 9580 -830
rect 9480 -950 9500 -880
rect 9560 -950 9580 -880
rect 9480 -1000 9580 -950
rect 9480 -1060 9500 -1000
rect 9560 -1060 9580 -1000
rect 9310 -1100 9410 -1080
rect 9310 -1160 9330 -1100
rect 9390 -1160 9410 -1100
rect 9310 -1180 9410 -1160
rect 9140 -1260 9160 -1200
rect 9220 -1260 9240 -1200
rect 9140 -1270 9240 -1260
rect 9480 -1200 9580 -1060
rect 9820 -770 9920 -750
rect 9820 -830 9840 -770
rect 9900 -830 9920 -770
rect 9820 -880 9920 -830
rect 9820 -950 9840 -880
rect 9900 -950 9920 -880
rect 9820 -1000 9920 -950
rect 9820 -1060 9840 -1000
rect 9900 -1060 9920 -1000
rect 9650 -1100 9750 -1080
rect 9650 -1160 9670 -1100
rect 9730 -1160 9750 -1100
rect 9650 -1180 9750 -1160
rect 9480 -1260 9500 -1200
rect 9560 -1260 9580 -1200
rect 9480 -1270 9580 -1260
rect 9820 -1200 9920 -1060
rect 10160 -770 10260 -750
rect 10160 -830 10180 -770
rect 10240 -830 10260 -770
rect 10160 -880 10260 -830
rect 10160 -950 10180 -880
rect 10240 -950 10260 -880
rect 10160 -1000 10260 -950
rect 10160 -1060 10180 -1000
rect 10240 -1060 10260 -1000
rect 9990 -1100 10090 -1080
rect 9990 -1160 10010 -1100
rect 10070 -1160 10090 -1100
rect 9990 -1180 10090 -1160
rect 9820 -1260 9840 -1200
rect 9900 -1260 9920 -1200
rect 9820 -1270 9920 -1260
rect 10160 -1200 10260 -1060
rect 10500 -770 10600 -750
rect 10500 -830 10520 -770
rect 10580 -830 10600 -770
rect 10500 -880 10600 -830
rect 10500 -950 10520 -880
rect 10580 -950 10600 -880
rect 10500 -1000 10600 -950
rect 10500 -1060 10520 -1000
rect 10580 -1060 10600 -1000
rect 10330 -1100 10430 -1080
rect 10330 -1160 10350 -1100
rect 10410 -1160 10430 -1100
rect 10330 -1180 10430 -1160
rect 10160 -1260 10180 -1200
rect 10240 -1260 10260 -1200
rect 10160 -1270 10260 -1260
rect 10500 -1200 10600 -1060
rect 10840 -770 10940 -750
rect 10840 -830 10860 -770
rect 10920 -830 10940 -770
rect 10840 -880 10940 -830
rect 10840 -950 10860 -880
rect 10920 -950 10940 -880
rect 10840 -1000 10940 -950
rect 10840 -1060 10860 -1000
rect 10920 -1060 10940 -1000
rect 10670 -1100 10770 -1080
rect 10670 -1160 10690 -1100
rect 10750 -1160 10770 -1100
rect 10670 -1180 10770 -1160
rect 10500 -1260 10520 -1200
rect 10580 -1260 10600 -1200
rect 10500 -1270 10600 -1260
rect 10840 -1200 10940 -1060
rect 11180 -770 11280 -750
rect 11180 -830 11200 -770
rect 11260 -830 11280 -770
rect 11180 -880 11280 -830
rect 11180 -950 11200 -880
rect 11260 -950 11280 -880
rect 11180 -1000 11280 -950
rect 11180 -1060 11200 -1000
rect 11260 -1060 11280 -1000
rect 11010 -1100 11110 -1080
rect 11010 -1160 11030 -1100
rect 11090 -1160 11110 -1100
rect 11010 -1180 11110 -1160
rect 10840 -1260 10860 -1200
rect 10920 -1260 10940 -1200
rect 10840 -1270 10940 -1260
rect 11180 -1200 11280 -1060
rect 11520 -770 11620 -750
rect 11520 -830 11540 -770
rect 11600 -830 11620 -770
rect 11520 -880 11620 -830
rect 11520 -950 11540 -880
rect 11600 -950 11620 -880
rect 11520 -1000 11620 -950
rect 11520 -1060 11540 -1000
rect 11600 -1060 11620 -1000
rect 11350 -1100 11450 -1080
rect 11350 -1160 11370 -1100
rect 11430 -1160 11450 -1100
rect 11350 -1180 11450 -1160
rect 11180 -1260 11200 -1200
rect 11260 -1260 11280 -1200
rect 11180 -1270 11280 -1260
rect 11520 -1200 11620 -1060
rect 11860 -770 11960 -750
rect 11860 -830 11880 -770
rect 11940 -830 11960 -770
rect 11860 -880 11960 -830
rect 11860 -950 11880 -880
rect 11940 -950 11960 -880
rect 11860 -1000 11960 -950
rect 11860 -1060 11880 -1000
rect 11940 -1060 11960 -1000
rect 11690 -1100 11790 -1080
rect 11690 -1160 11710 -1100
rect 11770 -1160 11790 -1100
rect 11690 -1180 11790 -1160
rect 11520 -1260 11540 -1200
rect 11600 -1260 11620 -1200
rect 11520 -1270 11620 -1260
rect 11860 -1200 11960 -1060
rect 12200 -770 12300 -750
rect 12200 -830 12220 -770
rect 12280 -830 12300 -770
rect 12200 -880 12300 -830
rect 12200 -950 12220 -880
rect 12280 -950 12300 -880
rect 12200 -1000 12300 -950
rect 12200 -1060 12220 -1000
rect 12280 -1060 12300 -1000
rect 12030 -1100 12130 -1080
rect 12030 -1160 12050 -1100
rect 12110 -1160 12130 -1100
rect 12030 -1180 12130 -1160
rect 11860 -1260 11880 -1200
rect 11940 -1260 11960 -1200
rect 11860 -1270 11960 -1260
rect 12200 -1200 12300 -1060
rect 12540 -770 12640 -750
rect 12540 -830 12560 -770
rect 12620 -830 12640 -770
rect 12540 -880 12640 -830
rect 12540 -950 12560 -880
rect 12620 -950 12640 -880
rect 12540 -1000 12640 -950
rect 12540 -1060 12560 -1000
rect 12620 -1060 12640 -1000
rect 12370 -1100 12470 -1080
rect 12370 -1160 12390 -1100
rect 12450 -1160 12470 -1100
rect 12370 -1180 12470 -1160
rect 12200 -1260 12220 -1200
rect 12280 -1260 12300 -1200
rect 12200 -1270 12300 -1260
rect 12540 -1200 12640 -1060
rect 12880 -770 12980 -750
rect 12880 -830 12900 -770
rect 12960 -830 12980 -770
rect 12880 -880 12980 -830
rect 12880 -950 12900 -880
rect 12960 -950 12980 -880
rect 12880 -1000 12980 -950
rect 12880 -1060 12900 -1000
rect 12960 -1060 12980 -1000
rect 12710 -1100 12810 -1080
rect 12710 -1160 12730 -1100
rect 12790 -1160 12810 -1100
rect 12710 -1180 12810 -1160
rect 12540 -1260 12560 -1200
rect 12620 -1260 12640 -1200
rect 12540 -1270 12640 -1260
rect 12880 -1200 12980 -1060
rect 13220 -770 13320 -750
rect 13220 -830 13240 -770
rect 13300 -830 13320 -770
rect 13220 -880 13320 -830
rect 13220 -950 13240 -880
rect 13300 -950 13320 -880
rect 13220 -1000 13320 -950
rect 13220 -1060 13240 -1000
rect 13300 -1060 13320 -1000
rect 13050 -1100 13150 -1080
rect 13050 -1160 13070 -1100
rect 13130 -1160 13150 -1100
rect 13050 -1180 13150 -1160
rect 12880 -1260 12900 -1200
rect 12960 -1260 12980 -1200
rect 12880 -1270 12980 -1260
rect 13220 -1200 13320 -1060
rect 13560 -770 13660 -750
rect 13560 -830 13580 -770
rect 13640 -830 13660 -770
rect 13560 -880 13660 -830
rect 13560 -950 13580 -880
rect 13640 -950 13660 -880
rect 13560 -1000 13660 -950
rect 13560 -1060 13580 -1000
rect 13640 -1060 13660 -1000
rect 13390 -1100 13490 -1080
rect 13390 -1160 13410 -1100
rect 13470 -1160 13490 -1100
rect 13390 -1180 13490 -1160
rect 13220 -1260 13240 -1200
rect 13300 -1260 13320 -1200
rect 13220 -1270 13320 -1260
rect 13560 -1200 13660 -1060
rect 13900 -770 14000 -750
rect 13900 -830 13920 -770
rect 13980 -830 14000 -770
rect 13900 -880 14000 -830
rect 13900 -950 13920 -880
rect 13980 -950 14000 -880
rect 13900 -1000 14000 -950
rect 13900 -1060 13920 -1000
rect 13980 -1060 14000 -1000
rect 13730 -1100 13830 -1080
rect 13730 -1160 13750 -1100
rect 13810 -1160 13830 -1100
rect 13730 -1180 13830 -1160
rect 13560 -1260 13580 -1200
rect 13640 -1260 13660 -1200
rect 13560 -1270 13660 -1260
rect 13900 -1200 14000 -1060
rect 14240 -770 14340 -750
rect 14240 -830 14260 -770
rect 14320 -830 14340 -770
rect 14240 -880 14340 -830
rect 14240 -950 14260 -880
rect 14320 -950 14340 -880
rect 14240 -1000 14340 -950
rect 14240 -1060 14260 -1000
rect 14320 -1060 14340 -1000
rect 14070 -1100 14170 -1080
rect 14070 -1160 14090 -1100
rect 14150 -1160 14170 -1100
rect 14070 -1180 14170 -1160
rect 13900 -1260 13920 -1200
rect 13980 -1260 14000 -1200
rect 13900 -1270 14000 -1260
rect 14240 -1200 14340 -1060
rect 14580 -770 14680 -750
rect 14580 -830 14600 -770
rect 14660 -830 14680 -770
rect 14580 -880 14680 -830
rect 14580 -950 14600 -880
rect 14660 -950 14680 -880
rect 14580 -1000 14680 -950
rect 14580 -1060 14600 -1000
rect 14660 -1060 14680 -1000
rect 14410 -1100 14510 -1080
rect 14410 -1160 14430 -1100
rect 14490 -1160 14510 -1100
rect 14410 -1180 14510 -1160
rect 14240 -1260 14260 -1200
rect 14320 -1260 14340 -1200
rect 14240 -1270 14340 -1260
rect 14580 -1200 14680 -1060
rect 14920 -770 15020 -750
rect 14920 -830 14940 -770
rect 15000 -830 15020 -770
rect 14920 -880 15020 -830
rect 14920 -950 14940 -880
rect 15000 -950 15020 -880
rect 14920 -1000 15020 -950
rect 14920 -1060 14940 -1000
rect 15000 -1060 15020 -1000
rect 14750 -1100 14850 -1080
rect 14750 -1160 14770 -1100
rect 14830 -1160 14850 -1100
rect 14750 -1180 14850 -1160
rect 14580 -1260 14600 -1200
rect 14660 -1260 14680 -1200
rect 14580 -1270 14680 -1260
rect 14920 -1200 15020 -1060
rect 15260 -770 15360 -750
rect 15260 -830 15280 -770
rect 15340 -830 15360 -770
rect 15260 -880 15360 -830
rect 15260 -950 15280 -880
rect 15340 -950 15360 -880
rect 15260 -1000 15360 -950
rect 15260 -1060 15280 -1000
rect 15340 -1060 15360 -1000
rect 15090 -1100 15190 -1080
rect 15090 -1160 15110 -1100
rect 15170 -1160 15190 -1100
rect 15090 -1180 15190 -1160
rect 14920 -1260 14940 -1200
rect 15000 -1260 15020 -1200
rect 14920 -1270 15020 -1260
rect 15260 -1200 15360 -1060
rect 15600 -770 15700 -750
rect 15600 -830 15620 -770
rect 15680 -830 15700 -770
rect 15600 -880 15700 -830
rect 15600 -950 15620 -880
rect 15680 -950 15700 -880
rect 15600 -1000 15700 -950
rect 15600 -1060 15620 -1000
rect 15680 -1060 15700 -1000
rect 15430 -1100 15530 -1080
rect 15430 -1160 15450 -1100
rect 15510 -1160 15530 -1100
rect 15430 -1180 15530 -1160
rect 15260 -1260 15280 -1200
rect 15340 -1260 15360 -1200
rect 15260 -1270 15360 -1260
rect 15600 -1200 15700 -1060
rect 15940 -770 16040 -750
rect 15940 -830 15960 -770
rect 16020 -830 16040 -770
rect 15940 -880 16040 -830
rect 15940 -950 15960 -880
rect 16020 -950 16040 -880
rect 15940 -1000 16040 -950
rect 15940 -1060 15960 -1000
rect 16020 -1060 16040 -1000
rect 15770 -1100 15870 -1080
rect 15770 -1160 15790 -1100
rect 15850 -1160 15870 -1100
rect 15770 -1180 15870 -1160
rect 15600 -1260 15620 -1200
rect 15680 -1260 15700 -1200
rect 15600 -1270 15700 -1260
rect 15940 -1200 16040 -1060
rect 16280 -770 16380 -750
rect 16280 -830 16300 -770
rect 16360 -830 16380 -770
rect 16280 -880 16380 -830
rect 16280 -950 16300 -880
rect 16360 -950 16380 -880
rect 16280 -1000 16380 -950
rect 16280 -1060 16300 -1000
rect 16360 -1060 16380 -1000
rect 16110 -1100 16210 -1080
rect 16110 -1160 16130 -1100
rect 16190 -1160 16210 -1100
rect 16110 -1180 16210 -1160
rect 15940 -1260 15960 -1200
rect 16020 -1260 16040 -1200
rect 15940 -1270 16040 -1260
rect 16280 -1200 16380 -1060
rect 16620 -770 16720 -750
rect 16620 -830 16640 -770
rect 16700 -830 16720 -770
rect 16620 -880 16720 -830
rect 16620 -950 16640 -880
rect 16700 -950 16720 -880
rect 16620 -1000 16720 -950
rect 16620 -1060 16640 -1000
rect 16700 -1060 16720 -1000
rect 16450 -1100 16550 -1080
rect 16450 -1160 16470 -1100
rect 16530 -1160 16550 -1100
rect 16450 -1180 16550 -1160
rect 16280 -1260 16300 -1200
rect 16360 -1260 16380 -1200
rect 16280 -1270 16380 -1260
rect 16620 -1200 16720 -1060
rect 16960 -770 17060 -750
rect 16960 -830 16980 -770
rect 17040 -830 17060 -770
rect 16960 -880 17060 -830
rect 16960 -950 16980 -880
rect 17040 -950 17060 -880
rect 16960 -1000 17060 -950
rect 16960 -1060 16980 -1000
rect 17040 -1060 17060 -1000
rect 16790 -1100 16890 -1080
rect 16790 -1160 16810 -1100
rect 16870 -1160 16890 -1100
rect 16790 -1180 16890 -1160
rect 16620 -1260 16640 -1200
rect 16700 -1260 16720 -1200
rect 16620 -1270 16720 -1260
rect 16960 -1200 17060 -1060
rect 17300 -770 17400 -750
rect 17300 -830 17320 -770
rect 17380 -830 17400 -770
rect 17300 -880 17400 -830
rect 17300 -950 17320 -880
rect 17380 -950 17400 -880
rect 17300 -1000 17400 -950
rect 17300 -1060 17320 -1000
rect 17380 -1060 17400 -1000
rect 17130 -1100 17230 -1080
rect 17130 -1160 17150 -1100
rect 17210 -1160 17230 -1100
rect 17130 -1180 17230 -1160
rect 16960 -1260 16980 -1200
rect 17040 -1260 17060 -1200
rect 16960 -1270 17060 -1260
rect 17300 -1200 17400 -1060
rect 17640 -770 17740 -750
rect 17640 -830 17660 -770
rect 17720 -830 17740 -770
rect 17640 -880 17740 -830
rect 17640 -950 17660 -880
rect 17720 -950 17740 -880
rect 17640 -1000 17740 -950
rect 17640 -1060 17660 -1000
rect 17720 -1060 17740 -1000
rect 17470 -1100 17570 -1080
rect 17470 -1160 17490 -1100
rect 17550 -1160 17570 -1100
rect 17470 -1180 17570 -1160
rect 17300 -1260 17320 -1200
rect 17380 -1260 17400 -1200
rect 17300 -1270 17400 -1260
rect 17640 -1200 17740 -1060
rect 17980 -770 18080 -750
rect 17980 -830 18000 -770
rect 18060 -830 18080 -770
rect 17980 -880 18080 -830
rect 17980 -950 18000 -880
rect 18060 -950 18080 -880
rect 17980 -1000 18080 -950
rect 17980 -1060 18000 -1000
rect 18060 -1060 18080 -1000
rect 17810 -1100 17910 -1080
rect 17810 -1160 17830 -1100
rect 17890 -1160 17910 -1100
rect 17810 -1180 17910 -1160
rect 17640 -1260 17660 -1200
rect 17720 -1260 17740 -1200
rect 17640 -1270 17740 -1260
rect 17980 -1200 18080 -1060
rect 18320 -770 18420 -750
rect 18320 -830 18340 -770
rect 18400 -830 18420 -770
rect 18320 -880 18420 -830
rect 18320 -950 18340 -880
rect 18400 -950 18420 -880
rect 18320 -1000 18420 -950
rect 18320 -1060 18340 -1000
rect 18400 -1060 18420 -1000
rect 18150 -1100 18250 -1080
rect 18150 -1160 18170 -1100
rect 18230 -1160 18250 -1100
rect 18150 -1180 18250 -1160
rect 17980 -1260 18000 -1200
rect 18060 -1260 18080 -1200
rect 17980 -1270 18080 -1260
rect 18320 -1200 18420 -1060
rect 18660 -770 18760 -750
rect 18660 -830 18680 -770
rect 18740 -830 18760 -770
rect 18660 -880 18760 -830
rect 18660 -950 18680 -880
rect 18740 -950 18760 -880
rect 18660 -1000 18760 -950
rect 18660 -1060 18680 -1000
rect 18740 -1060 18760 -1000
rect 18490 -1100 18590 -1080
rect 18490 -1160 18510 -1100
rect 18570 -1160 18590 -1100
rect 18490 -1180 18590 -1160
rect 18320 -1260 18340 -1200
rect 18400 -1260 18420 -1200
rect 18320 -1270 18420 -1260
rect 18660 -1200 18760 -1060
rect 19000 -770 19100 -750
rect 19000 -830 19020 -770
rect 19080 -830 19100 -770
rect 19000 -880 19100 -830
rect 19000 -950 19020 -880
rect 19080 -950 19100 -880
rect 19000 -1000 19100 -950
rect 19000 -1060 19020 -1000
rect 19080 -1060 19100 -1000
rect 18830 -1100 18930 -1080
rect 18830 -1160 18850 -1100
rect 18910 -1160 18930 -1100
rect 18830 -1180 18930 -1160
rect 18660 -1260 18680 -1200
rect 18740 -1260 18760 -1200
rect 18660 -1270 18760 -1260
rect 19000 -1200 19100 -1060
rect 19340 -770 19440 -750
rect 19340 -830 19360 -770
rect 19420 -830 19440 -770
rect 19340 -880 19440 -830
rect 19340 -950 19360 -880
rect 19420 -950 19440 -880
rect 19340 -1000 19440 -950
rect 19340 -1060 19360 -1000
rect 19420 -1060 19440 -1000
rect 19170 -1100 19270 -1080
rect 19170 -1160 19190 -1100
rect 19250 -1160 19270 -1100
rect 19170 -1180 19270 -1160
rect 19000 -1260 19020 -1200
rect 19080 -1260 19100 -1200
rect 19000 -1270 19100 -1260
rect 19340 -1200 19440 -1060
rect 19680 -770 19780 -750
rect 19680 -830 19700 -770
rect 19760 -830 19780 -770
rect 19680 -880 19780 -830
rect 19680 -950 19700 -880
rect 19760 -950 19780 -880
rect 19680 -1000 19780 -950
rect 19680 -1060 19700 -1000
rect 19760 -1060 19780 -1000
rect 19510 -1100 19610 -1080
rect 19510 -1160 19530 -1100
rect 19590 -1160 19610 -1100
rect 19510 -1180 19610 -1160
rect 19340 -1260 19360 -1200
rect 19420 -1260 19440 -1200
rect 19340 -1270 19440 -1260
rect 19680 -1200 19780 -1060
rect 20020 -770 20120 -750
rect 20020 -830 20040 -770
rect 20100 -830 20120 -770
rect 20020 -880 20120 -830
rect 20020 -950 20040 -880
rect 20100 -950 20120 -880
rect 20020 -1000 20120 -950
rect 20020 -1060 20040 -1000
rect 20100 -1060 20120 -1000
rect 19850 -1100 19950 -1080
rect 19850 -1160 19870 -1100
rect 19930 -1160 19950 -1100
rect 19850 -1180 19950 -1160
rect 19680 -1260 19700 -1200
rect 19760 -1260 19780 -1200
rect 19680 -1270 19780 -1260
rect 20020 -1200 20120 -1060
rect 20360 -770 20460 -750
rect 20360 -830 20380 -770
rect 20440 -830 20460 -770
rect 20360 -880 20460 -830
rect 20360 -950 20380 -880
rect 20440 -950 20460 -880
rect 20360 -1000 20460 -950
rect 20360 -1060 20380 -1000
rect 20440 -1060 20460 -1000
rect 20190 -1100 20290 -1080
rect 20190 -1160 20210 -1100
rect 20270 -1160 20290 -1100
rect 20190 -1180 20290 -1160
rect 20020 -1260 20040 -1200
rect 20100 -1260 20120 -1200
rect 20020 -1270 20120 -1260
rect 20360 -1200 20460 -1060
rect 20700 -770 20800 -750
rect 20700 -830 20720 -770
rect 20780 -830 20800 -770
rect 20700 -880 20800 -830
rect 20700 -950 20720 -880
rect 20780 -950 20800 -880
rect 20700 -1000 20800 -950
rect 20700 -1060 20720 -1000
rect 20780 -1060 20800 -1000
rect 20530 -1100 20630 -1080
rect 20530 -1160 20550 -1100
rect 20610 -1160 20630 -1100
rect 20530 -1180 20630 -1160
rect 20360 -1260 20380 -1200
rect 20440 -1260 20460 -1200
rect 20360 -1270 20460 -1260
rect 20700 -1200 20800 -1060
rect 21040 -770 21140 -750
rect 21040 -830 21060 -770
rect 21120 -830 21140 -770
rect 21040 -880 21140 -830
rect 21040 -950 21060 -880
rect 21120 -950 21140 -880
rect 21040 -1000 21140 -950
rect 21040 -1060 21060 -1000
rect 21120 -1060 21140 -1000
rect 20870 -1100 20970 -1080
rect 20870 -1160 20890 -1100
rect 20950 -1160 20970 -1100
rect 20870 -1180 20970 -1160
rect 20700 -1260 20720 -1200
rect 20780 -1260 20800 -1200
rect 20700 -1270 20800 -1260
rect 21040 -1200 21140 -1060
rect 21380 -770 21480 -750
rect 21380 -830 21400 -770
rect 21460 -830 21480 -770
rect 21380 -880 21480 -830
rect 21380 -950 21400 -880
rect 21460 -950 21480 -880
rect 21380 -1000 21480 -950
rect 21380 -1060 21400 -1000
rect 21460 -1060 21480 -1000
rect 21210 -1100 21310 -1080
rect 21210 -1160 21230 -1100
rect 21290 -1160 21310 -1100
rect 21210 -1180 21310 -1160
rect 21040 -1260 21060 -1200
rect 21120 -1260 21140 -1200
rect 21040 -1270 21140 -1260
rect 21380 -1200 21480 -1060
rect 21720 -770 21820 -750
rect 21720 -830 21740 -770
rect 21800 -830 21820 -770
rect 21720 -880 21820 -830
rect 21720 -950 21740 -880
rect 21800 -950 21820 -880
rect 21720 -1000 21820 -950
rect 21720 -1060 21740 -1000
rect 21800 -1060 21820 -1000
rect 21550 -1100 21650 -1080
rect 21550 -1160 21570 -1100
rect 21630 -1160 21650 -1100
rect 21550 -1180 21650 -1160
rect 21380 -1260 21400 -1200
rect 21460 -1260 21480 -1200
rect 21380 -1270 21480 -1260
rect 21720 -1200 21820 -1060
rect 22060 -770 22160 -750
rect 22060 -830 22080 -770
rect 22140 -830 22160 -770
rect 22060 -880 22160 -830
rect 22060 -950 22080 -880
rect 22140 -950 22160 -880
rect 22060 -1000 22160 -950
rect 22060 -1060 22080 -1000
rect 22140 -1060 22160 -1000
rect 21890 -1100 21990 -1080
rect 21890 -1160 21910 -1100
rect 21970 -1160 21990 -1100
rect 21890 -1180 21990 -1160
rect 21720 -1260 21740 -1200
rect 21800 -1260 21820 -1200
rect 21720 -1270 21820 -1260
rect 22060 -1200 22160 -1060
rect 22400 -770 22500 -750
rect 22400 -830 22420 -770
rect 22480 -830 22500 -770
rect 22400 -880 22500 -830
rect 22400 -950 22420 -880
rect 22480 -950 22500 -880
rect 22400 -1000 22500 -950
rect 22400 -1060 22420 -1000
rect 22480 -1060 22500 -1000
rect 22230 -1100 22330 -1080
rect 22230 -1160 22250 -1100
rect 22310 -1160 22330 -1100
rect 22230 -1180 22330 -1160
rect 22060 -1260 22080 -1200
rect 22140 -1260 22160 -1200
rect 22060 -1270 22160 -1260
rect 22400 -1200 22500 -1060
rect 22740 -770 22840 -750
rect 22740 -830 22760 -770
rect 22820 -830 22840 -770
rect 22740 -880 22840 -830
rect 22740 -950 22760 -880
rect 22820 -950 22840 -880
rect 22740 -1000 22840 -950
rect 22740 -1060 22760 -1000
rect 22820 -1060 22840 -1000
rect 22570 -1100 22670 -1080
rect 22570 -1160 22590 -1100
rect 22650 -1160 22670 -1100
rect 22570 -1180 22670 -1160
rect 22400 -1260 22420 -1200
rect 22480 -1260 22500 -1200
rect 22400 -1270 22500 -1260
rect 22740 -1200 22840 -1060
rect 23080 -770 23180 -750
rect 23080 -830 23100 -770
rect 23160 -830 23180 -770
rect 23080 -880 23180 -830
rect 23080 -950 23100 -880
rect 23160 -950 23180 -880
rect 23080 -1000 23180 -950
rect 23080 -1060 23100 -1000
rect 23160 -1060 23180 -1000
rect 22910 -1100 23010 -1080
rect 22910 -1160 22930 -1100
rect 22990 -1160 23010 -1100
rect 22910 -1180 23010 -1160
rect 22740 -1260 22760 -1200
rect 22820 -1260 22840 -1200
rect 22740 -1270 22840 -1260
rect 23080 -1200 23180 -1060
rect 23420 -770 23520 -750
rect 23420 -830 23440 -770
rect 23500 -830 23520 -770
rect 23420 -880 23520 -830
rect 23420 -950 23440 -880
rect 23500 -950 23520 -880
rect 23420 -1000 23520 -950
rect 23420 -1060 23440 -1000
rect 23500 -1060 23520 -1000
rect 23250 -1100 23350 -1080
rect 23250 -1160 23270 -1100
rect 23330 -1160 23350 -1100
rect 23250 -1180 23350 -1160
rect 23080 -1260 23100 -1200
rect 23160 -1260 23180 -1200
rect 23080 -1270 23180 -1260
rect 23420 -1200 23520 -1060
rect 23760 -770 23860 -750
rect 23760 -830 23780 -770
rect 23840 -830 23860 -770
rect 23760 -880 23860 -830
rect 23760 -950 23780 -880
rect 23840 -950 23860 -880
rect 23760 -1000 23860 -950
rect 23760 -1060 23780 -1000
rect 23840 -1060 23860 -1000
rect 23590 -1100 23690 -1080
rect 23590 -1160 23610 -1100
rect 23670 -1160 23690 -1100
rect 23590 -1180 23690 -1160
rect 23420 -1260 23440 -1200
rect 23500 -1260 23520 -1200
rect 23420 -1270 23520 -1260
rect 23760 -1200 23860 -1060
rect 24100 -770 24200 -750
rect 24100 -830 24120 -770
rect 24180 -830 24200 -770
rect 24100 -880 24200 -830
rect 24100 -950 24120 -880
rect 24180 -950 24200 -880
rect 24100 -1000 24200 -950
rect 24100 -1060 24120 -1000
rect 24180 -1060 24200 -1000
rect 23930 -1100 24030 -1080
rect 23930 -1160 23950 -1100
rect 24010 -1160 24030 -1100
rect 23930 -1180 24030 -1160
rect 23760 -1260 23780 -1200
rect 23840 -1260 23860 -1200
rect 23760 -1270 23860 -1260
rect 24100 -1200 24200 -1060
rect 24440 -770 24540 -750
rect 24440 -830 24460 -770
rect 24520 -830 24540 -770
rect 24440 -880 24540 -830
rect 24440 -950 24460 -880
rect 24520 -950 24540 -880
rect 24440 -1000 24540 -950
rect 24440 -1060 24460 -1000
rect 24520 -1060 24540 -1000
rect 24270 -1100 24370 -1080
rect 24270 -1160 24290 -1100
rect 24350 -1160 24370 -1100
rect 24270 -1180 24370 -1160
rect 24100 -1260 24120 -1200
rect 24180 -1260 24200 -1200
rect 24100 -1270 24200 -1260
rect 24440 -1200 24540 -1060
rect 24780 -770 24880 -750
rect 24780 -830 24800 -770
rect 24860 -830 24880 -770
rect 24780 -880 24880 -830
rect 24780 -950 24800 -880
rect 24860 -950 24880 -880
rect 24780 -1000 24880 -950
rect 24780 -1060 24800 -1000
rect 24860 -1060 24880 -1000
rect 24610 -1100 24710 -1080
rect 24610 -1160 24630 -1100
rect 24690 -1160 24710 -1100
rect 24610 -1180 24710 -1160
rect 24440 -1260 24460 -1200
rect 24520 -1260 24540 -1200
rect 24440 -1270 24540 -1260
rect 24780 -1200 24880 -1060
rect 25120 -770 25220 -750
rect 25120 -830 25140 -770
rect 25200 -830 25220 -770
rect 25120 -880 25220 -830
rect 25120 -950 25140 -880
rect 25200 -950 25220 -880
rect 25120 -1000 25220 -950
rect 25120 -1060 25140 -1000
rect 25200 -1060 25220 -1000
rect 24950 -1100 25050 -1080
rect 24950 -1160 24970 -1100
rect 25030 -1160 25050 -1100
rect 24950 -1180 25050 -1160
rect 24780 -1260 24800 -1200
rect 24860 -1260 24880 -1200
rect 24780 -1270 24880 -1260
rect 25120 -1200 25220 -1060
rect 25460 -770 25560 -750
rect 25460 -830 25480 -770
rect 25540 -830 25560 -770
rect 25460 -880 25560 -830
rect 25460 -950 25480 -880
rect 25540 -950 25560 -880
rect 25460 -1000 25560 -950
rect 25460 -1060 25480 -1000
rect 25540 -1060 25560 -1000
rect 25290 -1100 25390 -1080
rect 25290 -1160 25310 -1100
rect 25370 -1160 25390 -1100
rect 25290 -1180 25390 -1160
rect 25120 -1260 25140 -1200
rect 25200 -1260 25220 -1200
rect 25120 -1270 25220 -1260
rect 25460 -1200 25560 -1060
rect 25800 -770 25900 -750
rect 25800 -830 25820 -770
rect 25880 -830 25900 -770
rect 25800 -880 25900 -830
rect 25800 -950 25820 -880
rect 25880 -950 25900 -880
rect 25800 -1000 25900 -950
rect 25800 -1060 25820 -1000
rect 25880 -1060 25900 -1000
rect 25630 -1100 25730 -1080
rect 25630 -1160 25650 -1100
rect 25710 -1160 25730 -1100
rect 25630 -1180 25730 -1160
rect 25460 -1260 25480 -1200
rect 25540 -1260 25560 -1200
rect 25460 -1270 25560 -1260
rect 25800 -1200 25900 -1060
rect 26140 -770 26240 -750
rect 26140 -830 26160 -770
rect 26220 -830 26240 -770
rect 26140 -880 26240 -830
rect 26140 -950 26160 -880
rect 26220 -950 26240 -880
rect 26140 -1000 26240 -950
rect 26140 -1060 26160 -1000
rect 26220 -1060 26240 -1000
rect 25970 -1100 26070 -1080
rect 25970 -1160 25990 -1100
rect 26050 -1160 26070 -1100
rect 25970 -1180 26070 -1160
rect 25800 -1260 25820 -1200
rect 25880 -1260 25900 -1200
rect 25800 -1270 25900 -1260
rect 26140 -1200 26240 -1060
rect 26480 -770 26580 -750
rect 26480 -830 26500 -770
rect 26560 -830 26580 -770
rect 26480 -880 26580 -830
rect 26480 -950 26500 -880
rect 26560 -950 26580 -880
rect 26480 -1000 26580 -950
rect 26480 -1060 26500 -1000
rect 26560 -1060 26580 -1000
rect 26310 -1100 26410 -1080
rect 26310 -1160 26330 -1100
rect 26390 -1160 26410 -1100
rect 26310 -1180 26410 -1160
rect 26140 -1260 26160 -1200
rect 26220 -1260 26240 -1200
rect 26140 -1270 26240 -1260
rect 26480 -1200 26580 -1060
rect 26820 -770 26920 -750
rect 26820 -830 26840 -770
rect 26900 -830 26920 -770
rect 26820 -880 26920 -830
rect 26820 -950 26840 -880
rect 26900 -950 26920 -880
rect 26820 -1000 26920 -950
rect 26820 -1060 26840 -1000
rect 26900 -1060 26920 -1000
rect 26650 -1100 26750 -1080
rect 26650 -1160 26670 -1100
rect 26730 -1160 26750 -1100
rect 26650 -1180 26750 -1160
rect 26480 -1260 26500 -1200
rect 26560 -1260 26580 -1200
rect 26480 -1270 26580 -1260
rect 26820 -1200 26920 -1060
rect 27160 -770 27260 -750
rect 27160 -830 27180 -770
rect 27240 -830 27260 -770
rect 27160 -880 27260 -830
rect 27160 -950 27180 -880
rect 27240 -950 27260 -880
rect 27160 -1000 27260 -950
rect 27160 -1060 27180 -1000
rect 27240 -1060 27260 -1000
rect 26990 -1100 27090 -1080
rect 26990 -1160 27010 -1100
rect 27070 -1160 27090 -1100
rect 26990 -1180 27090 -1160
rect 26820 -1260 26840 -1200
rect 26900 -1260 26920 -1200
rect 26820 -1270 26920 -1260
rect 27160 -1200 27260 -1060
rect 27500 -770 27600 -750
rect 27500 -830 27520 -770
rect 27580 -830 27600 -770
rect 27500 -880 27600 -830
rect 27500 -950 27520 -880
rect 27580 -950 27600 -880
rect 27500 -1000 27600 -950
rect 27500 -1060 27520 -1000
rect 27580 -1060 27600 -1000
rect 27330 -1100 27430 -1080
rect 27330 -1160 27350 -1100
rect 27410 -1160 27430 -1100
rect 27330 -1180 27430 -1160
rect 27160 -1260 27180 -1200
rect 27240 -1260 27260 -1200
rect 27160 -1270 27260 -1260
rect 27500 -1200 27600 -1060
rect 27840 -770 27940 -750
rect 27840 -830 27860 -770
rect 27920 -830 27940 -770
rect 27840 -880 27940 -830
rect 27840 -950 27860 -880
rect 27920 -950 27940 -880
rect 27840 -1000 27940 -950
rect 27840 -1060 27860 -1000
rect 27920 -1060 27940 -1000
rect 27670 -1100 27770 -1080
rect 27670 -1160 27690 -1100
rect 27750 -1160 27770 -1100
rect 27670 -1180 27770 -1160
rect 27500 -1260 27520 -1200
rect 27580 -1260 27600 -1200
rect 27500 -1270 27600 -1260
rect 27840 -1200 27940 -1060
rect 28180 -770 28280 -750
rect 28180 -830 28200 -770
rect 28260 -830 28280 -770
rect 28180 -880 28280 -830
rect 28180 -950 28200 -880
rect 28260 -950 28280 -880
rect 28180 -1000 28280 -950
rect 28180 -1060 28200 -1000
rect 28260 -1060 28280 -1000
rect 28010 -1100 28110 -1080
rect 28010 -1160 28030 -1100
rect 28090 -1160 28110 -1100
rect 28010 -1180 28110 -1160
rect 27840 -1260 27860 -1200
rect 27920 -1260 27940 -1200
rect 27840 -1270 27940 -1260
rect 28180 -1200 28280 -1060
rect 28520 -770 28620 -750
rect 28520 -830 28540 -770
rect 28600 -830 28620 -770
rect 28520 -880 28620 -830
rect 28520 -950 28540 -880
rect 28600 -950 28620 -880
rect 28520 -1000 28620 -950
rect 28520 -1060 28540 -1000
rect 28600 -1060 28620 -1000
rect 28350 -1100 28450 -1080
rect 28350 -1160 28370 -1100
rect 28430 -1160 28450 -1100
rect 28350 -1180 28450 -1160
rect 28180 -1260 28200 -1200
rect 28260 -1260 28280 -1200
rect 28180 -1270 28280 -1260
rect 28520 -1200 28620 -1060
rect 28860 -770 28960 -750
rect 28860 -830 28880 -770
rect 28940 -830 28960 -770
rect 28860 -880 28960 -830
rect 28860 -950 28880 -880
rect 28940 -950 28960 -880
rect 28860 -1000 28960 -950
rect 28860 -1060 28880 -1000
rect 28940 -1060 28960 -1000
rect 28690 -1100 28790 -1080
rect 28690 -1160 28710 -1100
rect 28770 -1160 28790 -1100
rect 28690 -1180 28790 -1160
rect 28520 -1260 28540 -1200
rect 28600 -1260 28620 -1200
rect 28520 -1270 28620 -1260
rect 28860 -1200 28960 -1060
rect 29200 -770 29300 -750
rect 29200 -830 29220 -770
rect 29280 -830 29300 -770
rect 29200 -880 29300 -830
rect 29200 -950 29220 -880
rect 29280 -950 29300 -880
rect 29200 -1000 29300 -950
rect 29200 -1060 29220 -1000
rect 29280 -1060 29300 -1000
rect 29030 -1100 29130 -1080
rect 29030 -1160 29050 -1100
rect 29110 -1160 29130 -1100
rect 29030 -1180 29130 -1160
rect 28860 -1260 28880 -1200
rect 28940 -1260 28960 -1200
rect 28860 -1270 28960 -1260
rect 29200 -1200 29300 -1060
rect 29540 -770 29640 -750
rect 29540 -830 29560 -770
rect 29620 -830 29640 -770
rect 29540 -880 29640 -830
rect 29540 -950 29560 -880
rect 29620 -950 29640 -880
rect 29540 -1000 29640 -950
rect 29540 -1060 29560 -1000
rect 29620 -1060 29640 -1000
rect 29370 -1100 29470 -1080
rect 29370 -1160 29390 -1100
rect 29450 -1160 29470 -1100
rect 29370 -1180 29470 -1160
rect 29200 -1260 29220 -1200
rect 29280 -1260 29300 -1200
rect 29200 -1270 29300 -1260
rect 29540 -1200 29640 -1060
rect 29880 -770 29980 -750
rect 29880 -830 29900 -770
rect 29960 -830 29980 -770
rect 29880 -880 29980 -830
rect 29880 -950 29900 -880
rect 29960 -950 29980 -880
rect 29880 -1000 29980 -950
rect 29880 -1060 29900 -1000
rect 29960 -1060 29980 -1000
rect 29710 -1100 29810 -1080
rect 29710 -1160 29730 -1100
rect 29790 -1160 29810 -1100
rect 29710 -1180 29810 -1160
rect 29540 -1260 29560 -1200
rect 29620 -1260 29640 -1200
rect 29540 -1270 29640 -1260
rect 29880 -1200 29980 -1060
rect 30220 -770 30320 -750
rect 30220 -830 30240 -770
rect 30300 -830 30320 -770
rect 30220 -880 30320 -830
rect 30220 -950 30240 -880
rect 30300 -950 30320 -880
rect 30220 -1000 30320 -950
rect 30220 -1060 30240 -1000
rect 30300 -1060 30320 -1000
rect 30050 -1100 30150 -1080
rect 30050 -1160 30070 -1100
rect 30130 -1160 30150 -1100
rect 30050 -1180 30150 -1160
rect 29880 -1260 29900 -1200
rect 29960 -1260 29980 -1200
rect 29880 -1270 29980 -1260
rect 30220 -1200 30320 -1060
rect 30560 -770 30660 -750
rect 30560 -830 30580 -770
rect 30640 -830 30660 -770
rect 30560 -880 30660 -830
rect 30560 -950 30580 -880
rect 30640 -950 30660 -880
rect 30560 -1000 30660 -950
rect 30560 -1060 30580 -1000
rect 30640 -1060 30660 -1000
rect 30390 -1100 30490 -1080
rect 30390 -1160 30410 -1100
rect 30470 -1160 30490 -1100
rect 30390 -1180 30490 -1160
rect 30220 -1260 30240 -1200
rect 30300 -1260 30320 -1200
rect 30220 -1270 30320 -1260
rect 30560 -1200 30660 -1060
rect 30900 -770 31000 -750
rect 30900 -830 30920 -770
rect 30980 -830 31000 -770
rect 30900 -880 31000 -830
rect 30900 -950 30920 -880
rect 30980 -950 31000 -880
rect 30900 -1000 31000 -950
rect 30900 -1060 30920 -1000
rect 30980 -1060 31000 -1000
rect 30730 -1100 30830 -1080
rect 30730 -1160 30750 -1100
rect 30810 -1160 30830 -1100
rect 30730 -1180 30830 -1160
rect 30560 -1260 30580 -1200
rect 30640 -1260 30660 -1200
rect 30560 -1270 30660 -1260
rect 30900 -1200 31000 -1060
rect 31240 -770 31340 -750
rect 31240 -830 31260 -770
rect 31320 -830 31340 -770
rect 31240 -880 31340 -830
rect 31240 -950 31260 -880
rect 31320 -950 31340 -880
rect 31240 -1000 31340 -950
rect 31240 -1060 31260 -1000
rect 31320 -1060 31340 -1000
rect 31070 -1100 31170 -1080
rect 31070 -1160 31090 -1100
rect 31150 -1160 31170 -1100
rect 31070 -1180 31170 -1160
rect 30900 -1260 30920 -1200
rect 30980 -1260 31000 -1200
rect 30900 -1270 31000 -1260
rect 31240 -1200 31340 -1060
rect 31580 -770 31680 -750
rect 31580 -830 31600 -770
rect 31660 -830 31680 -770
rect 31580 -880 31680 -830
rect 31580 -950 31600 -880
rect 31660 -950 31680 -880
rect 31580 -1000 31680 -950
rect 31580 -1060 31600 -1000
rect 31660 -1060 31680 -1000
rect 31410 -1100 31510 -1080
rect 31410 -1160 31430 -1100
rect 31490 -1160 31510 -1100
rect 31410 -1180 31510 -1160
rect 31240 -1260 31260 -1200
rect 31320 -1260 31340 -1200
rect 31240 -1270 31340 -1260
rect 31580 -1200 31680 -1060
rect 31920 -770 32020 -750
rect 31920 -830 31940 -770
rect 32000 -830 32020 -770
rect 31920 -880 32020 -830
rect 31920 -950 31940 -880
rect 32000 -950 32020 -880
rect 31920 -1000 32020 -950
rect 31920 -1060 31940 -1000
rect 32000 -1060 32020 -1000
rect 31750 -1100 31850 -1080
rect 31750 -1160 31770 -1100
rect 31830 -1160 31850 -1100
rect 31750 -1180 31850 -1160
rect 31580 -1260 31600 -1200
rect 31660 -1260 31680 -1200
rect 31580 -1270 31680 -1260
rect 31920 -1200 32020 -1060
rect 32260 -770 32360 -750
rect 32260 -830 32280 -770
rect 32340 -830 32360 -770
rect 32260 -880 32360 -830
rect 32260 -950 32280 -880
rect 32340 -950 32360 -880
rect 32260 -1000 32360 -950
rect 32260 -1060 32280 -1000
rect 32340 -1060 32360 -1000
rect 32090 -1100 32190 -1080
rect 32090 -1160 32110 -1100
rect 32170 -1160 32190 -1100
rect 32090 -1180 32190 -1160
rect 31920 -1260 31940 -1200
rect 32000 -1260 32020 -1200
rect 31920 -1270 32020 -1260
rect 32260 -1200 32360 -1060
rect 32600 -770 32700 -750
rect 32600 -830 32620 -770
rect 32680 -830 32700 -770
rect 32600 -880 32700 -830
rect 32600 -950 32620 -880
rect 32680 -950 32700 -880
rect 32600 -1000 32700 -950
rect 32600 -1060 32620 -1000
rect 32680 -1060 32700 -1000
rect 32430 -1100 32530 -1080
rect 32430 -1160 32450 -1100
rect 32510 -1160 32530 -1100
rect 32430 -1180 32530 -1160
rect 32260 -1260 32280 -1200
rect 32340 -1260 32360 -1200
rect 32260 -1270 32360 -1260
rect 32600 -1200 32700 -1060
rect 32940 -770 33040 -750
rect 32940 -830 32960 -770
rect 33020 -830 33040 -770
rect 32940 -880 33040 -830
rect 32940 -950 32960 -880
rect 33020 -950 33040 -880
rect 32940 -1000 33040 -950
rect 32940 -1060 32960 -1000
rect 33020 -1060 33040 -1000
rect 32770 -1100 32870 -1080
rect 32770 -1160 32790 -1100
rect 32850 -1160 32870 -1100
rect 32770 -1180 32870 -1160
rect 32600 -1260 32620 -1200
rect 32680 -1260 32700 -1200
rect 32600 -1270 32700 -1260
rect 32940 -1200 33040 -1060
rect 33280 -770 33380 -750
rect 33280 -830 33300 -770
rect 33360 -830 33380 -770
rect 33280 -880 33380 -830
rect 33280 -950 33300 -880
rect 33360 -950 33380 -880
rect 33280 -1000 33380 -950
rect 33280 -1060 33300 -1000
rect 33360 -1060 33380 -1000
rect 33110 -1100 33210 -1080
rect 33110 -1160 33130 -1100
rect 33190 -1160 33210 -1100
rect 33110 -1180 33210 -1160
rect 32940 -1260 32960 -1200
rect 33020 -1260 33040 -1200
rect 32940 -1270 33040 -1260
rect 33280 -1200 33380 -1060
rect 33620 -770 33720 -750
rect 33620 -830 33640 -770
rect 33700 -830 33720 -770
rect 33620 -880 33720 -830
rect 33620 -950 33640 -880
rect 33700 -950 33720 -880
rect 33620 -1000 33720 -950
rect 33620 -1060 33640 -1000
rect 33700 -1060 33720 -1000
rect 33450 -1100 33550 -1080
rect 33450 -1160 33470 -1100
rect 33530 -1160 33550 -1100
rect 33450 -1180 33550 -1160
rect 33280 -1260 33300 -1200
rect 33360 -1260 33380 -1200
rect 33280 -1270 33380 -1260
rect 33620 -1200 33720 -1060
rect 33960 -770 34060 -750
rect 33960 -830 33980 -770
rect 34040 -830 34060 -770
rect 33960 -880 34060 -830
rect 33960 -950 33980 -880
rect 34040 -950 34060 -880
rect 33960 -1000 34060 -950
rect 33960 -1060 33980 -1000
rect 34040 -1060 34060 -1000
rect 33790 -1100 33890 -1080
rect 33790 -1160 33810 -1100
rect 33870 -1160 33890 -1100
rect 33790 -1180 33890 -1160
rect 33620 -1260 33640 -1200
rect 33700 -1260 33720 -1200
rect 33620 -1270 33720 -1260
rect 33960 -1200 34060 -1060
rect 34300 -770 34400 -750
rect 34300 -830 34320 -770
rect 34380 -830 34400 -770
rect 34300 -880 34400 -830
rect 34300 -950 34320 -880
rect 34380 -950 34400 -880
rect 34300 -1000 34400 -950
rect 34300 -1060 34320 -1000
rect 34380 -1060 34400 -1000
rect 34130 -1100 34230 -1080
rect 34130 -1160 34150 -1100
rect 34210 -1160 34230 -1100
rect 34130 -1180 34230 -1160
rect 33960 -1260 33980 -1200
rect 34040 -1260 34060 -1200
rect 33960 -1270 34060 -1260
rect 34300 -1200 34400 -1060
rect 34640 -770 34740 -750
rect 34640 -830 34660 -770
rect 34720 -830 34740 -770
rect 34640 -880 34740 -830
rect 34640 -950 34660 -880
rect 34720 -950 34740 -880
rect 34640 -1000 34740 -950
rect 34640 -1060 34660 -1000
rect 34720 -1060 34740 -1000
rect 34470 -1100 34570 -1080
rect 34470 -1160 34490 -1100
rect 34550 -1160 34570 -1100
rect 34470 -1180 34570 -1160
rect 34300 -1260 34320 -1200
rect 34380 -1260 34400 -1200
rect 34300 -1270 34400 -1260
rect 34640 -1200 34740 -1060
rect 34980 -770 35080 -750
rect 34980 -830 35000 -770
rect 35060 -830 35080 -770
rect 34980 -880 35080 -830
rect 34980 -950 35000 -880
rect 35060 -950 35080 -880
rect 34980 -1000 35080 -950
rect 34980 -1060 35000 -1000
rect 35060 -1060 35080 -1000
rect 34810 -1100 34910 -1080
rect 34810 -1160 34830 -1100
rect 34890 -1160 34910 -1100
rect 34810 -1180 34910 -1160
rect 34640 -1260 34660 -1200
rect 34720 -1260 34740 -1200
rect 34640 -1270 34740 -1260
rect 34980 -1200 35080 -1060
rect 35320 -770 35420 -750
rect 35320 -830 35340 -770
rect 35400 -830 35420 -770
rect 35320 -880 35420 -830
rect 35320 -950 35340 -880
rect 35400 -950 35420 -880
rect 35320 -1000 35420 -950
rect 35320 -1060 35340 -1000
rect 35400 -1060 35420 -1000
rect 35150 -1100 35250 -1080
rect 35150 -1160 35170 -1100
rect 35230 -1160 35250 -1100
rect 35150 -1180 35250 -1160
rect 34980 -1260 35000 -1200
rect 35060 -1260 35080 -1200
rect 34980 -1270 35080 -1260
rect 35320 -1200 35420 -1060
rect 35660 -770 35760 -750
rect 35660 -830 35680 -770
rect 35740 -830 35760 -770
rect 35660 -880 35760 -830
rect 35660 -950 35680 -880
rect 35740 -950 35760 -880
rect 35660 -1000 35760 -950
rect 35660 -1060 35680 -1000
rect 35740 -1060 35760 -1000
rect 35490 -1100 35590 -1080
rect 35490 -1160 35510 -1100
rect 35570 -1160 35590 -1100
rect 35490 -1180 35590 -1160
rect 35320 -1260 35340 -1200
rect 35400 -1260 35420 -1200
rect 35320 -1270 35420 -1260
rect 35660 -1200 35760 -1060
rect 36000 -770 36100 -750
rect 36000 -830 36020 -770
rect 36080 -830 36100 -770
rect 36000 -880 36100 -830
rect 36000 -950 36020 -880
rect 36080 -950 36100 -880
rect 36000 -1000 36100 -950
rect 36000 -1060 36020 -1000
rect 36080 -1060 36100 -1000
rect 35830 -1100 35930 -1080
rect 35830 -1160 35850 -1100
rect 35910 -1160 35930 -1100
rect 35830 -1180 35930 -1160
rect 35660 -1260 35680 -1200
rect 35740 -1260 35760 -1200
rect 35660 -1270 35760 -1260
rect 36000 -1200 36100 -1060
rect 36340 -770 36440 -750
rect 36340 -830 36360 -770
rect 36420 -830 36440 -770
rect 36340 -880 36440 -830
rect 36340 -950 36360 -880
rect 36420 -950 36440 -880
rect 36340 -1000 36440 -950
rect 36340 -1060 36360 -1000
rect 36420 -1060 36440 -1000
rect 36170 -1100 36270 -1080
rect 36170 -1160 36190 -1100
rect 36250 -1160 36270 -1100
rect 36170 -1180 36270 -1160
rect 36000 -1260 36020 -1200
rect 36080 -1260 36100 -1200
rect 36000 -1270 36100 -1260
rect 36340 -1200 36440 -1060
rect 36680 -770 36780 -750
rect 36680 -830 36700 -770
rect 36760 -830 36780 -770
rect 36680 -880 36780 -830
rect 36680 -950 36700 -880
rect 36760 -950 36780 -880
rect 36680 -1000 36780 -950
rect 36680 -1060 36700 -1000
rect 36760 -1060 36780 -1000
rect 36510 -1100 36610 -1080
rect 36510 -1160 36530 -1100
rect 36590 -1160 36610 -1100
rect 36510 -1180 36610 -1160
rect 36340 -1260 36360 -1200
rect 36420 -1260 36440 -1200
rect 36340 -1270 36440 -1260
rect 36680 -1200 36780 -1060
rect 37020 -770 37120 -750
rect 37020 -830 37040 -770
rect 37100 -830 37120 -770
rect 37020 -880 37120 -830
rect 37020 -950 37040 -880
rect 37100 -950 37120 -880
rect 37020 -1000 37120 -950
rect 37020 -1060 37040 -1000
rect 37100 -1060 37120 -1000
rect 36850 -1100 36950 -1080
rect 36850 -1160 36870 -1100
rect 36930 -1160 36950 -1100
rect 36850 -1180 36950 -1160
rect 36680 -1260 36700 -1200
rect 36760 -1260 36780 -1200
rect 36680 -1270 36780 -1260
rect 37020 -1200 37120 -1060
rect 37360 -770 37460 -750
rect 37360 -830 37380 -770
rect 37440 -830 37460 -770
rect 37360 -880 37460 -830
rect 37360 -950 37380 -880
rect 37440 -950 37460 -880
rect 37360 -1000 37460 -950
rect 37360 -1060 37380 -1000
rect 37440 -1060 37460 -1000
rect 37190 -1100 37290 -1080
rect 37190 -1160 37210 -1100
rect 37270 -1160 37290 -1100
rect 37190 -1180 37290 -1160
rect 37020 -1260 37040 -1200
rect 37100 -1260 37120 -1200
rect 37020 -1270 37120 -1260
rect 37360 -1200 37460 -1060
rect 37700 -770 37800 -750
rect 37700 -830 37720 -770
rect 37780 -830 37800 -770
rect 37700 -880 37800 -830
rect 37700 -950 37720 -880
rect 37780 -950 37800 -880
rect 37700 -1000 37800 -950
rect 37700 -1060 37720 -1000
rect 37780 -1060 37800 -1000
rect 37530 -1100 37630 -1080
rect 37530 -1160 37550 -1100
rect 37610 -1160 37630 -1100
rect 37530 -1180 37630 -1160
rect 37360 -1260 37380 -1200
rect 37440 -1260 37460 -1200
rect 37360 -1270 37460 -1260
rect 37700 -1200 37800 -1060
rect 38040 -770 38140 -750
rect 38040 -830 38060 -770
rect 38120 -830 38140 -770
rect 38040 -880 38140 -830
rect 38040 -950 38060 -880
rect 38120 -950 38140 -880
rect 38040 -1000 38140 -950
rect 38040 -1060 38060 -1000
rect 38120 -1060 38140 -1000
rect 37870 -1100 37970 -1080
rect 37870 -1160 37890 -1100
rect 37950 -1160 37970 -1100
rect 37870 -1180 37970 -1160
rect 37700 -1260 37720 -1200
rect 37780 -1260 37800 -1200
rect 37700 -1270 37800 -1260
rect 38040 -1200 38140 -1060
rect 38380 -770 38480 -750
rect 38380 -830 38400 -770
rect 38460 -830 38480 -770
rect 38380 -880 38480 -830
rect 38380 -950 38400 -880
rect 38460 -950 38480 -880
rect 38380 -1000 38480 -950
rect 38380 -1060 38400 -1000
rect 38460 -1060 38480 -1000
rect 38210 -1100 38310 -1080
rect 38210 -1160 38230 -1100
rect 38290 -1160 38310 -1100
rect 38210 -1180 38310 -1160
rect 38040 -1260 38060 -1200
rect 38120 -1260 38140 -1200
rect 38040 -1270 38140 -1260
rect 38380 -1200 38480 -1060
rect 38720 -770 38820 -750
rect 38720 -830 38740 -770
rect 38800 -830 38820 -770
rect 38720 -880 38820 -830
rect 38720 -950 38740 -880
rect 38800 -950 38820 -880
rect 38720 -1000 38820 -950
rect 38720 -1060 38740 -1000
rect 38800 -1060 38820 -1000
rect 38550 -1100 38650 -1080
rect 38550 -1160 38570 -1100
rect 38630 -1160 38650 -1100
rect 38550 -1180 38650 -1160
rect 38380 -1260 38400 -1200
rect 38460 -1260 38480 -1200
rect 38380 -1270 38480 -1260
rect 38720 -1200 38820 -1060
rect 39060 -770 39160 -750
rect 39060 -830 39080 -770
rect 39140 -830 39160 -770
rect 39060 -880 39160 -830
rect 39060 -950 39080 -880
rect 39140 -950 39160 -880
rect 39060 -1000 39160 -950
rect 39060 -1060 39080 -1000
rect 39140 -1060 39160 -1000
rect 38890 -1100 38990 -1080
rect 38890 -1160 38910 -1100
rect 38970 -1160 38990 -1100
rect 38890 -1180 38990 -1160
rect 38720 -1260 38740 -1200
rect 38800 -1260 38820 -1200
rect 38720 -1270 38820 -1260
rect 39060 -1200 39160 -1060
rect 39400 -770 39500 -750
rect 39400 -830 39420 -770
rect 39480 -830 39500 -770
rect 39400 -880 39500 -830
rect 39400 -950 39420 -880
rect 39480 -950 39500 -880
rect 39400 -1000 39500 -950
rect 39400 -1060 39420 -1000
rect 39480 -1060 39500 -1000
rect 39230 -1100 39330 -1080
rect 39230 -1160 39250 -1100
rect 39310 -1160 39330 -1100
rect 39230 -1180 39330 -1160
rect 39060 -1260 39080 -1200
rect 39140 -1260 39160 -1200
rect 39060 -1270 39160 -1260
rect 39400 -1200 39500 -1060
rect 39740 -770 39840 -750
rect 39740 -830 39760 -770
rect 39820 -830 39840 -770
rect 39740 -880 39840 -830
rect 39740 -950 39760 -880
rect 39820 -950 39840 -880
rect 39740 -1000 39840 -950
rect 39740 -1060 39760 -1000
rect 39820 -1060 39840 -1000
rect 39570 -1100 39670 -1080
rect 39570 -1160 39590 -1100
rect 39650 -1160 39670 -1100
rect 39570 -1180 39670 -1160
rect 39400 -1260 39420 -1200
rect 39480 -1260 39500 -1200
rect 39400 -1270 39500 -1260
rect 39740 -1200 39840 -1060
rect 40080 -770 40180 -750
rect 40080 -830 40100 -770
rect 40160 -830 40180 -770
rect 40080 -880 40180 -830
rect 40080 -950 40100 -880
rect 40160 -950 40180 -880
rect 40080 -1000 40180 -950
rect 40080 -1060 40100 -1000
rect 40160 -1060 40180 -1000
rect 39910 -1100 40010 -1080
rect 39910 -1160 39930 -1100
rect 39990 -1160 40010 -1100
rect 39910 -1180 40010 -1160
rect 39740 -1260 39760 -1200
rect 39820 -1260 39840 -1200
rect 39740 -1270 39840 -1260
rect 40080 -1200 40180 -1060
rect 40420 -770 40520 -750
rect 40420 -830 40440 -770
rect 40500 -830 40520 -770
rect 40420 -880 40520 -830
rect 40420 -950 40440 -880
rect 40500 -950 40520 -880
rect 40420 -1000 40520 -950
rect 40420 -1060 40440 -1000
rect 40500 -1060 40520 -1000
rect 40250 -1100 40350 -1080
rect 40250 -1160 40270 -1100
rect 40330 -1160 40350 -1100
rect 40250 -1180 40350 -1160
rect 40080 -1260 40100 -1200
rect 40160 -1260 40180 -1200
rect 40080 -1270 40180 -1260
rect 40420 -1200 40520 -1060
rect 40760 -770 40860 -750
rect 40760 -830 40780 -770
rect 40840 -830 40860 -770
rect 40760 -880 40860 -830
rect 40760 -950 40780 -880
rect 40840 -950 40860 -880
rect 40760 -1000 40860 -950
rect 40760 -1060 40780 -1000
rect 40840 -1060 40860 -1000
rect 40590 -1100 40690 -1080
rect 40590 -1160 40610 -1100
rect 40670 -1160 40690 -1100
rect 40590 -1180 40690 -1160
rect 40420 -1260 40440 -1200
rect 40500 -1260 40520 -1200
rect 40420 -1270 40520 -1260
rect 40760 -1200 40860 -1060
rect 41100 -770 41200 -750
rect 41100 -830 41120 -770
rect 41180 -830 41200 -770
rect 41100 -880 41200 -830
rect 41100 -950 41120 -880
rect 41180 -950 41200 -880
rect 41100 -1000 41200 -950
rect 41100 -1060 41120 -1000
rect 41180 -1060 41200 -1000
rect 40930 -1100 41030 -1080
rect 40930 -1160 40950 -1100
rect 41010 -1160 41030 -1100
rect 40930 -1180 41030 -1160
rect 40760 -1260 40780 -1200
rect 40840 -1260 40860 -1200
rect 40760 -1270 40860 -1260
rect 41100 -1200 41200 -1060
rect 41440 -770 41540 -750
rect 41440 -830 41460 -770
rect 41520 -830 41540 -770
rect 41440 -880 41540 -830
rect 41440 -950 41460 -880
rect 41520 -950 41540 -880
rect 41440 -1000 41540 -950
rect 41440 -1060 41460 -1000
rect 41520 -1060 41540 -1000
rect 41270 -1100 41370 -1080
rect 41270 -1160 41290 -1100
rect 41350 -1160 41370 -1100
rect 41270 -1180 41370 -1160
rect 41100 -1260 41120 -1200
rect 41180 -1260 41200 -1200
rect 41100 -1270 41200 -1260
rect 41440 -1200 41540 -1060
rect 41780 -770 41880 -750
rect 41780 -830 41800 -770
rect 41860 -830 41880 -770
rect 41780 -880 41880 -830
rect 41780 -950 41800 -880
rect 41860 -950 41880 -880
rect 41780 -1000 41880 -950
rect 41780 -1060 41800 -1000
rect 41860 -1060 41880 -1000
rect 41610 -1100 41710 -1080
rect 41610 -1160 41630 -1100
rect 41690 -1160 41710 -1100
rect 41610 -1180 41710 -1160
rect 41440 -1260 41460 -1200
rect 41520 -1260 41540 -1200
rect 41440 -1270 41540 -1260
rect 41780 -1200 41880 -1060
rect 42120 -770 42220 -750
rect 42120 -830 42140 -770
rect 42200 -830 42220 -770
rect 42120 -880 42220 -830
rect 42120 -950 42140 -880
rect 42200 -950 42220 -880
rect 42120 -1000 42220 -950
rect 42120 -1060 42140 -1000
rect 42200 -1060 42220 -1000
rect 41950 -1100 42050 -1080
rect 41950 -1160 41970 -1100
rect 42030 -1160 42050 -1100
rect 41950 -1180 42050 -1160
rect 41780 -1260 41800 -1200
rect 41860 -1260 41880 -1200
rect 41780 -1270 41880 -1260
rect 42120 -1200 42220 -1060
rect 42460 -770 42560 -750
rect 42460 -830 42480 -770
rect 42540 -830 42560 -770
rect 42460 -880 42560 -830
rect 42460 -950 42480 -880
rect 42540 -950 42560 -880
rect 42460 -1000 42560 -950
rect 42460 -1060 42480 -1000
rect 42540 -1060 42560 -1000
rect 42290 -1100 42390 -1080
rect 42290 -1160 42310 -1100
rect 42370 -1160 42390 -1100
rect 42290 -1180 42390 -1160
rect 42120 -1260 42140 -1200
rect 42200 -1260 42220 -1200
rect 42120 -1270 42220 -1260
rect 42460 -1200 42560 -1060
rect 42800 -770 42900 -750
rect 42800 -830 42820 -770
rect 42880 -830 42900 -770
rect 42800 -880 42900 -830
rect 42800 -950 42820 -880
rect 42880 -950 42900 -880
rect 42800 -1000 42900 -950
rect 42800 -1060 42820 -1000
rect 42880 -1060 42900 -1000
rect 42630 -1100 42730 -1080
rect 42630 -1160 42650 -1100
rect 42710 -1160 42730 -1100
rect 42630 -1180 42730 -1160
rect 42460 -1260 42480 -1200
rect 42540 -1260 42560 -1200
rect 42460 -1270 42560 -1260
rect 42800 -1200 42900 -1060
rect 43140 -770 43240 -750
rect 43140 -830 43160 -770
rect 43220 -830 43240 -770
rect 43140 -880 43240 -830
rect 43140 -950 43160 -880
rect 43220 -950 43240 -880
rect 43140 -1000 43240 -950
rect 43140 -1060 43160 -1000
rect 43220 -1060 43240 -1000
rect 42970 -1100 43070 -1080
rect 42970 -1160 42990 -1100
rect 43050 -1160 43070 -1100
rect 42970 -1180 43070 -1160
rect 42800 -1260 42820 -1200
rect 42880 -1260 42900 -1200
rect 42800 -1270 42900 -1260
rect 43140 -1200 43240 -1060
rect 43480 -770 43580 -750
rect 43480 -830 43500 -770
rect 43560 -830 43580 -770
rect 43480 -880 43580 -830
rect 43480 -950 43500 -880
rect 43560 -950 43580 -880
rect 43480 -1000 43580 -950
rect 43480 -1060 43500 -1000
rect 43560 -1060 43580 -1000
rect 43310 -1100 43410 -1080
rect 43310 -1160 43330 -1100
rect 43390 -1160 43410 -1100
rect 43310 -1180 43410 -1160
rect 43140 -1260 43160 -1200
rect 43220 -1260 43240 -1200
rect 43140 -1270 43240 -1260
rect 43480 -1200 43580 -1060
rect 43820 -770 43920 -750
rect 43820 -830 43840 -770
rect 43900 -830 43920 -770
rect 43820 -880 43920 -830
rect 43820 -950 43840 -880
rect 43900 -950 43920 -880
rect 43820 -1000 43920 -950
rect 43820 -1060 43840 -1000
rect 43900 -1060 43920 -1000
rect 43650 -1100 43750 -1080
rect 43650 -1160 43670 -1100
rect 43730 -1160 43750 -1100
rect 43650 -1180 43750 -1160
rect 43480 -1260 43500 -1200
rect 43560 -1260 43580 -1200
rect 43480 -1270 43580 -1260
rect 43820 -1200 43920 -1060
rect 44160 -770 44260 -750
rect 44160 -830 44180 -770
rect 44240 -830 44260 -770
rect 44160 -880 44260 -830
rect 44160 -950 44180 -880
rect 44240 -950 44260 -880
rect 44160 -1000 44260 -950
rect 44160 -1060 44180 -1000
rect 44240 -1060 44260 -1000
rect 43990 -1100 44090 -1080
rect 43990 -1160 44010 -1100
rect 44070 -1160 44090 -1100
rect 43990 -1180 44090 -1160
rect 43820 -1260 43840 -1200
rect 43900 -1260 43920 -1200
rect 43820 -1270 43920 -1260
rect 44160 -1200 44260 -1060
rect 44500 -770 44600 -750
rect 44500 -830 44520 -770
rect 44580 -830 44600 -770
rect 44500 -880 44600 -830
rect 44500 -950 44520 -880
rect 44580 -950 44600 -880
rect 44500 -1000 44600 -950
rect 44500 -1060 44520 -1000
rect 44580 -1060 44600 -1000
rect 44330 -1100 44430 -1080
rect 44330 -1160 44350 -1100
rect 44410 -1160 44430 -1100
rect 44330 -1180 44430 -1160
rect 44160 -1260 44180 -1200
rect 44240 -1260 44260 -1200
rect 44160 -1270 44260 -1260
rect 44500 -1200 44600 -1060
rect 44840 -770 44940 -750
rect 44840 -830 44860 -770
rect 44920 -830 44940 -770
rect 44840 -880 44940 -830
rect 44840 -950 44860 -880
rect 44920 -950 44940 -880
rect 44840 -1000 44940 -950
rect 44840 -1060 44860 -1000
rect 44920 -1060 44940 -1000
rect 44670 -1100 44770 -1080
rect 44670 -1160 44690 -1100
rect 44750 -1160 44770 -1100
rect 44670 -1180 44770 -1160
rect 44500 -1260 44520 -1200
rect 44580 -1260 44600 -1200
rect 44500 -1270 44600 -1260
rect 44840 -1200 44940 -1060
rect 45180 -770 45280 -750
rect 45180 -830 45200 -770
rect 45260 -830 45280 -770
rect 45180 -880 45280 -830
rect 45180 -950 45200 -880
rect 45260 -950 45280 -880
rect 45180 -1000 45280 -950
rect 45180 -1060 45200 -1000
rect 45260 -1060 45280 -1000
rect 45010 -1100 45110 -1080
rect 45010 -1160 45030 -1100
rect 45090 -1160 45110 -1100
rect 45010 -1180 45110 -1160
rect 44840 -1260 44860 -1200
rect 44920 -1260 44940 -1200
rect 44840 -1270 44940 -1260
rect 45180 -1200 45280 -1060
rect 45520 -770 45620 -750
rect 45520 -830 45540 -770
rect 45600 -830 45620 -770
rect 45520 -880 45620 -830
rect 45520 -950 45540 -880
rect 45600 -950 45620 -880
rect 45520 -1000 45620 -950
rect 45520 -1060 45540 -1000
rect 45600 -1060 45620 -1000
rect 45350 -1100 45450 -1080
rect 45350 -1160 45370 -1100
rect 45430 -1160 45450 -1100
rect 45350 -1180 45450 -1160
rect 45180 -1260 45200 -1200
rect 45260 -1260 45280 -1200
rect 45180 -1270 45280 -1260
rect 45520 -1200 45620 -1060
rect 45860 -770 45960 -750
rect 45860 -830 45880 -770
rect 45940 -830 45960 -770
rect 45860 -880 45960 -830
rect 45860 -950 45880 -880
rect 45940 -950 45960 -880
rect 45860 -1000 45960 -950
rect 45860 -1060 45880 -1000
rect 45940 -1060 45960 -1000
rect 45690 -1100 45790 -1080
rect 45690 -1160 45710 -1100
rect 45770 -1160 45790 -1100
rect 45690 -1180 45790 -1160
rect 45520 -1260 45540 -1200
rect 45600 -1260 45620 -1200
rect 45520 -1270 45620 -1260
rect 45860 -1200 45960 -1060
rect 46200 -770 46300 -750
rect 46200 -830 46220 -770
rect 46280 -830 46300 -770
rect 46200 -880 46300 -830
rect 46200 -950 46220 -880
rect 46280 -950 46300 -880
rect 46200 -1000 46300 -950
rect 46200 -1060 46220 -1000
rect 46280 -1060 46300 -1000
rect 46030 -1100 46130 -1080
rect 46030 -1160 46050 -1100
rect 46110 -1160 46130 -1100
rect 46030 -1180 46130 -1160
rect 45860 -1260 45880 -1200
rect 45940 -1260 45960 -1200
rect 45860 -1270 45960 -1260
rect 46200 -1200 46300 -1060
rect 46540 -770 46640 -750
rect 46540 -830 46560 -770
rect 46620 -830 46640 -770
rect 46540 -880 46640 -830
rect 46540 -950 46560 -880
rect 46620 -950 46640 -880
rect 46540 -1000 46640 -950
rect 46540 -1060 46560 -1000
rect 46620 -1060 46640 -1000
rect 46370 -1100 46470 -1080
rect 46370 -1160 46390 -1100
rect 46450 -1160 46470 -1100
rect 46370 -1180 46470 -1160
rect 46200 -1260 46220 -1200
rect 46280 -1260 46300 -1200
rect 46200 -1270 46300 -1260
rect 46540 -1200 46640 -1060
rect 46880 -770 46980 -750
rect 46880 -830 46900 -770
rect 46960 -830 46980 -770
rect 46880 -880 46980 -830
rect 46880 -950 46900 -880
rect 46960 -950 46980 -880
rect 46880 -1000 46980 -950
rect 46880 -1060 46900 -1000
rect 46960 -1060 46980 -1000
rect 46710 -1100 46810 -1080
rect 46710 -1160 46730 -1100
rect 46790 -1160 46810 -1100
rect 46710 -1180 46810 -1160
rect 46540 -1260 46560 -1200
rect 46620 -1260 46640 -1200
rect 46540 -1270 46640 -1260
rect 46880 -1200 46980 -1060
rect 47220 -770 47320 -750
rect 47220 -830 47240 -770
rect 47300 -830 47320 -770
rect 47220 -880 47320 -830
rect 47220 -950 47240 -880
rect 47300 -950 47320 -880
rect 47220 -1000 47320 -950
rect 47220 -1060 47240 -1000
rect 47300 -1060 47320 -1000
rect 47050 -1100 47150 -1080
rect 47050 -1160 47070 -1100
rect 47130 -1160 47150 -1100
rect 47050 -1180 47150 -1160
rect 46880 -1260 46900 -1200
rect 46960 -1260 46980 -1200
rect 46880 -1270 46980 -1260
rect 47220 -1200 47320 -1060
rect 47560 -770 47660 -750
rect 47560 -830 47580 -770
rect 47640 -830 47660 -770
rect 47560 -880 47660 -830
rect 47560 -950 47580 -880
rect 47640 -950 47660 -880
rect 47560 -1000 47660 -950
rect 47560 -1060 47580 -1000
rect 47640 -1060 47660 -1000
rect 47390 -1100 47490 -1080
rect 47390 -1160 47410 -1100
rect 47470 -1160 47490 -1100
rect 47390 -1180 47490 -1160
rect 47220 -1260 47240 -1200
rect 47300 -1260 47320 -1200
rect 47220 -1270 47320 -1260
rect 47560 -1200 47660 -1060
rect 47900 -770 48000 -750
rect 47900 -830 47920 -770
rect 47980 -830 48000 -770
rect 47900 -880 48000 -830
rect 47900 -950 47920 -880
rect 47980 -950 48000 -880
rect 47900 -1000 48000 -950
rect 47900 -1060 47920 -1000
rect 47980 -1060 48000 -1000
rect 47730 -1100 47830 -1080
rect 47730 -1160 47750 -1100
rect 47810 -1160 47830 -1100
rect 47730 -1180 47830 -1160
rect 47560 -1260 47580 -1200
rect 47640 -1260 47660 -1200
rect 47560 -1270 47660 -1260
rect 47900 -1200 48000 -1060
rect 48240 -770 48340 -750
rect 48240 -830 48260 -770
rect 48320 -830 48340 -770
rect 48240 -880 48340 -830
rect 48240 -950 48260 -880
rect 48320 -950 48340 -880
rect 48240 -1000 48340 -950
rect 48240 -1060 48260 -1000
rect 48320 -1060 48340 -1000
rect 48070 -1100 48170 -1080
rect 48070 -1160 48090 -1100
rect 48150 -1160 48170 -1100
rect 48070 -1180 48170 -1160
rect 47900 -1260 47920 -1200
rect 47980 -1260 48000 -1200
rect 47900 -1270 48000 -1260
rect 48240 -1200 48340 -1060
rect 48580 -770 48680 -750
rect 48580 -830 48600 -770
rect 48660 -830 48680 -770
rect 48580 -880 48680 -830
rect 48580 -950 48600 -880
rect 48660 -950 48680 -880
rect 48580 -1000 48680 -950
rect 48580 -1060 48600 -1000
rect 48660 -1060 48680 -1000
rect 48410 -1100 48510 -1080
rect 48410 -1160 48430 -1100
rect 48490 -1160 48510 -1100
rect 48410 -1180 48510 -1160
rect 48240 -1260 48260 -1200
rect 48320 -1260 48340 -1200
rect 48240 -1270 48340 -1260
rect 48580 -1200 48680 -1060
rect 48920 -770 49020 -750
rect 48920 -830 48940 -770
rect 49000 -830 49020 -770
rect 48920 -880 49020 -830
rect 48920 -950 48940 -880
rect 49000 -950 49020 -880
rect 48920 -1000 49020 -950
rect 48920 -1060 48940 -1000
rect 49000 -1060 49020 -1000
rect 48750 -1100 48850 -1080
rect 48750 -1160 48770 -1100
rect 48830 -1160 48850 -1100
rect 48750 -1180 48850 -1160
rect 48580 -1260 48600 -1200
rect 48660 -1260 48680 -1200
rect 48580 -1270 48680 -1260
rect 48920 -1200 49020 -1060
rect 49260 -770 49360 -750
rect 49260 -830 49280 -770
rect 49340 -830 49360 -770
rect 49260 -880 49360 -830
rect 49260 -950 49280 -880
rect 49340 -950 49360 -880
rect 49260 -1000 49360 -950
rect 49260 -1060 49280 -1000
rect 49340 -1060 49360 -1000
rect 49090 -1100 49190 -1080
rect 49090 -1160 49110 -1100
rect 49170 -1160 49190 -1100
rect 49090 -1180 49190 -1160
rect 48920 -1260 48940 -1200
rect 49000 -1260 49020 -1200
rect 48920 -1270 49020 -1260
rect 49260 -1200 49360 -1060
rect 49600 -770 49700 -750
rect 49600 -830 49620 -770
rect 49680 -830 49700 -770
rect 49600 -880 49700 -830
rect 49600 -950 49620 -880
rect 49680 -950 49700 -880
rect 49600 -1000 49700 -950
rect 49600 -1060 49620 -1000
rect 49680 -1060 49700 -1000
rect 49430 -1100 49530 -1080
rect 49430 -1160 49450 -1100
rect 49510 -1160 49530 -1100
rect 49430 -1180 49530 -1160
rect 49260 -1260 49280 -1200
rect 49340 -1260 49360 -1200
rect 49260 -1270 49360 -1260
rect 49600 -1200 49700 -1060
rect 49940 -770 50040 -750
rect 49940 -830 49960 -770
rect 50020 -830 50040 -770
rect 49940 -880 50040 -830
rect 49940 -950 49960 -880
rect 50020 -950 50040 -880
rect 49940 -1000 50040 -950
rect 49940 -1060 49960 -1000
rect 50020 -1060 50040 -1000
rect 49770 -1100 49870 -1080
rect 49770 -1160 49790 -1100
rect 49850 -1160 49870 -1100
rect 49770 -1180 49870 -1160
rect 49600 -1260 49620 -1200
rect 49680 -1260 49700 -1200
rect 49600 -1270 49700 -1260
rect 49940 -1200 50040 -1060
rect 50280 -770 50380 -750
rect 50280 -830 50300 -770
rect 50360 -830 50380 -770
rect 50280 -880 50380 -830
rect 50280 -950 50300 -880
rect 50360 -950 50380 -880
rect 50280 -1000 50380 -950
rect 50280 -1060 50300 -1000
rect 50360 -1060 50380 -1000
rect 50110 -1100 50210 -1080
rect 50110 -1160 50130 -1100
rect 50190 -1160 50210 -1100
rect 50110 -1180 50210 -1160
rect 49940 -1260 49960 -1200
rect 50020 -1260 50040 -1200
rect 49940 -1270 50040 -1260
rect 50280 -1200 50380 -1060
rect 50620 -770 50720 -750
rect 50620 -830 50640 -770
rect 50700 -830 50720 -770
rect 50620 -880 50720 -830
rect 50620 -950 50640 -880
rect 50700 -950 50720 -880
rect 50620 -1000 50720 -950
rect 50620 -1060 50640 -1000
rect 50700 -1060 50720 -1000
rect 50450 -1100 50550 -1080
rect 50450 -1160 50470 -1100
rect 50530 -1160 50550 -1100
rect 50450 -1180 50550 -1160
rect 50280 -1260 50300 -1200
rect 50360 -1260 50380 -1200
rect 50280 -1270 50380 -1260
rect 50620 -1200 50720 -1060
rect 50960 -770 51060 -750
rect 50960 -830 50980 -770
rect 51040 -830 51060 -770
rect 50960 -880 51060 -830
rect 50960 -950 50980 -880
rect 51040 -950 51060 -880
rect 50960 -1000 51060 -950
rect 50960 -1060 50980 -1000
rect 51040 -1060 51060 -1000
rect 50790 -1100 50890 -1080
rect 50790 -1160 50810 -1100
rect 50870 -1160 50890 -1100
rect 50790 -1180 50890 -1160
rect 50620 -1260 50640 -1200
rect 50700 -1260 50720 -1200
rect 50620 -1270 50720 -1260
rect 50960 -1200 51060 -1060
rect 51300 -770 51400 -750
rect 51300 -830 51320 -770
rect 51380 -830 51400 -770
rect 51300 -880 51400 -830
rect 51300 -950 51320 -880
rect 51380 -950 51400 -880
rect 51300 -1000 51400 -950
rect 51300 -1060 51320 -1000
rect 51380 -1060 51400 -1000
rect 51130 -1100 51230 -1080
rect 51130 -1160 51150 -1100
rect 51210 -1160 51230 -1100
rect 51130 -1180 51230 -1160
rect 50960 -1260 50980 -1200
rect 51040 -1260 51060 -1200
rect 50960 -1270 51060 -1260
rect 51300 -1200 51400 -1060
rect 51640 -770 51740 -750
rect 51640 -830 51660 -770
rect 51720 -830 51740 -770
rect 51640 -880 51740 -830
rect 51640 -950 51660 -880
rect 51720 -950 51740 -880
rect 51640 -1000 51740 -950
rect 51640 -1060 51660 -1000
rect 51720 -1060 51740 -1000
rect 51470 -1100 51570 -1080
rect 51470 -1160 51490 -1100
rect 51550 -1160 51570 -1100
rect 51470 -1180 51570 -1160
rect 51300 -1260 51320 -1200
rect 51380 -1260 51400 -1200
rect 51300 -1270 51400 -1260
rect 51640 -1200 51740 -1060
rect 51980 -770 52080 -750
rect 51980 -830 52000 -770
rect 52060 -830 52080 -770
rect 51980 -880 52080 -830
rect 51980 -950 52000 -880
rect 52060 -950 52080 -880
rect 51980 -1000 52080 -950
rect 51980 -1060 52000 -1000
rect 52060 -1060 52080 -1000
rect 51810 -1100 51910 -1080
rect 51810 -1160 51830 -1100
rect 51890 -1160 51910 -1100
rect 51810 -1180 51910 -1160
rect 51640 -1260 51660 -1200
rect 51720 -1260 51740 -1200
rect 51640 -1270 51740 -1260
rect 51980 -1200 52080 -1060
rect 52320 -770 52420 -750
rect 52320 -830 52340 -770
rect 52400 -830 52420 -770
rect 52320 -880 52420 -830
rect 52320 -950 52340 -880
rect 52400 -950 52420 -880
rect 52320 -1000 52420 -950
rect 52320 -1060 52340 -1000
rect 52400 -1060 52420 -1000
rect 52150 -1100 52250 -1080
rect 52150 -1160 52170 -1100
rect 52230 -1160 52250 -1100
rect 52150 -1180 52250 -1160
rect 51980 -1260 52000 -1200
rect 52060 -1260 52080 -1200
rect 51980 -1270 52080 -1260
rect 52320 -1200 52420 -1060
rect 52660 -770 52760 -750
rect 52660 -830 52680 -770
rect 52740 -830 52760 -770
rect 52660 -880 52760 -830
rect 52660 -950 52680 -880
rect 52740 -950 52760 -880
rect 52660 -1000 52760 -950
rect 52660 -1060 52680 -1000
rect 52740 -1060 52760 -1000
rect 52490 -1100 52590 -1080
rect 52490 -1160 52510 -1100
rect 52570 -1160 52590 -1100
rect 52490 -1180 52590 -1160
rect 52320 -1260 52340 -1200
rect 52400 -1260 52420 -1200
rect 52320 -1270 52420 -1260
rect 52660 -1200 52760 -1060
rect 53000 -770 53100 -750
rect 53000 -830 53020 -770
rect 53080 -830 53100 -770
rect 53000 -880 53100 -830
rect 53000 -950 53020 -880
rect 53080 -950 53100 -880
rect 53000 -1000 53100 -950
rect 53000 -1060 53020 -1000
rect 53080 -1060 53100 -1000
rect 52830 -1100 52930 -1080
rect 52830 -1160 52850 -1100
rect 52910 -1160 52930 -1100
rect 52830 -1180 52930 -1160
rect 52660 -1260 52680 -1200
rect 52740 -1260 52760 -1200
rect 52660 -1270 52760 -1260
rect 53000 -1200 53100 -1060
rect 53340 -770 53440 -750
rect 53340 -830 53360 -770
rect 53420 -830 53440 -770
rect 53340 -880 53440 -830
rect 53340 -950 53360 -880
rect 53420 -950 53440 -880
rect 53340 -1000 53440 -950
rect 53340 -1060 53360 -1000
rect 53420 -1060 53440 -1000
rect 53170 -1100 53270 -1080
rect 53170 -1160 53190 -1100
rect 53250 -1160 53270 -1100
rect 53170 -1180 53270 -1160
rect 53000 -1260 53020 -1200
rect 53080 -1260 53100 -1200
rect 53000 -1270 53100 -1260
rect 53340 -1200 53440 -1060
rect 53680 -770 53780 -750
rect 53680 -830 53700 -770
rect 53760 -830 53780 -770
rect 53680 -880 53780 -830
rect 53680 -950 53700 -880
rect 53760 -950 53780 -880
rect 53680 -1000 53780 -950
rect 53680 -1060 53700 -1000
rect 53760 -1060 53780 -1000
rect 53510 -1100 53610 -1080
rect 53510 -1160 53530 -1100
rect 53590 -1160 53610 -1100
rect 53510 -1180 53610 -1160
rect 53340 -1260 53360 -1200
rect 53420 -1260 53440 -1200
rect 53340 -1270 53440 -1260
rect 53680 -1200 53780 -1060
rect 54020 -770 54120 -750
rect 54020 -830 54040 -770
rect 54100 -830 54120 -770
rect 54020 -880 54120 -830
rect 54020 -950 54040 -880
rect 54100 -950 54120 -880
rect 54020 -1000 54120 -950
rect 54020 -1060 54040 -1000
rect 54100 -1060 54120 -1000
rect 53850 -1100 53950 -1080
rect 53850 -1160 53870 -1100
rect 53930 -1160 53950 -1100
rect 53850 -1180 53950 -1160
rect 53680 -1260 53700 -1200
rect 53760 -1260 53780 -1200
rect 53680 -1270 53780 -1260
rect 54020 -1200 54120 -1060
rect 54360 -770 54460 -750
rect 54360 -830 54380 -770
rect 54440 -830 54460 -770
rect 54360 -880 54460 -830
rect 54360 -950 54380 -880
rect 54440 -950 54460 -880
rect 54360 -1000 54460 -950
rect 54360 -1060 54380 -1000
rect 54440 -1060 54460 -1000
rect 54190 -1100 54290 -1080
rect 54190 -1160 54210 -1100
rect 54270 -1160 54290 -1100
rect 54190 -1180 54290 -1160
rect 54020 -1260 54040 -1200
rect 54100 -1260 54120 -1200
rect 54020 -1270 54120 -1260
rect 54360 -1200 54460 -1060
rect 54700 -770 54800 -750
rect 54700 -830 54720 -770
rect 54780 -830 54800 -770
rect 54700 -880 54800 -830
rect 54700 -950 54720 -880
rect 54780 -950 54800 -880
rect 54700 -1000 54800 -950
rect 54700 -1060 54720 -1000
rect 54780 -1060 54800 -1000
rect 54530 -1100 54630 -1080
rect 54530 -1160 54550 -1100
rect 54610 -1160 54630 -1100
rect 54530 -1180 54630 -1160
rect 54360 -1260 54380 -1200
rect 54440 -1260 54460 -1200
rect 54360 -1270 54460 -1260
rect 54700 -1200 54800 -1060
rect 55040 -770 55140 -750
rect 55040 -830 55060 -770
rect 55120 -830 55140 -770
rect 55040 -880 55140 -830
rect 55040 -950 55060 -880
rect 55120 -950 55140 -880
rect 55040 -1000 55140 -950
rect 55040 -1060 55060 -1000
rect 55120 -1060 55140 -1000
rect 54870 -1100 54970 -1080
rect 54870 -1160 54890 -1100
rect 54950 -1160 54970 -1100
rect 54870 -1180 54970 -1160
rect 54700 -1260 54720 -1200
rect 54780 -1260 54800 -1200
rect 54700 -1270 54800 -1260
rect 55040 -1200 55140 -1060
rect 55380 -770 55480 -750
rect 55380 -830 55400 -770
rect 55460 -830 55480 -770
rect 55380 -880 55480 -830
rect 55380 -950 55400 -880
rect 55460 -950 55480 -880
rect 55380 -1000 55480 -950
rect 55380 -1060 55400 -1000
rect 55460 -1060 55480 -1000
rect 55210 -1100 55310 -1080
rect 55210 -1160 55230 -1100
rect 55290 -1160 55310 -1100
rect 55210 -1180 55310 -1160
rect 55040 -1260 55060 -1200
rect 55120 -1260 55140 -1200
rect 55040 -1270 55140 -1260
rect 55380 -1200 55480 -1060
rect 55720 -770 55820 -750
rect 55720 -830 55740 -770
rect 55800 -830 55820 -770
rect 55720 -880 55820 -830
rect 55720 -950 55740 -880
rect 55800 -950 55820 -880
rect 55720 -1000 55820 -950
rect 55720 -1060 55740 -1000
rect 55800 -1060 55820 -1000
rect 55550 -1100 55650 -1080
rect 55550 -1160 55570 -1100
rect 55630 -1160 55650 -1100
rect 55550 -1180 55650 -1160
rect 55380 -1260 55400 -1200
rect 55460 -1260 55480 -1200
rect 55380 -1270 55480 -1260
rect 55720 -1200 55820 -1060
rect 56060 -770 56160 -750
rect 56060 -830 56080 -770
rect 56140 -830 56160 -770
rect 56060 -880 56160 -830
rect 56060 -950 56080 -880
rect 56140 -950 56160 -880
rect 56060 -1000 56160 -950
rect 56060 -1060 56080 -1000
rect 56140 -1060 56160 -1000
rect 55890 -1100 55990 -1080
rect 55890 -1160 55910 -1100
rect 55970 -1160 55990 -1100
rect 55890 -1180 55990 -1160
rect 55720 -1260 55740 -1200
rect 55800 -1260 55820 -1200
rect 55720 -1270 55820 -1260
rect 56060 -1200 56160 -1060
rect 56400 -770 56500 -750
rect 56400 -830 56420 -770
rect 56480 -830 56500 -770
rect 56400 -880 56500 -830
rect 56400 -950 56420 -880
rect 56480 -950 56500 -880
rect 56400 -1000 56500 -950
rect 56400 -1060 56420 -1000
rect 56480 -1060 56500 -1000
rect 56230 -1100 56330 -1080
rect 56230 -1160 56250 -1100
rect 56310 -1160 56330 -1100
rect 56230 -1180 56330 -1160
rect 56060 -1260 56080 -1200
rect 56140 -1260 56160 -1200
rect 56060 -1270 56160 -1260
rect 56400 -1200 56500 -1060
rect 56740 -770 56840 -750
rect 56740 -830 56760 -770
rect 56820 -830 56840 -770
rect 56740 -880 56840 -830
rect 56740 -950 56760 -880
rect 56820 -950 56840 -880
rect 56740 -1000 56840 -950
rect 56740 -1060 56760 -1000
rect 56820 -1060 56840 -1000
rect 56570 -1100 56670 -1080
rect 56570 -1160 56590 -1100
rect 56650 -1160 56670 -1100
rect 56570 -1180 56670 -1160
rect 56400 -1260 56420 -1200
rect 56480 -1260 56500 -1200
rect 56400 -1270 56500 -1260
rect 56740 -1200 56840 -1060
rect 57080 -770 57180 -750
rect 57080 -830 57100 -770
rect 57160 -830 57180 -770
rect 57080 -880 57180 -830
rect 57080 -950 57100 -880
rect 57160 -950 57180 -880
rect 57080 -1000 57180 -950
rect 57080 -1060 57100 -1000
rect 57160 -1060 57180 -1000
rect 56910 -1100 57010 -1080
rect 56910 -1160 56930 -1100
rect 56990 -1160 57010 -1100
rect 56910 -1180 57010 -1160
rect 56740 -1260 56760 -1200
rect 56820 -1260 56840 -1200
rect 56740 -1270 56840 -1260
rect 57080 -1200 57180 -1060
rect 57420 -770 57520 -750
rect 57420 -830 57440 -770
rect 57500 -830 57520 -770
rect 57420 -880 57520 -830
rect 57420 -950 57440 -880
rect 57500 -950 57520 -880
rect 57420 -1000 57520 -950
rect 57420 -1060 57440 -1000
rect 57500 -1060 57520 -1000
rect 57250 -1100 57350 -1080
rect 57250 -1160 57270 -1100
rect 57330 -1160 57350 -1100
rect 57250 -1180 57350 -1160
rect 57080 -1260 57100 -1200
rect 57160 -1260 57180 -1200
rect 57080 -1270 57180 -1260
rect 57420 -1200 57520 -1060
rect 57760 -770 57860 -750
rect 57760 -830 57780 -770
rect 57840 -830 57860 -770
rect 57760 -880 57860 -830
rect 57760 -950 57780 -880
rect 57840 -950 57860 -880
rect 57760 -1000 57860 -950
rect 57760 -1060 57780 -1000
rect 57840 -1060 57860 -1000
rect 57590 -1100 57690 -1080
rect 57590 -1160 57610 -1100
rect 57670 -1160 57690 -1100
rect 57590 -1180 57690 -1160
rect 57420 -1260 57440 -1200
rect 57500 -1260 57520 -1200
rect 57420 -1270 57520 -1260
rect 57760 -1200 57860 -1060
rect 58100 -770 58200 -750
rect 58100 -830 58120 -770
rect 58180 -830 58200 -770
rect 58100 -880 58200 -830
rect 58100 -950 58120 -880
rect 58180 -950 58200 -880
rect 58100 -1000 58200 -950
rect 58100 -1060 58120 -1000
rect 58180 -1060 58200 -1000
rect 57930 -1100 58030 -1080
rect 57930 -1160 57950 -1100
rect 58010 -1160 58030 -1100
rect 57930 -1180 58030 -1160
rect 57760 -1260 57780 -1200
rect 57840 -1260 57860 -1200
rect 57760 -1270 57860 -1260
rect 58100 -1200 58200 -1060
rect 58440 -770 58540 -750
rect 58440 -830 58460 -770
rect 58520 -830 58540 -770
rect 58440 -880 58540 -830
rect 58440 -950 58460 -880
rect 58520 -950 58540 -880
rect 58440 -1000 58540 -950
rect 58440 -1060 58460 -1000
rect 58520 -1060 58540 -1000
rect 58270 -1100 58370 -1080
rect 58270 -1160 58290 -1100
rect 58350 -1160 58370 -1100
rect 58270 -1180 58370 -1160
rect 58100 -1260 58120 -1200
rect 58180 -1260 58200 -1200
rect 58100 -1270 58200 -1260
rect 58440 -1200 58540 -1060
rect 58780 -770 58880 -750
rect 58780 -830 58800 -770
rect 58860 -830 58880 -770
rect 58780 -880 58880 -830
rect 58780 -950 58800 -880
rect 58860 -950 58880 -880
rect 58780 -1000 58880 -950
rect 58780 -1060 58800 -1000
rect 58860 -1060 58880 -1000
rect 58610 -1100 58710 -1080
rect 58610 -1160 58630 -1100
rect 58690 -1160 58710 -1100
rect 58610 -1180 58710 -1160
rect 58440 -1260 58460 -1200
rect 58520 -1260 58540 -1200
rect 58440 -1270 58540 -1260
rect 58780 -1200 58880 -1060
rect 59120 -770 59220 -750
rect 59120 -830 59140 -770
rect 59200 -830 59220 -770
rect 59120 -880 59220 -830
rect 59120 -950 59140 -880
rect 59200 -950 59220 -880
rect 59120 -1000 59220 -950
rect 59120 -1060 59140 -1000
rect 59200 -1060 59220 -1000
rect 58950 -1100 59050 -1080
rect 58950 -1160 58970 -1100
rect 59030 -1160 59050 -1100
rect 58950 -1180 59050 -1160
rect 58780 -1260 58800 -1200
rect 58860 -1260 58880 -1200
rect 58780 -1270 58880 -1260
rect 59120 -1200 59220 -1060
rect 59460 -770 59560 -750
rect 59460 -830 59480 -770
rect 59540 -830 59560 -770
rect 59460 -880 59560 -830
rect 59460 -950 59480 -880
rect 59540 -950 59560 -880
rect 59460 -1000 59560 -950
rect 59460 -1060 59480 -1000
rect 59540 -1060 59560 -1000
rect 59290 -1100 59390 -1080
rect 59290 -1160 59310 -1100
rect 59370 -1160 59390 -1100
rect 59290 -1180 59390 -1160
rect 59120 -1260 59140 -1200
rect 59200 -1260 59220 -1200
rect 59120 -1270 59220 -1260
rect 59460 -1200 59560 -1060
rect 59800 -770 59900 -750
rect 59800 -830 59820 -770
rect 59880 -830 59900 -770
rect 59800 -880 59900 -830
rect 59800 -950 59820 -880
rect 59880 -950 59900 -880
rect 59800 -1000 59900 -950
rect 59800 -1060 59820 -1000
rect 59880 -1060 59900 -1000
rect 59630 -1100 59730 -1080
rect 59630 -1160 59650 -1100
rect 59710 -1160 59730 -1100
rect 59630 -1180 59730 -1160
rect 59460 -1260 59480 -1200
rect 59540 -1260 59560 -1200
rect 59460 -1270 59560 -1260
rect 59800 -1200 59900 -1060
rect 60140 -770 60240 -750
rect 60140 -830 60160 -770
rect 60220 -830 60240 -770
rect 60140 -880 60240 -830
rect 60140 -950 60160 -880
rect 60220 -950 60240 -880
rect 60140 -1000 60240 -950
rect 60140 -1060 60160 -1000
rect 60220 -1060 60240 -1000
rect 59970 -1100 60070 -1080
rect 59970 -1160 59990 -1100
rect 60050 -1160 60070 -1100
rect 59970 -1180 60070 -1160
rect 59800 -1260 59820 -1200
rect 59880 -1260 59900 -1200
rect 59800 -1270 59900 -1260
rect 60140 -1200 60240 -1060
rect 60480 -770 60580 -750
rect 60480 -830 60500 -770
rect 60560 -830 60580 -770
rect 60480 -880 60580 -830
rect 60480 -950 60500 -880
rect 60560 -950 60580 -880
rect 60480 -1000 60580 -950
rect 60480 -1060 60500 -1000
rect 60560 -1060 60580 -1000
rect 60310 -1100 60410 -1080
rect 60310 -1160 60330 -1100
rect 60390 -1160 60410 -1100
rect 60310 -1180 60410 -1160
rect 60140 -1260 60160 -1200
rect 60220 -1260 60240 -1200
rect 60140 -1270 60240 -1260
rect 60480 -1200 60580 -1060
rect 60820 -770 60920 -750
rect 60820 -830 60840 -770
rect 60900 -830 60920 -770
rect 60820 -880 60920 -830
rect 60820 -950 60840 -880
rect 60900 -950 60920 -880
rect 60820 -1000 60920 -950
rect 60820 -1060 60840 -1000
rect 60900 -1060 60920 -1000
rect 60650 -1100 60750 -1080
rect 60650 -1160 60670 -1100
rect 60730 -1160 60750 -1100
rect 60650 -1180 60750 -1160
rect 60480 -1260 60500 -1200
rect 60560 -1260 60580 -1200
rect 60480 -1270 60580 -1260
rect 60820 -1200 60920 -1060
rect 61160 -770 61260 -750
rect 61160 -830 61180 -770
rect 61240 -830 61260 -770
rect 61160 -880 61260 -830
rect 61160 -950 61180 -880
rect 61240 -950 61260 -880
rect 61160 -1000 61260 -950
rect 61160 -1060 61180 -1000
rect 61240 -1060 61260 -1000
rect 60990 -1100 61090 -1080
rect 60990 -1160 61010 -1100
rect 61070 -1160 61090 -1100
rect 60990 -1180 61090 -1160
rect 60820 -1260 60840 -1200
rect 60900 -1260 60920 -1200
rect 60820 -1270 60920 -1260
rect 61160 -1200 61260 -1060
rect 61500 -770 61600 -750
rect 61500 -830 61520 -770
rect 61580 -830 61600 -770
rect 61500 -880 61600 -830
rect 61500 -950 61520 -880
rect 61580 -950 61600 -880
rect 61500 -1000 61600 -950
rect 61500 -1060 61520 -1000
rect 61580 -1060 61600 -1000
rect 61330 -1100 61430 -1080
rect 61330 -1160 61350 -1100
rect 61410 -1160 61430 -1100
rect 61330 -1180 61430 -1160
rect 61160 -1260 61180 -1200
rect 61240 -1260 61260 -1200
rect 61160 -1270 61260 -1260
rect 61500 -1200 61600 -1060
rect 61840 -770 61940 -750
rect 61840 -830 61860 -770
rect 61920 -830 61940 -770
rect 61840 -880 61940 -830
rect 61840 -950 61860 -880
rect 61920 -950 61940 -880
rect 61840 -1000 61940 -950
rect 61840 -1060 61860 -1000
rect 61920 -1060 61940 -1000
rect 61670 -1100 61770 -1080
rect 61670 -1160 61690 -1100
rect 61750 -1160 61770 -1100
rect 61670 -1180 61770 -1160
rect 61500 -1260 61520 -1200
rect 61580 -1260 61600 -1200
rect 61500 -1270 61600 -1260
rect 61840 -1200 61940 -1060
rect 62180 -770 62280 -750
rect 62180 -830 62200 -770
rect 62260 -830 62280 -770
rect 62180 -880 62280 -830
rect 62180 -950 62200 -880
rect 62260 -950 62280 -880
rect 62180 -1000 62280 -950
rect 62180 -1060 62200 -1000
rect 62260 -1060 62280 -1000
rect 62010 -1100 62110 -1080
rect 62010 -1160 62030 -1100
rect 62090 -1160 62110 -1100
rect 62010 -1180 62110 -1160
rect 61840 -1260 61860 -1200
rect 61920 -1260 61940 -1200
rect 61840 -1270 61940 -1260
rect 62180 -1200 62280 -1060
rect 62520 -770 62620 -750
rect 62520 -830 62540 -770
rect 62600 -830 62620 -770
rect 62520 -880 62620 -830
rect 62520 -950 62540 -880
rect 62600 -950 62620 -880
rect 62520 -1000 62620 -950
rect 62520 -1060 62540 -1000
rect 62600 -1060 62620 -1000
rect 62350 -1100 62450 -1080
rect 62350 -1160 62370 -1100
rect 62430 -1160 62450 -1100
rect 62350 -1180 62450 -1160
rect 62180 -1260 62200 -1200
rect 62260 -1260 62280 -1200
rect 62180 -1270 62280 -1260
rect 62520 -1200 62620 -1060
rect 62860 -770 62960 -750
rect 62860 -830 62880 -770
rect 62940 -830 62960 -770
rect 62860 -880 62960 -830
rect 62860 -950 62880 -880
rect 62940 -950 62960 -880
rect 62860 -1000 62960 -950
rect 62860 -1060 62880 -1000
rect 62940 -1060 62960 -1000
rect 62690 -1100 62790 -1080
rect 62690 -1160 62710 -1100
rect 62770 -1160 62790 -1100
rect 62690 -1180 62790 -1160
rect 62520 -1260 62540 -1200
rect 62600 -1260 62620 -1200
rect 62520 -1270 62620 -1260
rect 62860 -1200 62960 -1060
rect 63200 -770 63300 -750
rect 63200 -830 63220 -770
rect 63280 -830 63300 -770
rect 63200 -880 63300 -830
rect 63200 -950 63220 -880
rect 63280 -950 63300 -880
rect 63200 -1000 63300 -950
rect 63200 -1060 63220 -1000
rect 63280 -1060 63300 -1000
rect 63030 -1100 63130 -1080
rect 63030 -1160 63050 -1100
rect 63110 -1160 63130 -1100
rect 63030 -1180 63130 -1160
rect 62860 -1260 62880 -1200
rect 62940 -1260 62960 -1200
rect 62860 -1270 62960 -1260
rect 63200 -1200 63300 -1060
rect 63540 -770 63640 -750
rect 63540 -830 63560 -770
rect 63620 -830 63640 -770
rect 63540 -880 63640 -830
rect 63540 -950 63560 -880
rect 63620 -950 63640 -880
rect 63540 -1000 63640 -950
rect 63540 -1060 63560 -1000
rect 63620 -1060 63640 -1000
rect 63370 -1100 63470 -1080
rect 63370 -1160 63390 -1100
rect 63450 -1160 63470 -1100
rect 63370 -1180 63470 -1160
rect 63200 -1260 63220 -1200
rect 63280 -1260 63300 -1200
rect 63200 -1270 63300 -1260
rect 63540 -1200 63640 -1060
rect 63880 -770 63980 -750
rect 63880 -830 63900 -770
rect 63960 -830 63980 -770
rect 63880 -880 63980 -830
rect 63880 -950 63900 -880
rect 63960 -950 63980 -880
rect 63880 -1000 63980 -950
rect 63880 -1060 63900 -1000
rect 63960 -1060 63980 -1000
rect 63710 -1100 63810 -1080
rect 63710 -1160 63730 -1100
rect 63790 -1160 63810 -1100
rect 63710 -1180 63810 -1160
rect 63540 -1260 63560 -1200
rect 63620 -1260 63640 -1200
rect 63540 -1270 63640 -1260
rect 63880 -1200 63980 -1060
rect 64220 -770 64320 -750
rect 64220 -830 64240 -770
rect 64300 -830 64320 -770
rect 64220 -880 64320 -830
rect 64220 -950 64240 -880
rect 64300 -950 64320 -880
rect 64220 -1000 64320 -950
rect 64220 -1060 64240 -1000
rect 64300 -1060 64320 -1000
rect 64050 -1100 64150 -1080
rect 64050 -1160 64070 -1100
rect 64130 -1160 64150 -1100
rect 64050 -1180 64150 -1160
rect 63880 -1260 63900 -1200
rect 63960 -1260 63980 -1200
rect 63880 -1270 63980 -1260
rect 64220 -1200 64320 -1060
rect 64560 -770 64660 -750
rect 64560 -830 64580 -770
rect 64640 -830 64660 -770
rect 64560 -880 64660 -830
rect 64560 -950 64580 -880
rect 64640 -950 64660 -880
rect 64560 -1000 64660 -950
rect 64560 -1060 64580 -1000
rect 64640 -1060 64660 -1000
rect 64390 -1100 64490 -1080
rect 64390 -1160 64410 -1100
rect 64470 -1160 64490 -1100
rect 64390 -1180 64490 -1160
rect 64220 -1260 64240 -1200
rect 64300 -1260 64320 -1200
rect 64220 -1270 64320 -1260
rect 64560 -1200 64660 -1060
rect 64900 -770 65000 -750
rect 64900 -830 64920 -770
rect 64980 -830 65000 -770
rect 64900 -880 65000 -830
rect 64900 -950 64920 -880
rect 64980 -950 65000 -880
rect 64900 -1000 65000 -950
rect 64900 -1060 64920 -1000
rect 64980 -1060 65000 -1000
rect 64730 -1100 64830 -1080
rect 64730 -1160 64750 -1100
rect 64810 -1160 64830 -1100
rect 64730 -1180 64830 -1160
rect 64560 -1260 64580 -1200
rect 64640 -1260 64660 -1200
rect 64560 -1270 64660 -1260
rect 64900 -1200 65000 -1060
rect 65240 -770 65340 -750
rect 65240 -830 65260 -770
rect 65320 -830 65340 -770
rect 65240 -880 65340 -830
rect 65240 -950 65260 -880
rect 65320 -950 65340 -880
rect 65240 -1000 65340 -950
rect 65240 -1060 65260 -1000
rect 65320 -1060 65340 -1000
rect 65070 -1100 65170 -1080
rect 65070 -1160 65090 -1100
rect 65150 -1160 65170 -1100
rect 65070 -1180 65170 -1160
rect 64900 -1260 64920 -1200
rect 64980 -1260 65000 -1200
rect 64900 -1270 65000 -1260
rect 65240 -1200 65340 -1060
rect 65580 -770 65680 -750
rect 65580 -830 65600 -770
rect 65660 -830 65680 -770
rect 65580 -880 65680 -830
rect 65580 -950 65600 -880
rect 65660 -950 65680 -880
rect 65580 -1000 65680 -950
rect 65580 -1060 65600 -1000
rect 65660 -1060 65680 -1000
rect 65410 -1100 65510 -1080
rect 65410 -1160 65430 -1100
rect 65490 -1160 65510 -1100
rect 65410 -1180 65510 -1160
rect 65240 -1260 65260 -1200
rect 65320 -1260 65340 -1200
rect 65240 -1270 65340 -1260
rect 65580 -1200 65680 -1060
rect 65920 -770 66020 -750
rect 65920 -830 65940 -770
rect 66000 -830 66020 -770
rect 65920 -880 66020 -830
rect 65920 -950 65940 -880
rect 66000 -950 66020 -880
rect 65920 -1000 66020 -950
rect 65920 -1060 65940 -1000
rect 66000 -1060 66020 -1000
rect 65750 -1100 65850 -1080
rect 65750 -1160 65770 -1100
rect 65830 -1160 65850 -1100
rect 65750 -1180 65850 -1160
rect 65580 -1260 65600 -1200
rect 65660 -1260 65680 -1200
rect 65580 -1270 65680 -1260
rect 65920 -1200 66020 -1060
rect 66260 -770 66360 -750
rect 66260 -830 66280 -770
rect 66340 -830 66360 -770
rect 66260 -880 66360 -830
rect 66260 -950 66280 -880
rect 66340 -950 66360 -880
rect 66260 -1000 66360 -950
rect 66260 -1060 66280 -1000
rect 66340 -1060 66360 -1000
rect 66090 -1100 66190 -1080
rect 66090 -1160 66110 -1100
rect 66170 -1160 66190 -1100
rect 66090 -1180 66190 -1160
rect 65920 -1260 65940 -1200
rect 66000 -1260 66020 -1200
rect 65920 -1270 66020 -1260
rect 66260 -1200 66360 -1060
rect 66600 -770 66700 -750
rect 66600 -830 66620 -770
rect 66680 -830 66700 -770
rect 66600 -880 66700 -830
rect 66600 -950 66620 -880
rect 66680 -950 66700 -880
rect 66600 -1000 66700 -950
rect 66600 -1060 66620 -1000
rect 66680 -1060 66700 -1000
rect 66430 -1100 66530 -1080
rect 66430 -1160 66450 -1100
rect 66510 -1160 66530 -1100
rect 66430 -1180 66530 -1160
rect 66260 -1260 66280 -1200
rect 66340 -1260 66360 -1200
rect 66260 -1270 66360 -1260
rect 66600 -1200 66700 -1060
rect 66940 -770 67040 -750
rect 66940 -830 66960 -770
rect 67020 -830 67040 -770
rect 66940 -880 67040 -830
rect 66940 -950 66960 -880
rect 67020 -950 67040 -880
rect 66940 -1000 67040 -950
rect 66940 -1060 66960 -1000
rect 67020 -1060 67040 -1000
rect 66770 -1100 66870 -1080
rect 66770 -1160 66790 -1100
rect 66850 -1160 66870 -1100
rect 66770 -1180 66870 -1160
rect 66600 -1260 66620 -1200
rect 66680 -1260 66700 -1200
rect 66600 -1270 66700 -1260
rect 66940 -1200 67040 -1060
rect 67280 -770 67380 -750
rect 67280 -830 67300 -770
rect 67360 -830 67380 -770
rect 67280 -880 67380 -830
rect 67280 -950 67300 -880
rect 67360 -950 67380 -880
rect 67280 -1000 67380 -950
rect 67280 -1060 67300 -1000
rect 67360 -1060 67380 -1000
rect 67110 -1100 67210 -1080
rect 67110 -1160 67130 -1100
rect 67190 -1160 67210 -1100
rect 67110 -1180 67210 -1160
rect 66940 -1260 66960 -1200
rect 67020 -1260 67040 -1200
rect 66940 -1270 67040 -1260
rect 67280 -1200 67380 -1060
rect 67620 -770 67720 -750
rect 67620 -830 67640 -770
rect 67700 -830 67720 -770
rect 67620 -880 67720 -830
rect 67620 -950 67640 -880
rect 67700 -950 67720 -880
rect 67620 -1000 67720 -950
rect 67620 -1060 67640 -1000
rect 67700 -1060 67720 -1000
rect 67450 -1100 67550 -1080
rect 67450 -1160 67470 -1100
rect 67530 -1160 67550 -1100
rect 67450 -1180 67550 -1160
rect 67280 -1260 67300 -1200
rect 67360 -1260 67380 -1200
rect 67280 -1270 67380 -1260
rect 67620 -1200 67720 -1060
rect 67960 -770 68060 -750
rect 67960 -830 67980 -770
rect 68040 -830 68060 -770
rect 67960 -880 68060 -830
rect 67960 -950 67980 -880
rect 68040 -950 68060 -880
rect 67960 -1000 68060 -950
rect 67960 -1060 67980 -1000
rect 68040 -1060 68060 -1000
rect 67790 -1100 67890 -1080
rect 67790 -1160 67810 -1100
rect 67870 -1160 67890 -1100
rect 67790 -1180 67890 -1160
rect 67620 -1260 67640 -1200
rect 67700 -1260 67720 -1200
rect 67620 -1270 67720 -1260
rect 67960 -1200 68060 -1060
rect 68300 -770 68400 -750
rect 68300 -830 68320 -770
rect 68380 -830 68400 -770
rect 68300 -880 68400 -830
rect 68300 -950 68320 -880
rect 68380 -950 68400 -880
rect 68300 -1000 68400 -950
rect 68300 -1060 68320 -1000
rect 68380 -1060 68400 -1000
rect 68130 -1100 68230 -1080
rect 68130 -1160 68150 -1100
rect 68210 -1160 68230 -1100
rect 68130 -1180 68230 -1160
rect 67960 -1260 67980 -1200
rect 68040 -1260 68060 -1200
rect 67960 -1270 68060 -1260
rect 68300 -1200 68400 -1060
rect 68640 -770 68740 -750
rect 68640 -830 68660 -770
rect 68720 -830 68740 -770
rect 68640 -880 68740 -830
rect 68640 -950 68660 -880
rect 68720 -950 68740 -880
rect 68640 -1000 68740 -950
rect 68640 -1060 68660 -1000
rect 68720 -1060 68740 -1000
rect 68470 -1100 68570 -1080
rect 68470 -1160 68490 -1100
rect 68550 -1160 68570 -1100
rect 68470 -1180 68570 -1160
rect 68300 -1260 68320 -1200
rect 68380 -1260 68400 -1200
rect 68300 -1270 68400 -1260
rect 68640 -1200 68740 -1060
rect 68980 -770 69080 -750
rect 68980 -830 69000 -770
rect 69060 -830 69080 -770
rect 68980 -880 69080 -830
rect 68980 -950 69000 -880
rect 69060 -950 69080 -880
rect 68980 -1000 69080 -950
rect 68980 -1060 69000 -1000
rect 69060 -1060 69080 -1000
rect 68810 -1100 68910 -1080
rect 68810 -1160 68830 -1100
rect 68890 -1160 68910 -1100
rect 68810 -1180 68910 -1160
rect 68640 -1260 68660 -1200
rect 68720 -1260 68740 -1200
rect 68640 -1270 68740 -1260
rect 68980 -1200 69080 -1060
rect 69320 -770 69420 -750
rect 69320 -830 69340 -770
rect 69400 -830 69420 -770
rect 69320 -880 69420 -830
rect 69320 -950 69340 -880
rect 69400 -950 69420 -880
rect 69320 -1000 69420 -950
rect 69320 -1060 69340 -1000
rect 69400 -1060 69420 -1000
rect 69150 -1100 69250 -1080
rect 69150 -1160 69170 -1100
rect 69230 -1160 69250 -1100
rect 69150 -1180 69250 -1160
rect 68980 -1260 69000 -1200
rect 69060 -1260 69080 -1200
rect 68980 -1270 69080 -1260
rect 69320 -1200 69420 -1060
rect 69660 -770 69760 -750
rect 69660 -830 69680 -770
rect 69740 -830 69760 -770
rect 69660 -880 69760 -830
rect 69660 -950 69680 -880
rect 69740 -950 69760 -880
rect 69660 -1000 69760 -950
rect 69660 -1060 69680 -1000
rect 69740 -1060 69760 -1000
rect 69490 -1100 69590 -1080
rect 69490 -1160 69510 -1100
rect 69570 -1160 69590 -1100
rect 69490 -1180 69590 -1160
rect 69320 -1260 69340 -1200
rect 69400 -1260 69420 -1200
rect 69320 -1270 69420 -1260
rect 69660 -1200 69760 -1060
rect 70000 -770 70100 -750
rect 70000 -830 70020 -770
rect 70080 -830 70100 -770
rect 70000 -880 70100 -830
rect 70000 -950 70020 -880
rect 70080 -950 70100 -880
rect 70000 -1000 70100 -950
rect 70000 -1060 70020 -1000
rect 70080 -1060 70100 -1000
rect 69830 -1100 69930 -1080
rect 69830 -1160 69850 -1100
rect 69910 -1160 69930 -1100
rect 69830 -1180 69930 -1160
rect 69660 -1260 69680 -1200
rect 69740 -1260 69760 -1200
rect 69660 -1270 69760 -1260
rect 70000 -1200 70100 -1060
rect 70340 -770 70440 -750
rect 70340 -830 70360 -770
rect 70420 -830 70440 -770
rect 70340 -880 70440 -830
rect 70340 -950 70360 -880
rect 70420 -950 70440 -880
rect 70340 -1000 70440 -950
rect 70340 -1060 70360 -1000
rect 70420 -1060 70440 -1000
rect 70170 -1100 70270 -1080
rect 70170 -1160 70190 -1100
rect 70250 -1160 70270 -1100
rect 70170 -1180 70270 -1160
rect 70000 -1260 70020 -1200
rect 70080 -1260 70100 -1200
rect 70000 -1270 70100 -1260
rect 70340 -1200 70440 -1060
rect 70680 -770 70780 -750
rect 70680 -830 70700 -770
rect 70760 -830 70780 -770
rect 70680 -880 70780 -830
rect 70680 -950 70700 -880
rect 70760 -950 70780 -880
rect 70680 -1000 70780 -950
rect 70680 -1060 70700 -1000
rect 70760 -1060 70780 -1000
rect 70510 -1100 70610 -1080
rect 70510 -1160 70530 -1100
rect 70590 -1160 70610 -1100
rect 70510 -1180 70610 -1160
rect 70340 -1260 70360 -1200
rect 70420 -1260 70440 -1200
rect 70340 -1270 70440 -1260
rect 70680 -1200 70780 -1060
rect 71020 -770 71120 -750
rect 71020 -830 71040 -770
rect 71100 -830 71120 -770
rect 71020 -880 71120 -830
rect 71020 -950 71040 -880
rect 71100 -950 71120 -880
rect 71020 -1000 71120 -950
rect 71020 -1060 71040 -1000
rect 71100 -1060 71120 -1000
rect 70850 -1100 70950 -1080
rect 70850 -1160 70870 -1100
rect 70930 -1160 70950 -1100
rect 70850 -1180 70950 -1160
rect 70680 -1260 70700 -1200
rect 70760 -1260 70780 -1200
rect 70680 -1270 70780 -1260
rect 71020 -1200 71120 -1060
rect 71360 -770 71460 -750
rect 71360 -830 71380 -770
rect 71440 -830 71460 -770
rect 71360 -880 71460 -830
rect 71360 -950 71380 -880
rect 71440 -950 71460 -880
rect 71360 -1000 71460 -950
rect 71360 -1060 71380 -1000
rect 71440 -1060 71460 -1000
rect 71190 -1100 71290 -1080
rect 71190 -1160 71210 -1100
rect 71270 -1160 71290 -1100
rect 71190 -1180 71290 -1160
rect 71020 -1260 71040 -1200
rect 71100 -1260 71120 -1200
rect 71020 -1270 71120 -1260
rect 71360 -1200 71460 -1060
rect 71700 -770 71800 -750
rect 71700 -830 71720 -770
rect 71780 -830 71800 -770
rect 71700 -880 71800 -830
rect 71700 -950 71720 -880
rect 71780 -950 71800 -880
rect 71700 -1000 71800 -950
rect 71700 -1060 71720 -1000
rect 71780 -1060 71800 -1000
rect 71530 -1100 71630 -1080
rect 71530 -1160 71550 -1100
rect 71610 -1160 71630 -1100
rect 71530 -1180 71630 -1160
rect 71360 -1260 71380 -1200
rect 71440 -1260 71460 -1200
rect 71360 -1270 71460 -1260
rect 71700 -1200 71800 -1060
rect 72040 -770 72140 -750
rect 72040 -830 72060 -770
rect 72120 -830 72140 -770
rect 72040 -880 72140 -830
rect 72040 -950 72060 -880
rect 72120 -950 72140 -880
rect 72040 -1000 72140 -950
rect 72040 -1060 72060 -1000
rect 72120 -1060 72140 -1000
rect 71870 -1100 71970 -1080
rect 71870 -1160 71890 -1100
rect 71950 -1160 71970 -1100
rect 71870 -1180 71970 -1160
rect 71700 -1260 71720 -1200
rect 71780 -1260 71800 -1200
rect 71700 -1270 71800 -1260
rect 72040 -1200 72140 -1060
rect 72380 -770 72480 -750
rect 72380 -830 72400 -770
rect 72460 -830 72480 -770
rect 72380 -880 72480 -830
rect 72380 -950 72400 -880
rect 72460 -950 72480 -880
rect 72380 -1000 72480 -950
rect 72380 -1060 72400 -1000
rect 72460 -1060 72480 -1000
rect 72210 -1100 72310 -1080
rect 72210 -1160 72230 -1100
rect 72290 -1160 72310 -1100
rect 72210 -1180 72310 -1160
rect 72040 -1260 72060 -1200
rect 72120 -1260 72140 -1200
rect 72040 -1270 72140 -1260
rect 72380 -1200 72480 -1060
rect 72720 -770 72820 -750
rect 72720 -830 72740 -770
rect 72800 -830 72820 -770
rect 72720 -880 72820 -830
rect 72720 -950 72740 -880
rect 72800 -950 72820 -880
rect 72720 -1000 72820 -950
rect 72720 -1060 72740 -1000
rect 72800 -1060 72820 -1000
rect 72550 -1100 72650 -1080
rect 72550 -1160 72570 -1100
rect 72630 -1160 72650 -1100
rect 72550 -1180 72650 -1160
rect 72380 -1260 72400 -1200
rect 72460 -1260 72480 -1200
rect 72380 -1270 72480 -1260
rect 72720 -1200 72820 -1060
rect 73060 -770 73160 -750
rect 73060 -830 73080 -770
rect 73140 -830 73160 -770
rect 73060 -880 73160 -830
rect 73060 -950 73080 -880
rect 73140 -950 73160 -880
rect 73060 -1000 73160 -950
rect 73060 -1060 73080 -1000
rect 73140 -1060 73160 -1000
rect 72890 -1100 72990 -1080
rect 72890 -1160 72910 -1100
rect 72970 -1160 72990 -1100
rect 72890 -1180 72990 -1160
rect 72720 -1260 72740 -1200
rect 72800 -1260 72820 -1200
rect 72720 -1270 72820 -1260
rect 73060 -1200 73160 -1060
rect 73400 -770 73500 -750
rect 73400 -830 73420 -770
rect 73480 -830 73500 -770
rect 73400 -880 73500 -830
rect 73400 -950 73420 -880
rect 73480 -950 73500 -880
rect 73400 -1000 73500 -950
rect 73400 -1060 73420 -1000
rect 73480 -1060 73500 -1000
rect 73230 -1100 73330 -1080
rect 73230 -1160 73250 -1100
rect 73310 -1160 73330 -1100
rect 73230 -1180 73330 -1160
rect 73060 -1260 73080 -1200
rect 73140 -1260 73160 -1200
rect 73060 -1270 73160 -1260
rect 73400 -1200 73500 -1060
rect 73740 -770 73840 -750
rect 73740 -830 73760 -770
rect 73820 -830 73840 -770
rect 73740 -880 73840 -830
rect 73740 -950 73760 -880
rect 73820 -950 73840 -880
rect 73740 -1000 73840 -950
rect 73740 -1060 73760 -1000
rect 73820 -1060 73840 -1000
rect 73570 -1100 73670 -1080
rect 73570 -1160 73590 -1100
rect 73650 -1160 73670 -1100
rect 73570 -1180 73670 -1160
rect 73400 -1260 73420 -1200
rect 73480 -1260 73500 -1200
rect 73400 -1270 73500 -1260
rect 73740 -1200 73840 -1060
rect 74080 -770 74180 -750
rect 74080 -830 74100 -770
rect 74160 -830 74180 -770
rect 74080 -880 74180 -830
rect 74080 -950 74100 -880
rect 74160 -950 74180 -880
rect 74080 -1000 74180 -950
rect 74080 -1060 74100 -1000
rect 74160 -1060 74180 -1000
rect 73910 -1100 74010 -1080
rect 73910 -1160 73930 -1100
rect 73990 -1160 74010 -1100
rect 73910 -1180 74010 -1160
rect 73740 -1260 73760 -1200
rect 73820 -1260 73840 -1200
rect 73740 -1270 73840 -1260
rect 74080 -1200 74180 -1060
rect 74420 -770 74520 -750
rect 74420 -830 74440 -770
rect 74500 -830 74520 -770
rect 74420 -880 74520 -830
rect 74420 -950 74440 -880
rect 74500 -950 74520 -880
rect 74420 -1000 74520 -950
rect 74420 -1060 74440 -1000
rect 74500 -1060 74520 -1000
rect 74250 -1100 74350 -1080
rect 74250 -1160 74270 -1100
rect 74330 -1160 74350 -1100
rect 74250 -1180 74350 -1160
rect 74080 -1260 74100 -1200
rect 74160 -1260 74180 -1200
rect 74080 -1270 74180 -1260
rect 74420 -1200 74520 -1060
rect 74760 -770 74860 -750
rect 74760 -830 74780 -770
rect 74840 -830 74860 -770
rect 74760 -880 74860 -830
rect 74760 -950 74780 -880
rect 74840 -950 74860 -880
rect 74760 -1000 74860 -950
rect 74760 -1060 74780 -1000
rect 74840 -1060 74860 -1000
rect 74590 -1100 74690 -1080
rect 74590 -1160 74610 -1100
rect 74670 -1160 74690 -1100
rect 74590 -1180 74690 -1160
rect 74420 -1260 74440 -1200
rect 74500 -1260 74520 -1200
rect 74420 -1270 74520 -1260
rect 74760 -1200 74860 -1060
rect 75100 -770 75200 -750
rect 75100 -830 75120 -770
rect 75180 -830 75200 -770
rect 75100 -880 75200 -830
rect 75100 -950 75120 -880
rect 75180 -950 75200 -880
rect 75100 -1000 75200 -950
rect 75100 -1060 75120 -1000
rect 75180 -1060 75200 -1000
rect 74930 -1100 75030 -1080
rect 74930 -1160 74950 -1100
rect 75010 -1160 75030 -1100
rect 74930 -1180 75030 -1160
rect 74760 -1260 74780 -1200
rect 74840 -1260 74860 -1200
rect 74760 -1270 74860 -1260
rect 75100 -1200 75200 -1060
rect 75440 -770 75540 -750
rect 75440 -830 75460 -770
rect 75520 -830 75540 -770
rect 75440 -880 75540 -830
rect 75440 -950 75460 -880
rect 75520 -950 75540 -880
rect 75440 -1000 75540 -950
rect 75440 -1060 75460 -1000
rect 75520 -1060 75540 -1000
rect 75270 -1100 75370 -1080
rect 75270 -1160 75290 -1100
rect 75350 -1160 75370 -1100
rect 75270 -1180 75370 -1160
rect 75100 -1260 75120 -1200
rect 75180 -1260 75200 -1200
rect 75100 -1270 75200 -1260
rect 75440 -1200 75540 -1060
rect 75780 -770 75880 -750
rect 75780 -830 75800 -770
rect 75860 -830 75880 -770
rect 75780 -880 75880 -830
rect 75780 -950 75800 -880
rect 75860 -950 75880 -880
rect 75780 -1000 75880 -950
rect 75780 -1060 75800 -1000
rect 75860 -1060 75880 -1000
rect 75610 -1100 75710 -1080
rect 75610 -1160 75630 -1100
rect 75690 -1160 75710 -1100
rect 75610 -1180 75710 -1160
rect 75440 -1260 75460 -1200
rect 75520 -1260 75540 -1200
rect 75440 -1270 75540 -1260
rect 75780 -1200 75880 -1060
rect 76120 -770 76220 -750
rect 76120 -830 76140 -770
rect 76200 -830 76220 -770
rect 76120 -880 76220 -830
rect 76120 -950 76140 -880
rect 76200 -950 76220 -880
rect 76120 -1000 76220 -950
rect 76120 -1060 76140 -1000
rect 76200 -1060 76220 -1000
rect 75950 -1100 76050 -1080
rect 75950 -1160 75970 -1100
rect 76030 -1160 76050 -1100
rect 75950 -1180 76050 -1160
rect 75780 -1260 75800 -1200
rect 75860 -1260 75880 -1200
rect 75780 -1270 75880 -1260
rect 76120 -1200 76220 -1060
rect 76460 -770 76560 -750
rect 76460 -830 76480 -770
rect 76540 -830 76560 -770
rect 76460 -880 76560 -830
rect 76460 -950 76480 -880
rect 76540 -950 76560 -880
rect 76460 -1000 76560 -950
rect 76460 -1060 76480 -1000
rect 76540 -1060 76560 -1000
rect 76290 -1100 76390 -1080
rect 76290 -1160 76310 -1100
rect 76370 -1160 76390 -1100
rect 76290 -1180 76390 -1160
rect 76120 -1260 76140 -1200
rect 76200 -1260 76220 -1200
rect 76120 -1270 76220 -1260
rect 76460 -1200 76560 -1060
rect 76800 -770 76900 -750
rect 76800 -830 76820 -770
rect 76880 -830 76900 -770
rect 76800 -880 76900 -830
rect 76800 -950 76820 -880
rect 76880 -950 76900 -880
rect 76800 -1000 76900 -950
rect 76800 -1060 76820 -1000
rect 76880 -1060 76900 -1000
rect 76630 -1100 76730 -1080
rect 76630 -1160 76650 -1100
rect 76710 -1160 76730 -1100
rect 76630 -1180 76730 -1160
rect 76460 -1260 76480 -1200
rect 76540 -1260 76560 -1200
rect 76460 -1270 76560 -1260
rect 76800 -1200 76900 -1060
rect 77140 -770 77240 -750
rect 77140 -830 77160 -770
rect 77220 -830 77240 -770
rect 77140 -880 77240 -830
rect 77140 -950 77160 -880
rect 77220 -950 77240 -880
rect 77140 -1000 77240 -950
rect 77140 -1060 77160 -1000
rect 77220 -1060 77240 -1000
rect 76970 -1100 77070 -1080
rect 76970 -1160 76990 -1100
rect 77050 -1160 77070 -1100
rect 76970 -1180 77070 -1160
rect 76800 -1260 76820 -1200
rect 76880 -1260 76900 -1200
rect 76800 -1270 76900 -1260
rect 77140 -1200 77240 -1060
rect 77480 -770 77580 -750
rect 77480 -830 77500 -770
rect 77560 -830 77580 -770
rect 77480 -880 77580 -830
rect 77480 -950 77500 -880
rect 77560 -950 77580 -880
rect 77480 -1000 77580 -950
rect 77480 -1060 77500 -1000
rect 77560 -1060 77580 -1000
rect 77310 -1100 77410 -1080
rect 77310 -1160 77330 -1100
rect 77390 -1160 77410 -1100
rect 77310 -1180 77410 -1160
rect 77140 -1260 77160 -1200
rect 77220 -1260 77240 -1200
rect 77140 -1270 77240 -1260
rect 77480 -1200 77580 -1060
rect 77820 -770 77920 -750
rect 77820 -830 77840 -770
rect 77900 -830 77920 -770
rect 77820 -880 77920 -830
rect 77820 -950 77840 -880
rect 77900 -950 77920 -880
rect 77820 -1000 77920 -950
rect 77820 -1060 77840 -1000
rect 77900 -1060 77920 -1000
rect 77650 -1100 77750 -1080
rect 77650 -1160 77670 -1100
rect 77730 -1160 77750 -1100
rect 77650 -1180 77750 -1160
rect 77480 -1260 77500 -1200
rect 77560 -1260 77580 -1200
rect 77480 -1270 77580 -1260
rect 77820 -1200 77920 -1060
rect 78160 -770 78260 -750
rect 78160 -830 78180 -770
rect 78240 -830 78260 -770
rect 78160 -880 78260 -830
rect 78160 -950 78180 -880
rect 78240 -950 78260 -880
rect 78160 -1000 78260 -950
rect 78160 -1060 78180 -1000
rect 78240 -1060 78260 -1000
rect 77990 -1100 78090 -1080
rect 77990 -1160 78010 -1100
rect 78070 -1160 78090 -1100
rect 77990 -1180 78090 -1160
rect 77820 -1260 77840 -1200
rect 77900 -1260 77920 -1200
rect 77820 -1270 77920 -1260
rect 78160 -1200 78260 -1060
rect 78500 -770 78600 -750
rect 78500 -830 78520 -770
rect 78580 -830 78600 -770
rect 78500 -880 78600 -830
rect 78500 -950 78520 -880
rect 78580 -950 78600 -880
rect 78500 -1000 78600 -950
rect 78500 -1060 78520 -1000
rect 78580 -1060 78600 -1000
rect 78330 -1100 78430 -1080
rect 78330 -1160 78350 -1100
rect 78410 -1160 78430 -1100
rect 78330 -1180 78430 -1160
rect 78160 -1260 78180 -1200
rect 78240 -1260 78260 -1200
rect 78160 -1270 78260 -1260
rect 78500 -1200 78600 -1060
rect 78840 -770 78940 -750
rect 78840 -830 78860 -770
rect 78920 -830 78940 -770
rect 78840 -880 78940 -830
rect 78840 -950 78860 -880
rect 78920 -950 78940 -880
rect 78840 -1000 78940 -950
rect 78840 -1060 78860 -1000
rect 78920 -1060 78940 -1000
rect 78670 -1100 78770 -1080
rect 78670 -1160 78690 -1100
rect 78750 -1160 78770 -1100
rect 78670 -1180 78770 -1160
rect 78500 -1260 78520 -1200
rect 78580 -1260 78600 -1200
rect 78500 -1270 78600 -1260
rect 78840 -1200 78940 -1060
rect 79180 -770 79280 -750
rect 79180 -830 79200 -770
rect 79260 -830 79280 -770
rect 79180 -880 79280 -830
rect 79180 -950 79200 -880
rect 79260 -950 79280 -880
rect 79180 -1000 79280 -950
rect 79180 -1060 79200 -1000
rect 79260 -1060 79280 -1000
rect 79010 -1100 79110 -1080
rect 79010 -1160 79030 -1100
rect 79090 -1160 79110 -1100
rect 79010 -1180 79110 -1160
rect 78840 -1260 78860 -1200
rect 78920 -1260 78940 -1200
rect 78840 -1270 78940 -1260
rect 79180 -1200 79280 -1060
rect 79520 -770 79620 -750
rect 79520 -830 79540 -770
rect 79600 -830 79620 -770
rect 79520 -880 79620 -830
rect 79520 -950 79540 -880
rect 79600 -950 79620 -880
rect 79520 -1000 79620 -950
rect 79520 -1060 79540 -1000
rect 79600 -1060 79620 -1000
rect 79350 -1100 79450 -1080
rect 79350 -1160 79370 -1100
rect 79430 -1160 79450 -1100
rect 79350 -1180 79450 -1160
rect 79180 -1260 79200 -1200
rect 79260 -1260 79280 -1200
rect 79180 -1270 79280 -1260
rect 79520 -1200 79620 -1060
rect 79860 -770 79960 -750
rect 79860 -830 79880 -770
rect 79940 -830 79960 -770
rect 79860 -880 79960 -830
rect 79860 -950 79880 -880
rect 79940 -950 79960 -880
rect 79860 -1000 79960 -950
rect 79860 -1060 79880 -1000
rect 79940 -1060 79960 -1000
rect 79690 -1100 79790 -1080
rect 79690 -1160 79710 -1100
rect 79770 -1160 79790 -1100
rect 79690 -1180 79790 -1160
rect 79520 -1260 79540 -1200
rect 79600 -1260 79620 -1200
rect 79520 -1270 79620 -1260
rect 79860 -1200 79960 -1060
rect 80200 -770 80300 -750
rect 80200 -830 80220 -770
rect 80280 -830 80300 -770
rect 80200 -880 80300 -830
rect 80200 -950 80220 -880
rect 80280 -950 80300 -880
rect 80200 -1000 80300 -950
rect 80200 -1060 80220 -1000
rect 80280 -1060 80300 -1000
rect 80030 -1100 80130 -1080
rect 80030 -1160 80050 -1100
rect 80110 -1160 80130 -1100
rect 80030 -1180 80130 -1160
rect 79860 -1260 79880 -1200
rect 79940 -1260 79960 -1200
rect 79860 -1270 79960 -1260
rect 80200 -1200 80300 -1060
rect 80540 -770 80640 -750
rect 80540 -830 80560 -770
rect 80620 -830 80640 -770
rect 80540 -880 80640 -830
rect 80540 -950 80560 -880
rect 80620 -950 80640 -880
rect 80540 -1000 80640 -950
rect 80540 -1060 80560 -1000
rect 80620 -1060 80640 -1000
rect 80370 -1100 80470 -1080
rect 80370 -1160 80390 -1100
rect 80450 -1160 80470 -1100
rect 80370 -1180 80470 -1160
rect 80200 -1260 80220 -1200
rect 80280 -1260 80300 -1200
rect 80200 -1270 80300 -1260
rect 80540 -1200 80640 -1060
rect 80880 -770 80980 -750
rect 80880 -830 80900 -770
rect 80960 -830 80980 -770
rect 80880 -880 80980 -830
rect 80880 -950 80900 -880
rect 80960 -950 80980 -880
rect 80880 -1000 80980 -950
rect 80880 -1060 80900 -1000
rect 80960 -1060 80980 -1000
rect 80710 -1100 80810 -1080
rect 80710 -1160 80730 -1100
rect 80790 -1160 80810 -1100
rect 80710 -1180 80810 -1160
rect 80540 -1260 80560 -1200
rect 80620 -1260 80640 -1200
rect 80540 -1270 80640 -1260
rect 80880 -1200 80980 -1060
rect 81220 -770 81320 -750
rect 81220 -830 81240 -770
rect 81300 -830 81320 -770
rect 81220 -880 81320 -830
rect 81220 -950 81240 -880
rect 81300 -950 81320 -880
rect 81220 -1000 81320 -950
rect 81220 -1060 81240 -1000
rect 81300 -1060 81320 -1000
rect 81050 -1100 81150 -1080
rect 81050 -1160 81070 -1100
rect 81130 -1160 81150 -1100
rect 81050 -1180 81150 -1160
rect 80880 -1260 80900 -1200
rect 80960 -1260 80980 -1200
rect 80880 -1270 80980 -1260
rect 81220 -1200 81320 -1060
rect 81560 -770 81660 -750
rect 81560 -830 81580 -770
rect 81640 -830 81660 -770
rect 81560 -880 81660 -830
rect 81560 -950 81580 -880
rect 81640 -950 81660 -880
rect 81560 -1000 81660 -950
rect 81560 -1060 81580 -1000
rect 81640 -1060 81660 -1000
rect 81390 -1100 81490 -1080
rect 81390 -1160 81410 -1100
rect 81470 -1160 81490 -1100
rect 81390 -1180 81490 -1160
rect 81220 -1260 81240 -1200
rect 81300 -1260 81320 -1200
rect 81220 -1270 81320 -1260
rect 81560 -1200 81660 -1060
rect 81900 -770 82000 -750
rect 81900 -830 81920 -770
rect 81980 -830 82000 -770
rect 81900 -880 82000 -830
rect 81900 -950 81920 -880
rect 81980 -950 82000 -880
rect 81900 -1000 82000 -950
rect 81900 -1060 81920 -1000
rect 81980 -1060 82000 -1000
rect 81730 -1100 81830 -1080
rect 81730 -1160 81750 -1100
rect 81810 -1160 81830 -1100
rect 81730 -1180 81830 -1160
rect 81560 -1260 81580 -1200
rect 81640 -1260 81660 -1200
rect 81560 -1270 81660 -1260
rect 81900 -1200 82000 -1060
rect 82240 -770 82340 -750
rect 82240 -830 82260 -770
rect 82320 -830 82340 -770
rect 82240 -880 82340 -830
rect 82240 -950 82260 -880
rect 82320 -950 82340 -880
rect 82240 -1000 82340 -950
rect 82240 -1060 82260 -1000
rect 82320 -1060 82340 -1000
rect 82070 -1100 82170 -1080
rect 82070 -1160 82090 -1100
rect 82150 -1160 82170 -1100
rect 82070 -1180 82170 -1160
rect 81900 -1260 81920 -1200
rect 81980 -1260 82000 -1200
rect 81900 -1270 82000 -1260
rect 82240 -1200 82340 -1060
rect 82580 -770 82680 -750
rect 82580 -830 82600 -770
rect 82660 -830 82680 -770
rect 82580 -880 82680 -830
rect 82580 -950 82600 -880
rect 82660 -950 82680 -880
rect 82580 -1000 82680 -950
rect 82580 -1060 82600 -1000
rect 82660 -1060 82680 -1000
rect 82410 -1100 82510 -1080
rect 82410 -1160 82430 -1100
rect 82490 -1160 82510 -1100
rect 82410 -1180 82510 -1160
rect 82240 -1260 82260 -1200
rect 82320 -1260 82340 -1200
rect 82240 -1270 82340 -1260
rect 82580 -1200 82680 -1060
rect 82920 -770 83020 -750
rect 82920 -830 82940 -770
rect 83000 -830 83020 -770
rect 82920 -880 83020 -830
rect 82920 -950 82940 -880
rect 83000 -950 83020 -880
rect 82920 -1000 83020 -950
rect 82920 -1060 82940 -1000
rect 83000 -1060 83020 -1000
rect 82750 -1100 82850 -1080
rect 82750 -1160 82770 -1100
rect 82830 -1160 82850 -1100
rect 82750 -1180 82850 -1160
rect 82580 -1260 82600 -1200
rect 82660 -1260 82680 -1200
rect 82580 -1270 82680 -1260
rect 82920 -1200 83020 -1060
rect 83260 -770 83360 -750
rect 83260 -830 83280 -770
rect 83340 -830 83360 -770
rect 83260 -880 83360 -830
rect 83260 -950 83280 -880
rect 83340 -950 83360 -880
rect 83260 -1000 83360 -950
rect 83260 -1060 83280 -1000
rect 83340 -1060 83360 -1000
rect 83090 -1100 83190 -1080
rect 83090 -1160 83110 -1100
rect 83170 -1160 83190 -1100
rect 83090 -1180 83190 -1160
rect 82920 -1260 82940 -1200
rect 83000 -1260 83020 -1200
rect 82920 -1270 83020 -1260
rect 83260 -1200 83360 -1060
rect 83600 -770 83700 -750
rect 83600 -830 83620 -770
rect 83680 -830 83700 -770
rect 83600 -880 83700 -830
rect 83600 -950 83620 -880
rect 83680 -950 83700 -880
rect 83600 -1000 83700 -950
rect 83600 -1060 83620 -1000
rect 83680 -1060 83700 -1000
rect 83430 -1100 83530 -1080
rect 83430 -1160 83450 -1100
rect 83510 -1160 83530 -1100
rect 83430 -1180 83530 -1160
rect 83260 -1260 83280 -1200
rect 83340 -1260 83360 -1200
rect 83260 -1270 83360 -1260
rect 83600 -1200 83700 -1060
rect 83940 -770 84040 -750
rect 83940 -830 83960 -770
rect 84020 -830 84040 -770
rect 83940 -880 84040 -830
rect 83940 -950 83960 -880
rect 84020 -950 84040 -880
rect 83940 -1000 84040 -950
rect 83940 -1060 83960 -1000
rect 84020 -1060 84040 -1000
rect 83770 -1100 83870 -1080
rect 83770 -1160 83790 -1100
rect 83850 -1160 83870 -1100
rect 83770 -1180 83870 -1160
rect 83600 -1260 83620 -1200
rect 83680 -1260 83700 -1200
rect 83600 -1270 83700 -1260
rect 83940 -1200 84040 -1060
rect 84280 -770 84380 -750
rect 84280 -830 84300 -770
rect 84360 -830 84380 -770
rect 84280 -880 84380 -830
rect 84280 -950 84300 -880
rect 84360 -950 84380 -880
rect 84280 -1000 84380 -950
rect 84280 -1060 84300 -1000
rect 84360 -1060 84380 -1000
rect 84110 -1100 84210 -1080
rect 84110 -1160 84130 -1100
rect 84190 -1160 84210 -1100
rect 84110 -1180 84210 -1160
rect 83940 -1260 83960 -1200
rect 84020 -1260 84040 -1200
rect 83940 -1270 84040 -1260
rect 84280 -1200 84380 -1060
rect 84620 -770 84720 -750
rect 84620 -830 84640 -770
rect 84700 -830 84720 -770
rect 84620 -880 84720 -830
rect 84620 -950 84640 -880
rect 84700 -950 84720 -880
rect 84620 -1000 84720 -950
rect 84620 -1060 84640 -1000
rect 84700 -1060 84720 -1000
rect 84450 -1100 84550 -1080
rect 84450 -1160 84470 -1100
rect 84530 -1160 84550 -1100
rect 84450 -1180 84550 -1160
rect 84280 -1260 84300 -1200
rect 84360 -1260 84380 -1200
rect 84280 -1270 84380 -1260
rect 84620 -1200 84720 -1060
rect 84960 -770 85060 -750
rect 84960 -830 84980 -770
rect 85040 -830 85060 -770
rect 84960 -880 85060 -830
rect 84960 -950 84980 -880
rect 85040 -950 85060 -880
rect 84960 -1000 85060 -950
rect 84960 -1060 84980 -1000
rect 85040 -1060 85060 -1000
rect 84790 -1100 84890 -1080
rect 84790 -1160 84810 -1100
rect 84870 -1160 84890 -1100
rect 84790 -1180 84890 -1160
rect 84620 -1260 84640 -1200
rect 84700 -1260 84720 -1200
rect 84620 -1270 84720 -1260
rect 84960 -1200 85060 -1060
rect 85300 -770 85400 -750
rect 85300 -830 85320 -770
rect 85380 -830 85400 -770
rect 85300 -880 85400 -830
rect 85300 -950 85320 -880
rect 85380 -950 85400 -880
rect 85300 -1000 85400 -950
rect 85300 -1060 85320 -1000
rect 85380 -1060 85400 -1000
rect 85130 -1100 85230 -1080
rect 85130 -1160 85150 -1100
rect 85210 -1160 85230 -1100
rect 85130 -1180 85230 -1160
rect 84960 -1260 84980 -1200
rect 85040 -1260 85060 -1200
rect 84960 -1270 85060 -1260
rect 85300 -1200 85400 -1060
rect 85640 -770 85740 -750
rect 85640 -830 85660 -770
rect 85720 -830 85740 -770
rect 85640 -880 85740 -830
rect 85640 -950 85660 -880
rect 85720 -950 85740 -880
rect 85640 -1000 85740 -950
rect 85640 -1060 85660 -1000
rect 85720 -1060 85740 -1000
rect 85470 -1100 85570 -1080
rect 85470 -1160 85490 -1100
rect 85550 -1160 85570 -1100
rect 85470 -1180 85570 -1160
rect 85300 -1260 85320 -1200
rect 85380 -1260 85400 -1200
rect 85300 -1270 85400 -1260
rect 85640 -1200 85740 -1060
rect 85980 -770 86080 -750
rect 85980 -830 86000 -770
rect 86060 -830 86080 -770
rect 85980 -880 86080 -830
rect 85980 -950 86000 -880
rect 86060 -950 86080 -880
rect 85980 -1000 86080 -950
rect 85980 -1060 86000 -1000
rect 86060 -1060 86080 -1000
rect 85810 -1100 85910 -1080
rect 85810 -1160 85830 -1100
rect 85890 -1160 85910 -1100
rect 85810 -1180 85910 -1160
rect 85640 -1260 85660 -1200
rect 85720 -1260 85740 -1200
rect 85640 -1270 85740 -1260
rect 85980 -1200 86080 -1060
rect 86320 -770 86420 -750
rect 86320 -830 86340 -770
rect 86400 -830 86420 -770
rect 86320 -880 86420 -830
rect 86320 -950 86340 -880
rect 86400 -950 86420 -880
rect 86320 -1000 86420 -950
rect 86320 -1060 86340 -1000
rect 86400 -1060 86420 -1000
rect 86150 -1100 86250 -1080
rect 86150 -1160 86170 -1100
rect 86230 -1160 86250 -1100
rect 86150 -1180 86250 -1160
rect 85980 -1260 86000 -1200
rect 86060 -1260 86080 -1200
rect 85980 -1270 86080 -1260
rect 86320 -1200 86420 -1060
rect 86660 -770 86760 -750
rect 86660 -830 86680 -770
rect 86740 -830 86760 -770
rect 86660 -880 86760 -830
rect 86660 -950 86680 -880
rect 86740 -950 86760 -880
rect 86660 -1000 86760 -950
rect 86660 -1060 86680 -1000
rect 86740 -1060 86760 -1000
rect 86490 -1100 86590 -1080
rect 86490 -1160 86510 -1100
rect 86570 -1160 86590 -1100
rect 86490 -1180 86590 -1160
rect 86320 -1260 86340 -1200
rect 86400 -1260 86420 -1200
rect 86320 -1270 86420 -1260
rect 86660 -1200 86760 -1060
rect 87000 -770 87100 -750
rect 87000 -830 87020 -770
rect 87080 -830 87100 -770
rect 87000 -880 87100 -830
rect 87000 -950 87020 -880
rect 87080 -950 87100 -880
rect 87000 -1000 87100 -950
rect 87000 -1060 87020 -1000
rect 87080 -1060 87100 -1000
rect 86830 -1100 86930 -1080
rect 86830 -1160 86850 -1100
rect 86910 -1160 86930 -1100
rect 86830 -1180 86930 -1160
rect 86660 -1260 86680 -1200
rect 86740 -1260 86760 -1200
rect 86660 -1270 86760 -1260
rect 87000 -1200 87100 -1060
rect 87170 -1100 87270 -1080
rect 87170 -1160 87190 -1100
rect 87250 -1160 87270 -1100
rect 87170 -1180 87270 -1160
rect 87000 -1260 87020 -1200
rect 87080 -1260 87100 -1200
rect 87000 -1270 87100 -1260
rect 130 -1300 230 -1280
rect 130 -1360 150 -1300
rect 210 -1360 230 -1300
rect 130 -1380 230 -1360
rect 470 -1300 570 -1280
rect 470 -1360 490 -1300
rect 550 -1360 570 -1300
rect 470 -1380 570 -1360
rect 810 -1300 910 -1280
rect 810 -1360 830 -1300
rect 890 -1360 910 -1300
rect 810 -1380 910 -1360
rect 1150 -1300 1250 -1280
rect 1150 -1360 1170 -1300
rect 1230 -1360 1250 -1300
rect 1150 -1380 1250 -1360
rect 1490 -1300 1590 -1280
rect 1490 -1360 1510 -1300
rect 1570 -1360 1590 -1300
rect 1490 -1380 1590 -1360
rect 1830 -1300 1930 -1280
rect 1830 -1360 1850 -1300
rect 1910 -1360 1930 -1300
rect 1830 -1380 1930 -1360
rect 2170 -1300 2270 -1280
rect 2170 -1360 2190 -1300
rect 2250 -1360 2270 -1300
rect 2170 -1380 2270 -1360
rect 2510 -1300 2610 -1280
rect 2510 -1360 2530 -1300
rect 2590 -1360 2610 -1300
rect 2510 -1380 2610 -1360
rect 2850 -1300 2950 -1280
rect 2850 -1360 2870 -1300
rect 2930 -1360 2950 -1300
rect 2850 -1380 2950 -1360
rect 3190 -1300 3290 -1280
rect 3190 -1360 3210 -1300
rect 3270 -1360 3290 -1300
rect 3190 -1380 3290 -1360
rect 3530 -1300 3630 -1280
rect 3530 -1360 3550 -1300
rect 3610 -1360 3630 -1300
rect 3530 -1380 3630 -1360
rect 3870 -1300 3970 -1280
rect 3870 -1360 3890 -1300
rect 3950 -1360 3970 -1300
rect 3870 -1380 3970 -1360
rect 4210 -1300 4310 -1280
rect 4210 -1360 4230 -1300
rect 4290 -1360 4310 -1300
rect 4210 -1380 4310 -1360
rect 4550 -1300 4650 -1280
rect 4550 -1360 4570 -1300
rect 4630 -1360 4650 -1300
rect 4550 -1380 4650 -1360
rect 4890 -1300 4990 -1280
rect 4890 -1360 4910 -1300
rect 4970 -1360 4990 -1300
rect 4890 -1380 4990 -1360
rect 5230 -1300 5330 -1280
rect 5230 -1360 5250 -1300
rect 5310 -1360 5330 -1300
rect 5230 -1380 5330 -1360
rect 5570 -1300 5670 -1280
rect 5570 -1360 5590 -1300
rect 5650 -1360 5670 -1300
rect 5570 -1380 5670 -1360
rect 5910 -1300 6010 -1280
rect 5910 -1360 5930 -1300
rect 5990 -1360 6010 -1300
rect 5910 -1380 6010 -1360
rect 6250 -1300 6350 -1280
rect 6250 -1360 6270 -1300
rect 6330 -1360 6350 -1300
rect 6250 -1380 6350 -1360
rect 6590 -1300 6690 -1280
rect 6590 -1360 6610 -1300
rect 6670 -1360 6690 -1300
rect 6590 -1380 6690 -1360
rect 6930 -1300 7030 -1280
rect 6930 -1360 6950 -1300
rect 7010 -1360 7030 -1300
rect 6930 -1380 7030 -1360
rect 7270 -1300 7370 -1280
rect 7270 -1360 7290 -1300
rect 7350 -1360 7370 -1300
rect 7270 -1380 7370 -1360
rect 7610 -1300 7710 -1280
rect 7610 -1360 7630 -1300
rect 7690 -1360 7710 -1300
rect 7610 -1380 7710 -1360
rect 7950 -1300 8050 -1280
rect 7950 -1360 7970 -1300
rect 8030 -1360 8050 -1300
rect 7950 -1380 8050 -1360
rect 8290 -1300 8390 -1280
rect 8290 -1360 8310 -1300
rect 8370 -1360 8390 -1300
rect 8290 -1380 8390 -1360
rect 8630 -1300 8730 -1280
rect 8630 -1360 8650 -1300
rect 8710 -1360 8730 -1300
rect 8630 -1380 8730 -1360
rect 8970 -1300 9070 -1280
rect 8970 -1360 8990 -1300
rect 9050 -1360 9070 -1300
rect 8970 -1380 9070 -1360
rect 9310 -1300 9410 -1280
rect 9310 -1360 9330 -1300
rect 9390 -1360 9410 -1300
rect 9310 -1380 9410 -1360
rect 9650 -1300 9750 -1280
rect 9650 -1360 9670 -1300
rect 9730 -1360 9750 -1300
rect 9650 -1380 9750 -1360
rect 9990 -1300 10090 -1280
rect 9990 -1360 10010 -1300
rect 10070 -1360 10090 -1300
rect 9990 -1380 10090 -1360
rect 10330 -1300 10430 -1280
rect 10330 -1360 10350 -1300
rect 10410 -1360 10430 -1300
rect 10330 -1380 10430 -1360
rect 10670 -1300 10770 -1280
rect 10670 -1360 10690 -1300
rect 10750 -1360 10770 -1300
rect 10670 -1380 10770 -1360
rect 11010 -1300 11110 -1280
rect 11010 -1360 11030 -1300
rect 11090 -1360 11110 -1300
rect 11010 -1380 11110 -1360
rect 11350 -1300 11450 -1280
rect 11350 -1360 11370 -1300
rect 11430 -1360 11450 -1300
rect 11350 -1380 11450 -1360
rect 11690 -1300 11790 -1280
rect 11690 -1360 11710 -1300
rect 11770 -1360 11790 -1300
rect 11690 -1380 11790 -1360
rect 12030 -1300 12130 -1280
rect 12030 -1360 12050 -1300
rect 12110 -1360 12130 -1300
rect 12030 -1380 12130 -1360
rect 12370 -1300 12470 -1280
rect 12370 -1360 12390 -1300
rect 12450 -1360 12470 -1300
rect 12370 -1380 12470 -1360
rect 12710 -1300 12810 -1280
rect 12710 -1360 12730 -1300
rect 12790 -1360 12810 -1300
rect 12710 -1380 12810 -1360
rect 13050 -1300 13150 -1280
rect 13050 -1360 13070 -1300
rect 13130 -1360 13150 -1300
rect 13050 -1380 13150 -1360
rect 13390 -1300 13490 -1280
rect 13390 -1360 13410 -1300
rect 13470 -1360 13490 -1300
rect 13390 -1380 13490 -1360
rect 13730 -1300 13830 -1280
rect 13730 -1360 13750 -1300
rect 13810 -1360 13830 -1300
rect 13730 -1380 13830 -1360
rect 14070 -1300 14170 -1280
rect 14070 -1360 14090 -1300
rect 14150 -1360 14170 -1300
rect 14070 -1380 14170 -1360
rect 14410 -1300 14510 -1280
rect 14410 -1360 14430 -1300
rect 14490 -1360 14510 -1300
rect 14410 -1380 14510 -1360
rect 14750 -1300 14850 -1280
rect 14750 -1360 14770 -1300
rect 14830 -1360 14850 -1300
rect 14750 -1380 14850 -1360
rect 15090 -1300 15190 -1280
rect 15090 -1360 15110 -1300
rect 15170 -1360 15190 -1300
rect 15090 -1380 15190 -1360
rect 15430 -1300 15530 -1280
rect 15430 -1360 15450 -1300
rect 15510 -1360 15530 -1300
rect 15430 -1380 15530 -1360
rect 15770 -1300 15870 -1280
rect 15770 -1360 15790 -1300
rect 15850 -1360 15870 -1300
rect 15770 -1380 15870 -1360
rect 16110 -1300 16210 -1280
rect 16110 -1360 16130 -1300
rect 16190 -1360 16210 -1300
rect 16110 -1380 16210 -1360
rect 16450 -1300 16550 -1280
rect 16450 -1360 16470 -1300
rect 16530 -1360 16550 -1300
rect 16450 -1380 16550 -1360
rect 16790 -1300 16890 -1280
rect 16790 -1360 16810 -1300
rect 16870 -1360 16890 -1300
rect 16790 -1380 16890 -1360
rect 17130 -1300 17230 -1280
rect 17130 -1360 17150 -1300
rect 17210 -1360 17230 -1300
rect 17130 -1380 17230 -1360
rect 17470 -1300 17570 -1280
rect 17470 -1360 17490 -1300
rect 17550 -1360 17570 -1300
rect 17470 -1380 17570 -1360
rect 17810 -1300 17910 -1280
rect 17810 -1360 17830 -1300
rect 17890 -1360 17910 -1300
rect 17810 -1380 17910 -1360
rect 18150 -1300 18250 -1280
rect 18150 -1360 18170 -1300
rect 18230 -1360 18250 -1300
rect 18150 -1380 18250 -1360
rect 18490 -1300 18590 -1280
rect 18490 -1360 18510 -1300
rect 18570 -1360 18590 -1300
rect 18490 -1380 18590 -1360
rect 18830 -1300 18930 -1280
rect 18830 -1360 18850 -1300
rect 18910 -1360 18930 -1300
rect 18830 -1380 18930 -1360
rect 19170 -1300 19270 -1280
rect 19170 -1360 19190 -1300
rect 19250 -1360 19270 -1300
rect 19170 -1380 19270 -1360
rect 19510 -1300 19610 -1280
rect 19510 -1360 19530 -1300
rect 19590 -1360 19610 -1300
rect 19510 -1380 19610 -1360
rect 19850 -1300 19950 -1280
rect 19850 -1360 19870 -1300
rect 19930 -1360 19950 -1300
rect 19850 -1380 19950 -1360
rect 20190 -1300 20290 -1280
rect 20190 -1360 20210 -1300
rect 20270 -1360 20290 -1300
rect 20190 -1380 20290 -1360
rect 20530 -1300 20630 -1280
rect 20530 -1360 20550 -1300
rect 20610 -1360 20630 -1300
rect 20530 -1380 20630 -1360
rect 20870 -1300 20970 -1280
rect 20870 -1360 20890 -1300
rect 20950 -1360 20970 -1300
rect 20870 -1380 20970 -1360
rect 21210 -1300 21310 -1280
rect 21210 -1360 21230 -1300
rect 21290 -1360 21310 -1300
rect 21210 -1380 21310 -1360
rect 21550 -1300 21650 -1280
rect 21550 -1360 21570 -1300
rect 21630 -1360 21650 -1300
rect 21550 -1380 21650 -1360
rect 21890 -1300 21990 -1280
rect 21890 -1360 21910 -1300
rect 21970 -1360 21990 -1300
rect 21890 -1380 21990 -1360
rect 22230 -1300 22330 -1280
rect 22230 -1360 22250 -1300
rect 22310 -1360 22330 -1300
rect 22230 -1380 22330 -1360
rect 22570 -1300 22670 -1280
rect 22570 -1360 22590 -1300
rect 22650 -1360 22670 -1300
rect 22570 -1380 22670 -1360
rect 22910 -1300 23010 -1280
rect 22910 -1360 22930 -1300
rect 22990 -1360 23010 -1300
rect 22910 -1380 23010 -1360
rect 23250 -1300 23350 -1280
rect 23250 -1360 23270 -1300
rect 23330 -1360 23350 -1300
rect 23250 -1380 23350 -1360
rect 23590 -1300 23690 -1280
rect 23590 -1360 23610 -1300
rect 23670 -1360 23690 -1300
rect 23590 -1380 23690 -1360
rect 23930 -1300 24030 -1280
rect 23930 -1360 23950 -1300
rect 24010 -1360 24030 -1300
rect 23930 -1380 24030 -1360
rect 24270 -1300 24370 -1280
rect 24270 -1360 24290 -1300
rect 24350 -1360 24370 -1300
rect 24270 -1380 24370 -1360
rect 24610 -1300 24710 -1280
rect 24610 -1360 24630 -1300
rect 24690 -1360 24710 -1300
rect 24610 -1380 24710 -1360
rect 24950 -1300 25050 -1280
rect 24950 -1360 24970 -1300
rect 25030 -1360 25050 -1300
rect 24950 -1380 25050 -1360
rect 25290 -1300 25390 -1280
rect 25290 -1360 25310 -1300
rect 25370 -1360 25390 -1300
rect 25290 -1380 25390 -1360
rect 25630 -1300 25730 -1280
rect 25630 -1360 25650 -1300
rect 25710 -1360 25730 -1300
rect 25630 -1380 25730 -1360
rect 25970 -1300 26070 -1280
rect 25970 -1360 25990 -1300
rect 26050 -1360 26070 -1300
rect 25970 -1380 26070 -1360
rect 26310 -1300 26410 -1280
rect 26310 -1360 26330 -1300
rect 26390 -1360 26410 -1300
rect 26310 -1380 26410 -1360
rect 26650 -1300 26750 -1280
rect 26650 -1360 26670 -1300
rect 26730 -1360 26750 -1300
rect 26650 -1380 26750 -1360
rect 26990 -1300 27090 -1280
rect 26990 -1360 27010 -1300
rect 27070 -1360 27090 -1300
rect 26990 -1380 27090 -1360
rect 27330 -1300 27430 -1280
rect 27330 -1360 27350 -1300
rect 27410 -1360 27430 -1300
rect 27330 -1380 27430 -1360
rect 27670 -1300 27770 -1280
rect 27670 -1360 27690 -1300
rect 27750 -1360 27770 -1300
rect 27670 -1380 27770 -1360
rect 28010 -1300 28110 -1280
rect 28010 -1360 28030 -1300
rect 28090 -1360 28110 -1300
rect 28010 -1380 28110 -1360
rect 28350 -1300 28450 -1280
rect 28350 -1360 28370 -1300
rect 28430 -1360 28450 -1300
rect 28350 -1380 28450 -1360
rect 28690 -1300 28790 -1280
rect 28690 -1360 28710 -1300
rect 28770 -1360 28790 -1300
rect 28690 -1380 28790 -1360
rect 29030 -1300 29130 -1280
rect 29030 -1360 29050 -1300
rect 29110 -1360 29130 -1300
rect 29030 -1380 29130 -1360
rect 29370 -1300 29470 -1280
rect 29370 -1360 29390 -1300
rect 29450 -1360 29470 -1300
rect 29370 -1380 29470 -1360
rect 29710 -1300 29810 -1280
rect 29710 -1360 29730 -1300
rect 29790 -1360 29810 -1300
rect 29710 -1380 29810 -1360
rect 30050 -1300 30150 -1280
rect 30050 -1360 30070 -1300
rect 30130 -1360 30150 -1300
rect 30050 -1380 30150 -1360
rect 30390 -1300 30490 -1280
rect 30390 -1360 30410 -1300
rect 30470 -1360 30490 -1300
rect 30390 -1380 30490 -1360
rect 30730 -1300 30830 -1280
rect 30730 -1360 30750 -1300
rect 30810 -1360 30830 -1300
rect 30730 -1380 30830 -1360
rect 31070 -1300 31170 -1280
rect 31070 -1360 31090 -1300
rect 31150 -1360 31170 -1300
rect 31070 -1380 31170 -1360
rect 31410 -1300 31510 -1280
rect 31410 -1360 31430 -1300
rect 31490 -1360 31510 -1300
rect 31410 -1380 31510 -1360
rect 31750 -1300 31850 -1280
rect 31750 -1360 31770 -1300
rect 31830 -1360 31850 -1300
rect 31750 -1380 31850 -1360
rect 32090 -1300 32190 -1280
rect 32090 -1360 32110 -1300
rect 32170 -1360 32190 -1300
rect 32090 -1380 32190 -1360
rect 32430 -1300 32530 -1280
rect 32430 -1360 32450 -1300
rect 32510 -1360 32530 -1300
rect 32430 -1380 32530 -1360
rect 32770 -1300 32870 -1280
rect 32770 -1360 32790 -1300
rect 32850 -1360 32870 -1300
rect 32770 -1380 32870 -1360
rect 33110 -1300 33210 -1280
rect 33110 -1360 33130 -1300
rect 33190 -1360 33210 -1300
rect 33110 -1380 33210 -1360
rect 33450 -1300 33550 -1280
rect 33450 -1360 33470 -1300
rect 33530 -1360 33550 -1300
rect 33450 -1380 33550 -1360
rect 33790 -1300 33890 -1280
rect 33790 -1360 33810 -1300
rect 33870 -1360 33890 -1300
rect 33790 -1380 33890 -1360
rect 34130 -1300 34230 -1280
rect 34130 -1360 34150 -1300
rect 34210 -1360 34230 -1300
rect 34130 -1380 34230 -1360
rect 34470 -1300 34570 -1280
rect 34470 -1360 34490 -1300
rect 34550 -1360 34570 -1300
rect 34470 -1380 34570 -1360
rect 34810 -1300 34910 -1280
rect 34810 -1360 34830 -1300
rect 34890 -1360 34910 -1300
rect 34810 -1380 34910 -1360
rect 35150 -1300 35250 -1280
rect 35150 -1360 35170 -1300
rect 35230 -1360 35250 -1300
rect 35150 -1380 35250 -1360
rect 35490 -1300 35590 -1280
rect 35490 -1360 35510 -1300
rect 35570 -1360 35590 -1300
rect 35490 -1380 35590 -1360
rect 35830 -1300 35930 -1280
rect 35830 -1360 35850 -1300
rect 35910 -1360 35930 -1300
rect 35830 -1380 35930 -1360
rect 36170 -1300 36270 -1280
rect 36170 -1360 36190 -1300
rect 36250 -1360 36270 -1300
rect 36170 -1380 36270 -1360
rect 36510 -1300 36610 -1280
rect 36510 -1360 36530 -1300
rect 36590 -1360 36610 -1300
rect 36510 -1380 36610 -1360
rect 36850 -1300 36950 -1280
rect 36850 -1360 36870 -1300
rect 36930 -1360 36950 -1300
rect 36850 -1380 36950 -1360
rect 37190 -1300 37290 -1280
rect 37190 -1360 37210 -1300
rect 37270 -1360 37290 -1300
rect 37190 -1380 37290 -1360
rect 37530 -1300 37630 -1280
rect 37530 -1360 37550 -1300
rect 37610 -1360 37630 -1300
rect 37530 -1380 37630 -1360
rect 37870 -1300 37970 -1280
rect 37870 -1360 37890 -1300
rect 37950 -1360 37970 -1300
rect 37870 -1380 37970 -1360
rect 38210 -1300 38310 -1280
rect 38210 -1360 38230 -1300
rect 38290 -1360 38310 -1300
rect 38210 -1380 38310 -1360
rect 38550 -1300 38650 -1280
rect 38550 -1360 38570 -1300
rect 38630 -1360 38650 -1300
rect 38550 -1380 38650 -1360
rect 38890 -1300 38990 -1280
rect 38890 -1360 38910 -1300
rect 38970 -1360 38990 -1300
rect 38890 -1380 38990 -1360
rect 39230 -1300 39330 -1280
rect 39230 -1360 39250 -1300
rect 39310 -1360 39330 -1300
rect 39230 -1380 39330 -1360
rect 39570 -1300 39670 -1280
rect 39570 -1360 39590 -1300
rect 39650 -1360 39670 -1300
rect 39570 -1380 39670 -1360
rect 39910 -1300 40010 -1280
rect 39910 -1360 39930 -1300
rect 39990 -1360 40010 -1300
rect 39910 -1380 40010 -1360
rect 40250 -1300 40350 -1280
rect 40250 -1360 40270 -1300
rect 40330 -1360 40350 -1300
rect 40250 -1380 40350 -1360
rect 40590 -1300 40690 -1280
rect 40590 -1360 40610 -1300
rect 40670 -1360 40690 -1300
rect 40590 -1380 40690 -1360
rect 40930 -1300 41030 -1280
rect 40930 -1360 40950 -1300
rect 41010 -1360 41030 -1300
rect 40930 -1380 41030 -1360
rect 41270 -1300 41370 -1280
rect 41270 -1360 41290 -1300
rect 41350 -1360 41370 -1300
rect 41270 -1380 41370 -1360
rect 41610 -1300 41710 -1280
rect 41610 -1360 41630 -1300
rect 41690 -1360 41710 -1300
rect 41610 -1380 41710 -1360
rect 41950 -1300 42050 -1280
rect 41950 -1360 41970 -1300
rect 42030 -1360 42050 -1300
rect 41950 -1380 42050 -1360
rect 42290 -1300 42390 -1280
rect 42290 -1360 42310 -1300
rect 42370 -1360 42390 -1300
rect 42290 -1380 42390 -1360
rect 42630 -1300 42730 -1280
rect 42630 -1360 42650 -1300
rect 42710 -1360 42730 -1300
rect 42630 -1380 42730 -1360
rect 42970 -1300 43070 -1280
rect 42970 -1360 42990 -1300
rect 43050 -1360 43070 -1300
rect 42970 -1380 43070 -1360
rect 43310 -1300 43410 -1280
rect 43310 -1360 43330 -1300
rect 43390 -1360 43410 -1300
rect 43310 -1380 43410 -1360
rect 43650 -1300 43750 -1280
rect 43650 -1360 43670 -1300
rect 43730 -1360 43750 -1300
rect 43650 -1380 43750 -1360
rect 43990 -1300 44090 -1280
rect 43990 -1360 44010 -1300
rect 44070 -1360 44090 -1300
rect 43990 -1380 44090 -1360
rect 44330 -1300 44430 -1280
rect 44330 -1360 44350 -1300
rect 44410 -1360 44430 -1300
rect 44330 -1380 44430 -1360
rect 44670 -1300 44770 -1280
rect 44670 -1360 44690 -1300
rect 44750 -1360 44770 -1300
rect 44670 -1380 44770 -1360
rect 45010 -1300 45110 -1280
rect 45010 -1360 45030 -1300
rect 45090 -1360 45110 -1300
rect 45010 -1380 45110 -1360
rect 45350 -1300 45450 -1280
rect 45350 -1360 45370 -1300
rect 45430 -1360 45450 -1300
rect 45350 -1380 45450 -1360
rect 45690 -1300 45790 -1280
rect 45690 -1360 45710 -1300
rect 45770 -1360 45790 -1300
rect 45690 -1380 45790 -1360
rect 46030 -1300 46130 -1280
rect 46030 -1360 46050 -1300
rect 46110 -1360 46130 -1300
rect 46030 -1380 46130 -1360
rect 46370 -1300 46470 -1280
rect 46370 -1360 46390 -1300
rect 46450 -1360 46470 -1300
rect 46370 -1380 46470 -1360
rect 46710 -1300 46810 -1280
rect 46710 -1360 46730 -1300
rect 46790 -1360 46810 -1300
rect 46710 -1380 46810 -1360
rect 47050 -1300 47150 -1280
rect 47050 -1360 47070 -1300
rect 47130 -1360 47150 -1300
rect 47050 -1380 47150 -1360
rect 47390 -1300 47490 -1280
rect 47390 -1360 47410 -1300
rect 47470 -1360 47490 -1300
rect 47390 -1380 47490 -1360
rect 47730 -1300 47830 -1280
rect 47730 -1360 47750 -1300
rect 47810 -1360 47830 -1300
rect 47730 -1380 47830 -1360
rect 48070 -1300 48170 -1280
rect 48070 -1360 48090 -1300
rect 48150 -1360 48170 -1300
rect 48070 -1380 48170 -1360
rect 48410 -1300 48510 -1280
rect 48410 -1360 48430 -1300
rect 48490 -1360 48510 -1300
rect 48410 -1380 48510 -1360
rect 48750 -1300 48850 -1280
rect 48750 -1360 48770 -1300
rect 48830 -1360 48850 -1300
rect 48750 -1380 48850 -1360
rect 49090 -1300 49190 -1280
rect 49090 -1360 49110 -1300
rect 49170 -1360 49190 -1300
rect 49090 -1380 49190 -1360
rect 49430 -1300 49530 -1280
rect 49430 -1360 49450 -1300
rect 49510 -1360 49530 -1300
rect 49430 -1380 49530 -1360
rect 49770 -1300 49870 -1280
rect 49770 -1360 49790 -1300
rect 49850 -1360 49870 -1300
rect 49770 -1380 49870 -1360
rect 50110 -1300 50210 -1280
rect 50110 -1360 50130 -1300
rect 50190 -1360 50210 -1300
rect 50110 -1380 50210 -1360
rect 50450 -1300 50550 -1280
rect 50450 -1360 50470 -1300
rect 50530 -1360 50550 -1300
rect 50450 -1380 50550 -1360
rect 50790 -1300 50890 -1280
rect 50790 -1360 50810 -1300
rect 50870 -1360 50890 -1300
rect 50790 -1380 50890 -1360
rect 51130 -1300 51230 -1280
rect 51130 -1360 51150 -1300
rect 51210 -1360 51230 -1300
rect 51130 -1380 51230 -1360
rect 51470 -1300 51570 -1280
rect 51470 -1360 51490 -1300
rect 51550 -1360 51570 -1300
rect 51470 -1380 51570 -1360
rect 51810 -1300 51910 -1280
rect 51810 -1360 51830 -1300
rect 51890 -1360 51910 -1300
rect 51810 -1380 51910 -1360
rect 52150 -1300 52250 -1280
rect 52150 -1360 52170 -1300
rect 52230 -1360 52250 -1300
rect 52150 -1380 52250 -1360
rect 52490 -1300 52590 -1280
rect 52490 -1360 52510 -1300
rect 52570 -1360 52590 -1300
rect 52490 -1380 52590 -1360
rect 52830 -1300 52930 -1280
rect 52830 -1360 52850 -1300
rect 52910 -1360 52930 -1300
rect 52830 -1380 52930 -1360
rect 53170 -1300 53270 -1280
rect 53170 -1360 53190 -1300
rect 53250 -1360 53270 -1300
rect 53170 -1380 53270 -1360
rect 53510 -1300 53610 -1280
rect 53510 -1360 53530 -1300
rect 53590 -1360 53610 -1300
rect 53510 -1380 53610 -1360
rect 53850 -1300 53950 -1280
rect 53850 -1360 53870 -1300
rect 53930 -1360 53950 -1300
rect 53850 -1380 53950 -1360
rect 54190 -1300 54290 -1280
rect 54190 -1360 54210 -1300
rect 54270 -1360 54290 -1300
rect 54190 -1380 54290 -1360
rect 54530 -1300 54630 -1280
rect 54530 -1360 54550 -1300
rect 54610 -1360 54630 -1300
rect 54530 -1380 54630 -1360
rect 54870 -1300 54970 -1280
rect 54870 -1360 54890 -1300
rect 54950 -1360 54970 -1300
rect 54870 -1380 54970 -1360
rect 55210 -1300 55310 -1280
rect 55210 -1360 55230 -1300
rect 55290 -1360 55310 -1300
rect 55210 -1380 55310 -1360
rect 55550 -1300 55650 -1280
rect 55550 -1360 55570 -1300
rect 55630 -1360 55650 -1300
rect 55550 -1380 55650 -1360
rect 55890 -1300 55990 -1280
rect 55890 -1360 55910 -1300
rect 55970 -1360 55990 -1300
rect 55890 -1380 55990 -1360
rect 56230 -1300 56330 -1280
rect 56230 -1360 56250 -1300
rect 56310 -1360 56330 -1300
rect 56230 -1380 56330 -1360
rect 56570 -1300 56670 -1280
rect 56570 -1360 56590 -1300
rect 56650 -1360 56670 -1300
rect 56570 -1380 56670 -1360
rect 56910 -1300 57010 -1280
rect 56910 -1360 56930 -1300
rect 56990 -1360 57010 -1300
rect 56910 -1380 57010 -1360
rect 57250 -1300 57350 -1280
rect 57250 -1360 57270 -1300
rect 57330 -1360 57350 -1300
rect 57250 -1380 57350 -1360
rect 57590 -1300 57690 -1280
rect 57590 -1360 57610 -1300
rect 57670 -1360 57690 -1300
rect 57590 -1380 57690 -1360
rect 57930 -1300 58030 -1280
rect 57930 -1360 57950 -1300
rect 58010 -1360 58030 -1300
rect 57930 -1380 58030 -1360
rect 58270 -1300 58370 -1280
rect 58270 -1360 58290 -1300
rect 58350 -1360 58370 -1300
rect 58270 -1380 58370 -1360
rect 58610 -1300 58710 -1280
rect 58610 -1360 58630 -1300
rect 58690 -1360 58710 -1300
rect 58610 -1380 58710 -1360
rect 58950 -1300 59050 -1280
rect 58950 -1360 58970 -1300
rect 59030 -1360 59050 -1300
rect 58950 -1380 59050 -1360
rect 59290 -1300 59390 -1280
rect 59290 -1360 59310 -1300
rect 59370 -1360 59390 -1300
rect 59290 -1380 59390 -1360
rect 59630 -1300 59730 -1280
rect 59630 -1360 59650 -1300
rect 59710 -1360 59730 -1300
rect 59630 -1380 59730 -1360
rect 59970 -1300 60070 -1280
rect 59970 -1360 59990 -1300
rect 60050 -1360 60070 -1300
rect 59970 -1380 60070 -1360
rect 60310 -1300 60410 -1280
rect 60310 -1360 60330 -1300
rect 60390 -1360 60410 -1300
rect 60310 -1380 60410 -1360
rect 60650 -1300 60750 -1280
rect 60650 -1360 60670 -1300
rect 60730 -1360 60750 -1300
rect 60650 -1380 60750 -1360
rect 60990 -1300 61090 -1280
rect 60990 -1360 61010 -1300
rect 61070 -1360 61090 -1300
rect 60990 -1380 61090 -1360
rect 61330 -1300 61430 -1280
rect 61330 -1360 61350 -1300
rect 61410 -1360 61430 -1300
rect 61330 -1380 61430 -1360
rect 61670 -1300 61770 -1280
rect 61670 -1360 61690 -1300
rect 61750 -1360 61770 -1300
rect 61670 -1380 61770 -1360
rect 62010 -1300 62110 -1280
rect 62010 -1360 62030 -1300
rect 62090 -1360 62110 -1300
rect 62010 -1380 62110 -1360
rect 62350 -1300 62450 -1280
rect 62350 -1360 62370 -1300
rect 62430 -1360 62450 -1300
rect 62350 -1380 62450 -1360
rect 62690 -1300 62790 -1280
rect 62690 -1360 62710 -1300
rect 62770 -1360 62790 -1300
rect 62690 -1380 62790 -1360
rect 63030 -1300 63130 -1280
rect 63030 -1360 63050 -1300
rect 63110 -1360 63130 -1300
rect 63030 -1380 63130 -1360
rect 63370 -1300 63470 -1280
rect 63370 -1360 63390 -1300
rect 63450 -1360 63470 -1300
rect 63370 -1380 63470 -1360
rect 63710 -1300 63810 -1280
rect 63710 -1360 63730 -1300
rect 63790 -1360 63810 -1300
rect 63710 -1380 63810 -1360
rect 64050 -1300 64150 -1280
rect 64050 -1360 64070 -1300
rect 64130 -1360 64150 -1300
rect 64050 -1380 64150 -1360
rect 64390 -1300 64490 -1280
rect 64390 -1360 64410 -1300
rect 64470 -1360 64490 -1300
rect 64390 -1380 64490 -1360
rect 64730 -1300 64830 -1280
rect 64730 -1360 64750 -1300
rect 64810 -1360 64830 -1300
rect 64730 -1380 64830 -1360
rect 65070 -1300 65170 -1280
rect 65070 -1360 65090 -1300
rect 65150 -1360 65170 -1300
rect 65070 -1380 65170 -1360
rect 65410 -1300 65510 -1280
rect 65410 -1360 65430 -1300
rect 65490 -1360 65510 -1300
rect 65410 -1380 65510 -1360
rect 65750 -1300 65850 -1280
rect 65750 -1360 65770 -1300
rect 65830 -1360 65850 -1300
rect 65750 -1380 65850 -1360
rect 66090 -1300 66190 -1280
rect 66090 -1360 66110 -1300
rect 66170 -1360 66190 -1300
rect 66090 -1380 66190 -1360
rect 66430 -1300 66530 -1280
rect 66430 -1360 66450 -1300
rect 66510 -1360 66530 -1300
rect 66430 -1380 66530 -1360
rect 66770 -1300 66870 -1280
rect 66770 -1360 66790 -1300
rect 66850 -1360 66870 -1300
rect 66770 -1380 66870 -1360
rect 67110 -1300 67210 -1280
rect 67110 -1360 67130 -1300
rect 67190 -1360 67210 -1300
rect 67110 -1380 67210 -1360
rect 67450 -1300 67550 -1280
rect 67450 -1360 67470 -1300
rect 67530 -1360 67550 -1300
rect 67450 -1380 67550 -1360
rect 67790 -1300 67890 -1280
rect 67790 -1360 67810 -1300
rect 67870 -1360 67890 -1300
rect 67790 -1380 67890 -1360
rect 68130 -1300 68230 -1280
rect 68130 -1360 68150 -1300
rect 68210 -1360 68230 -1300
rect 68130 -1380 68230 -1360
rect 68470 -1300 68570 -1280
rect 68470 -1360 68490 -1300
rect 68550 -1360 68570 -1300
rect 68470 -1380 68570 -1360
rect 68810 -1300 68910 -1280
rect 68810 -1360 68830 -1300
rect 68890 -1360 68910 -1300
rect 68810 -1380 68910 -1360
rect 69150 -1300 69250 -1280
rect 69150 -1360 69170 -1300
rect 69230 -1360 69250 -1300
rect 69150 -1380 69250 -1360
rect 69490 -1300 69590 -1280
rect 69490 -1360 69510 -1300
rect 69570 -1360 69590 -1300
rect 69490 -1380 69590 -1360
rect 69830 -1300 69930 -1280
rect 69830 -1360 69850 -1300
rect 69910 -1360 69930 -1300
rect 69830 -1380 69930 -1360
rect 70170 -1300 70270 -1280
rect 70170 -1360 70190 -1300
rect 70250 -1360 70270 -1300
rect 70170 -1380 70270 -1360
rect 70510 -1300 70610 -1280
rect 70510 -1360 70530 -1300
rect 70590 -1360 70610 -1300
rect 70510 -1380 70610 -1360
rect 70850 -1300 70950 -1280
rect 70850 -1360 70870 -1300
rect 70930 -1360 70950 -1300
rect 70850 -1380 70950 -1360
rect 71190 -1300 71290 -1280
rect 71190 -1360 71210 -1300
rect 71270 -1360 71290 -1300
rect 71190 -1380 71290 -1360
rect 71530 -1300 71630 -1280
rect 71530 -1360 71550 -1300
rect 71610 -1360 71630 -1300
rect 71530 -1380 71630 -1360
rect 71870 -1300 71970 -1280
rect 71870 -1360 71890 -1300
rect 71950 -1360 71970 -1300
rect 71870 -1380 71970 -1360
rect 72210 -1300 72310 -1280
rect 72210 -1360 72230 -1300
rect 72290 -1360 72310 -1300
rect 72210 -1380 72310 -1360
rect 72550 -1300 72650 -1280
rect 72550 -1360 72570 -1300
rect 72630 -1360 72650 -1300
rect 72550 -1380 72650 -1360
rect 72890 -1300 72990 -1280
rect 72890 -1360 72910 -1300
rect 72970 -1360 72990 -1300
rect 72890 -1380 72990 -1360
rect 73230 -1300 73330 -1280
rect 73230 -1360 73250 -1300
rect 73310 -1360 73330 -1300
rect 73230 -1380 73330 -1360
rect 73570 -1300 73670 -1280
rect 73570 -1360 73590 -1300
rect 73650 -1360 73670 -1300
rect 73570 -1380 73670 -1360
rect 73910 -1300 74010 -1280
rect 73910 -1360 73930 -1300
rect 73990 -1360 74010 -1300
rect 73910 -1380 74010 -1360
rect 74250 -1300 74350 -1280
rect 74250 -1360 74270 -1300
rect 74330 -1360 74350 -1300
rect 74250 -1380 74350 -1360
rect 74590 -1300 74690 -1280
rect 74590 -1360 74610 -1300
rect 74670 -1360 74690 -1300
rect 74590 -1380 74690 -1360
rect 74930 -1300 75030 -1280
rect 74930 -1360 74950 -1300
rect 75010 -1360 75030 -1300
rect 74930 -1380 75030 -1360
rect 75270 -1300 75370 -1280
rect 75270 -1360 75290 -1300
rect 75350 -1360 75370 -1300
rect 75270 -1380 75370 -1360
rect 75610 -1300 75710 -1280
rect 75610 -1360 75630 -1300
rect 75690 -1360 75710 -1300
rect 75610 -1380 75710 -1360
rect 75950 -1300 76050 -1280
rect 75950 -1360 75970 -1300
rect 76030 -1360 76050 -1300
rect 75950 -1380 76050 -1360
rect 76290 -1300 76390 -1280
rect 76290 -1360 76310 -1300
rect 76370 -1360 76390 -1300
rect 76290 -1380 76390 -1360
rect 76630 -1300 76730 -1280
rect 76630 -1360 76650 -1300
rect 76710 -1360 76730 -1300
rect 76630 -1380 76730 -1360
rect 76970 -1300 77070 -1280
rect 76970 -1360 76990 -1300
rect 77050 -1360 77070 -1300
rect 76970 -1380 77070 -1360
rect 77310 -1300 77410 -1280
rect 77310 -1360 77330 -1300
rect 77390 -1360 77410 -1300
rect 77310 -1380 77410 -1360
rect 77650 -1300 77750 -1280
rect 77650 -1360 77670 -1300
rect 77730 -1360 77750 -1300
rect 77650 -1380 77750 -1360
rect 77990 -1300 78090 -1280
rect 77990 -1360 78010 -1300
rect 78070 -1360 78090 -1300
rect 77990 -1380 78090 -1360
rect 78330 -1300 78430 -1280
rect 78330 -1360 78350 -1300
rect 78410 -1360 78430 -1300
rect 78330 -1380 78430 -1360
rect 78670 -1300 78770 -1280
rect 78670 -1360 78690 -1300
rect 78750 -1360 78770 -1300
rect 78670 -1380 78770 -1360
rect 79010 -1300 79110 -1280
rect 79010 -1360 79030 -1300
rect 79090 -1360 79110 -1300
rect 79010 -1380 79110 -1360
rect 79350 -1300 79450 -1280
rect 79350 -1360 79370 -1300
rect 79430 -1360 79450 -1300
rect 79350 -1380 79450 -1360
rect 79690 -1300 79790 -1280
rect 79690 -1360 79710 -1300
rect 79770 -1360 79790 -1300
rect 79690 -1380 79790 -1360
rect 80030 -1300 80130 -1280
rect 80030 -1360 80050 -1300
rect 80110 -1360 80130 -1300
rect 80030 -1380 80130 -1360
rect 80370 -1300 80470 -1280
rect 80370 -1360 80390 -1300
rect 80450 -1360 80470 -1300
rect 80370 -1380 80470 -1360
rect 80710 -1300 80810 -1280
rect 80710 -1360 80730 -1300
rect 80790 -1360 80810 -1300
rect 80710 -1380 80810 -1360
rect 81050 -1300 81150 -1280
rect 81050 -1360 81070 -1300
rect 81130 -1360 81150 -1300
rect 81050 -1380 81150 -1360
rect 81390 -1300 81490 -1280
rect 81390 -1360 81410 -1300
rect 81470 -1360 81490 -1300
rect 81390 -1380 81490 -1360
rect 81730 -1300 81830 -1280
rect 81730 -1360 81750 -1300
rect 81810 -1360 81830 -1300
rect 81730 -1380 81830 -1360
rect 82070 -1300 82170 -1280
rect 82070 -1360 82090 -1300
rect 82150 -1360 82170 -1300
rect 82070 -1380 82170 -1360
rect 82410 -1300 82510 -1280
rect 82410 -1360 82430 -1300
rect 82490 -1360 82510 -1300
rect 82410 -1380 82510 -1360
rect 82750 -1300 82850 -1280
rect 82750 -1360 82770 -1300
rect 82830 -1360 82850 -1300
rect 82750 -1380 82850 -1360
rect 83090 -1300 83190 -1280
rect 83090 -1360 83110 -1300
rect 83170 -1360 83190 -1300
rect 83090 -1380 83190 -1360
rect 83430 -1300 83530 -1280
rect 83430 -1360 83450 -1300
rect 83510 -1360 83530 -1300
rect 83430 -1380 83530 -1360
rect 83770 -1300 83870 -1280
rect 83770 -1360 83790 -1300
rect 83850 -1360 83870 -1300
rect 83770 -1380 83870 -1360
rect 84110 -1300 84210 -1280
rect 84110 -1360 84130 -1300
rect 84190 -1360 84210 -1300
rect 84110 -1380 84210 -1360
rect 84450 -1300 84550 -1280
rect 84450 -1360 84470 -1300
rect 84530 -1360 84550 -1300
rect 84450 -1380 84550 -1360
rect 84790 -1300 84890 -1280
rect 84790 -1360 84810 -1300
rect 84870 -1360 84890 -1300
rect 84790 -1380 84890 -1360
rect 85130 -1300 85230 -1280
rect 85130 -1360 85150 -1300
rect 85210 -1360 85230 -1300
rect 85130 -1380 85230 -1360
rect 85470 -1300 85570 -1280
rect 85470 -1360 85490 -1300
rect 85550 -1360 85570 -1300
rect 85470 -1380 85570 -1360
rect 85810 -1300 85910 -1280
rect 85810 -1360 85830 -1300
rect 85890 -1360 85910 -1300
rect 85810 -1380 85910 -1360
rect 86150 -1300 86250 -1280
rect 86150 -1360 86170 -1300
rect 86230 -1360 86250 -1300
rect 86150 -1380 86250 -1360
rect 86490 -1300 86590 -1280
rect 86490 -1360 86510 -1300
rect 86570 -1360 86590 -1300
rect 86490 -1380 86590 -1360
rect 86830 -1300 86930 -1280
rect 86830 -1360 86850 -1300
rect 86910 -1360 86930 -1300
rect 86830 -1380 86930 -1360
rect 87170 -1300 87270 -1280
rect 87170 -1360 87190 -1300
rect 87250 -1360 87270 -1300
rect 87170 -1380 87270 -1360
rect 770 -1470 970 -1440
rect 770 -1540 830 -1470
rect 910 -1540 970 -1470
rect 770 -1570 970 -1540
rect 4940 -1470 5140 -1440
rect 4940 -1540 5000 -1470
rect 5080 -1540 5140 -1470
rect 4940 -1570 5140 -1540
rect 8970 -1470 9170 -1440
rect 8970 -1540 9030 -1470
rect 9110 -1540 9170 -1470
rect 8970 -1570 9170 -1540
rect 13000 -1470 13200 -1440
rect 13000 -1540 13060 -1470
rect 13140 -1540 13200 -1470
rect 13000 -1570 13200 -1540
rect 17040 -1470 17240 -1440
rect 17040 -1540 17100 -1470
rect 17180 -1540 17240 -1470
rect 17040 -1570 17240 -1540
rect 21140 -1470 21340 -1440
rect 21140 -1540 21200 -1470
rect 21280 -1540 21340 -1470
rect 21140 -1570 21340 -1540
rect 25250 -1470 25450 -1440
rect 25250 -1540 25310 -1470
rect 25390 -1540 25450 -1470
rect 25250 -1570 25450 -1540
rect 29350 -1470 29550 -1440
rect 29350 -1540 29410 -1470
rect 29490 -1540 29550 -1470
rect 29350 -1570 29550 -1540
rect 33380 -1470 33580 -1440
rect 33380 -1540 33440 -1470
rect 33520 -1540 33580 -1470
rect 33380 -1570 33580 -1540
rect 37490 -1470 37690 -1440
rect 37490 -1540 37550 -1470
rect 37630 -1540 37690 -1470
rect 37490 -1570 37690 -1540
rect 41590 -1470 41790 -1440
rect 41590 -1540 41650 -1470
rect 41730 -1540 41790 -1470
rect 41590 -1570 41790 -1540
rect 47040 -1470 47240 -1440
rect 47040 -1540 47100 -1470
rect 47180 -1540 47240 -1470
rect 47040 -1570 47240 -1540
rect 51120 -1470 51320 -1440
rect 51120 -1540 51180 -1470
rect 51260 -1540 51320 -1470
rect 51120 -1570 51320 -1540
rect 55230 -1470 55430 -1440
rect 55230 -1540 55290 -1470
rect 55370 -1540 55430 -1470
rect 55230 -1570 55430 -1540
rect 59260 -1470 59460 -1440
rect 59260 -1540 59320 -1470
rect 59400 -1540 59460 -1470
rect 59260 -1570 59460 -1540
rect 63360 -1470 63560 -1440
rect 63360 -1540 63420 -1470
rect 63500 -1540 63560 -1470
rect 63360 -1570 63560 -1540
rect 67470 -1470 67670 -1440
rect 67470 -1540 67530 -1470
rect 67610 -1540 67670 -1470
rect 67470 -1570 67670 -1540
rect 71500 -1470 71700 -1440
rect 71500 -1540 71560 -1470
rect 71640 -1540 71700 -1470
rect 71500 -1570 71700 -1540
rect 75750 -1470 75950 -1440
rect 75750 -1540 75810 -1470
rect 75890 -1540 75950 -1470
rect 75750 -1570 75950 -1540
rect 79710 -1470 79910 -1440
rect 79710 -1540 79770 -1470
rect 79850 -1540 79910 -1470
rect 79710 -1570 79910 -1540
rect 83890 -1470 84090 -1440
rect 83890 -1540 83950 -1470
rect 84030 -1540 84090 -1470
rect 83890 -1570 84090 -1540
rect 86450 -1474 86648 -1444
rect 86450 -1544 86508 -1474
rect 86588 -1544 86648 -1474
rect 86450 -1572 86648 -1544
<< via1 >>
rect 1300 650 1390 710
rect 790 520 870 590
rect 2170 520 2250 590
rect 3550 520 3630 590
rect 6390 630 6490 690
rect 5210 520 5290 590
rect 8040 520 8120 590
rect 10800 520 10880 590
rect 13430 520 13510 590
rect 16470 520 16550 590
rect 20540 520 20620 590
rect 24680 520 24760 590
rect 28760 520 28840 590
rect 32910 520 32990 590
rect 36780 520 36860 590
rect 40920 520 41000 590
rect 44910 520 44990 590
rect 48990 520 49070 590
rect 53080 520 53160 590
rect 57240 520 57320 590
rect 30 350 90 410
rect 450 350 510 410
rect 790 350 850 410
rect 1130 350 1190 410
rect 1520 350 1580 410
rect 1860 350 1920 410
rect 2200 350 2260 410
rect 2540 350 2600 410
rect 2880 350 2940 410
rect 3220 350 3280 410
rect 3560 350 3620 410
rect 3900 350 3960 410
rect 4240 350 4300 410
rect 4540 350 4600 410
rect 4880 350 4940 410
rect 5220 350 5280 410
rect 5560 350 5620 410
rect 5900 350 5960 410
rect 6240 350 6300 410
rect 6580 350 6640 410
rect 6920 350 6980 410
rect 7260 350 7320 410
rect 7600 350 7660 410
rect 7940 350 8000 410
rect 8280 350 8340 410
rect 8620 350 8680 410
rect 8960 350 9020 410
rect 9300 350 9360 410
rect 9640 350 9700 410
rect 9980 350 10040 410
rect 10320 350 10380 410
rect 10660 350 10720 410
rect 11000 350 11060 410
rect 11340 350 11400 410
rect 11680 350 11740 410
rect 12020 350 12080 410
rect 12360 350 12420 410
rect 12700 350 12760 410
rect 13040 350 13100 410
rect 13380 350 13440 410
rect 13720 350 13780 410
rect 14060 350 14120 410
rect 14400 350 14460 410
rect 14740 350 14800 410
rect 15080 350 15140 410
rect 15420 350 15480 410
rect 15720 350 15780 410
rect 16060 350 16120 410
rect 16400 350 16460 410
rect 16740 350 16800 410
rect 17080 350 17140 410
rect 17420 350 17480 410
rect 17760 350 17820 410
rect 18100 350 18160 410
rect 18440 350 18500 410
rect 18780 350 18840 410
rect 19120 350 19180 410
rect 19460 350 19520 410
rect 19800 350 19860 410
rect 20140 350 20200 410
rect 20480 350 20540 410
rect 20820 350 20880 410
rect 21160 350 21220 410
rect 21500 350 21560 410
rect 21840 350 21900 410
rect 22180 350 22240 410
rect 22520 350 22580 410
rect 22860 350 22920 410
rect 23200 350 23260 410
rect 23540 350 23600 410
rect 23880 350 23940 410
rect 24220 350 24280 410
rect 24560 350 24620 410
rect 24900 350 24960 410
rect 25240 350 25300 410
rect 25580 350 25640 410
rect 25920 350 25980 410
rect 26260 350 26320 410
rect 26600 350 26660 410
rect 26940 350 27000 410
rect 27280 350 27340 410
rect 27620 350 27680 410
rect 27960 350 28020 410
rect 28300 350 28360 410
rect 28640 350 28700 410
rect 28980 350 29040 410
rect 29320 350 29380 410
rect 29660 350 29720 410
rect 30000 350 30060 410
rect 30340 350 30400 410
rect 30680 350 30740 410
rect 31020 350 31080 410
rect 31360 350 31420 410
rect 31700 350 31760 410
rect 32040 350 32100 410
rect 32380 350 32440 410
rect 32720 350 32780 410
rect 33060 350 33120 410
rect 33400 350 33460 410
rect 33740 350 33800 410
rect 34080 350 34140 410
rect 34420 350 34480 410
rect 34760 350 34820 410
rect 35100 350 35160 410
rect 35440 350 35500 410
rect 35780 350 35840 410
rect 36120 350 36180 410
rect 36460 350 36520 410
rect 36800 350 36860 410
rect 37140 350 37200 410
rect 37480 350 37540 410
rect 37820 350 37880 410
rect 38160 350 38220 410
rect 38500 350 38560 410
rect 38840 350 38900 410
rect 39180 350 39240 410
rect 39520 350 39580 410
rect 39860 350 39920 410
rect 40200 350 40260 410
rect 40540 350 40600 410
rect 40880 350 40940 410
rect 41220 350 41280 410
rect 41560 350 41620 410
rect 41900 350 41960 410
rect 42240 350 42300 410
rect 42580 350 42640 410
rect 42920 350 42980 410
rect 43260 350 43320 410
rect 43600 350 43660 410
rect 43940 350 44000 410
rect 44280 350 44340 410
rect 44620 350 44680 410
rect 44960 350 45020 410
rect 45300 350 45360 410
rect 45640 350 45700 410
rect 45980 350 46040 410
rect 46320 350 46380 410
rect 46660 350 46720 410
rect 47000 350 47060 410
rect 47340 350 47400 410
rect 47680 350 47740 410
rect 48020 350 48080 410
rect 48360 350 48420 410
rect 48700 350 48760 410
rect 49040 350 49100 410
rect 49380 350 49440 410
rect 49720 350 49780 410
rect 50060 350 50120 410
rect 50400 350 50460 410
rect 50740 350 50800 410
rect 51080 350 51140 410
rect 51420 350 51480 410
rect 51760 350 51820 410
rect 52100 350 52160 410
rect 52440 350 52500 410
rect 52780 350 52840 410
rect 53120 350 53180 410
rect 53460 350 53520 410
rect 53800 350 53860 410
rect 54140 350 54200 410
rect 54480 350 54540 410
rect 54820 350 54880 410
rect 55160 350 55220 410
rect 55500 350 55560 410
rect 55840 350 55900 410
rect 56180 350 56240 410
rect 56520 350 56580 410
rect 56860 350 56920 410
rect 57200 350 57260 410
rect 57540 350 57600 410
rect 57880 350 57940 410
rect 58220 350 58280 410
rect 58560 350 58620 410
rect 58900 350 58960 410
rect 59240 350 59300 410
rect 70 30 130 110
rect 30 -120 90 -60
rect 620 130 680 200
rect 450 20 510 80
rect 960 130 1020 200
rect 790 20 850 80
rect 1690 130 1750 200
rect 1130 20 1190 80
rect 1520 20 1580 80
rect 2030 130 2090 200
rect 1860 20 1920 80
rect 2370 130 2430 200
rect 2200 20 2260 80
rect 2710 130 2770 200
rect 2540 20 2600 80
rect 3050 130 3110 200
rect 2880 20 2940 80
rect 3390 130 3450 200
rect 3220 20 3280 80
rect 3730 130 3790 200
rect 3560 20 3620 80
rect 4070 130 4130 200
rect 3900 20 3960 80
rect 4710 130 4770 200
rect 4240 20 4300 80
rect 4540 20 4600 80
rect 5050 130 5110 200
rect 4880 20 4940 80
rect 5390 130 5450 200
rect 5220 20 5280 80
rect 5730 130 5790 200
rect 5560 20 5620 80
rect 6070 130 6130 200
rect 5900 20 5960 80
rect 6410 130 6470 200
rect 6240 20 6300 80
rect 6750 130 6810 200
rect 6580 20 6640 80
rect 7090 130 7150 200
rect 6920 20 6980 80
rect 7430 130 7490 200
rect 7260 20 7320 80
rect 7770 130 7830 200
rect 7600 20 7660 80
rect 8110 130 8170 200
rect 7940 20 8000 80
rect 8450 130 8510 200
rect 8280 20 8340 80
rect 8790 130 8850 200
rect 8620 20 8680 80
rect 9130 130 9190 200
rect 8960 20 9020 80
rect 9470 130 9530 200
rect 9300 20 9360 80
rect 9810 130 9870 200
rect 9640 20 9700 80
rect 10150 130 10210 200
rect 9980 20 10040 80
rect 10490 130 10550 200
rect 10320 20 10380 80
rect 10830 130 10890 200
rect 10660 20 10720 80
rect 11170 130 11230 200
rect 11000 20 11060 80
rect 11510 130 11570 200
rect 11340 20 11400 80
rect 11850 130 11910 200
rect 11680 20 11740 80
rect 12190 130 12250 200
rect 12020 20 12080 80
rect 12530 130 12590 200
rect 12360 20 12420 80
rect 12870 130 12930 200
rect 12700 20 12760 80
rect 13210 130 13270 200
rect 13040 20 13100 80
rect 13550 130 13610 200
rect 13380 20 13440 80
rect 13890 130 13950 200
rect 13720 20 13780 80
rect 14230 130 14290 200
rect 14060 20 14120 80
rect 14570 130 14630 200
rect 14400 20 14460 80
rect 14910 130 14970 200
rect 14740 20 14800 80
rect 15250 130 15310 200
rect 15080 20 15140 80
rect 15890 130 15950 200
rect 15420 20 15480 80
rect 15720 20 15780 80
rect 16230 130 16290 200
rect 16060 20 16120 80
rect 16570 130 16630 200
rect 16400 20 16460 80
rect 16910 130 16970 200
rect 16740 20 16800 80
rect 17250 130 17310 200
rect 17080 20 17140 80
rect 17590 130 17650 200
rect 17420 20 17480 80
rect 17930 130 17990 200
rect 17760 20 17820 80
rect 18270 130 18330 200
rect 18100 20 18160 80
rect 18610 130 18670 200
rect 18440 20 18500 80
rect 18950 130 19010 200
rect 18780 20 18840 80
rect 19290 130 19350 200
rect 19120 20 19180 80
rect 19630 130 19690 200
rect 19460 20 19520 80
rect 19970 130 20030 200
rect 19800 20 19860 80
rect 20310 130 20370 200
rect 20140 20 20200 80
rect 20650 130 20710 200
rect 20480 20 20540 80
rect 20990 130 21050 200
rect 20820 20 20880 80
rect 21330 130 21390 200
rect 21160 20 21220 80
rect 21670 130 21730 200
rect 21500 20 21560 80
rect 22010 130 22070 200
rect 21840 20 21900 80
rect 22350 130 22410 200
rect 22180 20 22240 80
rect 22690 130 22750 200
rect 22520 20 22580 80
rect 23030 130 23090 200
rect 22860 20 22920 80
rect 23370 130 23430 200
rect 23200 20 23260 80
rect 23710 130 23770 200
rect 23540 20 23600 80
rect 24050 130 24110 200
rect 23880 20 23940 80
rect 24390 130 24450 200
rect 24220 20 24280 80
rect 24730 130 24790 200
rect 24560 20 24620 80
rect 25070 130 25130 200
rect 24900 20 24960 80
rect 25410 130 25470 200
rect 25240 20 25300 80
rect 25750 130 25810 200
rect 25580 20 25640 80
rect 26090 130 26150 200
rect 25920 20 25980 80
rect 26430 130 26490 200
rect 26260 20 26320 80
rect 26770 130 26830 200
rect 26600 20 26660 80
rect 27110 130 27170 200
rect 26940 20 27000 80
rect 27450 130 27510 200
rect 27280 20 27340 80
rect 27790 130 27850 200
rect 27620 20 27680 80
rect 28130 130 28190 200
rect 27960 20 28020 80
rect 28470 130 28530 200
rect 28300 20 28360 80
rect 28810 130 28870 200
rect 28640 20 28700 80
rect 29150 130 29210 200
rect 28980 20 29040 80
rect 29490 130 29550 200
rect 29320 20 29380 80
rect 29830 130 29890 200
rect 29660 20 29720 80
rect 30170 130 30230 200
rect 30000 20 30060 80
rect 30510 130 30570 200
rect 30340 20 30400 80
rect 30850 130 30910 200
rect 30680 20 30740 80
rect 31190 130 31250 200
rect 31020 20 31080 80
rect 31530 130 31590 200
rect 31360 20 31420 80
rect 31870 130 31930 200
rect 31700 20 31760 80
rect 32210 130 32270 200
rect 32040 20 32100 80
rect 32550 130 32610 200
rect 32380 20 32440 80
rect 32890 130 32950 200
rect 32720 20 32780 80
rect 33230 130 33290 200
rect 33060 20 33120 80
rect 33570 130 33630 200
rect 33400 20 33460 80
rect 33910 130 33970 200
rect 33740 20 33800 80
rect 34250 130 34310 200
rect 34080 20 34140 80
rect 34590 130 34650 200
rect 34420 20 34480 80
rect 34930 130 34990 200
rect 34760 20 34820 80
rect 35270 130 35330 200
rect 35100 20 35160 80
rect 35610 130 35670 200
rect 35440 20 35500 80
rect 35950 130 36010 200
rect 35780 20 35840 80
rect 36290 130 36350 200
rect 36120 20 36180 80
rect 36630 130 36690 200
rect 36460 20 36520 80
rect 36970 130 37030 200
rect 36800 20 36860 80
rect 37310 130 37370 200
rect 37140 20 37200 80
rect 37650 130 37710 200
rect 37480 20 37540 80
rect 37990 130 38050 200
rect 37820 20 37880 80
rect 38330 130 38390 200
rect 38160 20 38220 80
rect 38670 130 38730 200
rect 38500 20 38560 80
rect 39010 130 39070 200
rect 38840 20 38900 80
rect 39350 130 39410 200
rect 39180 20 39240 80
rect 39690 130 39750 200
rect 39520 20 39580 80
rect 40030 130 40090 200
rect 39860 20 39920 80
rect 40370 130 40430 200
rect 40200 20 40260 80
rect 40710 130 40770 200
rect 40540 20 40600 80
rect 41050 130 41110 200
rect 40880 20 40940 80
rect 41390 130 41450 200
rect 41220 20 41280 80
rect 41730 130 41790 200
rect 41560 20 41620 80
rect 42070 130 42130 200
rect 41900 20 41960 80
rect 42410 130 42470 200
rect 42240 20 42300 80
rect 42750 130 42810 200
rect 42580 20 42640 80
rect 43090 130 43150 200
rect 42920 20 42980 80
rect 43430 130 43490 200
rect 43260 20 43320 80
rect 43770 130 43830 200
rect 43600 20 43660 80
rect 44110 130 44170 200
rect 43940 20 44000 80
rect 44450 130 44510 200
rect 44280 20 44340 80
rect 44790 130 44850 200
rect 44620 20 44680 80
rect 45130 130 45190 200
rect 44960 20 45020 80
rect 45470 130 45530 200
rect 45300 20 45360 80
rect 45810 130 45870 200
rect 45640 20 45700 80
rect 46150 130 46210 200
rect 45980 20 46040 80
rect 46490 130 46550 200
rect 46320 20 46380 80
rect 46830 130 46890 200
rect 46660 20 46720 80
rect 47170 130 47230 200
rect 47000 20 47060 80
rect 47510 130 47570 200
rect 47340 20 47400 80
rect 47850 130 47910 200
rect 47680 20 47740 80
rect 48190 130 48250 200
rect 48020 20 48080 80
rect 48530 130 48590 200
rect 48360 20 48420 80
rect 48870 130 48930 200
rect 48700 20 48760 80
rect 49210 130 49270 200
rect 49040 20 49100 80
rect 49550 130 49610 200
rect 49380 20 49440 80
rect 49890 130 49950 200
rect 49720 20 49780 80
rect 50230 130 50290 200
rect 50060 20 50120 80
rect 50570 130 50630 200
rect 50400 20 50460 80
rect 50910 130 50970 200
rect 50740 20 50800 80
rect 51250 130 51310 200
rect 51080 20 51140 80
rect 51590 130 51650 200
rect 51420 20 51480 80
rect 51930 130 51990 200
rect 51760 20 51820 80
rect 52270 130 52330 200
rect 52100 20 52160 80
rect 52610 130 52670 200
rect 52440 20 52500 80
rect 52950 130 53010 200
rect 52780 20 52840 80
rect 53290 130 53350 200
rect 53120 20 53180 80
rect 53630 130 53690 200
rect 53460 20 53520 80
rect 53970 130 54030 200
rect 53800 20 53860 80
rect 54310 130 54370 200
rect 54140 20 54200 80
rect 54650 130 54710 200
rect 54480 20 54540 80
rect 54990 130 55050 200
rect 54820 20 54880 80
rect 55330 130 55390 200
rect 55160 20 55220 80
rect 55670 130 55730 200
rect 55500 20 55560 80
rect 56010 130 56070 200
rect 55840 20 55900 80
rect 56350 130 56410 200
rect 56180 20 56240 80
rect 56690 130 56750 200
rect 56520 20 56580 80
rect 57030 130 57090 200
rect 56860 20 56920 80
rect 57370 130 57430 200
rect 57200 20 57260 80
rect 57710 130 57770 200
rect 57540 20 57600 80
rect 58050 130 58110 200
rect 57880 20 57940 80
rect 58390 130 58450 200
rect 58220 20 58280 80
rect 58730 130 58790 200
rect 58560 20 58620 80
rect 59070 130 59130 200
rect 58900 20 58960 80
rect 59240 20 59300 80
rect 200 -120 260 -60
rect 530 -120 600 -60
rect 700 -120 770 -60
rect 870 -120 940 -60
rect 1040 -120 1110 -60
rect 1600 -120 1670 -60
rect 1770 -120 1840 -60
rect 1940 -120 2010 -60
rect 2110 -120 2180 -60
rect 2280 -120 2350 -60
rect 2450 -120 2520 -60
rect 2620 -120 2690 -60
rect 2790 -120 2860 -60
rect 2960 -120 3030 -60
rect 3130 -120 3200 -60
rect 3300 -120 3370 -60
rect 3470 -120 3540 -60
rect 3640 -120 3710 -60
rect 3810 -120 3880 -60
rect 3980 -120 4050 -60
rect 4150 -120 4220 -60
rect 4620 -120 4690 -60
rect 4790 -120 4860 -60
rect 4960 -120 5030 -60
rect 5130 -120 5200 -60
rect 5300 -120 5370 -60
rect 5470 -120 5540 -60
rect 5640 -120 5710 -60
rect 5810 -120 5880 -60
rect 5980 -120 6050 -60
rect 6150 -120 6220 -60
rect 6320 -120 6390 -60
rect 6490 -120 6560 -60
rect 6660 -120 6730 -60
rect 6830 -120 6900 -60
rect 7000 -120 7070 -60
rect 7170 -120 7240 -60
rect 7340 -120 7410 -60
rect 7510 -120 7580 -60
rect 7680 -120 7750 -60
rect 7850 -120 7920 -60
rect 8020 -120 8090 -60
rect 8190 -120 8260 -60
rect 8360 -120 8430 -60
rect 8530 -120 8600 -60
rect 8700 -120 8770 -60
rect 8870 -120 8940 -60
rect 9040 -120 9110 -60
rect 9210 -120 9280 -60
rect 9380 -120 9450 -60
rect 9550 -120 9620 -60
rect 9720 -120 9790 -60
rect 9890 -120 9960 -60
rect 10060 -120 10130 -60
rect 10230 -120 10300 -60
rect 10400 -120 10470 -60
rect 10570 -120 10640 -60
rect 10740 -120 10810 -60
rect 10910 -120 10980 -60
rect 11080 -120 11150 -60
rect 11250 -120 11320 -60
rect 11420 -120 11490 -60
rect 11590 -120 11660 -60
rect 11760 -120 11830 -60
rect 11930 -120 12000 -60
rect 12100 -120 12170 -60
rect 12270 -120 12340 -60
rect 12440 -120 12510 -60
rect 12610 -120 12680 -60
rect 12780 -120 12850 -60
rect 12950 -120 13020 -60
rect 13120 -120 13190 -60
rect 13290 -120 13360 -60
rect 13460 -120 13530 -60
rect 13630 -120 13700 -60
rect 13800 -120 13870 -60
rect 13970 -120 14040 -60
rect 14140 -120 14210 -60
rect 14310 -120 14380 -60
rect 14480 -120 14550 -60
rect 14650 -120 14720 -60
rect 14820 -120 14890 -60
rect 14990 -120 15060 -60
rect 15160 -120 15230 -60
rect 15330 -120 15400 -60
rect 15800 -120 15870 -60
rect 15970 -120 16040 -60
rect 16140 -120 16210 -60
rect 16310 -120 16380 -60
rect 16480 -120 16550 -60
rect 16650 -120 16720 -60
rect 16820 -120 16890 -60
rect 16990 -120 17060 -60
rect 17160 -120 17230 -60
rect 17330 -120 17400 -60
rect 17500 -120 17570 -60
rect 17670 -120 17740 -60
rect 17840 -120 17910 -60
rect 18010 -120 18080 -60
rect 18180 -120 18250 -60
rect 18350 -120 18420 -60
rect 18520 -120 18590 -60
rect 18690 -120 18760 -60
rect 18860 -120 18930 -60
rect 19030 -120 19100 -60
rect 19200 -120 19270 -60
rect 19370 -120 19440 -60
rect 19540 -120 19610 -60
rect 19710 -120 19780 -60
rect 19880 -120 19950 -60
rect 20050 -120 20120 -60
rect 20220 -120 20290 -60
rect 20390 -120 20460 -60
rect 20560 -120 20630 -60
rect 20730 -120 20800 -60
rect 20900 -120 20970 -60
rect 21070 -120 21140 -60
rect 21240 -120 21310 -60
rect 21410 -120 21480 -60
rect 21580 -120 21650 -60
rect 21750 -120 21820 -60
rect 21920 -120 21990 -60
rect 22090 -120 22160 -60
rect 22260 -120 22330 -60
rect 22430 -120 22500 -60
rect 22600 -120 22670 -60
rect 22770 -120 22840 -60
rect 22940 -120 23010 -60
rect 23110 -120 23180 -60
rect 23280 -120 23350 -60
rect 23450 -120 23520 -60
rect 23620 -120 23690 -60
rect 23790 -120 23860 -60
rect 23960 -120 24030 -60
rect 24130 -120 24200 -60
rect 24300 -120 24370 -60
rect 24470 -120 24540 -60
rect 24640 -120 24710 -60
rect 24810 -120 24880 -60
rect 24980 -120 25050 -60
rect 25150 -120 25220 -60
rect 25320 -120 25390 -60
rect 25490 -120 25560 -60
rect 25660 -120 25730 -60
rect 25830 -120 25900 -60
rect 26000 -120 26070 -60
rect 26170 -120 26240 -60
rect 26340 -120 26410 -60
rect 26510 -120 26580 -60
rect 26680 -120 26750 -60
rect 26850 -120 26920 -60
rect 27020 -120 27090 -60
rect 27190 -120 27260 -60
rect 27360 -120 27430 -60
rect 27530 -120 27600 -60
rect 27700 -120 27770 -60
rect 27870 -120 27940 -60
rect 28040 -120 28110 -60
rect 28210 -120 28280 -60
rect 28380 -120 28450 -60
rect 28550 -120 28620 -60
rect 28720 -120 28790 -60
rect 28890 -120 28960 -60
rect 29060 -120 29130 -60
rect 29230 -120 29300 -60
rect 29400 -120 29470 -60
rect 29570 -120 29640 -60
rect 29740 -120 29810 -60
rect 29910 -120 29980 -60
rect 30080 -120 30150 -60
rect 30250 -120 30320 -60
rect 30420 -120 30490 -60
rect 30590 -120 30660 -60
rect 30760 -120 30830 -60
rect 30930 -120 31000 -60
rect 31100 -120 31170 -60
rect 31270 -120 31340 -60
rect 31440 -120 31510 -60
rect 31610 -120 31680 -60
rect 31780 -120 31850 -60
rect 31950 -120 32020 -60
rect 32120 -120 32190 -60
rect 32290 -120 32360 -60
rect 32460 -120 32530 -60
rect 32630 -120 32700 -60
rect 32800 -120 32870 -60
rect 32970 -120 33040 -60
rect 33140 -120 33210 -60
rect 33310 -120 33380 -60
rect 33480 -120 33550 -60
rect 33650 -120 33720 -60
rect 33820 -120 33890 -60
rect 33990 -120 34060 -60
rect 34160 -120 34230 -60
rect 34330 -120 34400 -60
rect 34500 -120 34570 -60
rect 34670 -120 34740 -60
rect 34840 -120 34910 -60
rect 35010 -120 35080 -60
rect 35180 -120 35250 -60
rect 35350 -120 35420 -60
rect 35520 -120 35590 -60
rect 35690 -120 35760 -60
rect 35860 -120 35930 -60
rect 36030 -120 36100 -60
rect 36200 -120 36270 -60
rect 36370 -120 36440 -60
rect 36540 -120 36610 -60
rect 36710 -120 36780 -60
rect 36880 -120 36950 -60
rect 37050 -120 37120 -60
rect 37220 -120 37290 -60
rect 37390 -120 37460 -60
rect 37560 -120 37630 -60
rect 37730 -120 37800 -60
rect 37900 -120 37970 -60
rect 38070 -120 38140 -60
rect 38240 -120 38310 -60
rect 38410 -120 38480 -60
rect 38580 -120 38650 -60
rect 38750 -120 38820 -60
rect 38920 -120 38990 -60
rect 39090 -120 39160 -60
rect 39260 -120 39330 -60
rect 39430 -120 39500 -60
rect 39600 -120 39670 -60
rect 39770 -120 39840 -60
rect 39940 -120 40010 -60
rect 40110 -120 40180 -60
rect 40280 -120 40350 -60
rect 40450 -120 40520 -60
rect 40620 -120 40690 -60
rect 40790 -120 40860 -60
rect 40960 -120 41030 -60
rect 41130 -120 41200 -60
rect 41300 -120 41370 -60
rect 41470 -120 41540 -60
rect 41640 -120 41710 -60
rect 41810 -120 41880 -60
rect 41980 -120 42050 -60
rect 42150 -120 42220 -60
rect 42320 -120 42390 -60
rect 42490 -120 42560 -60
rect 42660 -120 42730 -60
rect 42830 -120 42900 -60
rect 43000 -120 43070 -60
rect 43170 -120 43240 -60
rect 43340 -120 43410 -60
rect 43510 -120 43580 -60
rect 43680 -120 43750 -60
rect 43850 -120 43920 -60
rect 44020 -120 44090 -60
rect 44190 -120 44260 -60
rect 44360 -120 44430 -60
rect 44530 -120 44600 -60
rect 44700 -120 44770 -60
rect 44870 -120 44940 -60
rect 45040 -120 45110 -60
rect 45210 -120 45280 -60
rect 45380 -120 45450 -60
rect 45550 -120 45620 -60
rect 45720 -120 45790 -60
rect 45890 -120 45960 -60
rect 46060 -120 46130 -60
rect 46230 -120 46300 -60
rect 46400 -120 46470 -60
rect 46570 -120 46640 -60
rect 46740 -120 46810 -60
rect 46910 -120 46980 -60
rect 47080 -120 47150 -60
rect 47250 -120 47320 -60
rect 47420 -120 47490 -60
rect 47590 -120 47660 -60
rect 47760 -120 47830 -60
rect 47930 -120 48000 -60
rect 48100 -120 48170 -60
rect 48270 -120 48340 -60
rect 48440 -120 48510 -60
rect 48610 -120 48680 -60
rect 48780 -120 48850 -60
rect 48950 -120 49020 -60
rect 49120 -120 49190 -60
rect 49290 -120 49360 -60
rect 49460 -120 49530 -60
rect 49630 -120 49700 -60
rect 49800 -120 49870 -60
rect 49970 -120 50040 -60
rect 50140 -120 50210 -60
rect 50310 -120 50380 -60
rect 50480 -120 50550 -60
rect 50650 -120 50720 -60
rect 50820 -120 50890 -60
rect 50990 -120 51060 -60
rect 51160 -120 51230 -60
rect 51330 -120 51400 -60
rect 51500 -120 51570 -60
rect 51670 -120 51740 -60
rect 51840 -120 51910 -60
rect 52010 -120 52080 -60
rect 52180 -120 52250 -60
rect 52350 -120 52420 -60
rect 52520 -120 52590 -60
rect 52690 -120 52760 -60
rect 52860 -120 52930 -60
rect 53030 -120 53100 -60
rect 53200 -120 53270 -60
rect 53370 -120 53440 -60
rect 53540 -120 53610 -60
rect 53710 -120 53780 -60
rect 53880 -120 53950 -60
rect 54050 -120 54120 -60
rect 54220 -120 54290 -60
rect 54390 -120 54460 -60
rect 54560 -120 54630 -60
rect 54730 -120 54800 -60
rect 54900 -120 54970 -60
rect 55070 -120 55140 -60
rect 55240 -120 55310 -60
rect 55410 -120 55480 -60
rect 55580 -120 55650 -60
rect 55750 -120 55820 -60
rect 55920 -120 55990 -60
rect 56090 -120 56160 -60
rect 56260 -120 56330 -60
rect 56430 -120 56500 -60
rect 56600 -120 56670 -60
rect 56770 -120 56840 -60
rect 56940 -120 57010 -60
rect 57110 -120 57180 -60
rect 57280 -120 57350 -60
rect 57450 -120 57520 -60
rect 57620 -120 57690 -60
rect 57790 -120 57860 -60
rect 57960 -120 58030 -60
rect 58130 -120 58200 -60
rect 58300 -120 58370 -60
rect 58470 -120 58540 -60
rect 58640 -120 58710 -60
rect 58810 -120 58880 -60
rect 58980 -120 59050 -60
rect 59150 -120 59220 -60
rect 2120 -390 2350 -260
rect 5138 -398 5368 -268
rect 7624 -398 7854 -268
rect 9044 -398 9274 -268
rect 13668 -394 13898 -264
rect 16868 -394 17098 -264
rect 20424 -394 20654 -264
rect 25758 -394 25988 -264
rect 28602 -394 28832 -264
rect 32514 -394 32744 -264
rect 34670 -394 34900 -264
rect 37492 -394 37722 -264
rect 40692 -394 40922 -264
rect 45668 -394 45898 -264
rect 48868 -394 49098 -264
rect 51002 -394 51232 -264
rect 54558 -394 54788 -264
rect 57402 -394 57632 -264
rect 61314 -394 61544 -264
rect 64158 -394 64388 -264
rect 67714 -394 67944 -264
rect 70558 -394 70788 -264
rect 74468 -394 74698 -264
rect 78380 -394 78610 -264
rect 82292 -394 82522 -264
rect 86202 -394 86432 -264
rect 230 -590 300 -530
rect 400 -590 470 -530
rect 570 -590 640 -530
rect 740 -590 810 -530
rect 910 -590 980 -530
rect 1080 -590 1150 -530
rect 1250 -590 1320 -530
rect 1420 -590 1490 -530
rect 1590 -590 1660 -530
rect 1760 -590 1830 -530
rect 1930 -590 2000 -530
rect 2100 -590 2170 -530
rect 2270 -590 2340 -530
rect 2440 -590 2510 -530
rect 2610 -590 2680 -530
rect 2780 -590 2850 -530
rect 2950 -590 3020 -530
rect 3120 -590 3190 -530
rect 3290 -590 3360 -530
rect 3460 -590 3530 -530
rect 3630 -590 3700 -530
rect 3800 -590 3870 -530
rect 3970 -590 4040 -530
rect 4140 -590 4210 -530
rect 4310 -590 4380 -530
rect 4480 -590 4550 -530
rect 4650 -590 4720 -530
rect 4820 -590 4890 -530
rect 4990 -590 5060 -530
rect 5160 -590 5230 -530
rect 5330 -590 5400 -530
rect 5500 -590 5570 -530
rect 5670 -590 5740 -530
rect 5840 -590 5910 -530
rect 6010 -590 6080 -530
rect 6180 -590 6250 -530
rect 6350 -590 6420 -530
rect 6520 -590 6590 -530
rect 6690 -590 6760 -530
rect 6860 -590 6930 -530
rect 7030 -590 7100 -530
rect 7200 -590 7270 -530
rect 7370 -590 7440 -530
rect 7540 -590 7610 -530
rect 7710 -590 7780 -530
rect 7880 -590 7950 -530
rect 8050 -590 8120 -530
rect 8220 -590 8290 -530
rect 8390 -590 8460 -530
rect 8560 -590 8630 -530
rect 8730 -590 8800 -530
rect 8900 -590 8970 -530
rect 9070 -590 9140 -530
rect 9240 -590 9310 -530
rect 9410 -590 9480 -530
rect 9580 -590 9650 -530
rect 9750 -590 9820 -530
rect 9920 -590 9990 -530
rect 10090 -590 10160 -530
rect 10260 -590 10330 -530
rect 10430 -590 10500 -530
rect 10600 -590 10670 -530
rect 10770 -590 10840 -530
rect 10940 -590 11010 -530
rect 11110 -590 11180 -530
rect 11280 -590 11350 -530
rect 11450 -590 11520 -530
rect 11620 -590 11690 -530
rect 11790 -590 11860 -530
rect 11960 -590 12030 -530
rect 12130 -590 12200 -530
rect 12300 -590 12370 -530
rect 12470 -590 12540 -530
rect 12640 -590 12710 -530
rect 12810 -590 12880 -530
rect 12980 -590 13050 -530
rect 13150 -590 13220 -530
rect 13320 -590 13390 -530
rect 13490 -590 13560 -530
rect 13660 -590 13730 -530
rect 13830 -590 13900 -530
rect 14000 -590 14070 -530
rect 14170 -590 14240 -530
rect 14340 -590 14410 -530
rect 14510 -590 14580 -530
rect 14680 -590 14750 -530
rect 14850 -590 14920 -530
rect 15020 -590 15090 -530
rect 15190 -590 15260 -530
rect 15360 -590 15430 -530
rect 15530 -590 15600 -530
rect 15700 -590 15770 -530
rect 15870 -590 15940 -530
rect 16040 -590 16110 -530
rect 16210 -590 16280 -530
rect 16380 -590 16450 -530
rect 16550 -590 16620 -530
rect 16720 -590 16790 -530
rect 16890 -590 16960 -530
rect 17060 -590 17130 -530
rect 17230 -590 17300 -530
rect 17400 -590 17470 -530
rect 17570 -590 17640 -530
rect 17740 -590 17810 -530
rect 17910 -590 17980 -530
rect 18080 -590 18150 -530
rect 18250 -590 18320 -530
rect 18420 -590 18490 -530
rect 18590 -590 18660 -530
rect 18760 -590 18830 -530
rect 18930 -590 19000 -530
rect 19100 -590 19170 -530
rect 19270 -590 19340 -530
rect 19440 -590 19510 -530
rect 19610 -590 19680 -530
rect 19780 -590 19850 -530
rect 19950 -590 20020 -530
rect 20120 -590 20190 -530
rect 20290 -590 20360 -530
rect 20460 -590 20530 -530
rect 20630 -590 20700 -530
rect 20800 -590 20870 -530
rect 20970 -590 21040 -530
rect 21140 -590 21210 -530
rect 21310 -590 21380 -530
rect 21480 -590 21550 -530
rect 21650 -590 21720 -530
rect 21820 -590 21890 -530
rect 21990 -590 22060 -530
rect 22160 -590 22230 -530
rect 22330 -590 22400 -530
rect 22500 -590 22570 -530
rect 22670 -590 22740 -530
rect 22840 -590 22910 -530
rect 23010 -590 23080 -530
rect 23180 -590 23250 -530
rect 23350 -590 23420 -530
rect 23520 -590 23590 -530
rect 23690 -590 23760 -530
rect 23860 -590 23930 -530
rect 24030 -590 24100 -530
rect 24200 -590 24270 -530
rect 24370 -590 24440 -530
rect 24540 -590 24610 -530
rect 24710 -590 24780 -530
rect 24880 -590 24950 -530
rect 25050 -590 25120 -530
rect 25220 -590 25290 -530
rect 25390 -590 25460 -530
rect 25560 -590 25630 -530
rect 25730 -590 25800 -530
rect 25900 -590 25970 -530
rect 26070 -590 26140 -530
rect 26240 -590 26310 -530
rect 26410 -590 26480 -530
rect 26580 -590 26650 -530
rect 26750 -590 26820 -530
rect 26920 -590 26990 -530
rect 27090 -590 27160 -530
rect 27260 -590 27330 -530
rect 27430 -590 27500 -530
rect 27600 -590 27670 -530
rect 27770 -590 27840 -530
rect 27940 -590 28010 -530
rect 28110 -590 28180 -530
rect 28280 -590 28350 -530
rect 28450 -590 28520 -530
rect 28620 -590 28690 -530
rect 28790 -590 28860 -530
rect 28960 -590 29030 -530
rect 29130 -590 29200 -530
rect 29300 -590 29370 -530
rect 29470 -590 29540 -530
rect 29640 -590 29710 -530
rect 29810 -590 29880 -530
rect 29980 -590 30050 -530
rect 30150 -590 30220 -530
rect 30320 -590 30390 -530
rect 30490 -590 30560 -530
rect 30660 -590 30730 -530
rect 30830 -590 30900 -530
rect 31000 -590 31070 -530
rect 31170 -590 31240 -530
rect 31340 -590 31410 -530
rect 31510 -590 31580 -530
rect 31680 -590 31750 -530
rect 31850 -590 31920 -530
rect 32020 -590 32090 -530
rect 32190 -590 32260 -530
rect 32360 -590 32430 -530
rect 32530 -590 32600 -530
rect 32700 -590 32770 -530
rect 32870 -590 32940 -530
rect 33040 -590 33110 -530
rect 33210 -590 33280 -530
rect 33380 -590 33450 -530
rect 33550 -590 33620 -530
rect 33720 -590 33790 -530
rect 33890 -590 33960 -530
rect 34060 -590 34130 -530
rect 34230 -590 34300 -530
rect 34400 -590 34470 -530
rect 34570 -590 34640 -530
rect 34740 -590 34810 -530
rect 34910 -590 34980 -530
rect 35080 -590 35150 -530
rect 35250 -590 35320 -530
rect 35420 -590 35490 -530
rect 35590 -590 35660 -530
rect 35760 -590 35830 -530
rect 35930 -590 36000 -530
rect 36100 -590 36170 -530
rect 36270 -590 36340 -530
rect 36440 -590 36510 -530
rect 36610 -590 36680 -530
rect 36780 -590 36850 -530
rect 36950 -590 37020 -530
rect 37120 -590 37190 -530
rect 37290 -590 37360 -530
rect 37460 -590 37530 -530
rect 37630 -590 37700 -530
rect 37800 -590 37870 -530
rect 37970 -590 38040 -530
rect 38140 -590 38210 -530
rect 38310 -590 38380 -530
rect 38480 -590 38550 -530
rect 38650 -590 38720 -530
rect 38820 -590 38890 -530
rect 38990 -590 39060 -530
rect 39160 -590 39230 -530
rect 39330 -590 39400 -530
rect 39500 -590 39570 -530
rect 39670 -590 39740 -530
rect 39840 -590 39910 -530
rect 40010 -590 40080 -530
rect 40180 -590 40250 -530
rect 40350 -590 40420 -530
rect 40520 -590 40590 -530
rect 40690 -590 40760 -530
rect 40860 -590 40930 -530
rect 41030 -590 41100 -530
rect 41200 -590 41270 -530
rect 41370 -590 41440 -530
rect 41540 -590 41610 -530
rect 41710 -590 41780 -530
rect 41880 -590 41950 -530
rect 42050 -590 42120 -530
rect 42220 -590 42290 -530
rect 42390 -590 42460 -530
rect 42560 -590 42630 -530
rect 42730 -590 42800 -530
rect 42900 -590 42970 -530
rect 43070 -590 43140 -530
rect 43240 -590 43310 -530
rect 43410 -590 43480 -530
rect 43580 -590 43650 -530
rect 43750 -590 43820 -530
rect 43920 -590 43990 -530
rect 44090 -590 44160 -530
rect 44260 -590 44330 -530
rect 44430 -590 44500 -530
rect 44600 -590 44670 -530
rect 44770 -590 44840 -530
rect 44940 -590 45010 -530
rect 45110 -590 45180 -530
rect 45280 -590 45350 -530
rect 45450 -590 45520 -530
rect 45620 -590 45690 -530
rect 45790 -590 45860 -530
rect 45960 -590 46030 -530
rect 46130 -590 46200 -530
rect 46300 -590 46370 -530
rect 46470 -590 46540 -530
rect 46640 -590 46710 -530
rect 46810 -590 46880 -530
rect 46980 -590 47050 -530
rect 47150 -590 47220 -530
rect 47320 -590 47390 -530
rect 47490 -590 47560 -530
rect 47660 -590 47730 -530
rect 47830 -590 47900 -530
rect 48000 -590 48070 -530
rect 48170 -590 48240 -530
rect 48340 -590 48410 -530
rect 48510 -590 48580 -530
rect 48680 -590 48750 -530
rect 48850 -590 48920 -530
rect 49020 -590 49090 -530
rect 49190 -590 49260 -530
rect 49360 -590 49430 -530
rect 49530 -590 49600 -530
rect 49700 -590 49770 -530
rect 49870 -590 49940 -530
rect 50040 -590 50110 -530
rect 50210 -590 50280 -530
rect 50380 -590 50450 -530
rect 50550 -590 50620 -530
rect 50720 -590 50790 -530
rect 50890 -590 50960 -530
rect 51060 -590 51130 -530
rect 51230 -590 51300 -530
rect 51400 -590 51470 -530
rect 51570 -590 51640 -530
rect 51740 -590 51810 -530
rect 51910 -590 51980 -530
rect 52080 -590 52150 -530
rect 52250 -590 52320 -530
rect 52420 -590 52490 -530
rect 52590 -590 52660 -530
rect 52760 -590 52830 -530
rect 52930 -590 53000 -530
rect 53100 -590 53170 -530
rect 53270 -590 53340 -530
rect 53440 -590 53510 -530
rect 53610 -590 53680 -530
rect 53780 -590 53850 -530
rect 53950 -590 54020 -530
rect 54120 -590 54190 -530
rect 54290 -590 54360 -530
rect 54460 -590 54530 -530
rect 54630 -590 54700 -530
rect 54800 -590 54870 -530
rect 54970 -590 55040 -530
rect 55140 -590 55210 -530
rect 55310 -590 55380 -530
rect 55480 -590 55550 -530
rect 55650 -590 55720 -530
rect 55820 -590 55890 -530
rect 55990 -590 56060 -530
rect 56160 -590 56230 -530
rect 56330 -590 56400 -530
rect 56500 -590 56570 -530
rect 56670 -590 56740 -530
rect 56840 -590 56910 -530
rect 57010 -590 57080 -530
rect 57180 -590 57250 -530
rect 57350 -590 57420 -530
rect 57520 -590 57590 -530
rect 57690 -590 57760 -530
rect 57860 -590 57930 -530
rect 58030 -590 58100 -530
rect 58200 -590 58270 -530
rect 58370 -590 58440 -530
rect 58540 -590 58610 -530
rect 58710 -590 58780 -530
rect 58880 -590 58950 -530
rect 59050 -590 59120 -530
rect 59220 -590 59290 -530
rect 59390 -590 59460 -530
rect 59560 -590 59630 -530
rect 59730 -590 59800 -530
rect 59900 -590 59970 -530
rect 60070 -590 60140 -530
rect 60240 -590 60310 -530
rect 60410 -590 60480 -530
rect 60580 -590 60650 -530
rect 60750 -590 60820 -530
rect 60920 -590 60990 -530
rect 61090 -590 61160 -530
rect 61260 -590 61330 -530
rect 61430 -590 61500 -530
rect 61600 -590 61670 -530
rect 61770 -590 61840 -530
rect 61940 -590 62010 -530
rect 62110 -590 62180 -530
rect 62280 -590 62350 -530
rect 62450 -590 62520 -530
rect 62620 -590 62690 -530
rect 62790 -590 62860 -530
rect 62960 -590 63030 -530
rect 63130 -590 63200 -530
rect 63300 -590 63370 -530
rect 63470 -590 63540 -530
rect 63640 -590 63710 -530
rect 63810 -590 63880 -530
rect 63980 -590 64050 -530
rect 64150 -590 64220 -530
rect 64320 -590 64390 -530
rect 64490 -590 64560 -530
rect 64660 -590 64730 -530
rect 64830 -590 64900 -530
rect 65000 -590 65070 -530
rect 65170 -590 65240 -530
rect 65340 -590 65410 -530
rect 65510 -590 65580 -530
rect 65680 -590 65750 -530
rect 65850 -590 65920 -530
rect 66020 -590 66090 -530
rect 66190 -590 66260 -530
rect 66360 -590 66430 -530
rect 66530 -590 66600 -530
rect 66700 -590 66770 -530
rect 66870 -590 66940 -530
rect 67040 -590 67110 -530
rect 67210 -590 67280 -530
rect 67380 -590 67450 -530
rect 67550 -590 67620 -530
rect 67720 -590 67790 -530
rect 67890 -590 67960 -530
rect 68060 -590 68130 -530
rect 68230 -590 68300 -530
rect 68400 -590 68470 -530
rect 68570 -590 68640 -530
rect 68740 -590 68810 -530
rect 68910 -590 68980 -530
rect 69080 -590 69150 -530
rect 69250 -590 69320 -530
rect 69420 -590 69490 -530
rect 69590 -590 69660 -530
rect 69760 -590 69830 -530
rect 69930 -590 70000 -530
rect 70100 -590 70170 -530
rect 70270 -590 70340 -530
rect 70440 -590 70510 -530
rect 70610 -590 70680 -530
rect 70780 -590 70850 -530
rect 70950 -590 71020 -530
rect 71120 -590 71190 -530
rect 71290 -590 71360 -530
rect 71460 -590 71530 -530
rect 71630 -590 71700 -530
rect 71800 -590 71870 -530
rect 71970 -590 72040 -530
rect 72140 -590 72210 -530
rect 72310 -590 72380 -530
rect 72480 -590 72550 -530
rect 72650 -590 72720 -530
rect 72820 -590 72890 -530
rect 72990 -590 73060 -530
rect 73160 -590 73230 -530
rect 73330 -590 73400 -530
rect 73500 -590 73570 -530
rect 73670 -590 73740 -530
rect 73840 -590 73910 -530
rect 74010 -590 74080 -530
rect 74180 -590 74250 -530
rect 74350 -590 74420 -530
rect 74520 -590 74590 -530
rect 74690 -590 74760 -530
rect 74860 -590 74930 -530
rect 75030 -590 75100 -530
rect 75200 -590 75270 -530
rect 75370 -590 75440 -530
rect 75540 -590 75610 -530
rect 75710 -590 75780 -530
rect 75880 -590 75950 -530
rect 76050 -590 76120 -530
rect 76220 -590 76290 -530
rect 76390 -590 76460 -530
rect 76560 -590 76630 -530
rect 76730 -590 76800 -530
rect 76900 -590 76970 -530
rect 77070 -590 77140 -530
rect 77240 -590 77310 -530
rect 77410 -590 77480 -530
rect 77580 -590 77650 -530
rect 77750 -590 77820 -530
rect 77920 -590 77990 -530
rect 78090 -590 78160 -530
rect 78260 -590 78330 -530
rect 78430 -590 78500 -530
rect 78600 -590 78670 -530
rect 78770 -590 78840 -530
rect 78940 -590 79010 -530
rect 79110 -590 79180 -530
rect 79280 -590 79350 -530
rect 79450 -590 79520 -530
rect 79620 -590 79690 -530
rect 79790 -590 79860 -530
rect 79960 -590 80030 -530
rect 80130 -590 80200 -530
rect 80300 -590 80370 -530
rect 80470 -590 80540 -530
rect 80640 -590 80710 -530
rect 80810 -590 80880 -530
rect 80980 -590 81050 -530
rect 81150 -590 81220 -530
rect 81320 -590 81390 -530
rect 81490 -590 81560 -530
rect 81660 -590 81730 -530
rect 81830 -590 81900 -530
rect 82000 -590 82070 -530
rect 82170 -590 82240 -530
rect 82340 -590 82410 -530
rect 82510 -590 82580 -530
rect 82680 -590 82750 -530
rect 82850 -590 82920 -530
rect 83020 -590 83090 -530
rect 83190 -590 83260 -530
rect 83360 -590 83430 -530
rect 83530 -590 83600 -530
rect 83700 -590 83770 -530
rect 83870 -590 83940 -530
rect 84040 -590 84110 -530
rect 84210 -590 84280 -530
rect 84380 -590 84450 -530
rect 84550 -590 84620 -530
rect 84720 -590 84790 -530
rect 84890 -590 84960 -530
rect 85060 -590 85130 -530
rect 85230 -590 85300 -530
rect 85400 -590 85470 -530
rect 85570 -590 85640 -530
rect 85740 -590 85810 -530
rect 85910 -590 85980 -530
rect 86080 -590 86150 -530
rect 86250 -590 86320 -530
rect 86420 -590 86490 -530
rect 86590 -590 86660 -530
rect 86760 -590 86830 -530
rect 86930 -590 87000 -530
rect 87100 -590 87170 -530
rect 150 -730 210 -670
rect 490 -730 550 -670
rect 830 -730 890 -670
rect 1170 -730 1230 -670
rect 1510 -730 1570 -670
rect 1850 -730 1910 -670
rect 2190 -730 2250 -670
rect 2530 -730 2590 -670
rect 2870 -730 2930 -670
rect 3210 -730 3270 -670
rect 3550 -730 3610 -670
rect 3890 -730 3950 -670
rect 4230 -730 4290 -670
rect 4570 -730 4630 -670
rect 4910 -730 4970 -670
rect 5250 -730 5310 -670
rect 5590 -730 5650 -670
rect 5930 -730 5990 -670
rect 6270 -730 6330 -670
rect 6610 -730 6670 -670
rect 6950 -730 7010 -670
rect 7290 -730 7350 -670
rect 7630 -730 7690 -670
rect 7970 -730 8030 -670
rect 8310 -730 8370 -670
rect 8650 -730 8710 -670
rect 8990 -730 9050 -670
rect 9330 -730 9390 -670
rect 9670 -730 9730 -670
rect 10010 -730 10070 -670
rect 10350 -730 10410 -670
rect 10690 -730 10750 -670
rect 11030 -730 11090 -670
rect 11370 -730 11430 -670
rect 11710 -730 11770 -670
rect 12050 -730 12110 -670
rect 12390 -730 12450 -670
rect 12730 -730 12790 -670
rect 13070 -730 13130 -670
rect 13410 -730 13470 -670
rect 13750 -730 13810 -670
rect 14090 -730 14150 -670
rect 14430 -730 14490 -670
rect 14770 -730 14830 -670
rect 15110 -730 15170 -670
rect 15450 -730 15510 -670
rect 15790 -730 15850 -670
rect 16130 -730 16190 -670
rect 16470 -730 16530 -670
rect 16810 -730 16870 -670
rect 17150 -730 17210 -670
rect 17490 -730 17550 -670
rect 17830 -730 17890 -670
rect 18170 -730 18230 -670
rect 18510 -730 18570 -670
rect 18850 -730 18910 -670
rect 19190 -730 19250 -670
rect 19530 -730 19590 -670
rect 19870 -730 19930 -670
rect 20210 -730 20270 -670
rect 20550 -730 20610 -670
rect 20890 -730 20950 -670
rect 21230 -730 21290 -670
rect 21570 -730 21630 -670
rect 21910 -730 21970 -670
rect 22250 -730 22310 -670
rect 22590 -730 22650 -670
rect 22930 -730 22990 -670
rect 23270 -730 23330 -670
rect 23610 -730 23670 -670
rect 23950 -730 24010 -670
rect 24290 -730 24350 -670
rect 24630 -730 24690 -670
rect 24970 -730 25030 -670
rect 25310 -730 25370 -670
rect 25650 -730 25710 -670
rect 25990 -730 26050 -670
rect 26330 -730 26390 -670
rect 26670 -730 26730 -670
rect 27010 -730 27070 -670
rect 27350 -730 27410 -670
rect 27690 -730 27750 -670
rect 28030 -730 28090 -670
rect 28370 -730 28430 -670
rect 28710 -730 28770 -670
rect 29050 -730 29110 -670
rect 29390 -730 29450 -670
rect 29730 -730 29790 -670
rect 30070 -730 30130 -670
rect 30410 -730 30470 -670
rect 30750 -730 30810 -670
rect 31090 -730 31150 -670
rect 31430 -730 31490 -670
rect 31770 -730 31830 -670
rect 32110 -730 32170 -670
rect 32450 -730 32510 -670
rect 32790 -730 32850 -670
rect 33130 -730 33190 -670
rect 33470 -730 33530 -670
rect 33810 -730 33870 -670
rect 34150 -730 34210 -670
rect 34490 -730 34550 -670
rect 34830 -730 34890 -670
rect 35170 -730 35230 -670
rect 35510 -730 35570 -670
rect 35850 -730 35910 -670
rect 36190 -730 36250 -670
rect 36530 -730 36590 -670
rect 36870 -730 36930 -670
rect 37210 -730 37270 -670
rect 37550 -730 37610 -670
rect 37890 -730 37950 -670
rect 38230 -730 38290 -670
rect 38570 -730 38630 -670
rect 38910 -730 38970 -670
rect 39250 -730 39310 -670
rect 39590 -730 39650 -670
rect 39930 -730 39990 -670
rect 40270 -730 40330 -670
rect 40610 -730 40670 -670
rect 40950 -730 41010 -670
rect 41290 -730 41350 -670
rect 41630 -730 41690 -670
rect 41970 -730 42030 -670
rect 42310 -730 42370 -670
rect 42650 -730 42710 -670
rect 42990 -730 43050 -670
rect 43330 -730 43390 -670
rect 43670 -730 43730 -670
rect 44010 -730 44070 -670
rect 44350 -730 44410 -670
rect 44690 -730 44750 -670
rect 45030 -730 45090 -670
rect 45370 -730 45430 -670
rect 45710 -730 45770 -670
rect 46050 -730 46110 -670
rect 46390 -730 46450 -670
rect 46730 -730 46790 -670
rect 47070 -730 47130 -670
rect 47410 -730 47470 -670
rect 47750 -730 47810 -670
rect 48090 -730 48150 -670
rect 48430 -730 48490 -670
rect 48770 -730 48830 -670
rect 49110 -730 49170 -670
rect 49450 -730 49510 -670
rect 49790 -730 49850 -670
rect 50130 -730 50190 -670
rect 50470 -730 50530 -670
rect 50810 -730 50870 -670
rect 51150 -730 51210 -670
rect 51490 -730 51550 -670
rect 51830 -730 51890 -670
rect 52170 -730 52230 -670
rect 52510 -730 52570 -670
rect 52850 -730 52910 -670
rect 53190 -730 53250 -670
rect 53530 -730 53590 -670
rect 53870 -730 53930 -670
rect 54210 -730 54270 -670
rect 54550 -730 54610 -670
rect 54890 -730 54950 -670
rect 55230 -730 55290 -670
rect 55570 -730 55630 -670
rect 55910 -730 55970 -670
rect 56250 -730 56310 -670
rect 56590 -730 56650 -670
rect 56930 -730 56990 -670
rect 57270 -730 57330 -670
rect 57610 -730 57670 -670
rect 57950 -730 58010 -670
rect 58290 -730 58350 -670
rect 58630 -730 58690 -670
rect 58970 -730 59030 -670
rect 59310 -730 59370 -670
rect 59650 -730 59710 -670
rect 59990 -730 60050 -670
rect 60330 -730 60390 -670
rect 60670 -730 60730 -670
rect 61010 -730 61070 -670
rect 61350 -730 61410 -670
rect 61690 -730 61750 -670
rect 62030 -730 62090 -670
rect 62370 -730 62430 -670
rect 62710 -730 62770 -670
rect 63050 -730 63110 -670
rect 63390 -730 63450 -670
rect 63730 -730 63790 -670
rect 64070 -730 64130 -670
rect 64410 -730 64470 -670
rect 64750 -730 64810 -670
rect 65090 -730 65150 -670
rect 65430 -730 65490 -670
rect 65770 -730 65830 -670
rect 66110 -730 66170 -670
rect 66450 -730 66510 -670
rect 66790 -730 66850 -670
rect 67130 -730 67190 -670
rect 67470 -730 67530 -670
rect 67810 -730 67870 -670
rect 68150 -730 68210 -670
rect 68490 -730 68550 -670
rect 68830 -730 68890 -670
rect 69170 -730 69230 -670
rect 69510 -730 69570 -670
rect 69850 -730 69910 -670
rect 70190 -730 70250 -670
rect 70530 -730 70590 -670
rect 70870 -730 70930 -670
rect 71210 -730 71270 -670
rect 71550 -730 71610 -670
rect 71890 -730 71950 -670
rect 72230 -730 72290 -670
rect 72570 -730 72630 -670
rect 72910 -730 72970 -670
rect 73250 -730 73310 -670
rect 73590 -730 73650 -670
rect 73930 -730 73990 -670
rect 74270 -730 74330 -670
rect 74610 -730 74670 -670
rect 74950 -730 75010 -670
rect 75290 -730 75350 -670
rect 75630 -730 75690 -670
rect 75970 -730 76030 -670
rect 76310 -730 76370 -670
rect 76650 -730 76710 -670
rect 76990 -730 77050 -670
rect 77330 -730 77390 -670
rect 77670 -730 77730 -670
rect 78010 -730 78070 -670
rect 78350 -730 78410 -670
rect 78690 -730 78750 -670
rect 79030 -730 79090 -670
rect 79370 -730 79430 -670
rect 79710 -730 79770 -670
rect 80050 -730 80110 -670
rect 80390 -730 80450 -670
rect 80730 -730 80790 -670
rect 81070 -730 81130 -670
rect 81410 -730 81470 -670
rect 81750 -730 81810 -670
rect 82090 -730 82150 -670
rect 82430 -730 82490 -670
rect 82770 -730 82830 -670
rect 83110 -730 83170 -670
rect 83450 -730 83510 -670
rect 83790 -730 83850 -670
rect 84130 -730 84190 -670
rect 84470 -730 84530 -670
rect 84810 -730 84870 -670
rect 85150 -730 85210 -670
rect 85490 -730 85550 -670
rect 85830 -730 85890 -670
rect 86170 -730 86230 -670
rect 86510 -730 86570 -670
rect 86850 -730 86910 -670
rect 87190 -730 87250 -670
rect 320 -950 380 -880
rect 150 -1160 210 -1100
rect 660 -950 720 -880
rect 490 -1160 550 -1100
rect 1000 -950 1060 -880
rect 830 -1160 890 -1100
rect 1340 -950 1400 -880
rect 1170 -1160 1230 -1100
rect 1680 -950 1740 -880
rect 1510 -1160 1570 -1100
rect 2020 -950 2080 -880
rect 1850 -1160 1910 -1100
rect 2360 -950 2420 -880
rect 2190 -1160 2250 -1100
rect 2700 -950 2760 -880
rect 2530 -1160 2590 -1100
rect 3040 -950 3100 -880
rect 2870 -1160 2930 -1100
rect 3380 -950 3440 -880
rect 3210 -1160 3270 -1100
rect 3720 -950 3780 -880
rect 3550 -1160 3610 -1100
rect 4060 -950 4120 -880
rect 3890 -1160 3950 -1100
rect 4400 -950 4460 -880
rect 4230 -1160 4290 -1100
rect 4740 -950 4800 -880
rect 4570 -1160 4630 -1100
rect 5080 -950 5140 -880
rect 4910 -1160 4970 -1100
rect 5420 -950 5480 -880
rect 5250 -1160 5310 -1100
rect 5760 -950 5820 -880
rect 5590 -1160 5650 -1100
rect 6100 -950 6160 -880
rect 5930 -1160 5990 -1100
rect 6440 -950 6500 -880
rect 6270 -1160 6330 -1100
rect 6780 -950 6840 -880
rect 6610 -1160 6670 -1100
rect 7120 -950 7180 -880
rect 6950 -1160 7010 -1100
rect 7460 -950 7520 -880
rect 7290 -1160 7350 -1100
rect 7800 -950 7860 -880
rect 7630 -1160 7690 -1100
rect 8140 -950 8200 -880
rect 7970 -1160 8030 -1100
rect 8480 -950 8540 -880
rect 8310 -1160 8370 -1100
rect 8820 -950 8880 -880
rect 8650 -1160 8710 -1100
rect 9160 -950 9220 -880
rect 8990 -1160 9050 -1100
rect 9500 -950 9560 -880
rect 9330 -1160 9390 -1100
rect 9840 -950 9900 -880
rect 9670 -1160 9730 -1100
rect 10180 -950 10240 -880
rect 10010 -1160 10070 -1100
rect 10520 -950 10580 -880
rect 10350 -1160 10410 -1100
rect 10860 -950 10920 -880
rect 10690 -1160 10750 -1100
rect 11200 -950 11260 -880
rect 11030 -1160 11090 -1100
rect 11540 -950 11600 -880
rect 11370 -1160 11430 -1100
rect 11880 -950 11940 -880
rect 11710 -1160 11770 -1100
rect 12220 -950 12280 -880
rect 12050 -1160 12110 -1100
rect 12560 -950 12620 -880
rect 12390 -1160 12450 -1100
rect 12900 -950 12960 -880
rect 12730 -1160 12790 -1100
rect 13240 -950 13300 -880
rect 13070 -1160 13130 -1100
rect 13580 -950 13640 -880
rect 13410 -1160 13470 -1100
rect 13920 -950 13980 -880
rect 13750 -1160 13810 -1100
rect 14260 -950 14320 -880
rect 14090 -1160 14150 -1100
rect 14600 -950 14660 -880
rect 14430 -1160 14490 -1100
rect 14940 -950 15000 -880
rect 14770 -1160 14830 -1100
rect 15280 -950 15340 -880
rect 15110 -1160 15170 -1100
rect 15620 -950 15680 -880
rect 15450 -1160 15510 -1100
rect 15960 -950 16020 -880
rect 15790 -1160 15850 -1100
rect 16300 -950 16360 -880
rect 16130 -1160 16190 -1100
rect 16640 -950 16700 -880
rect 16470 -1160 16530 -1100
rect 16980 -950 17040 -880
rect 16810 -1160 16870 -1100
rect 17320 -950 17380 -880
rect 17150 -1160 17210 -1100
rect 17660 -950 17720 -880
rect 17490 -1160 17550 -1100
rect 18000 -950 18060 -880
rect 17830 -1160 17890 -1100
rect 18340 -950 18400 -880
rect 18170 -1160 18230 -1100
rect 18680 -950 18740 -880
rect 18510 -1160 18570 -1100
rect 19020 -950 19080 -880
rect 18850 -1160 18910 -1100
rect 19360 -950 19420 -880
rect 19190 -1160 19250 -1100
rect 19700 -950 19760 -880
rect 19530 -1160 19590 -1100
rect 20040 -950 20100 -880
rect 19870 -1160 19930 -1100
rect 20380 -950 20440 -880
rect 20210 -1160 20270 -1100
rect 20720 -950 20780 -880
rect 20550 -1160 20610 -1100
rect 21060 -950 21120 -880
rect 20890 -1160 20950 -1100
rect 21400 -950 21460 -880
rect 21230 -1160 21290 -1100
rect 21740 -950 21800 -880
rect 21570 -1160 21630 -1100
rect 22080 -950 22140 -880
rect 21910 -1160 21970 -1100
rect 22420 -950 22480 -880
rect 22250 -1160 22310 -1100
rect 22760 -950 22820 -880
rect 22590 -1160 22650 -1100
rect 23100 -950 23160 -880
rect 22930 -1160 22990 -1100
rect 23440 -950 23500 -880
rect 23270 -1160 23330 -1100
rect 23780 -950 23840 -880
rect 23610 -1160 23670 -1100
rect 24120 -950 24180 -880
rect 23950 -1160 24010 -1100
rect 24460 -950 24520 -880
rect 24290 -1160 24350 -1100
rect 24800 -950 24860 -880
rect 24630 -1160 24690 -1100
rect 25140 -950 25200 -880
rect 24970 -1160 25030 -1100
rect 25480 -950 25540 -880
rect 25310 -1160 25370 -1100
rect 25820 -950 25880 -880
rect 25650 -1160 25710 -1100
rect 26160 -950 26220 -880
rect 25990 -1160 26050 -1100
rect 26500 -950 26560 -880
rect 26330 -1160 26390 -1100
rect 26840 -950 26900 -880
rect 26670 -1160 26730 -1100
rect 27180 -950 27240 -880
rect 27010 -1160 27070 -1100
rect 27520 -950 27580 -880
rect 27350 -1160 27410 -1100
rect 27860 -950 27920 -880
rect 27690 -1160 27750 -1100
rect 28200 -950 28260 -880
rect 28030 -1160 28090 -1100
rect 28540 -950 28600 -880
rect 28370 -1160 28430 -1100
rect 28880 -950 28940 -880
rect 28710 -1160 28770 -1100
rect 29220 -950 29280 -880
rect 29050 -1160 29110 -1100
rect 29560 -950 29620 -880
rect 29390 -1160 29450 -1100
rect 29900 -950 29960 -880
rect 29730 -1160 29790 -1100
rect 30240 -950 30300 -880
rect 30070 -1160 30130 -1100
rect 30580 -950 30640 -880
rect 30410 -1160 30470 -1100
rect 30920 -950 30980 -880
rect 30750 -1160 30810 -1100
rect 31260 -950 31320 -880
rect 31090 -1160 31150 -1100
rect 31600 -950 31660 -880
rect 31430 -1160 31490 -1100
rect 31940 -950 32000 -880
rect 31770 -1160 31830 -1100
rect 32280 -950 32340 -880
rect 32110 -1160 32170 -1100
rect 32620 -950 32680 -880
rect 32450 -1160 32510 -1100
rect 32960 -950 33020 -880
rect 32790 -1160 32850 -1100
rect 33300 -950 33360 -880
rect 33130 -1160 33190 -1100
rect 33640 -950 33700 -880
rect 33470 -1160 33530 -1100
rect 33980 -950 34040 -880
rect 33810 -1160 33870 -1100
rect 34320 -950 34380 -880
rect 34150 -1160 34210 -1100
rect 34660 -950 34720 -880
rect 34490 -1160 34550 -1100
rect 35000 -950 35060 -880
rect 34830 -1160 34890 -1100
rect 35340 -950 35400 -880
rect 35170 -1160 35230 -1100
rect 35680 -950 35740 -880
rect 35510 -1160 35570 -1100
rect 36020 -950 36080 -880
rect 35850 -1160 35910 -1100
rect 36360 -950 36420 -880
rect 36190 -1160 36250 -1100
rect 36700 -950 36760 -880
rect 36530 -1160 36590 -1100
rect 37040 -950 37100 -880
rect 36870 -1160 36930 -1100
rect 37380 -950 37440 -880
rect 37210 -1160 37270 -1100
rect 37720 -950 37780 -880
rect 37550 -1160 37610 -1100
rect 38060 -950 38120 -880
rect 37890 -1160 37950 -1100
rect 38400 -950 38460 -880
rect 38230 -1160 38290 -1100
rect 38740 -950 38800 -880
rect 38570 -1160 38630 -1100
rect 39080 -950 39140 -880
rect 38910 -1160 38970 -1100
rect 39420 -950 39480 -880
rect 39250 -1160 39310 -1100
rect 39760 -950 39820 -880
rect 39590 -1160 39650 -1100
rect 40100 -950 40160 -880
rect 39930 -1160 39990 -1100
rect 40440 -950 40500 -880
rect 40270 -1160 40330 -1100
rect 40780 -950 40840 -880
rect 40610 -1160 40670 -1100
rect 41120 -950 41180 -880
rect 40950 -1160 41010 -1100
rect 41460 -950 41520 -880
rect 41290 -1160 41350 -1100
rect 41800 -950 41860 -880
rect 41630 -1160 41690 -1100
rect 42140 -950 42200 -880
rect 41970 -1160 42030 -1100
rect 42480 -950 42540 -880
rect 42310 -1160 42370 -1100
rect 42820 -950 42880 -880
rect 42650 -1160 42710 -1100
rect 43160 -950 43220 -880
rect 42990 -1160 43050 -1100
rect 43500 -950 43560 -880
rect 43330 -1160 43390 -1100
rect 43840 -950 43900 -880
rect 43670 -1160 43730 -1100
rect 44180 -950 44240 -880
rect 44010 -1160 44070 -1100
rect 44520 -950 44580 -880
rect 44350 -1160 44410 -1100
rect 44860 -950 44920 -880
rect 44690 -1160 44750 -1100
rect 45200 -950 45260 -880
rect 45030 -1160 45090 -1100
rect 45540 -950 45600 -880
rect 45370 -1160 45430 -1100
rect 45880 -950 45940 -880
rect 45710 -1160 45770 -1100
rect 46220 -950 46280 -880
rect 46050 -1160 46110 -1100
rect 46560 -950 46620 -880
rect 46390 -1160 46450 -1100
rect 46900 -950 46960 -880
rect 46730 -1160 46790 -1100
rect 47240 -950 47300 -880
rect 47070 -1160 47130 -1100
rect 47580 -950 47640 -880
rect 47410 -1160 47470 -1100
rect 47920 -950 47980 -880
rect 47750 -1160 47810 -1100
rect 48260 -950 48320 -880
rect 48090 -1160 48150 -1100
rect 48600 -950 48660 -880
rect 48430 -1160 48490 -1100
rect 48940 -950 49000 -880
rect 48770 -1160 48830 -1100
rect 49280 -950 49340 -880
rect 49110 -1160 49170 -1100
rect 49620 -950 49680 -880
rect 49450 -1160 49510 -1100
rect 49960 -950 50020 -880
rect 49790 -1160 49850 -1100
rect 50300 -950 50360 -880
rect 50130 -1160 50190 -1100
rect 50640 -950 50700 -880
rect 50470 -1160 50530 -1100
rect 50980 -950 51040 -880
rect 50810 -1160 50870 -1100
rect 51320 -950 51380 -880
rect 51150 -1160 51210 -1100
rect 51660 -950 51720 -880
rect 51490 -1160 51550 -1100
rect 52000 -950 52060 -880
rect 51830 -1160 51890 -1100
rect 52340 -950 52400 -880
rect 52170 -1160 52230 -1100
rect 52680 -950 52740 -880
rect 52510 -1160 52570 -1100
rect 53020 -950 53080 -880
rect 52850 -1160 52910 -1100
rect 53360 -950 53420 -880
rect 53190 -1160 53250 -1100
rect 53700 -950 53760 -880
rect 53530 -1160 53590 -1100
rect 54040 -950 54100 -880
rect 53870 -1160 53930 -1100
rect 54380 -950 54440 -880
rect 54210 -1160 54270 -1100
rect 54720 -950 54780 -880
rect 54550 -1160 54610 -1100
rect 55060 -950 55120 -880
rect 54890 -1160 54950 -1100
rect 55400 -950 55460 -880
rect 55230 -1160 55290 -1100
rect 55740 -950 55800 -880
rect 55570 -1160 55630 -1100
rect 56080 -950 56140 -880
rect 55910 -1160 55970 -1100
rect 56420 -950 56480 -880
rect 56250 -1160 56310 -1100
rect 56760 -950 56820 -880
rect 56590 -1160 56650 -1100
rect 57100 -950 57160 -880
rect 56930 -1160 56990 -1100
rect 57440 -950 57500 -880
rect 57270 -1160 57330 -1100
rect 57780 -950 57840 -880
rect 57610 -1160 57670 -1100
rect 58120 -950 58180 -880
rect 57950 -1160 58010 -1100
rect 58460 -950 58520 -880
rect 58290 -1160 58350 -1100
rect 58800 -950 58860 -880
rect 58630 -1160 58690 -1100
rect 59140 -950 59200 -880
rect 58970 -1160 59030 -1100
rect 59480 -950 59540 -880
rect 59310 -1160 59370 -1100
rect 59820 -950 59880 -880
rect 59650 -1160 59710 -1100
rect 60160 -950 60220 -880
rect 59990 -1160 60050 -1100
rect 60500 -950 60560 -880
rect 60330 -1160 60390 -1100
rect 60840 -950 60900 -880
rect 60670 -1160 60730 -1100
rect 61180 -950 61240 -880
rect 61010 -1160 61070 -1100
rect 61520 -950 61580 -880
rect 61350 -1160 61410 -1100
rect 61860 -950 61920 -880
rect 61690 -1160 61750 -1100
rect 62200 -950 62260 -880
rect 62030 -1160 62090 -1100
rect 62540 -950 62600 -880
rect 62370 -1160 62430 -1100
rect 62880 -950 62940 -880
rect 62710 -1160 62770 -1100
rect 63220 -950 63280 -880
rect 63050 -1160 63110 -1100
rect 63560 -950 63620 -880
rect 63390 -1160 63450 -1100
rect 63900 -950 63960 -880
rect 63730 -1160 63790 -1100
rect 64240 -950 64300 -880
rect 64070 -1160 64130 -1100
rect 64580 -950 64640 -880
rect 64410 -1160 64470 -1100
rect 64920 -950 64980 -880
rect 64750 -1160 64810 -1100
rect 65260 -950 65320 -880
rect 65090 -1160 65150 -1100
rect 65600 -950 65660 -880
rect 65430 -1160 65490 -1100
rect 65940 -950 66000 -880
rect 65770 -1160 65830 -1100
rect 66280 -950 66340 -880
rect 66110 -1160 66170 -1100
rect 66620 -950 66680 -880
rect 66450 -1160 66510 -1100
rect 66960 -950 67020 -880
rect 66790 -1160 66850 -1100
rect 67300 -950 67360 -880
rect 67130 -1160 67190 -1100
rect 67640 -950 67700 -880
rect 67470 -1160 67530 -1100
rect 67980 -950 68040 -880
rect 67810 -1160 67870 -1100
rect 68320 -950 68380 -880
rect 68150 -1160 68210 -1100
rect 68660 -950 68720 -880
rect 68490 -1160 68550 -1100
rect 69000 -950 69060 -880
rect 68830 -1160 68890 -1100
rect 69340 -950 69400 -880
rect 69170 -1160 69230 -1100
rect 69680 -950 69740 -880
rect 69510 -1160 69570 -1100
rect 70020 -950 70080 -880
rect 69850 -1160 69910 -1100
rect 70360 -950 70420 -880
rect 70190 -1160 70250 -1100
rect 70700 -950 70760 -880
rect 70530 -1160 70590 -1100
rect 71040 -950 71100 -880
rect 70870 -1160 70930 -1100
rect 71380 -950 71440 -880
rect 71210 -1160 71270 -1100
rect 71720 -950 71780 -880
rect 71550 -1160 71610 -1100
rect 72060 -950 72120 -880
rect 71890 -1160 71950 -1100
rect 72400 -950 72460 -880
rect 72230 -1160 72290 -1100
rect 72740 -950 72800 -880
rect 72570 -1160 72630 -1100
rect 73080 -950 73140 -880
rect 72910 -1160 72970 -1100
rect 73420 -950 73480 -880
rect 73250 -1160 73310 -1100
rect 73760 -950 73820 -880
rect 73590 -1160 73650 -1100
rect 74100 -950 74160 -880
rect 73930 -1160 73990 -1100
rect 74440 -950 74500 -880
rect 74270 -1160 74330 -1100
rect 74780 -950 74840 -880
rect 74610 -1160 74670 -1100
rect 75120 -950 75180 -880
rect 74950 -1160 75010 -1100
rect 75460 -950 75520 -880
rect 75290 -1160 75350 -1100
rect 75800 -950 75860 -880
rect 75630 -1160 75690 -1100
rect 76140 -950 76200 -880
rect 75970 -1160 76030 -1100
rect 76480 -950 76540 -880
rect 76310 -1160 76370 -1100
rect 76820 -950 76880 -880
rect 76650 -1160 76710 -1100
rect 77160 -950 77220 -880
rect 76990 -1160 77050 -1100
rect 77500 -950 77560 -880
rect 77330 -1160 77390 -1100
rect 77840 -950 77900 -880
rect 77670 -1160 77730 -1100
rect 78180 -950 78240 -880
rect 78010 -1160 78070 -1100
rect 78520 -950 78580 -880
rect 78350 -1160 78410 -1100
rect 78860 -950 78920 -880
rect 78690 -1160 78750 -1100
rect 79200 -950 79260 -880
rect 79030 -1160 79090 -1100
rect 79540 -950 79600 -880
rect 79370 -1160 79430 -1100
rect 79880 -950 79940 -880
rect 79710 -1160 79770 -1100
rect 80220 -950 80280 -880
rect 80050 -1160 80110 -1100
rect 80560 -950 80620 -880
rect 80390 -1160 80450 -1100
rect 80900 -950 80960 -880
rect 80730 -1160 80790 -1100
rect 81240 -950 81300 -880
rect 81070 -1160 81130 -1100
rect 81580 -950 81640 -880
rect 81410 -1160 81470 -1100
rect 81920 -950 81980 -880
rect 81750 -1160 81810 -1100
rect 82260 -950 82320 -880
rect 82090 -1160 82150 -1100
rect 82600 -950 82660 -880
rect 82430 -1160 82490 -1100
rect 82940 -950 83000 -880
rect 82770 -1160 82830 -1100
rect 83280 -950 83340 -880
rect 83110 -1160 83170 -1100
rect 83620 -950 83680 -880
rect 83450 -1160 83510 -1100
rect 83960 -950 84020 -880
rect 83790 -1160 83850 -1100
rect 84300 -950 84360 -880
rect 84130 -1160 84190 -1100
rect 84640 -950 84700 -880
rect 84470 -1160 84530 -1100
rect 84980 -950 85040 -880
rect 84810 -1160 84870 -1100
rect 85320 -950 85380 -880
rect 85150 -1160 85210 -1100
rect 85660 -950 85720 -880
rect 85490 -1160 85550 -1100
rect 86000 -950 86060 -880
rect 85830 -1160 85890 -1100
rect 86340 -950 86400 -880
rect 86170 -1160 86230 -1100
rect 86680 -950 86740 -880
rect 86510 -1160 86570 -1100
rect 87020 -950 87080 -880
rect 86850 -1160 86910 -1100
rect 87190 -1160 87250 -1100
rect 150 -1360 210 -1300
rect 490 -1360 550 -1300
rect 830 -1360 890 -1300
rect 1170 -1360 1230 -1300
rect 1510 -1360 1570 -1300
rect 1850 -1360 1910 -1300
rect 2190 -1360 2250 -1300
rect 2530 -1360 2590 -1300
rect 2870 -1360 2930 -1300
rect 3210 -1360 3270 -1300
rect 3550 -1360 3610 -1300
rect 3890 -1360 3950 -1300
rect 4230 -1360 4290 -1300
rect 4570 -1360 4630 -1300
rect 4910 -1360 4970 -1300
rect 5250 -1360 5310 -1300
rect 5590 -1360 5650 -1300
rect 5930 -1360 5990 -1300
rect 6270 -1360 6330 -1300
rect 6610 -1360 6670 -1300
rect 6950 -1360 7010 -1300
rect 7290 -1360 7350 -1300
rect 7630 -1360 7690 -1300
rect 7970 -1360 8030 -1300
rect 8310 -1360 8370 -1300
rect 8650 -1360 8710 -1300
rect 8990 -1360 9050 -1300
rect 9330 -1360 9390 -1300
rect 9670 -1360 9730 -1300
rect 10010 -1360 10070 -1300
rect 10350 -1360 10410 -1300
rect 10690 -1360 10750 -1300
rect 11030 -1360 11090 -1300
rect 11370 -1360 11430 -1300
rect 11710 -1360 11770 -1300
rect 12050 -1360 12110 -1300
rect 12390 -1360 12450 -1300
rect 12730 -1360 12790 -1300
rect 13070 -1360 13130 -1300
rect 13410 -1360 13470 -1300
rect 13750 -1360 13810 -1300
rect 14090 -1360 14150 -1300
rect 14430 -1360 14490 -1300
rect 14770 -1360 14830 -1300
rect 15110 -1360 15170 -1300
rect 15450 -1360 15510 -1300
rect 15790 -1360 15850 -1300
rect 16130 -1360 16190 -1300
rect 16470 -1360 16530 -1300
rect 16810 -1360 16870 -1300
rect 17150 -1360 17210 -1300
rect 17490 -1360 17550 -1300
rect 17830 -1360 17890 -1300
rect 18170 -1360 18230 -1300
rect 18510 -1360 18570 -1300
rect 18850 -1360 18910 -1300
rect 19190 -1360 19250 -1300
rect 19530 -1360 19590 -1300
rect 19870 -1360 19930 -1300
rect 20210 -1360 20270 -1300
rect 20550 -1360 20610 -1300
rect 20890 -1360 20950 -1300
rect 21230 -1360 21290 -1300
rect 21570 -1360 21630 -1300
rect 21910 -1360 21970 -1300
rect 22250 -1360 22310 -1300
rect 22590 -1360 22650 -1300
rect 22930 -1360 22990 -1300
rect 23270 -1360 23330 -1300
rect 23610 -1360 23670 -1300
rect 23950 -1360 24010 -1300
rect 24290 -1360 24350 -1300
rect 24630 -1360 24690 -1300
rect 24970 -1360 25030 -1300
rect 25310 -1360 25370 -1300
rect 25650 -1360 25710 -1300
rect 25990 -1360 26050 -1300
rect 26330 -1360 26390 -1300
rect 26670 -1360 26730 -1300
rect 27010 -1360 27070 -1300
rect 27350 -1360 27410 -1300
rect 27690 -1360 27750 -1300
rect 28030 -1360 28090 -1300
rect 28370 -1360 28430 -1300
rect 28710 -1360 28770 -1300
rect 29050 -1360 29110 -1300
rect 29390 -1360 29450 -1300
rect 29730 -1360 29790 -1300
rect 30070 -1360 30130 -1300
rect 30410 -1360 30470 -1300
rect 30750 -1360 30810 -1300
rect 31090 -1360 31150 -1300
rect 31430 -1360 31490 -1300
rect 31770 -1360 31830 -1300
rect 32110 -1360 32170 -1300
rect 32450 -1360 32510 -1300
rect 32790 -1360 32850 -1300
rect 33130 -1360 33190 -1300
rect 33470 -1360 33530 -1300
rect 33810 -1360 33870 -1300
rect 34150 -1360 34210 -1300
rect 34490 -1360 34550 -1300
rect 34830 -1360 34890 -1300
rect 35170 -1360 35230 -1300
rect 35510 -1360 35570 -1300
rect 35850 -1360 35910 -1300
rect 36190 -1360 36250 -1300
rect 36530 -1360 36590 -1300
rect 36870 -1360 36930 -1300
rect 37210 -1360 37270 -1300
rect 37550 -1360 37610 -1300
rect 37890 -1360 37950 -1300
rect 38230 -1360 38290 -1300
rect 38570 -1360 38630 -1300
rect 38910 -1360 38970 -1300
rect 39250 -1360 39310 -1300
rect 39590 -1360 39650 -1300
rect 39930 -1360 39990 -1300
rect 40270 -1360 40330 -1300
rect 40610 -1360 40670 -1300
rect 40950 -1360 41010 -1300
rect 41290 -1360 41350 -1300
rect 41630 -1360 41690 -1300
rect 41970 -1360 42030 -1300
rect 42310 -1360 42370 -1300
rect 42650 -1360 42710 -1300
rect 42990 -1360 43050 -1300
rect 43330 -1360 43390 -1300
rect 43670 -1360 43730 -1300
rect 44010 -1360 44070 -1300
rect 44350 -1360 44410 -1300
rect 44690 -1360 44750 -1300
rect 45030 -1360 45090 -1300
rect 45370 -1360 45430 -1300
rect 45710 -1360 45770 -1300
rect 46050 -1360 46110 -1300
rect 46390 -1360 46450 -1300
rect 46730 -1360 46790 -1300
rect 47070 -1360 47130 -1300
rect 47410 -1360 47470 -1300
rect 47750 -1360 47810 -1300
rect 48090 -1360 48150 -1300
rect 48430 -1360 48490 -1300
rect 48770 -1360 48830 -1300
rect 49110 -1360 49170 -1300
rect 49450 -1360 49510 -1300
rect 49790 -1360 49850 -1300
rect 50130 -1360 50190 -1300
rect 50470 -1360 50530 -1300
rect 50810 -1360 50870 -1300
rect 51150 -1360 51210 -1300
rect 51490 -1360 51550 -1300
rect 51830 -1360 51890 -1300
rect 52170 -1360 52230 -1300
rect 52510 -1360 52570 -1300
rect 52850 -1360 52910 -1300
rect 53190 -1360 53250 -1300
rect 53530 -1360 53590 -1300
rect 53870 -1360 53930 -1300
rect 54210 -1360 54270 -1300
rect 54550 -1360 54610 -1300
rect 54890 -1360 54950 -1300
rect 55230 -1360 55290 -1300
rect 55570 -1360 55630 -1300
rect 55910 -1360 55970 -1300
rect 56250 -1360 56310 -1300
rect 56590 -1360 56650 -1300
rect 56930 -1360 56990 -1300
rect 57270 -1360 57330 -1300
rect 57610 -1360 57670 -1300
rect 57950 -1360 58010 -1300
rect 58290 -1360 58350 -1300
rect 58630 -1360 58690 -1300
rect 58970 -1360 59030 -1300
rect 59310 -1360 59370 -1300
rect 59650 -1360 59710 -1300
rect 59990 -1360 60050 -1300
rect 60330 -1360 60390 -1300
rect 60670 -1360 60730 -1300
rect 61010 -1360 61070 -1300
rect 61350 -1360 61410 -1300
rect 61690 -1360 61750 -1300
rect 62030 -1360 62090 -1300
rect 62370 -1360 62430 -1300
rect 62710 -1360 62770 -1300
rect 63050 -1360 63110 -1300
rect 63390 -1360 63450 -1300
rect 63730 -1360 63790 -1300
rect 64070 -1360 64130 -1300
rect 64410 -1360 64470 -1300
rect 64750 -1360 64810 -1300
rect 65090 -1360 65150 -1300
rect 65430 -1360 65490 -1300
rect 65770 -1360 65830 -1300
rect 66110 -1360 66170 -1300
rect 66450 -1360 66510 -1300
rect 66790 -1360 66850 -1300
rect 67130 -1360 67190 -1300
rect 67470 -1360 67530 -1300
rect 67810 -1360 67870 -1300
rect 68150 -1360 68210 -1300
rect 68490 -1360 68550 -1300
rect 68830 -1360 68890 -1300
rect 69170 -1360 69230 -1300
rect 69510 -1360 69570 -1300
rect 69850 -1360 69910 -1300
rect 70190 -1360 70250 -1300
rect 70530 -1360 70590 -1300
rect 70870 -1360 70930 -1300
rect 71210 -1360 71270 -1300
rect 71550 -1360 71610 -1300
rect 71890 -1360 71950 -1300
rect 72230 -1360 72290 -1300
rect 72570 -1360 72630 -1300
rect 72910 -1360 72970 -1300
rect 73250 -1360 73310 -1300
rect 73590 -1360 73650 -1300
rect 73930 -1360 73990 -1300
rect 74270 -1360 74330 -1300
rect 74610 -1360 74670 -1300
rect 74950 -1360 75010 -1300
rect 75290 -1360 75350 -1300
rect 75630 -1360 75690 -1300
rect 75970 -1360 76030 -1300
rect 76310 -1360 76370 -1300
rect 76650 -1360 76710 -1300
rect 76990 -1360 77050 -1300
rect 77330 -1360 77390 -1300
rect 77670 -1360 77730 -1300
rect 78010 -1360 78070 -1300
rect 78350 -1360 78410 -1300
rect 78690 -1360 78750 -1300
rect 79030 -1360 79090 -1300
rect 79370 -1360 79430 -1300
rect 79710 -1360 79770 -1300
rect 80050 -1360 80110 -1300
rect 80390 -1360 80450 -1300
rect 80730 -1360 80790 -1300
rect 81070 -1360 81130 -1300
rect 81410 -1360 81470 -1300
rect 81750 -1360 81810 -1300
rect 82090 -1360 82150 -1300
rect 82430 -1360 82490 -1300
rect 82770 -1360 82830 -1300
rect 83110 -1360 83170 -1300
rect 83450 -1360 83510 -1300
rect 83790 -1360 83850 -1300
rect 84130 -1360 84190 -1300
rect 84470 -1360 84530 -1300
rect 84810 -1360 84870 -1300
rect 85150 -1360 85210 -1300
rect 85490 -1360 85550 -1300
rect 85830 -1360 85890 -1300
rect 86170 -1360 86230 -1300
rect 86510 -1360 86570 -1300
rect 86850 -1360 86910 -1300
rect 87190 -1360 87250 -1300
rect 830 -1540 910 -1470
rect 5000 -1540 5080 -1470
rect 9030 -1540 9110 -1470
rect 13060 -1540 13140 -1470
rect 17100 -1540 17180 -1470
rect 21200 -1540 21280 -1470
rect 25310 -1540 25390 -1470
rect 29410 -1540 29490 -1470
rect 33440 -1540 33520 -1470
rect 37550 -1540 37630 -1470
rect 41650 -1540 41730 -1470
rect 47100 -1540 47180 -1470
rect 51180 -1540 51260 -1470
rect 55290 -1540 55370 -1470
rect 59320 -1540 59400 -1470
rect 63420 -1540 63500 -1470
rect 67530 -1540 67610 -1470
rect 71560 -1540 71640 -1470
rect 75810 -1540 75890 -1470
rect 79770 -1540 79850 -1470
rect 83950 -1540 84030 -1470
rect 86508 -1544 86588 -1474
<< metal2 >>
rect 1280 710 1410 730
rect 1280 650 1300 710
rect 1390 650 1410 710
rect 1280 630 1410 650
rect 6370 690 6510 710
rect 6370 630 6390 690
rect 6490 630 6510 690
rect 730 590 930 620
rect 730 520 790 590
rect 870 520 930 590
rect 730 490 930 520
rect 2110 590 2310 620
rect 2110 520 2170 590
rect 2250 520 2310 590
rect 2110 490 2310 520
rect 3490 590 3690 620
rect 3490 520 3550 590
rect 3630 520 3690 590
rect 3490 490 3690 520
rect 5150 590 5350 620
rect 6370 610 6510 630
rect 5150 520 5210 590
rect 5290 520 5350 590
rect 5150 490 5350 520
rect 7980 590 8180 620
rect 7980 520 8040 590
rect 8120 520 8180 590
rect 7980 490 8180 520
rect 10740 590 10940 620
rect 10740 520 10800 590
rect 10880 520 10940 590
rect 10740 490 10940 520
rect 13370 590 13570 620
rect 13370 520 13430 590
rect 13510 520 13570 590
rect 13370 490 13570 520
rect 16410 590 16610 620
rect 16410 520 16470 590
rect 16550 520 16610 590
rect 16410 490 16610 520
rect 20480 590 20680 620
rect 20480 520 20540 590
rect 20620 520 20680 590
rect 20480 490 20680 520
rect 24620 590 24820 620
rect 24620 520 24680 590
rect 24760 520 24820 590
rect 24620 490 24820 520
rect 28700 590 28900 620
rect 28700 520 28760 590
rect 28840 520 28900 590
rect 28700 490 28900 520
rect 32850 590 33050 620
rect 32850 520 32910 590
rect 32990 520 33050 590
rect 32850 490 33050 520
rect 36720 590 36920 620
rect 36720 520 36780 590
rect 36860 520 36920 590
rect 36720 490 36920 520
rect 40860 590 41060 620
rect 40860 520 40920 590
rect 41000 520 41060 590
rect 40860 490 41060 520
rect 44850 590 45050 620
rect 44850 520 44910 590
rect 44990 520 45050 590
rect 44850 490 45050 520
rect 48930 590 49130 620
rect 48930 520 48990 590
rect 49070 520 49130 590
rect 48930 490 49130 520
rect 53020 590 53220 620
rect 53020 520 53080 590
rect 53160 520 53220 590
rect 53020 490 53220 520
rect 57180 590 57380 620
rect 57180 520 57240 590
rect 57320 520 57380 590
rect 57180 490 57380 520
rect 10 410 110 430
rect 10 350 30 410
rect 90 350 110 410
rect 10 330 110 350
rect 430 410 530 430
rect 770 410 870 430
rect 1110 410 1210 430
rect 1500 410 1600 430
rect 1840 410 1940 430
rect 2180 410 2280 430
rect 2520 410 2620 430
rect 2860 410 2960 430
rect 3200 410 3300 430
rect 3540 410 3640 430
rect 3880 410 3980 430
rect 4220 410 4320 430
rect 4520 410 4620 430
rect 4860 410 4960 430
rect 5200 410 5300 430
rect 5540 410 5640 430
rect 5880 410 5980 430
rect 6220 410 6320 430
rect 6560 410 6660 430
rect 6900 410 7000 430
rect 7240 410 7340 430
rect 7580 410 7680 430
rect 7920 410 8020 430
rect 8260 410 8360 430
rect 8600 410 8700 430
rect 8940 410 9040 430
rect 9280 410 9380 430
rect 9620 410 9720 430
rect 9960 410 10060 430
rect 10300 410 10400 430
rect 10640 410 10740 430
rect 10980 410 11080 430
rect 11320 410 11420 430
rect 11660 410 11760 430
rect 12000 410 12100 430
rect 12340 410 12440 430
rect 12680 410 12780 430
rect 13020 410 13120 430
rect 13360 410 13460 430
rect 13700 410 13800 430
rect 14040 410 14140 430
rect 14380 410 14480 430
rect 14720 410 14820 430
rect 15060 410 15160 430
rect 15400 410 15500 430
rect 15700 410 15800 430
rect 16040 410 16140 430
rect 16380 410 16480 430
rect 16720 410 16820 430
rect 17060 410 17160 430
rect 17400 410 17500 430
rect 17740 410 17840 430
rect 18080 410 18180 430
rect 18420 410 18520 430
rect 18760 410 18860 430
rect 19100 410 19200 430
rect 19440 410 19540 430
rect 19780 410 19880 430
rect 20120 410 20220 430
rect 20460 410 20560 430
rect 20800 410 20900 430
rect 21140 410 21240 430
rect 21480 410 21580 430
rect 21820 410 21920 430
rect 22160 410 22260 430
rect 22500 410 22600 430
rect 22840 410 22940 430
rect 23180 410 23280 430
rect 23520 410 23620 430
rect 23860 410 23960 430
rect 24200 410 24300 430
rect 24540 410 24640 430
rect 24880 410 24980 430
rect 25220 410 25320 430
rect 25560 410 25660 430
rect 25900 410 26000 430
rect 26240 410 26340 430
rect 26580 410 26680 430
rect 26920 410 27020 430
rect 27260 410 27360 430
rect 27600 410 27700 430
rect 27940 410 28040 430
rect 28280 410 28380 430
rect 28620 410 28720 430
rect 28960 410 29060 430
rect 29300 410 29400 430
rect 29640 410 29740 430
rect 29980 410 30080 430
rect 30320 410 30420 430
rect 30660 410 30760 430
rect 31000 410 31100 430
rect 31340 410 31440 430
rect 31680 410 31780 430
rect 32020 410 32120 430
rect 32360 410 32460 430
rect 32700 410 32800 430
rect 33040 410 33140 430
rect 33380 410 33480 430
rect 33720 410 33820 430
rect 34060 410 34160 430
rect 34400 410 34500 430
rect 34740 410 34840 430
rect 35080 410 35180 430
rect 35420 410 35520 430
rect 35760 410 35860 430
rect 36100 410 36200 430
rect 36440 410 36540 430
rect 36780 410 36880 430
rect 37120 410 37220 430
rect 37460 410 37560 430
rect 37800 410 37900 430
rect 38140 410 38240 430
rect 38480 410 38580 430
rect 38820 410 38920 430
rect 39160 410 39260 430
rect 39500 410 39600 430
rect 39840 410 39940 430
rect 40180 410 40280 430
rect 40520 410 40620 430
rect 40860 410 40960 430
rect 41200 410 41300 430
rect 41540 410 41640 430
rect 41880 410 41980 430
rect 42220 410 42320 430
rect 42560 410 42660 430
rect 42900 410 43000 430
rect 43240 410 43340 430
rect 43580 410 43680 430
rect 43920 410 44020 430
rect 44260 410 44360 430
rect 44600 410 44700 430
rect 44940 410 45040 430
rect 45280 410 45380 430
rect 45620 410 45720 430
rect 45960 410 46060 430
rect 46300 410 46400 430
rect 46640 410 46740 430
rect 46980 410 47080 430
rect 47320 410 47420 430
rect 47660 410 47760 430
rect 48000 410 48100 430
rect 48340 410 48440 430
rect 48680 410 48780 430
rect 49020 410 49120 430
rect 49360 410 49460 430
rect 49700 410 49800 430
rect 50040 410 50140 430
rect 50380 410 50480 430
rect 50720 410 50820 430
rect 51060 410 51160 430
rect 51400 410 51500 430
rect 51740 410 51840 430
rect 52080 410 52180 430
rect 52420 410 52520 430
rect 52760 410 52860 430
rect 53100 410 53200 430
rect 53440 410 53540 430
rect 53780 410 53880 430
rect 54120 410 54220 430
rect 54460 410 54560 430
rect 54800 410 54900 430
rect 55140 410 55240 430
rect 55480 410 55580 430
rect 55820 410 55920 430
rect 56160 410 56260 430
rect 56500 410 56600 430
rect 56840 410 56940 430
rect 57180 410 57280 430
rect 57520 410 57620 430
rect 57860 410 57960 430
rect 58200 410 58300 430
rect 58540 410 58640 430
rect 58880 410 58980 430
rect 59220 410 59320 430
rect 430 350 450 410
rect 510 350 790 410
rect 850 350 1130 410
rect 1190 350 1230 410
rect 1500 350 1520 410
rect 1580 350 1860 410
rect 1920 350 2200 410
rect 2260 350 2540 410
rect 2600 350 2880 410
rect 2940 350 3220 410
rect 3280 350 3560 410
rect 3620 350 3900 410
rect 3960 350 4240 410
rect 4300 350 4340 410
rect 4520 350 4540 410
rect 4600 350 4880 410
rect 4940 350 5220 410
rect 5280 350 5560 410
rect 5620 350 5900 410
rect 5960 350 6240 410
rect 6300 350 6580 410
rect 6640 350 6920 410
rect 6980 350 7260 410
rect 7320 350 7600 410
rect 7660 350 7940 410
rect 8000 350 8280 410
rect 8340 350 8620 410
rect 8680 350 8960 410
rect 9020 350 9300 410
rect 9360 350 9640 410
rect 9700 350 9980 410
rect 10040 350 10320 410
rect 10380 350 10660 410
rect 10720 350 11000 410
rect 11060 350 11340 410
rect 11400 350 11680 410
rect 11740 350 12020 410
rect 12080 350 12360 410
rect 12420 350 12700 410
rect 12760 350 13040 410
rect 13100 350 13380 410
rect 13440 350 13720 410
rect 13780 350 14060 410
rect 14120 350 14400 410
rect 14460 350 14740 410
rect 14800 350 15080 410
rect 15140 350 15420 410
rect 15480 350 15520 410
rect 15700 350 15720 410
rect 15780 350 16060 410
rect 16120 350 16400 410
rect 16460 350 16740 410
rect 16800 350 17080 410
rect 17140 350 17420 410
rect 17480 350 17760 410
rect 17820 350 18100 410
rect 18160 350 18440 410
rect 18500 350 18780 410
rect 18840 350 19120 410
rect 19180 350 19460 410
rect 19520 350 19800 410
rect 19860 350 20140 410
rect 20200 350 20480 410
rect 20540 350 20820 410
rect 20880 350 21160 410
rect 21220 350 21500 410
rect 21560 350 21840 410
rect 21900 350 22180 410
rect 22240 350 22520 410
rect 22580 350 22860 410
rect 22920 350 23200 410
rect 23260 350 23540 410
rect 23600 350 23880 410
rect 23940 350 24220 410
rect 24280 350 24560 410
rect 24620 350 24900 410
rect 24960 350 25240 410
rect 25300 350 25580 410
rect 25640 350 25920 410
rect 25980 350 26260 410
rect 26320 350 26600 410
rect 26660 350 26940 410
rect 27000 350 27280 410
rect 27340 350 27620 410
rect 27680 350 27960 410
rect 28020 350 28300 410
rect 28360 350 28640 410
rect 28700 350 28980 410
rect 29040 350 29320 410
rect 29380 350 29660 410
rect 29720 350 30000 410
rect 30060 350 30340 410
rect 30400 350 30680 410
rect 30740 350 31020 410
rect 31080 350 31360 410
rect 31420 350 31700 410
rect 31760 350 32040 410
rect 32100 350 32380 410
rect 32440 350 32720 410
rect 32780 350 33060 410
rect 33120 350 33400 410
rect 33460 350 33740 410
rect 33800 350 34080 410
rect 34140 350 34420 410
rect 34480 350 34760 410
rect 34820 350 35100 410
rect 35160 350 35440 410
rect 35500 350 35780 410
rect 35840 350 36120 410
rect 36180 350 36460 410
rect 36520 350 36800 410
rect 36860 350 37140 410
rect 37200 350 37480 410
rect 37540 350 37820 410
rect 37880 350 38160 410
rect 38220 350 38500 410
rect 38560 350 38840 410
rect 38900 350 39180 410
rect 39240 350 39520 410
rect 39580 350 39860 410
rect 39920 350 40200 410
rect 40260 350 40540 410
rect 40600 350 40880 410
rect 40940 350 41220 410
rect 41280 350 41560 410
rect 41620 350 41900 410
rect 41960 350 42240 410
rect 42300 350 42580 410
rect 42640 350 42920 410
rect 42980 350 43260 410
rect 43320 350 43600 410
rect 43660 350 43940 410
rect 44000 350 44280 410
rect 44340 350 44620 410
rect 44680 350 44960 410
rect 45020 350 45300 410
rect 45360 350 45640 410
rect 45700 350 45980 410
rect 46040 350 46320 410
rect 46380 350 46660 410
rect 46720 350 47000 410
rect 47060 350 47340 410
rect 47400 350 47680 410
rect 47740 350 48020 410
rect 48080 350 48360 410
rect 48420 350 48700 410
rect 48760 350 49040 410
rect 49100 350 49380 410
rect 49440 350 49720 410
rect 49780 350 50060 410
rect 50120 350 50400 410
rect 50460 350 50740 410
rect 50800 350 51080 410
rect 51140 350 51420 410
rect 51480 350 51760 410
rect 51820 350 52100 410
rect 52160 350 52440 410
rect 52500 350 52780 410
rect 52840 350 53120 410
rect 53180 350 53460 410
rect 53520 350 53800 410
rect 53860 350 54140 410
rect 54200 350 54480 410
rect 54540 350 54820 410
rect 54880 350 55160 410
rect 55220 350 55500 410
rect 55560 350 55840 410
rect 55900 350 56180 410
rect 56240 350 56520 410
rect 56580 350 56860 410
rect 56920 350 57200 410
rect 57260 350 57540 410
rect 57600 350 57880 410
rect 57940 350 58220 410
rect 58280 350 58560 410
rect 58620 350 58900 410
rect 58960 350 59240 410
rect 59300 350 59320 410
rect 430 330 530 350
rect 770 330 870 350
rect 1110 330 1210 350
rect 1500 330 1600 350
rect 1840 330 1940 350
rect 2180 330 2280 350
rect 2520 330 2620 350
rect 2860 330 2960 350
rect 3200 330 3300 350
rect 3540 330 3640 350
rect 3880 330 3980 350
rect 4220 330 4320 350
rect 4520 330 4620 350
rect 4860 330 4960 350
rect 5200 330 5300 350
rect 5540 330 5640 350
rect 5880 330 5980 350
rect 6220 330 6320 350
rect 6560 330 6660 350
rect 6900 330 7000 350
rect 7240 330 7340 350
rect 7580 330 7680 350
rect 7920 330 8020 350
rect 8260 330 8360 350
rect 8600 330 8700 350
rect 8940 330 9040 350
rect 9280 330 9380 350
rect 9620 330 9720 350
rect 9960 330 10060 350
rect 10300 330 10400 350
rect 10640 330 10740 350
rect 10980 330 11080 350
rect 11320 330 11420 350
rect 11660 330 11760 350
rect 12000 330 12100 350
rect 12340 330 12440 350
rect 12680 330 12780 350
rect 13020 330 13120 350
rect 13360 330 13460 350
rect 13700 330 13800 350
rect 14040 330 14140 350
rect 14380 330 14480 350
rect 14720 330 14820 350
rect 15060 330 15160 350
rect 15400 330 15500 350
rect 15700 330 15800 350
rect 16040 330 16140 350
rect 16380 330 16480 350
rect 16720 330 16820 350
rect 17060 330 17160 350
rect 17400 330 17500 350
rect 17740 330 17840 350
rect 18080 330 18180 350
rect 18420 330 18520 350
rect 18760 330 18860 350
rect 19100 330 19200 350
rect 19440 330 19540 350
rect 19780 330 19880 350
rect 20120 330 20220 350
rect 20460 330 20560 350
rect 20800 330 20900 350
rect 21140 330 21240 350
rect 21480 330 21580 350
rect 21820 330 21920 350
rect 22160 330 22260 350
rect 22500 330 22600 350
rect 22840 330 22940 350
rect 23180 330 23280 350
rect 23520 330 23620 350
rect 23860 330 23960 350
rect 24200 330 24300 350
rect 24540 330 24640 350
rect 24880 330 24980 350
rect 25220 330 25320 350
rect 25560 330 25660 350
rect 25900 330 26000 350
rect 26240 330 26340 350
rect 26580 330 26680 350
rect 26920 330 27020 350
rect 27260 330 27360 350
rect 27600 330 27700 350
rect 27940 330 28040 350
rect 28280 330 28380 350
rect 28620 330 28720 350
rect 28960 330 29060 350
rect 29300 330 29400 350
rect 29640 330 29740 350
rect 29980 330 30080 350
rect 30320 330 30420 350
rect 30660 330 30760 350
rect 31000 330 31100 350
rect 31340 330 31440 350
rect 31680 330 31780 350
rect 32020 330 32120 350
rect 32360 330 32460 350
rect 32700 330 32800 350
rect 33040 330 33140 350
rect 33380 330 33480 350
rect 33720 330 33820 350
rect 34060 330 34160 350
rect 34400 330 34500 350
rect 34740 330 34840 350
rect 35080 330 35180 350
rect 35420 330 35520 350
rect 35760 330 35860 350
rect 36100 330 36200 350
rect 36440 330 36540 350
rect 36780 330 36880 350
rect 37120 330 37220 350
rect 37460 330 37560 350
rect 37800 330 37900 350
rect 38140 330 38240 350
rect 38480 330 38580 350
rect 38820 330 38920 350
rect 39160 330 39260 350
rect 39500 330 39600 350
rect 39840 330 39940 350
rect 40180 330 40280 350
rect 40520 330 40620 350
rect 40860 330 40960 350
rect 41200 330 41300 350
rect 41540 330 41640 350
rect 41880 330 41980 350
rect 42220 330 42320 350
rect 42560 330 42660 350
rect 42900 330 43000 350
rect 43240 330 43340 350
rect 43580 330 43680 350
rect 43920 330 44020 350
rect 44260 330 44360 350
rect 44600 330 44700 350
rect 44940 330 45040 350
rect 45280 330 45380 350
rect 45620 330 45720 350
rect 45960 330 46060 350
rect 46300 330 46400 350
rect 46640 330 46740 350
rect 46980 330 47080 350
rect 47320 330 47420 350
rect 47660 330 47760 350
rect 48000 330 48100 350
rect 48340 330 48440 350
rect 48680 330 48780 350
rect 49020 330 49120 350
rect 49360 330 49460 350
rect 49700 330 49800 350
rect 50040 330 50140 350
rect 50380 330 50480 350
rect 50720 330 50820 350
rect 51060 330 51160 350
rect 51400 330 51500 350
rect 51740 330 51840 350
rect 52080 330 52180 350
rect 52420 330 52520 350
rect 52760 330 52860 350
rect 53100 330 53200 350
rect 53440 330 53540 350
rect 53780 330 53880 350
rect 54120 330 54220 350
rect 54460 330 54560 350
rect 54800 330 54900 350
rect 55140 330 55240 350
rect 55480 330 55580 350
rect 55820 330 55920 350
rect 56160 330 56260 350
rect 56500 330 56600 350
rect 56840 330 56940 350
rect 57180 330 57280 350
rect 57520 330 57620 350
rect 57860 330 57960 350
rect 58200 330 58300 350
rect 58540 330 58640 350
rect 58880 330 58980 350
rect 59220 330 59320 350
rect 610 200 690 210
rect 610 130 620 200
rect 680 130 690 200
rect -940 110 150 130
rect 610 120 690 130
rect 950 200 1030 210
rect 950 130 960 200
rect 1020 130 1030 200
rect 950 120 1030 130
rect 1680 200 1760 210
rect 1680 130 1690 200
rect 1750 130 1760 200
rect 1680 120 1760 130
rect 2020 200 2100 210
rect 2020 130 2030 200
rect 2090 130 2100 200
rect 2020 120 2100 130
rect 2360 200 2440 210
rect 2360 130 2370 200
rect 2430 130 2440 200
rect 2360 120 2440 130
rect 2700 200 2780 210
rect 2700 130 2710 200
rect 2770 130 2780 200
rect 2700 120 2780 130
rect 3040 200 3120 210
rect 3040 130 3050 200
rect 3110 130 3120 200
rect 3040 120 3120 130
rect 3380 200 3460 210
rect 3380 130 3390 200
rect 3450 130 3460 200
rect 3380 120 3460 130
rect 3720 200 3800 210
rect 3720 130 3730 200
rect 3790 130 3800 200
rect 3720 120 3800 130
rect 4060 200 4140 210
rect 4060 130 4070 200
rect 4130 130 4140 200
rect 4060 120 4140 130
rect 4700 200 4780 210
rect 4700 130 4710 200
rect 4770 130 4780 200
rect 4700 120 4780 130
rect 5040 200 5120 210
rect 5040 130 5050 200
rect 5110 130 5120 200
rect 5040 120 5120 130
rect 5380 200 5460 210
rect 5380 130 5390 200
rect 5450 130 5460 200
rect 5380 120 5460 130
rect 5720 200 5800 210
rect 5720 130 5730 200
rect 5790 130 5800 200
rect 5720 120 5800 130
rect 6060 200 6140 210
rect 6060 130 6070 200
rect 6130 130 6140 200
rect 6060 120 6140 130
rect 6400 200 6480 210
rect 6400 130 6410 200
rect 6470 130 6480 200
rect 6400 120 6480 130
rect 6740 200 6820 210
rect 6740 130 6750 200
rect 6810 130 6820 200
rect 6740 120 6820 130
rect 7080 200 7160 210
rect 7080 130 7090 200
rect 7150 130 7160 200
rect 7080 120 7160 130
rect 7420 200 7500 210
rect 7420 130 7430 200
rect 7490 130 7500 200
rect 7420 120 7500 130
rect 7760 200 7840 210
rect 7760 130 7770 200
rect 7830 130 7840 200
rect 7760 120 7840 130
rect 8100 200 8180 210
rect 8100 130 8110 200
rect 8170 130 8180 200
rect 8100 120 8180 130
rect 8440 200 8520 210
rect 8440 130 8450 200
rect 8510 130 8520 200
rect 8440 120 8520 130
rect 8780 200 8860 210
rect 8780 130 8790 200
rect 8850 130 8860 200
rect 8780 120 8860 130
rect 9120 200 9200 210
rect 9120 130 9130 200
rect 9190 130 9200 200
rect 9120 120 9200 130
rect 9460 200 9540 210
rect 9460 130 9470 200
rect 9530 130 9540 200
rect 9460 120 9540 130
rect 9800 200 9880 210
rect 9800 130 9810 200
rect 9870 130 9880 200
rect 9800 120 9880 130
rect 10140 200 10220 210
rect 10140 130 10150 200
rect 10210 130 10220 200
rect 10140 120 10220 130
rect 10480 200 10560 210
rect 10480 130 10490 200
rect 10550 130 10560 200
rect 10480 120 10560 130
rect 10820 200 10900 210
rect 10820 130 10830 200
rect 10890 130 10900 200
rect 10820 120 10900 130
rect 11160 200 11240 210
rect 11160 130 11170 200
rect 11230 130 11240 200
rect 11160 120 11240 130
rect 11500 200 11580 210
rect 11500 130 11510 200
rect 11570 130 11580 200
rect 11500 120 11580 130
rect 11840 200 11920 210
rect 11840 130 11850 200
rect 11910 130 11920 200
rect 11840 120 11920 130
rect 12180 200 12260 210
rect 12180 130 12190 200
rect 12250 130 12260 200
rect 12180 120 12260 130
rect 12520 200 12600 210
rect 12520 130 12530 200
rect 12590 130 12600 200
rect 12520 120 12600 130
rect 12860 200 12940 210
rect 12860 130 12870 200
rect 12930 130 12940 200
rect 12860 120 12940 130
rect 13200 200 13280 210
rect 13200 130 13210 200
rect 13270 130 13280 200
rect 13200 120 13280 130
rect 13540 200 13620 210
rect 13540 130 13550 200
rect 13610 130 13620 200
rect 13540 120 13620 130
rect 13880 200 13960 210
rect 13880 130 13890 200
rect 13950 130 13960 200
rect 13880 120 13960 130
rect 14220 200 14300 210
rect 14220 130 14230 200
rect 14290 130 14300 200
rect 14220 120 14300 130
rect 14560 200 14640 210
rect 14560 130 14570 200
rect 14630 130 14640 200
rect 14560 120 14640 130
rect 14900 200 14980 210
rect 14900 130 14910 200
rect 14970 130 14980 200
rect 14900 120 14980 130
rect 15240 200 15320 210
rect 15240 130 15250 200
rect 15310 130 15320 200
rect 15240 120 15320 130
rect 15880 200 15960 210
rect 15880 130 15890 200
rect 15950 130 15960 200
rect 15880 120 15960 130
rect 16220 200 16300 210
rect 16220 130 16230 200
rect 16290 130 16300 200
rect 16220 120 16300 130
rect 16560 200 16640 210
rect 16560 130 16570 200
rect 16630 130 16640 200
rect 16560 120 16640 130
rect 16900 200 16980 210
rect 16900 130 16910 200
rect 16970 130 16980 200
rect 16900 120 16980 130
rect 17240 200 17320 210
rect 17240 130 17250 200
rect 17310 130 17320 200
rect 17240 120 17320 130
rect 17580 200 17660 210
rect 17580 130 17590 200
rect 17650 130 17660 200
rect 17580 120 17660 130
rect 17920 200 18000 210
rect 17920 130 17930 200
rect 17990 130 18000 200
rect 17920 120 18000 130
rect 18260 200 18340 210
rect 18260 130 18270 200
rect 18330 130 18340 200
rect 18260 120 18340 130
rect 18600 200 18680 210
rect 18600 130 18610 200
rect 18670 130 18680 200
rect 18600 120 18680 130
rect 18940 200 19020 210
rect 18940 130 18950 200
rect 19010 130 19020 200
rect 18940 120 19020 130
rect 19280 200 19360 210
rect 19280 130 19290 200
rect 19350 130 19360 200
rect 19280 120 19360 130
rect 19620 200 19700 210
rect 19620 130 19630 200
rect 19690 130 19700 200
rect 19620 120 19700 130
rect 19960 200 20040 210
rect 19960 130 19970 200
rect 20030 130 20040 200
rect 19960 120 20040 130
rect 20300 200 20380 210
rect 20300 130 20310 200
rect 20370 130 20380 200
rect 20300 120 20380 130
rect 20640 200 20720 210
rect 20640 130 20650 200
rect 20710 130 20720 200
rect 20640 120 20720 130
rect 20980 200 21060 210
rect 20980 130 20990 200
rect 21050 130 21060 200
rect 20980 120 21060 130
rect 21320 200 21400 210
rect 21320 130 21330 200
rect 21390 130 21400 200
rect 21320 120 21400 130
rect 21660 200 21740 210
rect 21660 130 21670 200
rect 21730 130 21740 200
rect 21660 120 21740 130
rect 22000 200 22080 210
rect 22000 130 22010 200
rect 22070 130 22080 200
rect 22000 120 22080 130
rect 22340 200 22420 210
rect 22340 130 22350 200
rect 22410 130 22420 200
rect 22340 120 22420 130
rect 22680 200 22760 210
rect 22680 130 22690 200
rect 22750 130 22760 200
rect 22680 120 22760 130
rect 23020 200 23100 210
rect 23020 130 23030 200
rect 23090 130 23100 200
rect 23020 120 23100 130
rect 23360 200 23440 210
rect 23360 130 23370 200
rect 23430 130 23440 200
rect 23360 120 23440 130
rect 23700 200 23780 210
rect 23700 130 23710 200
rect 23770 130 23780 200
rect 23700 120 23780 130
rect 24040 200 24120 210
rect 24040 130 24050 200
rect 24110 130 24120 200
rect 24040 120 24120 130
rect 24380 200 24460 210
rect 24380 130 24390 200
rect 24450 130 24460 200
rect 24380 120 24460 130
rect 24720 200 24800 210
rect 24720 130 24730 200
rect 24790 130 24800 200
rect 24720 120 24800 130
rect 25060 200 25140 210
rect 25060 130 25070 200
rect 25130 130 25140 200
rect 25060 120 25140 130
rect 25400 200 25480 210
rect 25400 130 25410 200
rect 25470 130 25480 200
rect 25400 120 25480 130
rect 25740 200 25820 210
rect 25740 130 25750 200
rect 25810 130 25820 200
rect 25740 120 25820 130
rect 26080 200 26160 210
rect 26080 130 26090 200
rect 26150 130 26160 200
rect 26080 120 26160 130
rect 26420 200 26500 210
rect 26420 130 26430 200
rect 26490 130 26500 200
rect 26420 120 26500 130
rect 26760 200 26840 210
rect 26760 130 26770 200
rect 26830 130 26840 200
rect 26760 120 26840 130
rect 27100 200 27180 210
rect 27100 130 27110 200
rect 27170 130 27180 200
rect 27100 120 27180 130
rect 27440 200 27520 210
rect 27440 130 27450 200
rect 27510 130 27520 200
rect 27440 120 27520 130
rect 27780 200 27860 210
rect 27780 130 27790 200
rect 27850 130 27860 200
rect 27780 120 27860 130
rect 28120 200 28200 210
rect 28120 130 28130 200
rect 28190 130 28200 200
rect 28120 120 28200 130
rect 28460 200 28540 210
rect 28460 130 28470 200
rect 28530 130 28540 200
rect 28460 120 28540 130
rect 28800 200 28880 210
rect 28800 130 28810 200
rect 28870 130 28880 200
rect 28800 120 28880 130
rect 29140 200 29220 210
rect 29140 130 29150 200
rect 29210 130 29220 200
rect 29140 120 29220 130
rect 29480 200 29560 210
rect 29480 130 29490 200
rect 29550 130 29560 200
rect 29480 120 29560 130
rect 29820 200 29900 210
rect 29820 130 29830 200
rect 29890 130 29900 200
rect 29820 120 29900 130
rect 30160 200 30240 210
rect 30160 130 30170 200
rect 30230 130 30240 200
rect 30160 120 30240 130
rect 30500 200 30580 210
rect 30500 130 30510 200
rect 30570 130 30580 200
rect 30500 120 30580 130
rect 30840 200 30920 210
rect 30840 130 30850 200
rect 30910 130 30920 200
rect 30840 120 30920 130
rect 31180 200 31260 210
rect 31180 130 31190 200
rect 31250 130 31260 200
rect 31180 120 31260 130
rect 31520 200 31600 210
rect 31520 130 31530 200
rect 31590 130 31600 200
rect 31520 120 31600 130
rect 31860 200 31940 210
rect 31860 130 31870 200
rect 31930 130 31940 200
rect 31860 120 31940 130
rect 32200 200 32280 210
rect 32200 130 32210 200
rect 32270 130 32280 200
rect 32200 120 32280 130
rect 32540 200 32620 210
rect 32540 130 32550 200
rect 32610 130 32620 200
rect 32540 120 32620 130
rect 32880 200 32960 210
rect 32880 130 32890 200
rect 32950 130 32960 200
rect 32880 120 32960 130
rect 33220 200 33300 210
rect 33220 130 33230 200
rect 33290 130 33300 200
rect 33220 120 33300 130
rect 33560 200 33640 210
rect 33560 130 33570 200
rect 33630 130 33640 200
rect 33560 120 33640 130
rect 33900 200 33980 210
rect 33900 130 33910 200
rect 33970 130 33980 200
rect 33900 120 33980 130
rect 34240 200 34320 210
rect 34240 130 34250 200
rect 34310 130 34320 200
rect 34240 120 34320 130
rect 34580 200 34660 210
rect 34580 130 34590 200
rect 34650 130 34660 200
rect 34580 120 34660 130
rect 34920 200 35000 210
rect 34920 130 34930 200
rect 34990 130 35000 200
rect 34920 120 35000 130
rect 35260 200 35340 210
rect 35260 130 35270 200
rect 35330 130 35340 200
rect 35260 120 35340 130
rect 35600 200 35680 210
rect 35600 130 35610 200
rect 35670 130 35680 200
rect 35600 120 35680 130
rect 35940 200 36020 210
rect 35940 130 35950 200
rect 36010 130 36020 200
rect 35940 120 36020 130
rect 36280 200 36360 210
rect 36280 130 36290 200
rect 36350 130 36360 200
rect 36280 120 36360 130
rect 36620 200 36700 210
rect 36620 130 36630 200
rect 36690 130 36700 200
rect 36620 120 36700 130
rect 36960 200 37040 210
rect 36960 130 36970 200
rect 37030 130 37040 200
rect 36960 120 37040 130
rect 37300 200 37380 210
rect 37300 130 37310 200
rect 37370 130 37380 200
rect 37300 120 37380 130
rect 37640 200 37720 210
rect 37640 130 37650 200
rect 37710 130 37720 200
rect 37640 120 37720 130
rect 37980 200 38060 210
rect 37980 130 37990 200
rect 38050 130 38060 200
rect 37980 120 38060 130
rect 38320 200 38400 210
rect 38320 130 38330 200
rect 38390 130 38400 200
rect 38320 120 38400 130
rect 38660 200 38740 210
rect 38660 130 38670 200
rect 38730 130 38740 200
rect 38660 120 38740 130
rect 39000 200 39080 210
rect 39000 130 39010 200
rect 39070 130 39080 200
rect 39000 120 39080 130
rect 39340 200 39420 210
rect 39340 130 39350 200
rect 39410 130 39420 200
rect 39340 120 39420 130
rect 39680 200 39760 210
rect 39680 130 39690 200
rect 39750 130 39760 200
rect 39680 120 39760 130
rect 40020 200 40100 210
rect 40020 130 40030 200
rect 40090 130 40100 200
rect 40020 120 40100 130
rect 40360 200 40440 210
rect 40360 130 40370 200
rect 40430 130 40440 200
rect 40360 120 40440 130
rect 40700 200 40780 210
rect 40700 130 40710 200
rect 40770 130 40780 200
rect 40700 120 40780 130
rect 41040 200 41120 210
rect 41040 130 41050 200
rect 41110 130 41120 200
rect 41040 120 41120 130
rect 41380 200 41460 210
rect 41380 130 41390 200
rect 41450 130 41460 200
rect 41380 120 41460 130
rect 41720 200 41800 210
rect 41720 130 41730 200
rect 41790 130 41800 200
rect 41720 120 41800 130
rect 42060 200 42140 210
rect 42060 130 42070 200
rect 42130 130 42140 200
rect 42060 120 42140 130
rect 42400 200 42480 210
rect 42400 130 42410 200
rect 42470 130 42480 200
rect 42400 120 42480 130
rect 42740 200 42820 210
rect 42740 130 42750 200
rect 42810 130 42820 200
rect 42740 120 42820 130
rect 43080 200 43160 210
rect 43080 130 43090 200
rect 43150 130 43160 200
rect 43080 120 43160 130
rect 43420 200 43500 210
rect 43420 130 43430 200
rect 43490 130 43500 200
rect 43420 120 43500 130
rect 43760 200 43840 210
rect 43760 130 43770 200
rect 43830 130 43840 200
rect 43760 120 43840 130
rect 44100 200 44180 210
rect 44100 130 44110 200
rect 44170 130 44180 200
rect 44100 120 44180 130
rect 44440 200 44520 210
rect 44440 130 44450 200
rect 44510 130 44520 200
rect 44440 120 44520 130
rect 44780 200 44860 210
rect 44780 130 44790 200
rect 44850 130 44860 200
rect 44780 120 44860 130
rect 45120 200 45200 210
rect 45120 130 45130 200
rect 45190 130 45200 200
rect 45120 120 45200 130
rect 45460 200 45540 210
rect 45460 130 45470 200
rect 45530 130 45540 200
rect 45460 120 45540 130
rect 45800 200 45880 210
rect 45800 130 45810 200
rect 45870 130 45880 200
rect 45800 120 45880 130
rect 46140 200 46220 210
rect 46140 130 46150 200
rect 46210 130 46220 200
rect 46140 120 46220 130
rect 46480 200 46560 210
rect 46480 130 46490 200
rect 46550 130 46560 200
rect 46480 120 46560 130
rect 46820 200 46900 210
rect 46820 130 46830 200
rect 46890 130 46900 200
rect 46820 120 46900 130
rect 47160 200 47240 210
rect 47160 130 47170 200
rect 47230 130 47240 200
rect 47160 120 47240 130
rect 47500 200 47580 210
rect 47500 130 47510 200
rect 47570 130 47580 200
rect 47500 120 47580 130
rect 47840 200 47920 210
rect 47840 130 47850 200
rect 47910 130 47920 200
rect 47840 120 47920 130
rect 48180 200 48260 210
rect 48180 130 48190 200
rect 48250 130 48260 200
rect 48180 120 48260 130
rect 48520 200 48600 210
rect 48520 130 48530 200
rect 48590 130 48600 200
rect 48520 120 48600 130
rect 48860 200 48940 210
rect 48860 130 48870 200
rect 48930 130 48940 200
rect 48860 120 48940 130
rect 49200 200 49280 210
rect 49200 130 49210 200
rect 49270 130 49280 200
rect 49200 120 49280 130
rect 49540 200 49620 210
rect 49540 130 49550 200
rect 49610 130 49620 200
rect 49540 120 49620 130
rect 49880 200 49960 210
rect 49880 130 49890 200
rect 49950 130 49960 200
rect 49880 120 49960 130
rect 50220 200 50300 210
rect 50220 130 50230 200
rect 50290 130 50300 200
rect 50220 120 50300 130
rect 50560 200 50640 210
rect 50560 130 50570 200
rect 50630 130 50640 200
rect 50560 120 50640 130
rect 50900 200 50980 210
rect 50900 130 50910 200
rect 50970 130 50980 200
rect 50900 120 50980 130
rect 51240 200 51320 210
rect 51240 130 51250 200
rect 51310 130 51320 200
rect 51240 120 51320 130
rect 51580 200 51660 210
rect 51580 130 51590 200
rect 51650 130 51660 200
rect 51580 120 51660 130
rect 51920 200 52000 210
rect 51920 130 51930 200
rect 51990 130 52000 200
rect 51920 120 52000 130
rect 52260 200 52340 210
rect 52260 130 52270 200
rect 52330 130 52340 200
rect 52260 120 52340 130
rect 52600 200 52680 210
rect 52600 130 52610 200
rect 52670 130 52680 200
rect 52600 120 52680 130
rect 52940 200 53020 210
rect 52940 130 52950 200
rect 53010 130 53020 200
rect 52940 120 53020 130
rect 53280 200 53360 210
rect 53280 130 53290 200
rect 53350 130 53360 200
rect 53280 120 53360 130
rect 53620 200 53700 210
rect 53620 130 53630 200
rect 53690 130 53700 200
rect 53620 120 53700 130
rect 53960 200 54040 210
rect 53960 130 53970 200
rect 54030 130 54040 200
rect 53960 120 54040 130
rect 54300 200 54380 210
rect 54300 130 54310 200
rect 54370 130 54380 200
rect 54300 120 54380 130
rect 54640 200 54720 210
rect 54640 130 54650 200
rect 54710 130 54720 200
rect 54640 120 54720 130
rect 54980 200 55060 210
rect 54980 130 54990 200
rect 55050 130 55060 200
rect 54980 120 55060 130
rect 55320 200 55400 210
rect 55320 130 55330 200
rect 55390 130 55400 200
rect 55320 120 55400 130
rect 55660 200 55740 210
rect 55660 130 55670 200
rect 55730 130 55740 200
rect 55660 120 55740 130
rect 56000 200 56080 210
rect 56000 130 56010 200
rect 56070 130 56080 200
rect 56000 120 56080 130
rect 56340 200 56420 210
rect 56340 130 56350 200
rect 56410 130 56420 200
rect 56340 120 56420 130
rect 56680 200 56760 210
rect 56680 130 56690 200
rect 56750 130 56760 200
rect 56680 120 56760 130
rect 57020 200 57100 210
rect 57020 130 57030 200
rect 57090 130 57100 200
rect 57020 120 57100 130
rect 57360 200 57440 210
rect 57360 130 57370 200
rect 57430 130 57440 200
rect 57360 120 57440 130
rect 57700 200 57780 210
rect 57700 130 57710 200
rect 57770 130 57780 200
rect 57700 120 57780 130
rect 58040 200 58120 210
rect 58040 130 58050 200
rect 58110 130 58120 200
rect 58040 120 58120 130
rect 58380 200 58460 210
rect 58380 130 58390 200
rect 58450 130 58460 200
rect 58380 120 58460 130
rect 58720 200 58800 210
rect 58720 130 58730 200
rect 58790 130 58800 200
rect 58720 120 58800 130
rect 59060 200 59140 210
rect 59060 130 59070 200
rect 59130 130 59140 200
rect 59060 120 59140 130
rect -940 30 70 110
rect 130 30 150 110
rect -940 10 150 30
rect 430 80 530 100
rect 770 80 870 100
rect 1110 80 1210 100
rect 430 20 450 80
rect 510 20 790 80
rect 850 20 1130 80
rect 1190 20 1210 80
rect 430 0 530 20
rect 770 0 870 20
rect 1110 0 1210 20
rect 1500 80 1600 100
rect 1840 80 1940 100
rect 2180 80 2280 100
rect 2520 80 2620 100
rect 2860 80 2960 100
rect 3200 80 3300 100
rect 3540 80 3640 100
rect 3880 80 3980 100
rect 4220 80 4320 100
rect 1500 20 1520 80
rect 1580 20 1860 80
rect 1920 20 2200 80
rect 2260 20 2540 80
rect 2600 20 2880 80
rect 2940 20 3220 80
rect 3280 20 3560 80
rect 3620 20 3900 80
rect 3960 20 4240 80
rect 4300 20 4320 80
rect 1500 0 1600 20
rect 1840 0 1940 20
rect 2180 0 2280 20
rect 2520 0 2620 20
rect 2860 0 2960 20
rect 3200 0 3300 20
rect 3540 0 3640 20
rect 3880 0 3980 20
rect 4220 0 4320 20
rect 4520 80 4620 100
rect 4860 80 4960 100
rect 5200 80 5300 100
rect 5540 80 5640 100
rect 5880 80 5980 100
rect 6220 80 6320 100
rect 6560 80 6660 100
rect 6900 80 7000 100
rect 7240 80 7340 100
rect 7580 80 7680 100
rect 7920 80 8020 100
rect 8260 80 8360 100
rect 8600 80 8700 100
rect 8940 80 9040 100
rect 9280 80 9380 100
rect 9620 80 9720 100
rect 9960 80 10060 100
rect 10300 80 10400 100
rect 10640 80 10740 100
rect 10980 80 11080 100
rect 11320 80 11420 100
rect 11660 80 11760 100
rect 12000 80 12100 100
rect 12340 80 12440 100
rect 12680 80 12780 100
rect 13020 80 13120 100
rect 13360 80 13460 100
rect 13700 80 13800 100
rect 14040 80 14140 100
rect 14380 80 14480 100
rect 14720 80 14820 100
rect 15060 80 15160 100
rect 15400 80 15500 100
rect 4520 20 4540 80
rect 4600 20 4880 80
rect 4940 20 5220 80
rect 5280 20 5560 80
rect 5620 20 5900 80
rect 5960 20 6240 80
rect 6300 20 6580 80
rect 6640 20 6920 80
rect 6980 20 7260 80
rect 7320 20 7600 80
rect 7660 20 7940 80
rect 8000 20 8280 80
rect 8340 20 8620 80
rect 8680 20 8960 80
rect 9020 20 9300 80
rect 9360 20 9640 80
rect 9700 20 9980 80
rect 10040 20 10320 80
rect 10380 20 10660 80
rect 10720 20 11000 80
rect 11060 20 11340 80
rect 11400 20 11680 80
rect 11740 20 12020 80
rect 12080 20 12360 80
rect 12420 20 12700 80
rect 12760 20 13040 80
rect 13100 20 13380 80
rect 13440 20 13720 80
rect 13780 20 14060 80
rect 14120 20 14400 80
rect 14460 20 14740 80
rect 14800 20 15080 80
rect 15140 20 15420 80
rect 15480 20 15500 80
rect 4520 0 4620 20
rect 4860 0 4960 20
rect 5200 0 5300 20
rect 5540 0 5640 20
rect 5880 0 5980 20
rect 6220 0 6320 20
rect 6560 0 6660 20
rect 6900 0 7000 20
rect 7240 0 7340 20
rect 7580 0 7680 20
rect 7920 0 8020 20
rect 8260 0 8360 20
rect 8600 0 8700 20
rect 8940 0 9040 20
rect 9280 0 9380 20
rect 9620 0 9720 20
rect 9960 0 10060 20
rect 10300 0 10400 20
rect 10640 0 10740 20
rect 10980 0 11080 20
rect 11320 0 11420 20
rect 11660 0 11760 20
rect 12000 0 12100 20
rect 12340 0 12440 20
rect 12680 0 12780 20
rect 13020 0 13120 20
rect 13360 0 13460 20
rect 13700 0 13800 20
rect 14040 0 14140 20
rect 14380 0 14480 20
rect 14720 0 14820 20
rect 15060 0 15160 20
rect 15400 0 15500 20
rect 15700 80 15800 100
rect 16040 80 16140 100
rect 16380 80 16480 100
rect 16720 80 16820 100
rect 17060 80 17160 100
rect 17400 80 17500 100
rect 17740 80 17840 100
rect 18080 80 18180 100
rect 18420 80 18520 100
rect 18760 80 18860 100
rect 19100 80 19200 100
rect 19440 80 19540 100
rect 19780 80 19880 100
rect 20120 80 20220 100
rect 20460 80 20560 100
rect 20800 80 20900 100
rect 21140 80 21240 100
rect 21480 80 21580 100
rect 21820 80 21920 100
rect 22160 80 22260 100
rect 22500 80 22600 100
rect 22840 80 22940 100
rect 23180 80 23280 100
rect 23520 80 23620 100
rect 23860 80 23960 100
rect 24200 80 24300 100
rect 24540 80 24640 100
rect 24880 80 24980 100
rect 25220 80 25320 100
rect 25560 80 25660 100
rect 25900 80 26000 100
rect 26240 80 26340 100
rect 26580 80 26680 100
rect 26920 80 27020 100
rect 27260 80 27360 100
rect 27600 80 27700 100
rect 27940 80 28040 100
rect 28280 80 28380 100
rect 28620 80 28720 100
rect 28960 80 29060 100
rect 29300 80 29400 100
rect 29640 80 29740 100
rect 29980 80 30080 100
rect 30320 80 30420 100
rect 30660 80 30760 100
rect 31000 80 31100 100
rect 31340 80 31440 100
rect 31680 80 31780 100
rect 32020 80 32120 100
rect 32360 80 32460 100
rect 32700 80 32800 100
rect 33040 80 33140 100
rect 33380 80 33480 100
rect 33720 80 33820 100
rect 34060 80 34160 100
rect 34400 80 34500 100
rect 34740 80 34840 100
rect 35080 80 35180 100
rect 35420 80 35520 100
rect 35760 80 35860 100
rect 36100 80 36200 100
rect 36440 80 36540 100
rect 36780 80 36880 100
rect 37120 80 37220 100
rect 37460 80 37560 100
rect 37800 80 37900 100
rect 38140 80 38240 100
rect 38480 80 38580 100
rect 38820 80 38920 100
rect 39160 80 39260 100
rect 39500 80 39600 100
rect 39840 80 39940 100
rect 40180 80 40280 100
rect 40520 80 40620 100
rect 40860 80 40960 100
rect 41200 80 41300 100
rect 41540 80 41640 100
rect 41880 80 41980 100
rect 42220 80 42320 100
rect 42560 80 42660 100
rect 42900 80 43000 100
rect 43240 80 43340 100
rect 43580 80 43680 100
rect 43920 80 44020 100
rect 44260 80 44360 100
rect 44600 80 44700 100
rect 44940 80 45040 100
rect 45280 80 45380 100
rect 45620 80 45720 100
rect 45960 80 46060 100
rect 46300 80 46400 100
rect 46640 80 46740 100
rect 46980 80 47080 100
rect 47320 80 47420 100
rect 47660 80 47760 100
rect 48000 80 48100 100
rect 48340 80 48440 100
rect 48680 80 48780 100
rect 49020 80 49120 100
rect 49360 80 49460 100
rect 49700 80 49800 100
rect 50040 80 50140 100
rect 50380 80 50480 100
rect 50720 80 50820 100
rect 51060 80 51160 100
rect 51400 80 51500 100
rect 51740 80 51840 100
rect 52080 80 52180 100
rect 52420 80 52520 100
rect 52760 80 52860 100
rect 53100 80 53200 100
rect 53440 80 53540 100
rect 53780 80 53880 100
rect 54120 80 54220 100
rect 54460 80 54560 100
rect 54800 80 54900 100
rect 55140 80 55240 100
rect 55480 80 55580 100
rect 55820 80 55920 100
rect 56160 80 56260 100
rect 56500 80 56600 100
rect 56840 80 56940 100
rect 57180 80 57280 100
rect 57520 80 57620 100
rect 57860 80 57960 100
rect 58200 80 58300 100
rect 58540 80 58640 100
rect 58880 80 58980 100
rect 59220 80 59320 100
rect 15700 20 15720 80
rect 15780 20 16060 80
rect 16120 20 16400 80
rect 16460 20 16740 80
rect 16800 20 17080 80
rect 17140 20 17420 80
rect 17480 20 17760 80
rect 17820 20 18100 80
rect 18160 20 18440 80
rect 18500 20 18780 80
rect 18840 20 19120 80
rect 19180 20 19460 80
rect 19520 20 19800 80
rect 19860 20 20140 80
rect 20200 20 20480 80
rect 20540 20 20820 80
rect 20880 20 21160 80
rect 21220 20 21500 80
rect 21560 20 21840 80
rect 21900 20 22180 80
rect 22240 20 22520 80
rect 22580 20 22860 80
rect 22920 20 23200 80
rect 23260 20 23540 80
rect 23600 20 23880 80
rect 23940 20 24220 80
rect 24280 20 24560 80
rect 24620 20 24900 80
rect 24960 20 25240 80
rect 25300 20 25580 80
rect 25640 20 25920 80
rect 25980 20 26260 80
rect 26320 20 26600 80
rect 26660 20 26940 80
rect 27000 20 27280 80
rect 27340 20 27620 80
rect 27680 20 27960 80
rect 28020 20 28300 80
rect 28360 20 28640 80
rect 28700 20 28980 80
rect 29040 20 29320 80
rect 29380 20 29660 80
rect 29720 20 30000 80
rect 30060 20 30340 80
rect 30400 20 30680 80
rect 30740 20 31020 80
rect 31080 20 31360 80
rect 31420 20 31700 80
rect 31760 20 32040 80
rect 32100 20 32380 80
rect 32440 20 32720 80
rect 32780 20 33060 80
rect 33120 20 33400 80
rect 33460 20 33740 80
rect 33800 20 34080 80
rect 34140 20 34420 80
rect 34480 20 34760 80
rect 34820 20 35100 80
rect 35160 20 35440 80
rect 35500 20 35780 80
rect 35840 20 36120 80
rect 36180 20 36460 80
rect 36520 20 36800 80
rect 36860 20 37140 80
rect 37200 20 37480 80
rect 37540 20 37820 80
rect 37880 20 38160 80
rect 38220 20 38500 80
rect 38560 20 38840 80
rect 38900 20 39180 80
rect 39240 20 39520 80
rect 39580 20 39860 80
rect 39920 20 40200 80
rect 40260 20 40540 80
rect 40600 20 40880 80
rect 40940 20 41220 80
rect 41280 20 41560 80
rect 41620 20 41900 80
rect 41960 20 42240 80
rect 42300 20 42580 80
rect 42640 20 42920 80
rect 42980 20 43260 80
rect 43320 20 43600 80
rect 43660 20 43940 80
rect 44000 20 44280 80
rect 44340 20 44620 80
rect 44680 20 44960 80
rect 45020 20 45300 80
rect 45360 20 45640 80
rect 45700 20 45980 80
rect 46040 20 46320 80
rect 46380 20 46660 80
rect 46720 20 47000 80
rect 47060 20 47340 80
rect 47400 20 47680 80
rect 47740 20 48020 80
rect 48080 20 48360 80
rect 48420 20 48700 80
rect 48760 20 49040 80
rect 49100 20 49380 80
rect 49440 20 49720 80
rect 49780 20 50060 80
rect 50120 20 50400 80
rect 50460 20 50740 80
rect 50800 20 51080 80
rect 51140 20 51420 80
rect 51480 20 51760 80
rect 51820 20 52100 80
rect 52160 20 52440 80
rect 52500 20 52780 80
rect 52840 20 53120 80
rect 53180 20 53460 80
rect 53520 20 53800 80
rect 53860 20 54140 80
rect 54200 20 54480 80
rect 54540 20 54820 80
rect 54880 20 55160 80
rect 55220 20 55500 80
rect 55560 20 55840 80
rect 55900 20 56180 80
rect 56240 20 56520 80
rect 56580 20 56860 80
rect 56920 20 57200 80
rect 57260 20 57540 80
rect 57600 20 57880 80
rect 57940 20 58220 80
rect 58280 20 58560 80
rect 58620 20 58900 80
rect 58960 20 59240 80
rect 59300 20 59320 80
rect 15700 0 15800 20
rect 16040 0 16140 20
rect 16380 0 16480 20
rect 16720 0 16820 20
rect 17060 0 17160 20
rect 17400 0 17500 20
rect 17740 0 17840 20
rect 18080 0 18180 20
rect 18420 0 18520 20
rect 18760 0 18860 20
rect 19100 0 19200 20
rect 19440 0 19540 20
rect 19780 0 19880 20
rect 20120 0 20220 20
rect 20460 0 20560 20
rect 20800 0 20900 20
rect 21140 0 21240 20
rect 21480 0 21580 20
rect 21820 0 21920 20
rect 22160 0 22260 20
rect 22500 0 22600 20
rect 22840 0 22940 20
rect 23180 0 23280 20
rect 23520 0 23620 20
rect 23860 0 23960 20
rect 24200 0 24300 20
rect 24540 0 24640 20
rect 24880 0 24980 20
rect 25220 0 25320 20
rect 25560 0 25660 20
rect 25900 0 26000 20
rect 26240 0 26340 20
rect 26580 0 26680 20
rect 26920 0 27020 20
rect 27260 0 27360 20
rect 27600 0 27700 20
rect 27940 0 28040 20
rect 28280 0 28380 20
rect 28620 0 28720 20
rect 28960 0 29060 20
rect 29300 0 29400 20
rect 29640 0 29740 20
rect 29980 0 30080 20
rect 30320 0 30420 20
rect 30660 0 30760 20
rect 31000 0 31100 20
rect 31340 0 31440 20
rect 31680 0 31780 20
rect 32020 0 32120 20
rect 32360 0 32460 20
rect 32700 0 32800 20
rect 33040 0 33140 20
rect 33380 0 33480 20
rect 33720 0 33820 20
rect 34060 0 34160 20
rect 34400 0 34500 20
rect 34740 0 34840 20
rect 35080 0 35180 20
rect 35420 0 35520 20
rect 35760 0 35860 20
rect 36100 0 36200 20
rect 36440 0 36540 20
rect 36780 0 36880 20
rect 37120 0 37220 20
rect 37460 0 37560 20
rect 37800 0 37900 20
rect 38140 0 38240 20
rect 38480 0 38580 20
rect 38820 0 38920 20
rect 39160 0 39260 20
rect 39500 0 39600 20
rect 39840 0 39940 20
rect 40180 0 40280 20
rect 40520 0 40620 20
rect 40860 0 40960 20
rect 41200 0 41300 20
rect 41540 0 41640 20
rect 41880 0 41980 20
rect 42220 0 42320 20
rect 42560 0 42660 20
rect 42900 0 43000 20
rect 43240 0 43340 20
rect 43580 0 43680 20
rect 43920 0 44020 20
rect 44260 0 44360 20
rect 44600 0 44700 20
rect 44940 0 45040 20
rect 45280 0 45380 20
rect 45620 0 45720 20
rect 45960 0 46060 20
rect 46300 0 46400 20
rect 46640 0 46740 20
rect 46980 0 47080 20
rect 47320 0 47420 20
rect 47660 0 47760 20
rect 48000 0 48100 20
rect 48340 0 48440 20
rect 48680 0 48780 20
rect 49020 0 49120 20
rect 49360 0 49460 20
rect 49700 0 49800 20
rect 50040 0 50140 20
rect 50380 0 50480 20
rect 50720 0 50820 20
rect 51060 0 51160 20
rect 51400 0 51500 20
rect 51740 0 51840 20
rect 52080 0 52180 20
rect 52420 0 52520 20
rect 52760 0 52860 20
rect 53100 0 53200 20
rect 53440 0 53540 20
rect 53780 0 53880 20
rect 54120 0 54220 20
rect 54460 0 54560 20
rect 54800 0 54900 20
rect 55140 0 55240 20
rect 55480 0 55580 20
rect 55820 0 55920 20
rect 56160 0 56260 20
rect 56500 0 56600 20
rect 56840 0 56940 20
rect 57180 0 57280 20
rect 57520 0 57620 20
rect 57860 0 57960 20
rect 58200 0 58300 20
rect 58540 0 58640 20
rect 58880 0 58980 20
rect 59220 0 59320 20
rect 10 -60 110 -40
rect 10 -120 30 -60
rect 90 -120 110 -60
rect 10 -140 110 -120
rect 180 -60 1130 -40
rect 180 -120 200 -60
rect 260 -120 530 -60
rect 600 -120 700 -60
rect 770 -120 870 -60
rect 940 -120 1040 -60
rect 1110 -120 1130 -60
rect 180 -140 1130 -120
rect 1290 -50 4240 -40
rect 1290 -130 1300 -50
rect 1400 -60 4240 -50
rect 1400 -120 1600 -60
rect 1670 -120 1770 -60
rect 1840 -120 1940 -60
rect 2010 -120 2110 -60
rect 2180 -120 2280 -60
rect 2350 -120 2450 -60
rect 2520 -120 2620 -60
rect 2690 -120 2790 -60
rect 2860 -120 2960 -60
rect 3030 -120 3130 -60
rect 3200 -120 3300 -60
rect 3370 -120 3470 -60
rect 3540 -120 3640 -60
rect 3710 -120 3810 -60
rect 3880 -120 3980 -60
rect 4050 -120 4150 -60
rect 4220 -120 4240 -60
rect 1400 -130 4240 -120
rect 1290 -140 4240 -130
rect 4370 -50 15420 -40
rect 4370 -130 4380 -50
rect 4480 -60 15420 -50
rect 4480 -120 4620 -60
rect 4690 -120 4790 -60
rect 4860 -120 4960 -60
rect 5030 -120 5130 -60
rect 5200 -120 5300 -60
rect 5370 -120 5470 -60
rect 5540 -120 5640 -60
rect 5710 -120 5810 -60
rect 5880 -120 5980 -60
rect 6050 -120 6150 -60
rect 6220 -120 6320 -60
rect 6390 -120 6490 -60
rect 6560 -120 6660 -60
rect 6730 -120 6830 -60
rect 6900 -120 7000 -60
rect 7070 -120 7170 -60
rect 7240 -120 7340 -60
rect 7410 -120 7510 -60
rect 7580 -120 7680 -60
rect 7750 -120 7850 -60
rect 7920 -120 8020 -60
rect 8090 -120 8190 -60
rect 8260 -120 8360 -60
rect 8430 -120 8530 -60
rect 8600 -120 8700 -60
rect 8770 -120 8870 -60
rect 8940 -120 9040 -60
rect 9110 -120 9210 -60
rect 9280 -120 9380 -60
rect 9450 -120 9550 -60
rect 9620 -120 9720 -60
rect 9790 -120 9890 -60
rect 9960 -120 10060 -60
rect 10130 -120 10230 -60
rect 10300 -120 10400 -60
rect 10470 -120 10570 -60
rect 10640 -120 10740 -60
rect 10810 -120 10910 -60
rect 10980 -120 11080 -60
rect 11150 -120 11250 -60
rect 11320 -120 11420 -60
rect 11490 -120 11590 -60
rect 11660 -120 11760 -60
rect 11830 -120 11930 -60
rect 12000 -120 12100 -60
rect 12170 -120 12270 -60
rect 12340 -120 12440 -60
rect 12510 -120 12610 -60
rect 12680 -120 12780 -60
rect 12850 -120 12950 -60
rect 13020 -120 13120 -60
rect 13190 -120 13290 -60
rect 13360 -120 13460 -60
rect 13530 -120 13630 -60
rect 13700 -120 13800 -60
rect 13870 -120 13970 -60
rect 14040 -120 14140 -60
rect 14210 -120 14310 -60
rect 14380 -120 14480 -60
rect 14550 -120 14650 -60
rect 14720 -120 14820 -60
rect 14890 -120 14990 -60
rect 15060 -120 15160 -60
rect 15230 -120 15330 -60
rect 15400 -120 15420 -60
rect 4480 -130 15420 -120
rect 4370 -140 15420 -130
rect 15550 -50 59240 -40
rect 15550 -130 15560 -50
rect 15660 -60 59240 -50
rect 15660 -120 15800 -60
rect 15870 -120 15970 -60
rect 16040 -120 16140 -60
rect 16210 -120 16310 -60
rect 16380 -120 16480 -60
rect 16550 -120 16650 -60
rect 16720 -120 16820 -60
rect 16890 -120 16990 -60
rect 17060 -120 17160 -60
rect 17230 -120 17330 -60
rect 17400 -120 17500 -60
rect 17570 -120 17670 -60
rect 17740 -120 17840 -60
rect 17910 -120 18010 -60
rect 18080 -120 18180 -60
rect 18250 -120 18350 -60
rect 18420 -120 18520 -60
rect 18590 -120 18690 -60
rect 18760 -120 18860 -60
rect 18930 -120 19030 -60
rect 19100 -120 19200 -60
rect 19270 -120 19370 -60
rect 19440 -120 19540 -60
rect 19610 -120 19710 -60
rect 19780 -120 19880 -60
rect 19950 -120 20050 -60
rect 20120 -120 20220 -60
rect 20290 -120 20390 -60
rect 20460 -120 20560 -60
rect 20630 -120 20730 -60
rect 20800 -120 20900 -60
rect 20970 -120 21070 -60
rect 21140 -120 21240 -60
rect 21310 -120 21410 -60
rect 21480 -120 21580 -60
rect 21650 -120 21750 -60
rect 21820 -120 21920 -60
rect 21990 -120 22090 -60
rect 22160 -120 22260 -60
rect 22330 -120 22430 -60
rect 22500 -120 22600 -60
rect 22670 -120 22770 -60
rect 22840 -120 22940 -60
rect 23010 -120 23110 -60
rect 23180 -120 23280 -60
rect 23350 -120 23450 -60
rect 23520 -120 23620 -60
rect 23690 -120 23790 -60
rect 23860 -120 23960 -60
rect 24030 -120 24130 -60
rect 24200 -120 24300 -60
rect 24370 -120 24470 -60
rect 24540 -120 24640 -60
rect 24710 -120 24810 -60
rect 24880 -120 24980 -60
rect 25050 -120 25150 -60
rect 25220 -120 25320 -60
rect 25390 -120 25490 -60
rect 25560 -120 25660 -60
rect 25730 -120 25830 -60
rect 25900 -120 26000 -60
rect 26070 -120 26170 -60
rect 26240 -120 26340 -60
rect 26410 -120 26510 -60
rect 26580 -120 26680 -60
rect 26750 -120 26850 -60
rect 26920 -120 27020 -60
rect 27090 -120 27190 -60
rect 27260 -120 27360 -60
rect 27430 -120 27530 -60
rect 27600 -120 27700 -60
rect 27770 -120 27870 -60
rect 27940 -120 28040 -60
rect 28110 -120 28210 -60
rect 28280 -120 28380 -60
rect 28450 -120 28550 -60
rect 28620 -120 28720 -60
rect 28790 -120 28890 -60
rect 28960 -120 29060 -60
rect 29130 -120 29230 -60
rect 29300 -120 29400 -60
rect 29470 -120 29570 -60
rect 29640 -120 29740 -60
rect 29810 -120 29910 -60
rect 29980 -120 30080 -60
rect 30150 -120 30250 -60
rect 30320 -120 30420 -60
rect 30490 -120 30590 -60
rect 30660 -120 30760 -60
rect 30830 -120 30930 -60
rect 31000 -120 31100 -60
rect 31170 -120 31270 -60
rect 31340 -120 31440 -60
rect 31510 -120 31610 -60
rect 31680 -120 31780 -60
rect 31850 -120 31950 -60
rect 32020 -120 32120 -60
rect 32190 -120 32290 -60
rect 32360 -120 32460 -60
rect 32530 -120 32630 -60
rect 32700 -120 32800 -60
rect 32870 -120 32970 -60
rect 33040 -120 33140 -60
rect 33210 -120 33310 -60
rect 33380 -120 33480 -60
rect 33550 -120 33650 -60
rect 33720 -120 33820 -60
rect 33890 -120 33990 -60
rect 34060 -120 34160 -60
rect 34230 -120 34330 -60
rect 34400 -120 34500 -60
rect 34570 -120 34670 -60
rect 34740 -120 34840 -60
rect 34910 -120 35010 -60
rect 35080 -120 35180 -60
rect 35250 -120 35350 -60
rect 35420 -120 35520 -60
rect 35590 -120 35690 -60
rect 35760 -120 35860 -60
rect 35930 -120 36030 -60
rect 36100 -120 36200 -60
rect 36270 -120 36370 -60
rect 36440 -120 36540 -60
rect 36610 -120 36710 -60
rect 36780 -120 36880 -60
rect 36950 -120 37050 -60
rect 37120 -120 37220 -60
rect 37290 -120 37390 -60
rect 37460 -120 37560 -60
rect 37630 -120 37730 -60
rect 37800 -120 37900 -60
rect 37970 -120 38070 -60
rect 38140 -120 38240 -60
rect 38310 -120 38410 -60
rect 38480 -120 38580 -60
rect 38650 -120 38750 -60
rect 38820 -120 38920 -60
rect 38990 -120 39090 -60
rect 39160 -120 39260 -60
rect 39330 -120 39430 -60
rect 39500 -120 39600 -60
rect 39670 -120 39770 -60
rect 39840 -120 39940 -60
rect 40010 -120 40110 -60
rect 40180 -120 40280 -60
rect 40350 -120 40450 -60
rect 40520 -120 40620 -60
rect 40690 -120 40790 -60
rect 40860 -120 40960 -60
rect 41030 -120 41130 -60
rect 41200 -120 41300 -60
rect 41370 -120 41470 -60
rect 41540 -120 41640 -60
rect 41710 -120 41810 -60
rect 41880 -120 41980 -60
rect 42050 -120 42150 -60
rect 42220 -120 42320 -60
rect 42390 -120 42490 -60
rect 42560 -120 42660 -60
rect 42730 -120 42830 -60
rect 42900 -120 43000 -60
rect 43070 -120 43170 -60
rect 43240 -120 43340 -60
rect 43410 -120 43510 -60
rect 43580 -120 43680 -60
rect 43750 -120 43850 -60
rect 43920 -120 44020 -60
rect 44090 -120 44190 -60
rect 44260 -120 44360 -60
rect 44430 -120 44530 -60
rect 44600 -120 44700 -60
rect 44770 -120 44870 -60
rect 44940 -120 45040 -60
rect 45110 -120 45210 -60
rect 45280 -120 45380 -60
rect 45450 -120 45550 -60
rect 45620 -120 45720 -60
rect 45790 -120 45890 -60
rect 45960 -120 46060 -60
rect 46130 -120 46230 -60
rect 46300 -120 46400 -60
rect 46470 -120 46570 -60
rect 46640 -120 46740 -60
rect 46810 -120 46910 -60
rect 46980 -120 47080 -60
rect 47150 -120 47250 -60
rect 47320 -120 47420 -60
rect 47490 -120 47590 -60
rect 47660 -120 47760 -60
rect 47830 -120 47930 -60
rect 48000 -120 48100 -60
rect 48170 -120 48270 -60
rect 48340 -120 48440 -60
rect 48510 -120 48610 -60
rect 48680 -120 48780 -60
rect 48850 -120 48950 -60
rect 49020 -120 49120 -60
rect 49190 -120 49290 -60
rect 49360 -120 49460 -60
rect 49530 -120 49630 -60
rect 49700 -120 49800 -60
rect 49870 -120 49970 -60
rect 50040 -120 50140 -60
rect 50210 -120 50310 -60
rect 50380 -120 50480 -60
rect 50550 -120 50650 -60
rect 50720 -120 50820 -60
rect 50890 -120 50990 -60
rect 51060 -120 51160 -60
rect 51230 -120 51330 -60
rect 51400 -120 51500 -60
rect 51570 -120 51670 -60
rect 51740 -120 51840 -60
rect 51910 -120 52010 -60
rect 52080 -120 52180 -60
rect 52250 -120 52350 -60
rect 52420 -120 52520 -60
rect 52590 -120 52690 -60
rect 52760 -120 52860 -60
rect 52930 -120 53030 -60
rect 53100 -120 53200 -60
rect 53270 -120 53370 -60
rect 53440 -120 53540 -60
rect 53610 -120 53710 -60
rect 53780 -120 53880 -60
rect 53950 -120 54050 -60
rect 54120 -120 54220 -60
rect 54290 -120 54390 -60
rect 54460 -120 54560 -60
rect 54630 -120 54730 -60
rect 54800 -120 54900 -60
rect 54970 -120 55070 -60
rect 55140 -120 55240 -60
rect 55310 -120 55410 -60
rect 55480 -120 55580 -60
rect 55650 -120 55750 -60
rect 55820 -120 55920 -60
rect 55990 -120 56090 -60
rect 56160 -120 56260 -60
rect 56330 -120 56430 -60
rect 56500 -120 56600 -60
rect 56670 -120 56770 -60
rect 56840 -120 56940 -60
rect 57010 -120 57110 -60
rect 57180 -120 57280 -60
rect 57350 -120 57450 -60
rect 57520 -120 57620 -60
rect 57690 -120 57790 -60
rect 57860 -120 57960 -60
rect 58030 -120 58130 -60
rect 58200 -120 58300 -60
rect 58370 -120 58470 -60
rect 58540 -120 58640 -60
rect 58710 -120 58810 -60
rect 58880 -120 58980 -60
rect 59050 -120 59150 -60
rect 59220 -120 59240 -60
rect 15660 -130 59240 -120
rect 15550 -140 59240 -130
rect 2070 -260 2400 -240
rect 2070 -390 2120 -260
rect 2350 -390 2400 -260
rect 2070 -410 2400 -390
rect 5088 -268 5418 -248
rect 5088 -398 5138 -268
rect 5368 -398 5418 -268
rect 5088 -418 5418 -398
rect 7574 -268 7904 -248
rect 7574 -398 7624 -268
rect 7854 -398 7904 -268
rect 7574 -418 7904 -398
rect 8994 -268 9324 -248
rect 8994 -398 9044 -268
rect 9274 -398 9324 -268
rect 8994 -418 9324 -398
rect 13618 -264 13948 -244
rect 13618 -394 13668 -264
rect 13898 -394 13948 -264
rect 13618 -414 13948 -394
rect 16818 -264 17148 -244
rect 16818 -394 16868 -264
rect 17098 -394 17148 -264
rect 16818 -414 17148 -394
rect 20374 -264 20704 -244
rect 20374 -394 20424 -264
rect 20654 -394 20704 -264
rect 20374 -414 20704 -394
rect 25708 -264 26038 -244
rect 25708 -394 25758 -264
rect 25988 -394 26038 -264
rect 25708 -414 26038 -394
rect 28552 -264 28882 -244
rect 28552 -394 28602 -264
rect 28832 -394 28882 -264
rect 28552 -414 28882 -394
rect 32464 -264 32794 -244
rect 32464 -394 32514 -264
rect 32744 -394 32794 -264
rect 32464 -414 32794 -394
rect 34620 -264 34950 -244
rect 34620 -394 34670 -264
rect 34900 -394 34950 -264
rect 34620 -414 34950 -394
rect 37442 -264 37772 -244
rect 37442 -394 37492 -264
rect 37722 -394 37772 -264
rect 37442 -414 37772 -394
rect 40642 -264 40972 -244
rect 40642 -394 40692 -264
rect 40922 -394 40972 -264
rect 40642 -414 40972 -394
rect 45618 -264 45948 -244
rect 45618 -394 45668 -264
rect 45898 -394 45948 -264
rect 45618 -414 45948 -394
rect 48818 -264 49148 -244
rect 48818 -394 48868 -264
rect 49098 -394 49148 -264
rect 48818 -414 49148 -394
rect 50952 -264 51282 -244
rect 50952 -394 51002 -264
rect 51232 -394 51282 -264
rect 50952 -414 51282 -394
rect 54508 -264 54838 -244
rect 54508 -394 54558 -264
rect 54788 -394 54838 -264
rect 54508 -414 54838 -394
rect 57352 -264 57682 -244
rect 57352 -394 57402 -264
rect 57632 -394 57682 -264
rect 57352 -414 57682 -394
rect 61264 -264 61594 -244
rect 61264 -394 61314 -264
rect 61544 -394 61594 -264
rect 61264 -414 61594 -394
rect 64108 -264 64438 -244
rect 64108 -394 64158 -264
rect 64388 -394 64438 -264
rect 64108 -414 64438 -394
rect 67664 -264 67994 -244
rect 67664 -394 67714 -264
rect 67944 -394 67994 -264
rect 67664 -414 67994 -394
rect 70508 -264 70838 -244
rect 70508 -394 70558 -264
rect 70788 -394 70838 -264
rect 70508 -414 70838 -394
rect 74418 -264 74748 -244
rect 74418 -394 74468 -264
rect 74698 -394 74748 -264
rect 74418 -414 74748 -394
rect 78330 -264 78660 -244
rect 78330 -394 78380 -264
rect 78610 -394 78660 -264
rect 78330 -414 78660 -394
rect 82242 -264 82572 -244
rect 82242 -394 82292 -264
rect 82522 -394 82572 -264
rect 82242 -414 82572 -394
rect 86152 -264 86482 -244
rect 86152 -394 86202 -264
rect 86432 -394 86482 -264
rect 86152 -414 86482 -394
rect 15850 -460 16010 -450
rect 15850 -510 15930 -460
rect 210 -520 15930 -510
rect 16000 -510 16010 -460
rect 31150 -460 31310 -450
rect 31150 -510 31230 -460
rect 16000 -520 31230 -510
rect 31300 -510 31310 -460
rect 59030 -460 59190 -450
rect 59030 -510 59110 -460
rect 31300 -520 59110 -510
rect 59180 -510 59190 -460
rect 59180 -520 87250 -510
rect 210 -530 87250 -520
rect 210 -590 230 -530
rect 300 -590 400 -530
rect 470 -590 570 -530
rect 640 -590 740 -530
rect 810 -590 910 -530
rect 980 -590 1080 -530
rect 1150 -590 1250 -530
rect 1320 -590 1420 -530
rect 1490 -590 1590 -530
rect 1660 -590 1760 -530
rect 1830 -590 1930 -530
rect 2000 -590 2100 -530
rect 2170 -590 2270 -530
rect 2340 -590 2440 -530
rect 2510 -590 2610 -530
rect 2680 -590 2780 -530
rect 2850 -590 2950 -530
rect 3020 -590 3120 -530
rect 3190 -590 3290 -530
rect 3360 -590 3460 -530
rect 3530 -590 3630 -530
rect 3700 -590 3800 -530
rect 3870 -590 3970 -530
rect 4040 -590 4140 -530
rect 4210 -590 4310 -530
rect 4380 -590 4480 -530
rect 4550 -590 4650 -530
rect 4720 -590 4820 -530
rect 4890 -590 4990 -530
rect 5060 -590 5160 -530
rect 5230 -590 5330 -530
rect 5400 -590 5500 -530
rect 5570 -590 5670 -530
rect 5740 -590 5840 -530
rect 5910 -590 6010 -530
rect 6080 -590 6180 -530
rect 6250 -590 6350 -530
rect 6420 -590 6520 -530
rect 6590 -590 6690 -530
rect 6760 -590 6860 -530
rect 6930 -590 7030 -530
rect 7100 -590 7200 -530
rect 7270 -590 7370 -530
rect 7440 -590 7540 -530
rect 7610 -590 7710 -530
rect 7780 -590 7880 -530
rect 7950 -590 8050 -530
rect 8120 -590 8220 -530
rect 8290 -590 8390 -530
rect 8460 -590 8560 -530
rect 8630 -590 8730 -530
rect 8800 -590 8900 -530
rect 8970 -590 9070 -530
rect 9140 -590 9240 -530
rect 9310 -590 9410 -530
rect 9480 -590 9580 -530
rect 9650 -590 9750 -530
rect 9820 -590 9920 -530
rect 9990 -590 10090 -530
rect 10160 -590 10260 -530
rect 10330 -590 10430 -530
rect 10500 -590 10600 -530
rect 10670 -590 10770 -530
rect 10840 -590 10940 -530
rect 11010 -590 11110 -530
rect 11180 -590 11280 -530
rect 11350 -590 11450 -530
rect 11520 -590 11620 -530
rect 11690 -590 11790 -530
rect 11860 -590 11960 -530
rect 12030 -590 12130 -530
rect 12200 -590 12300 -530
rect 12370 -590 12470 -530
rect 12540 -590 12640 -530
rect 12710 -590 12810 -530
rect 12880 -590 12980 -530
rect 13050 -590 13150 -530
rect 13220 -590 13320 -530
rect 13390 -590 13490 -530
rect 13560 -590 13660 -530
rect 13730 -590 13830 -530
rect 13900 -590 14000 -530
rect 14070 -590 14170 -530
rect 14240 -590 14340 -530
rect 14410 -590 14510 -530
rect 14580 -590 14680 -530
rect 14750 -590 14850 -530
rect 14920 -590 15020 -530
rect 15090 -590 15190 -530
rect 15260 -590 15360 -530
rect 15430 -590 15530 -530
rect 15600 -590 15700 -530
rect 15770 -590 15870 -530
rect 15940 -590 16040 -530
rect 16110 -590 16210 -530
rect 16280 -590 16380 -530
rect 16450 -590 16550 -530
rect 16620 -590 16720 -530
rect 16790 -590 16890 -530
rect 16960 -590 17060 -530
rect 17130 -590 17230 -530
rect 17300 -590 17400 -530
rect 17470 -590 17570 -530
rect 17640 -590 17740 -530
rect 17810 -590 17910 -530
rect 17980 -590 18080 -530
rect 18150 -590 18250 -530
rect 18320 -590 18420 -530
rect 18490 -590 18590 -530
rect 18660 -590 18760 -530
rect 18830 -590 18930 -530
rect 19000 -590 19100 -530
rect 19170 -590 19270 -530
rect 19340 -590 19440 -530
rect 19510 -590 19610 -530
rect 19680 -590 19780 -530
rect 19850 -590 19950 -530
rect 20020 -590 20120 -530
rect 20190 -590 20290 -530
rect 20360 -590 20460 -530
rect 20530 -590 20630 -530
rect 20700 -590 20800 -530
rect 20870 -590 20970 -530
rect 21040 -590 21140 -530
rect 21210 -590 21310 -530
rect 21380 -590 21480 -530
rect 21550 -590 21650 -530
rect 21720 -590 21820 -530
rect 21890 -590 21990 -530
rect 22060 -590 22160 -530
rect 22230 -590 22330 -530
rect 22400 -590 22500 -530
rect 22570 -590 22670 -530
rect 22740 -590 22840 -530
rect 22910 -590 23010 -530
rect 23080 -590 23180 -530
rect 23250 -590 23350 -530
rect 23420 -590 23520 -530
rect 23590 -590 23690 -530
rect 23760 -590 23860 -530
rect 23930 -590 24030 -530
rect 24100 -590 24200 -530
rect 24270 -590 24370 -530
rect 24440 -590 24540 -530
rect 24610 -590 24710 -530
rect 24780 -590 24880 -530
rect 24950 -590 25050 -530
rect 25120 -590 25220 -530
rect 25290 -590 25390 -530
rect 25460 -590 25560 -530
rect 25630 -590 25730 -530
rect 25800 -590 25900 -530
rect 25970 -590 26070 -530
rect 26140 -590 26240 -530
rect 26310 -590 26410 -530
rect 26480 -590 26580 -530
rect 26650 -590 26750 -530
rect 26820 -590 26920 -530
rect 26990 -590 27090 -530
rect 27160 -590 27260 -530
rect 27330 -590 27430 -530
rect 27500 -590 27600 -530
rect 27670 -590 27770 -530
rect 27840 -590 27940 -530
rect 28010 -590 28110 -530
rect 28180 -590 28280 -530
rect 28350 -590 28450 -530
rect 28520 -590 28620 -530
rect 28690 -590 28790 -530
rect 28860 -590 28960 -530
rect 29030 -590 29130 -530
rect 29200 -590 29300 -530
rect 29370 -590 29470 -530
rect 29540 -590 29640 -530
rect 29710 -590 29810 -530
rect 29880 -590 29980 -530
rect 30050 -590 30150 -530
rect 30220 -590 30320 -530
rect 30390 -590 30490 -530
rect 30560 -590 30660 -530
rect 30730 -590 30830 -530
rect 30900 -590 31000 -530
rect 31070 -590 31170 -530
rect 31240 -590 31340 -530
rect 31410 -590 31510 -530
rect 31580 -590 31680 -530
rect 31750 -590 31850 -530
rect 31920 -590 32020 -530
rect 32090 -590 32190 -530
rect 32260 -590 32360 -530
rect 32430 -590 32530 -530
rect 32600 -590 32700 -530
rect 32770 -590 32870 -530
rect 32940 -590 33040 -530
rect 33110 -590 33210 -530
rect 33280 -590 33380 -530
rect 33450 -590 33550 -530
rect 33620 -590 33720 -530
rect 33790 -590 33890 -530
rect 33960 -590 34060 -530
rect 34130 -590 34230 -530
rect 34300 -590 34400 -530
rect 34470 -590 34570 -530
rect 34640 -590 34740 -530
rect 34810 -590 34910 -530
rect 34980 -590 35080 -530
rect 35150 -590 35250 -530
rect 35320 -590 35420 -530
rect 35490 -590 35590 -530
rect 35660 -590 35760 -530
rect 35830 -590 35930 -530
rect 36000 -590 36100 -530
rect 36170 -590 36270 -530
rect 36340 -590 36440 -530
rect 36510 -590 36610 -530
rect 36680 -590 36780 -530
rect 36850 -590 36950 -530
rect 37020 -590 37120 -530
rect 37190 -590 37290 -530
rect 37360 -590 37460 -530
rect 37530 -590 37630 -530
rect 37700 -590 37800 -530
rect 37870 -590 37970 -530
rect 38040 -590 38140 -530
rect 38210 -590 38310 -530
rect 38380 -590 38480 -530
rect 38550 -590 38650 -530
rect 38720 -590 38820 -530
rect 38890 -590 38990 -530
rect 39060 -590 39160 -530
rect 39230 -590 39330 -530
rect 39400 -590 39500 -530
rect 39570 -590 39670 -530
rect 39740 -590 39840 -530
rect 39910 -590 40010 -530
rect 40080 -590 40180 -530
rect 40250 -590 40350 -530
rect 40420 -590 40520 -530
rect 40590 -590 40690 -530
rect 40760 -590 40860 -530
rect 40930 -590 41030 -530
rect 41100 -590 41200 -530
rect 41270 -590 41370 -530
rect 41440 -590 41540 -530
rect 41610 -590 41710 -530
rect 41780 -590 41880 -530
rect 41950 -590 42050 -530
rect 42120 -590 42220 -530
rect 42290 -590 42390 -530
rect 42460 -590 42560 -530
rect 42630 -590 42730 -530
rect 42800 -590 42900 -530
rect 42970 -590 43070 -530
rect 43140 -590 43240 -530
rect 43310 -590 43410 -530
rect 43480 -590 43580 -530
rect 43650 -590 43750 -530
rect 43820 -590 43920 -530
rect 43990 -590 44090 -530
rect 44160 -590 44260 -530
rect 44330 -590 44430 -530
rect 44500 -590 44600 -530
rect 44670 -590 44770 -530
rect 44840 -590 44940 -530
rect 45010 -590 45110 -530
rect 45180 -590 45280 -530
rect 45350 -590 45450 -530
rect 45520 -590 45620 -530
rect 45690 -590 45790 -530
rect 45860 -590 45960 -530
rect 46030 -590 46130 -530
rect 46200 -590 46300 -530
rect 46370 -590 46470 -530
rect 46540 -590 46640 -530
rect 46710 -590 46810 -530
rect 46880 -590 46980 -530
rect 47050 -590 47150 -530
rect 47220 -590 47320 -530
rect 47390 -590 47490 -530
rect 47560 -590 47660 -530
rect 47730 -590 47830 -530
rect 47900 -590 48000 -530
rect 48070 -590 48170 -530
rect 48240 -590 48340 -530
rect 48410 -590 48510 -530
rect 48580 -590 48680 -530
rect 48750 -590 48850 -530
rect 48920 -590 49020 -530
rect 49090 -590 49190 -530
rect 49260 -590 49360 -530
rect 49430 -590 49530 -530
rect 49600 -590 49700 -530
rect 49770 -590 49870 -530
rect 49940 -590 50040 -530
rect 50110 -590 50210 -530
rect 50280 -590 50380 -530
rect 50450 -590 50550 -530
rect 50620 -590 50720 -530
rect 50790 -590 50890 -530
rect 50960 -590 51060 -530
rect 51130 -590 51230 -530
rect 51300 -590 51400 -530
rect 51470 -590 51570 -530
rect 51640 -590 51740 -530
rect 51810 -590 51910 -530
rect 51980 -590 52080 -530
rect 52150 -590 52250 -530
rect 52320 -590 52420 -530
rect 52490 -590 52590 -530
rect 52660 -590 52760 -530
rect 52830 -590 52930 -530
rect 53000 -590 53100 -530
rect 53170 -590 53270 -530
rect 53340 -590 53440 -530
rect 53510 -590 53610 -530
rect 53680 -590 53780 -530
rect 53850 -590 53950 -530
rect 54020 -590 54120 -530
rect 54190 -590 54290 -530
rect 54360 -590 54460 -530
rect 54530 -590 54630 -530
rect 54700 -590 54800 -530
rect 54870 -590 54970 -530
rect 55040 -590 55140 -530
rect 55210 -590 55310 -530
rect 55380 -590 55480 -530
rect 55550 -590 55650 -530
rect 55720 -590 55820 -530
rect 55890 -590 55990 -530
rect 56060 -590 56160 -530
rect 56230 -590 56330 -530
rect 56400 -590 56500 -530
rect 56570 -590 56670 -530
rect 56740 -590 56840 -530
rect 56910 -590 57010 -530
rect 57080 -590 57180 -530
rect 57250 -590 57350 -530
rect 57420 -590 57520 -530
rect 57590 -590 57690 -530
rect 57760 -590 57860 -530
rect 57930 -590 58030 -530
rect 58100 -590 58200 -530
rect 58270 -590 58370 -530
rect 58440 -590 58540 -530
rect 58610 -590 58710 -530
rect 58780 -590 58880 -530
rect 58950 -590 59050 -530
rect 59120 -590 59220 -530
rect 59290 -590 59390 -530
rect 59460 -590 59560 -530
rect 59630 -590 59730 -530
rect 59800 -590 59900 -530
rect 59970 -590 60070 -530
rect 60140 -590 60240 -530
rect 60310 -590 60410 -530
rect 60480 -590 60580 -530
rect 60650 -590 60750 -530
rect 60820 -590 60920 -530
rect 60990 -590 61090 -530
rect 61160 -590 61260 -530
rect 61330 -590 61430 -530
rect 61500 -590 61600 -530
rect 61670 -590 61770 -530
rect 61840 -590 61940 -530
rect 62010 -590 62110 -530
rect 62180 -590 62280 -530
rect 62350 -590 62450 -530
rect 62520 -590 62620 -530
rect 62690 -590 62790 -530
rect 62860 -590 62960 -530
rect 63030 -590 63130 -530
rect 63200 -590 63300 -530
rect 63370 -590 63470 -530
rect 63540 -590 63640 -530
rect 63710 -590 63810 -530
rect 63880 -590 63980 -530
rect 64050 -590 64150 -530
rect 64220 -590 64320 -530
rect 64390 -590 64490 -530
rect 64560 -590 64660 -530
rect 64730 -590 64830 -530
rect 64900 -590 65000 -530
rect 65070 -590 65170 -530
rect 65240 -590 65340 -530
rect 65410 -590 65510 -530
rect 65580 -590 65680 -530
rect 65750 -590 65850 -530
rect 65920 -590 66020 -530
rect 66090 -590 66190 -530
rect 66260 -590 66360 -530
rect 66430 -590 66530 -530
rect 66600 -590 66700 -530
rect 66770 -590 66870 -530
rect 66940 -590 67040 -530
rect 67110 -590 67210 -530
rect 67280 -590 67380 -530
rect 67450 -590 67550 -530
rect 67620 -590 67720 -530
rect 67790 -590 67890 -530
rect 67960 -590 68060 -530
rect 68130 -590 68230 -530
rect 68300 -590 68400 -530
rect 68470 -590 68570 -530
rect 68640 -590 68740 -530
rect 68810 -590 68910 -530
rect 68980 -590 69080 -530
rect 69150 -590 69250 -530
rect 69320 -590 69420 -530
rect 69490 -590 69590 -530
rect 69660 -590 69760 -530
rect 69830 -590 69930 -530
rect 70000 -590 70100 -530
rect 70170 -590 70270 -530
rect 70340 -590 70440 -530
rect 70510 -590 70610 -530
rect 70680 -590 70780 -530
rect 70850 -590 70950 -530
rect 71020 -590 71120 -530
rect 71190 -590 71290 -530
rect 71360 -590 71460 -530
rect 71530 -590 71630 -530
rect 71700 -590 71800 -530
rect 71870 -590 71970 -530
rect 72040 -590 72140 -530
rect 72210 -590 72310 -530
rect 72380 -590 72480 -530
rect 72550 -590 72650 -530
rect 72720 -590 72820 -530
rect 72890 -590 72990 -530
rect 73060 -590 73160 -530
rect 73230 -590 73330 -530
rect 73400 -590 73500 -530
rect 73570 -590 73670 -530
rect 73740 -590 73840 -530
rect 73910 -590 74010 -530
rect 74080 -590 74180 -530
rect 74250 -590 74350 -530
rect 74420 -590 74520 -530
rect 74590 -590 74690 -530
rect 74760 -590 74860 -530
rect 74930 -590 75030 -530
rect 75100 -590 75200 -530
rect 75270 -590 75370 -530
rect 75440 -590 75540 -530
rect 75610 -590 75710 -530
rect 75780 -590 75880 -530
rect 75950 -590 76050 -530
rect 76120 -590 76220 -530
rect 76290 -590 76390 -530
rect 76460 -590 76560 -530
rect 76630 -590 76730 -530
rect 76800 -590 76900 -530
rect 76970 -590 77070 -530
rect 77140 -590 77240 -530
rect 77310 -590 77410 -530
rect 77480 -590 77580 -530
rect 77650 -590 77750 -530
rect 77820 -590 77920 -530
rect 77990 -590 78090 -530
rect 78160 -590 78260 -530
rect 78330 -590 78430 -530
rect 78500 -590 78600 -530
rect 78670 -590 78770 -530
rect 78840 -590 78940 -530
rect 79010 -590 79110 -530
rect 79180 -590 79280 -530
rect 79350 -590 79450 -530
rect 79520 -590 79620 -530
rect 79690 -590 79790 -530
rect 79860 -590 79960 -530
rect 80030 -590 80130 -530
rect 80200 -590 80300 -530
rect 80370 -590 80470 -530
rect 80540 -590 80640 -530
rect 80710 -590 80810 -530
rect 80880 -590 80980 -530
rect 81050 -590 81150 -530
rect 81220 -590 81320 -530
rect 81390 -590 81490 -530
rect 81560 -590 81660 -530
rect 81730 -590 81830 -530
rect 81900 -590 82000 -530
rect 82070 -590 82170 -530
rect 82240 -590 82340 -530
rect 82410 -590 82510 -530
rect 82580 -590 82680 -530
rect 82750 -590 82850 -530
rect 82920 -590 83020 -530
rect 83090 -590 83190 -530
rect 83260 -590 83360 -530
rect 83430 -590 83530 -530
rect 83600 -590 83700 -530
rect 83770 -590 83870 -530
rect 83940 -590 84040 -530
rect 84110 -590 84210 -530
rect 84280 -590 84380 -530
rect 84450 -590 84550 -530
rect 84620 -590 84720 -530
rect 84790 -590 84890 -530
rect 84960 -590 85060 -530
rect 85130 -590 85230 -530
rect 85300 -590 85400 -530
rect 85470 -590 85570 -530
rect 85640 -590 85740 -530
rect 85810 -590 85910 -530
rect 85980 -590 86080 -530
rect 86150 -590 86250 -530
rect 86320 -590 86420 -530
rect 86490 -590 86590 -530
rect 86660 -590 86760 -530
rect 86830 -590 86930 -530
rect 87000 -590 87100 -530
rect 87170 -590 87250 -530
rect 210 -610 87250 -590
rect 130 -670 230 -650
rect 470 -670 570 -650
rect 810 -670 910 -650
rect 1150 -670 1250 -650
rect 1490 -670 1590 -650
rect 1830 -670 1930 -650
rect 2170 -670 2270 -650
rect 2510 -670 2610 -650
rect 2850 -670 2950 -650
rect 3190 -670 3290 -650
rect 3530 -670 3630 -650
rect 3870 -670 3970 -650
rect 4210 -670 4310 -650
rect 4550 -670 4650 -650
rect 4890 -670 4990 -650
rect 5230 -670 5330 -650
rect 5570 -670 5670 -650
rect 5910 -670 6010 -650
rect 6250 -670 6350 -650
rect 6590 -670 6690 -650
rect 6930 -670 7030 -650
rect 7270 -670 7370 -650
rect 7610 -670 7710 -650
rect 7950 -670 8050 -650
rect 8290 -670 8390 -650
rect 8630 -670 8730 -650
rect 8970 -670 9070 -650
rect 9310 -670 9410 -650
rect 9650 -670 9750 -650
rect 9990 -670 10090 -650
rect 10330 -670 10430 -650
rect 10670 -670 10770 -650
rect 11010 -670 11110 -650
rect 11350 -670 11450 -650
rect 11690 -670 11790 -650
rect 12030 -670 12130 -650
rect 12370 -670 12470 -650
rect 12710 -670 12810 -650
rect 13050 -670 13150 -650
rect 13390 -670 13490 -650
rect 13730 -670 13830 -650
rect 14070 -670 14170 -650
rect 14410 -670 14510 -650
rect 14750 -670 14850 -650
rect 15090 -670 15190 -650
rect 15430 -670 15530 -650
rect 15770 -670 15870 -650
rect 16110 -670 16210 -650
rect 16450 -670 16550 -650
rect 16790 -670 16890 -650
rect 17130 -670 17230 -650
rect 17470 -670 17570 -650
rect 17810 -670 17910 -650
rect 18150 -670 18250 -650
rect 18490 -670 18590 -650
rect 18830 -670 18930 -650
rect 19170 -670 19270 -650
rect 19510 -670 19610 -650
rect 19850 -670 19950 -650
rect 20190 -670 20290 -650
rect 20530 -670 20630 -650
rect 20870 -670 20970 -650
rect 21210 -670 21310 -650
rect 21550 -670 21650 -650
rect 21890 -670 21990 -650
rect 22230 -670 22330 -650
rect 22570 -670 22670 -650
rect 22910 -670 23010 -650
rect 23250 -670 23350 -650
rect 23590 -670 23690 -650
rect 23930 -670 24030 -650
rect 24270 -670 24370 -650
rect 24610 -670 24710 -650
rect 24950 -670 25050 -650
rect 25290 -670 25390 -650
rect 25630 -670 25730 -650
rect 25970 -670 26070 -650
rect 26310 -670 26410 -650
rect 26650 -670 26750 -650
rect 26990 -670 27090 -650
rect 27330 -670 27430 -650
rect 27670 -670 27770 -650
rect 28010 -670 28110 -650
rect 28350 -670 28450 -650
rect 28690 -670 28790 -650
rect 29030 -670 29130 -650
rect 29370 -670 29470 -650
rect 29710 -670 29810 -650
rect 30050 -670 30150 -650
rect 30390 -670 30490 -650
rect 30730 -670 30830 -650
rect 31070 -670 31170 -650
rect 31410 -670 31510 -650
rect 31750 -670 31850 -650
rect 32090 -670 32190 -650
rect 32430 -670 32530 -650
rect 32770 -670 32870 -650
rect 33110 -670 33210 -650
rect 33450 -670 33550 -650
rect 33790 -670 33890 -650
rect 34130 -670 34230 -650
rect 34470 -670 34570 -650
rect 34810 -670 34910 -650
rect 35150 -670 35250 -650
rect 35490 -670 35590 -650
rect 35830 -670 35930 -650
rect 36170 -670 36270 -650
rect 36510 -670 36610 -650
rect 36850 -670 36950 -650
rect 37190 -670 37290 -650
rect 37530 -670 37630 -650
rect 37870 -670 37970 -650
rect 38210 -670 38310 -650
rect 38550 -670 38650 -650
rect 38890 -670 38990 -650
rect 39230 -670 39330 -650
rect 39570 -670 39670 -650
rect 39910 -670 40010 -650
rect 40250 -670 40350 -650
rect 40590 -670 40690 -650
rect 40930 -670 41030 -650
rect 41270 -670 41370 -650
rect 41610 -670 41710 -650
rect 41950 -670 42050 -650
rect 42290 -670 42390 -650
rect 42630 -670 42730 -650
rect 42970 -670 43070 -650
rect 43310 -670 43410 -650
rect 43650 -670 43750 -650
rect 43990 -670 44090 -650
rect 44330 -670 44430 -650
rect 44670 -670 44770 -650
rect 45010 -670 45110 -650
rect 45350 -670 45450 -650
rect 45690 -670 45790 -650
rect 46030 -670 46130 -650
rect 46370 -670 46470 -650
rect 46710 -670 46810 -650
rect 47050 -670 47150 -650
rect 47390 -670 47490 -650
rect 47730 -670 47830 -650
rect 48070 -670 48170 -650
rect 48410 -670 48510 -650
rect 48750 -670 48850 -650
rect 49090 -670 49190 -650
rect 49430 -670 49530 -650
rect 49770 -670 49870 -650
rect 50110 -670 50210 -650
rect 50450 -670 50550 -650
rect 50790 -670 50890 -650
rect 51130 -670 51230 -650
rect 51470 -670 51570 -650
rect 51810 -670 51910 -650
rect 52150 -670 52250 -650
rect 52490 -670 52590 -650
rect 52830 -670 52930 -650
rect 53170 -670 53270 -650
rect 53510 -670 53610 -650
rect 53850 -670 53950 -650
rect 54190 -670 54290 -650
rect 54530 -670 54630 -650
rect 54870 -670 54970 -650
rect 55210 -670 55310 -650
rect 55550 -670 55650 -650
rect 55890 -670 55990 -650
rect 56230 -670 56330 -650
rect 56570 -670 56670 -650
rect 56910 -670 57010 -650
rect 57250 -670 57350 -650
rect 57590 -670 57690 -650
rect 57930 -670 58030 -650
rect 58270 -670 58370 -650
rect 58610 -670 58710 -650
rect 58950 -670 59050 -650
rect 59290 -670 59390 -650
rect 59630 -670 59730 -650
rect 59970 -670 60070 -650
rect 60310 -670 60410 -650
rect 60650 -670 60750 -650
rect 60990 -670 61090 -650
rect 61330 -670 61430 -650
rect 61670 -670 61770 -650
rect 62010 -670 62110 -650
rect 62350 -670 62450 -650
rect 62690 -670 62790 -650
rect 63030 -670 63130 -650
rect 63370 -670 63470 -650
rect 63710 -670 63810 -650
rect 64050 -670 64150 -650
rect 64390 -670 64490 -650
rect 64730 -670 64830 -650
rect 65070 -670 65170 -650
rect 65410 -670 65510 -650
rect 65750 -670 65850 -650
rect 66090 -670 66190 -650
rect 66430 -670 66530 -650
rect 66770 -670 66870 -650
rect 67110 -670 67210 -650
rect 67450 -670 67550 -650
rect 67790 -670 67890 -650
rect 68130 -670 68230 -650
rect 68470 -670 68570 -650
rect 68810 -670 68910 -650
rect 69150 -670 69250 -650
rect 69490 -670 69590 -650
rect 69830 -670 69930 -650
rect 70170 -670 70270 -650
rect 70510 -670 70610 -650
rect 70850 -670 70950 -650
rect 71190 -670 71290 -650
rect 71530 -670 71630 -650
rect 71870 -670 71970 -650
rect 72210 -670 72310 -650
rect 72550 -670 72650 -650
rect 72890 -670 72990 -650
rect 73230 -670 73330 -650
rect 73570 -670 73670 -650
rect 73910 -670 74010 -650
rect 74250 -670 74350 -650
rect 74590 -670 74690 -650
rect 74930 -670 75030 -650
rect 75270 -670 75370 -650
rect 75610 -670 75710 -650
rect 75950 -670 76050 -650
rect 76290 -670 76390 -650
rect 76630 -670 76730 -650
rect 76970 -670 77070 -650
rect 77310 -670 77410 -650
rect 77650 -670 77750 -650
rect 77990 -670 78090 -650
rect 78330 -670 78430 -650
rect 78670 -670 78770 -650
rect 79010 -670 79110 -650
rect 79350 -670 79450 -650
rect 79690 -670 79790 -650
rect 80030 -670 80130 -650
rect 80370 -670 80470 -650
rect 80710 -670 80810 -650
rect 81050 -670 81150 -650
rect 81390 -670 81490 -650
rect 81730 -670 81830 -650
rect 82070 -670 82170 -650
rect 82410 -670 82510 -650
rect 82750 -670 82850 -650
rect 83090 -670 83190 -650
rect 83430 -670 83530 -650
rect 83770 -670 83870 -650
rect 84110 -670 84210 -650
rect 84450 -670 84550 -650
rect 84790 -670 84890 -650
rect 85130 -670 85230 -650
rect 85470 -670 85570 -650
rect 85810 -670 85910 -650
rect 86150 -670 86250 -650
rect 86490 -670 86590 -650
rect 86830 -670 86930 -650
rect 87170 -670 87270 -650
rect 130 -730 150 -670
rect 210 -730 490 -670
rect 550 -730 830 -670
rect 890 -730 1170 -670
rect 1230 -730 1510 -670
rect 1570 -730 1850 -670
rect 1910 -730 2190 -670
rect 2250 -730 2530 -670
rect 2590 -730 2870 -670
rect 2930 -730 3210 -670
rect 3270 -730 3550 -670
rect 3610 -730 3890 -670
rect 3950 -730 4230 -670
rect 4290 -730 4570 -670
rect 4630 -730 4910 -670
rect 4970 -730 5250 -670
rect 5310 -730 5590 -670
rect 5650 -730 5930 -670
rect 5990 -730 6270 -670
rect 6330 -730 6610 -670
rect 6670 -730 6950 -670
rect 7010 -730 7290 -670
rect 7350 -730 7630 -670
rect 7690 -730 7970 -670
rect 8030 -730 8310 -670
rect 8370 -730 8650 -670
rect 8710 -730 8990 -670
rect 9050 -730 9330 -670
rect 9390 -730 9670 -670
rect 9730 -730 10010 -670
rect 10070 -730 10350 -670
rect 10410 -730 10690 -670
rect 10750 -730 11030 -670
rect 11090 -730 11370 -670
rect 11430 -730 11710 -670
rect 11770 -730 12050 -670
rect 12110 -730 12390 -670
rect 12450 -730 12730 -670
rect 12790 -730 13070 -670
rect 13130 -730 13410 -670
rect 13470 -730 13750 -670
rect 13810 -730 14090 -670
rect 14150 -730 14430 -670
rect 14490 -730 14770 -670
rect 14830 -730 15110 -670
rect 15170 -730 15450 -670
rect 15510 -730 15790 -670
rect 15850 -730 16130 -670
rect 16190 -730 16470 -670
rect 16530 -730 16810 -670
rect 16870 -730 17150 -670
rect 17210 -730 17490 -670
rect 17550 -730 17830 -670
rect 17890 -730 18170 -670
rect 18230 -730 18510 -670
rect 18570 -730 18850 -670
rect 18910 -730 19190 -670
rect 19250 -730 19530 -670
rect 19590 -730 19870 -670
rect 19930 -730 20210 -670
rect 20270 -730 20550 -670
rect 20610 -730 20890 -670
rect 20950 -730 21230 -670
rect 21290 -730 21570 -670
rect 21630 -730 21910 -670
rect 21970 -730 22250 -670
rect 22310 -730 22590 -670
rect 22650 -730 22930 -670
rect 22990 -730 23270 -670
rect 23330 -730 23610 -670
rect 23670 -730 23950 -670
rect 24010 -730 24290 -670
rect 24350 -730 24630 -670
rect 24690 -730 24970 -670
rect 25030 -730 25310 -670
rect 25370 -730 25650 -670
rect 25710 -730 25990 -670
rect 26050 -730 26330 -670
rect 26390 -730 26670 -670
rect 26730 -730 27010 -670
rect 27070 -730 27350 -670
rect 27410 -730 27690 -670
rect 27750 -730 28030 -670
rect 28090 -730 28370 -670
rect 28430 -730 28710 -670
rect 28770 -730 29050 -670
rect 29110 -730 29390 -670
rect 29450 -730 29730 -670
rect 29790 -730 30070 -670
rect 30130 -730 30410 -670
rect 30470 -730 30750 -670
rect 30810 -730 31090 -670
rect 31150 -730 31430 -670
rect 31490 -730 31770 -670
rect 31830 -730 32110 -670
rect 32170 -730 32450 -670
rect 32510 -730 32790 -670
rect 32850 -730 33130 -670
rect 33190 -730 33470 -670
rect 33530 -730 33810 -670
rect 33870 -730 34150 -670
rect 34210 -730 34490 -670
rect 34550 -730 34830 -670
rect 34890 -730 35170 -670
rect 35230 -730 35510 -670
rect 35570 -730 35850 -670
rect 35910 -730 36190 -670
rect 36250 -730 36530 -670
rect 36590 -730 36870 -670
rect 36930 -730 37210 -670
rect 37270 -730 37550 -670
rect 37610 -730 37890 -670
rect 37950 -730 38230 -670
rect 38290 -730 38570 -670
rect 38630 -730 38910 -670
rect 38970 -730 39250 -670
rect 39310 -730 39590 -670
rect 39650 -730 39930 -670
rect 39990 -730 40270 -670
rect 40330 -730 40610 -670
rect 40670 -730 40950 -670
rect 41010 -730 41290 -670
rect 41350 -730 41630 -670
rect 41690 -730 41970 -670
rect 42030 -730 42310 -670
rect 42370 -730 42650 -670
rect 42710 -730 42990 -670
rect 43050 -730 43330 -670
rect 43390 -730 43670 -670
rect 43730 -730 44010 -670
rect 44070 -730 44350 -670
rect 44410 -730 44690 -670
rect 44750 -730 45030 -670
rect 45090 -730 45370 -670
rect 45430 -730 45710 -670
rect 45770 -730 46050 -670
rect 46110 -730 46390 -670
rect 46450 -730 46730 -670
rect 46790 -730 47070 -670
rect 47130 -730 47410 -670
rect 47470 -730 47750 -670
rect 47810 -730 48090 -670
rect 48150 -730 48430 -670
rect 48490 -730 48770 -670
rect 48830 -730 49110 -670
rect 49170 -730 49450 -670
rect 49510 -730 49790 -670
rect 49850 -730 50130 -670
rect 50190 -730 50470 -670
rect 50530 -730 50810 -670
rect 50870 -730 51150 -670
rect 51210 -730 51490 -670
rect 51550 -730 51830 -670
rect 51890 -730 52170 -670
rect 52230 -730 52510 -670
rect 52570 -730 52850 -670
rect 52910 -730 53190 -670
rect 53250 -730 53530 -670
rect 53590 -730 53870 -670
rect 53930 -730 54210 -670
rect 54270 -730 54550 -670
rect 54610 -730 54890 -670
rect 54950 -730 55230 -670
rect 55290 -730 55570 -670
rect 55630 -730 55910 -670
rect 55970 -730 56250 -670
rect 56310 -730 56590 -670
rect 56650 -730 56930 -670
rect 56990 -730 57270 -670
rect 57330 -730 57610 -670
rect 57670 -730 57950 -670
rect 58010 -730 58290 -670
rect 58350 -730 58630 -670
rect 58690 -730 58970 -670
rect 59030 -730 59310 -670
rect 59370 -730 59650 -670
rect 59710 -730 59990 -670
rect 60050 -730 60330 -670
rect 60390 -730 60670 -670
rect 60730 -730 61010 -670
rect 61070 -730 61350 -670
rect 61410 -730 61690 -670
rect 61750 -730 62030 -670
rect 62090 -730 62370 -670
rect 62430 -730 62710 -670
rect 62770 -730 63050 -670
rect 63110 -730 63390 -670
rect 63450 -730 63730 -670
rect 63790 -730 64070 -670
rect 64130 -730 64410 -670
rect 64470 -730 64750 -670
rect 64810 -730 65090 -670
rect 65150 -730 65430 -670
rect 65490 -730 65770 -670
rect 65830 -730 66110 -670
rect 66170 -730 66450 -670
rect 66510 -730 66790 -670
rect 66850 -730 67130 -670
rect 67190 -730 67470 -670
rect 67530 -730 67810 -670
rect 67870 -730 68150 -670
rect 68210 -730 68490 -670
rect 68550 -730 68830 -670
rect 68890 -730 69170 -670
rect 69230 -730 69510 -670
rect 69570 -730 69850 -670
rect 69910 -730 70190 -670
rect 70250 -730 70530 -670
rect 70590 -730 70870 -670
rect 70930 -730 71210 -670
rect 71270 -730 71550 -670
rect 71610 -730 71890 -670
rect 71950 -730 72230 -670
rect 72290 -730 72570 -670
rect 72630 -730 72910 -670
rect 72970 -730 73250 -670
rect 73310 -730 73590 -670
rect 73650 -730 73930 -670
rect 73990 -730 74270 -670
rect 74330 -730 74610 -670
rect 74670 -730 74950 -670
rect 75010 -730 75290 -670
rect 75350 -730 75630 -670
rect 75690 -730 75970 -670
rect 76030 -730 76310 -670
rect 76370 -730 76650 -670
rect 76710 -730 76990 -670
rect 77050 -730 77330 -670
rect 77390 -730 77670 -670
rect 77730 -730 78010 -670
rect 78070 -730 78350 -670
rect 78410 -730 78690 -670
rect 78750 -730 79030 -670
rect 79090 -730 79370 -670
rect 79430 -730 79710 -670
rect 79770 -730 80050 -670
rect 80110 -730 80390 -670
rect 80450 -730 80730 -670
rect 80790 -730 81070 -670
rect 81130 -730 81410 -670
rect 81470 -730 81750 -670
rect 81810 -730 82090 -670
rect 82150 -730 82430 -670
rect 82490 -730 82770 -670
rect 82830 -730 83110 -670
rect 83170 -730 83450 -670
rect 83510 -730 83790 -670
rect 83850 -730 84130 -670
rect 84190 -730 84470 -670
rect 84530 -730 84810 -670
rect 84870 -730 85150 -670
rect 85210 -730 85490 -670
rect 85550 -730 85830 -670
rect 85890 -730 86170 -670
rect 86230 -730 86510 -670
rect 86570 -730 86850 -670
rect 86910 -730 87190 -670
rect 87250 -730 87290 -670
rect 130 -750 230 -730
rect 470 -750 570 -730
rect 810 -750 910 -730
rect 1150 -750 1250 -730
rect 1490 -750 1590 -730
rect 1830 -750 1930 -730
rect 2170 -750 2270 -730
rect 2510 -750 2610 -730
rect 2850 -750 2950 -730
rect 3190 -750 3290 -730
rect 3530 -750 3630 -730
rect 3870 -750 3970 -730
rect 4210 -750 4310 -730
rect 4550 -750 4650 -730
rect 4890 -750 4990 -730
rect 5230 -750 5330 -730
rect 5570 -750 5670 -730
rect 5910 -750 6010 -730
rect 6250 -750 6350 -730
rect 6590 -750 6690 -730
rect 6930 -750 7030 -730
rect 7270 -750 7370 -730
rect 7610 -750 7710 -730
rect 7950 -750 8050 -730
rect 8290 -750 8390 -730
rect 8630 -750 8730 -730
rect 8970 -750 9070 -730
rect 9310 -750 9410 -730
rect 9650 -750 9750 -730
rect 9990 -750 10090 -730
rect 10330 -750 10430 -730
rect 10670 -750 10770 -730
rect 11010 -750 11110 -730
rect 11350 -750 11450 -730
rect 11690 -750 11790 -730
rect 12030 -750 12130 -730
rect 12370 -750 12470 -730
rect 12710 -750 12810 -730
rect 13050 -750 13150 -730
rect 13390 -750 13490 -730
rect 13730 -750 13830 -730
rect 14070 -750 14170 -730
rect 14410 -750 14510 -730
rect 14750 -750 14850 -730
rect 15090 -750 15190 -730
rect 15430 -750 15530 -730
rect 15770 -750 15870 -730
rect 16110 -750 16210 -730
rect 16450 -750 16550 -730
rect 16790 -750 16890 -730
rect 17130 -750 17230 -730
rect 17470 -750 17570 -730
rect 17810 -750 17910 -730
rect 18150 -750 18250 -730
rect 18490 -750 18590 -730
rect 18830 -750 18930 -730
rect 19170 -750 19270 -730
rect 19510 -750 19610 -730
rect 19850 -750 19950 -730
rect 20190 -750 20290 -730
rect 20530 -750 20630 -730
rect 20870 -750 20970 -730
rect 21210 -750 21310 -730
rect 21550 -750 21650 -730
rect 21890 -750 21990 -730
rect 22230 -750 22330 -730
rect 22570 -750 22670 -730
rect 22910 -750 23010 -730
rect 23250 -750 23350 -730
rect 23590 -750 23690 -730
rect 23930 -750 24030 -730
rect 24270 -750 24370 -730
rect 24610 -750 24710 -730
rect 24950 -750 25050 -730
rect 25290 -750 25390 -730
rect 25630 -750 25730 -730
rect 25970 -750 26070 -730
rect 26310 -750 26410 -730
rect 26650 -750 26750 -730
rect 26990 -750 27090 -730
rect 27330 -750 27430 -730
rect 27670 -750 27770 -730
rect 28010 -750 28110 -730
rect 28350 -750 28450 -730
rect 28690 -750 28790 -730
rect 29030 -750 29130 -730
rect 29370 -750 29470 -730
rect 29710 -750 29810 -730
rect 30050 -750 30150 -730
rect 30390 -750 30490 -730
rect 30730 -750 30830 -730
rect 31070 -750 31170 -730
rect 31410 -750 31510 -730
rect 31750 -750 31850 -730
rect 32090 -750 32190 -730
rect 32430 -750 32530 -730
rect 32770 -750 32870 -730
rect 33110 -750 33210 -730
rect 33450 -750 33550 -730
rect 33790 -750 33890 -730
rect 34130 -750 34230 -730
rect 34470 -750 34570 -730
rect 34810 -750 34910 -730
rect 35150 -750 35250 -730
rect 35490 -750 35590 -730
rect 35830 -750 35930 -730
rect 36170 -750 36270 -730
rect 36510 -750 36610 -730
rect 36850 -750 36950 -730
rect 37190 -750 37290 -730
rect 37530 -750 37630 -730
rect 37870 -750 37970 -730
rect 38210 -750 38310 -730
rect 38550 -750 38650 -730
rect 38890 -750 38990 -730
rect 39230 -750 39330 -730
rect 39570 -750 39670 -730
rect 39910 -750 40010 -730
rect 40250 -750 40350 -730
rect 40590 -750 40690 -730
rect 40930 -750 41030 -730
rect 41270 -750 41370 -730
rect 41610 -750 41710 -730
rect 41950 -750 42050 -730
rect 42290 -750 42390 -730
rect 42630 -750 42730 -730
rect 42970 -750 43070 -730
rect 43310 -750 43410 -730
rect 43650 -750 43750 -730
rect 43990 -750 44090 -730
rect 44330 -750 44430 -730
rect 44670 -750 44770 -730
rect 45010 -750 45110 -730
rect 45350 -750 45450 -730
rect 45690 -750 45790 -730
rect 46030 -750 46130 -730
rect 46370 -750 46470 -730
rect 46710 -750 46810 -730
rect 47050 -750 47150 -730
rect 47390 -750 47490 -730
rect 47730 -750 47830 -730
rect 48070 -750 48170 -730
rect 48410 -750 48510 -730
rect 48750 -750 48850 -730
rect 49090 -750 49190 -730
rect 49430 -750 49530 -730
rect 49770 -750 49870 -730
rect 50110 -750 50210 -730
rect 50450 -750 50550 -730
rect 50790 -750 50890 -730
rect 51130 -750 51230 -730
rect 51470 -750 51570 -730
rect 51810 -750 51910 -730
rect 52150 -750 52250 -730
rect 52490 -750 52590 -730
rect 52830 -750 52930 -730
rect 53170 -750 53270 -730
rect 53510 -750 53610 -730
rect 53850 -750 53950 -730
rect 54190 -750 54290 -730
rect 54530 -750 54630 -730
rect 54870 -750 54970 -730
rect 55210 -750 55310 -730
rect 55550 -750 55650 -730
rect 55890 -750 55990 -730
rect 56230 -750 56330 -730
rect 56570 -750 56670 -730
rect 56910 -750 57010 -730
rect 57250 -750 57350 -730
rect 57590 -750 57690 -730
rect 57930 -750 58030 -730
rect 58270 -750 58370 -730
rect 58610 -750 58710 -730
rect 58950 -750 59050 -730
rect 59290 -750 59390 -730
rect 59630 -750 59730 -730
rect 59970 -750 60070 -730
rect 60310 -750 60410 -730
rect 60650 -750 60750 -730
rect 60990 -750 61090 -730
rect 61330 -750 61430 -730
rect 61670 -750 61770 -730
rect 62010 -750 62110 -730
rect 62350 -750 62450 -730
rect 62690 -750 62790 -730
rect 63030 -750 63130 -730
rect 63370 -750 63470 -730
rect 63710 -750 63810 -730
rect 64050 -750 64150 -730
rect 64390 -750 64490 -730
rect 64730 -750 64830 -730
rect 65070 -750 65170 -730
rect 65410 -750 65510 -730
rect 65750 -750 65850 -730
rect 66090 -750 66190 -730
rect 66430 -750 66530 -730
rect 66770 -750 66870 -730
rect 67110 -750 67210 -730
rect 67450 -750 67550 -730
rect 67790 -750 67890 -730
rect 68130 -750 68230 -730
rect 68470 -750 68570 -730
rect 68810 -750 68910 -730
rect 69150 -750 69250 -730
rect 69490 -750 69590 -730
rect 69830 -750 69930 -730
rect 70170 -750 70270 -730
rect 70510 -750 70610 -730
rect 70850 -750 70950 -730
rect 71190 -750 71290 -730
rect 71530 -750 71630 -730
rect 71870 -750 71970 -730
rect 72210 -750 72310 -730
rect 72550 -750 72650 -730
rect 72890 -750 72990 -730
rect 73230 -750 73330 -730
rect 73570 -750 73670 -730
rect 73910 -750 74010 -730
rect 74250 -750 74350 -730
rect 74590 -750 74690 -730
rect 74930 -750 75030 -730
rect 75270 -750 75370 -730
rect 75610 -750 75710 -730
rect 75950 -750 76050 -730
rect 76290 -750 76390 -730
rect 76630 -750 76730 -730
rect 76970 -750 77070 -730
rect 77310 -750 77410 -730
rect 77650 -750 77750 -730
rect 77990 -750 78090 -730
rect 78330 -750 78430 -730
rect 78670 -750 78770 -730
rect 79010 -750 79110 -730
rect 79350 -750 79450 -730
rect 79690 -750 79790 -730
rect 80030 -750 80130 -730
rect 80370 -750 80470 -730
rect 80710 -750 80810 -730
rect 81050 -750 81150 -730
rect 81390 -750 81490 -730
rect 81730 -750 81830 -730
rect 82070 -750 82170 -730
rect 82410 -750 82510 -730
rect 82750 -750 82850 -730
rect 83090 -750 83190 -730
rect 83430 -750 83530 -730
rect 83770 -750 83870 -730
rect 84110 -750 84210 -730
rect 84450 -750 84550 -730
rect 84790 -750 84890 -730
rect 85130 -750 85230 -730
rect 85470 -750 85570 -730
rect 85810 -750 85910 -730
rect 86150 -750 86250 -730
rect 86490 -750 86590 -730
rect 86830 -750 86930 -730
rect 87170 -750 87270 -730
rect 310 -880 390 -870
rect 310 -950 320 -880
rect 380 -950 390 -880
rect 310 -960 390 -950
rect 650 -880 730 -870
rect 650 -950 660 -880
rect 720 -950 730 -880
rect 650 -960 730 -950
rect 990 -880 1070 -870
rect 990 -950 1000 -880
rect 1060 -950 1070 -880
rect 990 -960 1070 -950
rect 1330 -880 1410 -870
rect 1330 -950 1340 -880
rect 1400 -950 1410 -880
rect 1330 -960 1410 -950
rect 1670 -880 1750 -870
rect 1670 -950 1680 -880
rect 1740 -950 1750 -880
rect 1670 -960 1750 -950
rect 2010 -880 2090 -870
rect 2010 -950 2020 -880
rect 2080 -950 2090 -880
rect 2010 -960 2090 -950
rect 2350 -880 2430 -870
rect 2350 -950 2360 -880
rect 2420 -950 2430 -880
rect 2350 -960 2430 -950
rect 2690 -880 2770 -870
rect 2690 -950 2700 -880
rect 2760 -950 2770 -880
rect 2690 -960 2770 -950
rect 3030 -880 3110 -870
rect 3030 -950 3040 -880
rect 3100 -950 3110 -880
rect 3030 -960 3110 -950
rect 3370 -880 3450 -870
rect 3370 -950 3380 -880
rect 3440 -950 3450 -880
rect 3370 -960 3450 -950
rect 3710 -880 3790 -870
rect 3710 -950 3720 -880
rect 3780 -950 3790 -880
rect 3710 -960 3790 -950
rect 4050 -880 4130 -870
rect 4050 -950 4060 -880
rect 4120 -950 4130 -880
rect 4050 -960 4130 -950
rect 4390 -880 4470 -870
rect 4390 -950 4400 -880
rect 4460 -950 4470 -880
rect 4390 -960 4470 -950
rect 4730 -880 4810 -870
rect 4730 -950 4740 -880
rect 4800 -950 4810 -880
rect 4730 -960 4810 -950
rect 5070 -880 5150 -870
rect 5070 -950 5080 -880
rect 5140 -950 5150 -880
rect 5070 -960 5150 -950
rect 5410 -880 5490 -870
rect 5410 -950 5420 -880
rect 5480 -950 5490 -880
rect 5410 -960 5490 -950
rect 5750 -880 5830 -870
rect 5750 -950 5760 -880
rect 5820 -950 5830 -880
rect 5750 -960 5830 -950
rect 6090 -880 6170 -870
rect 6090 -950 6100 -880
rect 6160 -950 6170 -880
rect 6090 -960 6170 -950
rect 6430 -880 6510 -870
rect 6430 -950 6440 -880
rect 6500 -950 6510 -880
rect 6430 -960 6510 -950
rect 6770 -880 6850 -870
rect 6770 -950 6780 -880
rect 6840 -950 6850 -880
rect 6770 -960 6850 -950
rect 7110 -880 7190 -870
rect 7110 -950 7120 -880
rect 7180 -950 7190 -880
rect 7110 -960 7190 -950
rect 7450 -880 7530 -870
rect 7450 -950 7460 -880
rect 7520 -950 7530 -880
rect 7450 -960 7530 -950
rect 7790 -880 7870 -870
rect 7790 -950 7800 -880
rect 7860 -950 7870 -880
rect 7790 -960 7870 -950
rect 8130 -880 8210 -870
rect 8130 -950 8140 -880
rect 8200 -950 8210 -880
rect 8130 -960 8210 -950
rect 8470 -880 8550 -870
rect 8470 -950 8480 -880
rect 8540 -950 8550 -880
rect 8470 -960 8550 -950
rect 8810 -880 8890 -870
rect 8810 -950 8820 -880
rect 8880 -950 8890 -880
rect 8810 -960 8890 -950
rect 9150 -880 9230 -870
rect 9150 -950 9160 -880
rect 9220 -950 9230 -880
rect 9150 -960 9230 -950
rect 9490 -880 9570 -870
rect 9490 -950 9500 -880
rect 9560 -950 9570 -880
rect 9490 -960 9570 -950
rect 9830 -880 9910 -870
rect 9830 -950 9840 -880
rect 9900 -950 9910 -880
rect 9830 -960 9910 -950
rect 10170 -880 10250 -870
rect 10170 -950 10180 -880
rect 10240 -950 10250 -880
rect 10170 -960 10250 -950
rect 10510 -880 10590 -870
rect 10510 -950 10520 -880
rect 10580 -950 10590 -880
rect 10510 -960 10590 -950
rect 10850 -880 10930 -870
rect 10850 -950 10860 -880
rect 10920 -950 10930 -880
rect 10850 -960 10930 -950
rect 11190 -880 11270 -870
rect 11190 -950 11200 -880
rect 11260 -950 11270 -880
rect 11190 -960 11270 -950
rect 11530 -880 11610 -870
rect 11530 -950 11540 -880
rect 11600 -950 11610 -880
rect 11530 -960 11610 -950
rect 11870 -880 11950 -870
rect 11870 -950 11880 -880
rect 11940 -950 11950 -880
rect 11870 -960 11950 -950
rect 12210 -880 12290 -870
rect 12210 -950 12220 -880
rect 12280 -950 12290 -880
rect 12210 -960 12290 -950
rect 12550 -880 12630 -870
rect 12550 -950 12560 -880
rect 12620 -950 12630 -880
rect 12550 -960 12630 -950
rect 12890 -880 12970 -870
rect 12890 -950 12900 -880
rect 12960 -950 12970 -880
rect 12890 -960 12970 -950
rect 13230 -880 13310 -870
rect 13230 -950 13240 -880
rect 13300 -950 13310 -880
rect 13230 -960 13310 -950
rect 13570 -880 13650 -870
rect 13570 -950 13580 -880
rect 13640 -950 13650 -880
rect 13570 -960 13650 -950
rect 13910 -880 13990 -870
rect 13910 -950 13920 -880
rect 13980 -950 13990 -880
rect 13910 -960 13990 -950
rect 14250 -880 14330 -870
rect 14250 -950 14260 -880
rect 14320 -950 14330 -880
rect 14250 -960 14330 -950
rect 14590 -880 14670 -870
rect 14590 -950 14600 -880
rect 14660 -950 14670 -880
rect 14590 -960 14670 -950
rect 14930 -880 15010 -870
rect 14930 -950 14940 -880
rect 15000 -950 15010 -880
rect 14930 -960 15010 -950
rect 15270 -880 15350 -870
rect 15270 -950 15280 -880
rect 15340 -950 15350 -880
rect 15270 -960 15350 -950
rect 15610 -880 15690 -870
rect 15610 -950 15620 -880
rect 15680 -950 15690 -880
rect 15610 -960 15690 -950
rect 15950 -880 16030 -870
rect 15950 -950 15960 -880
rect 16020 -950 16030 -880
rect 15950 -960 16030 -950
rect 16290 -880 16370 -870
rect 16290 -950 16300 -880
rect 16360 -950 16370 -880
rect 16290 -960 16370 -950
rect 16630 -880 16710 -870
rect 16630 -950 16640 -880
rect 16700 -950 16710 -880
rect 16630 -960 16710 -950
rect 16970 -880 17050 -870
rect 16970 -950 16980 -880
rect 17040 -950 17050 -880
rect 16970 -960 17050 -950
rect 17310 -880 17390 -870
rect 17310 -950 17320 -880
rect 17380 -950 17390 -880
rect 17310 -960 17390 -950
rect 17650 -880 17730 -870
rect 17650 -950 17660 -880
rect 17720 -950 17730 -880
rect 17650 -960 17730 -950
rect 17990 -880 18070 -870
rect 17990 -950 18000 -880
rect 18060 -950 18070 -880
rect 17990 -960 18070 -950
rect 18330 -880 18410 -870
rect 18330 -950 18340 -880
rect 18400 -950 18410 -880
rect 18330 -960 18410 -950
rect 18670 -880 18750 -870
rect 18670 -950 18680 -880
rect 18740 -950 18750 -880
rect 18670 -960 18750 -950
rect 19010 -880 19090 -870
rect 19010 -950 19020 -880
rect 19080 -950 19090 -880
rect 19010 -960 19090 -950
rect 19350 -880 19430 -870
rect 19350 -950 19360 -880
rect 19420 -950 19430 -880
rect 19350 -960 19430 -950
rect 19690 -880 19770 -870
rect 19690 -950 19700 -880
rect 19760 -950 19770 -880
rect 19690 -960 19770 -950
rect 20030 -880 20110 -870
rect 20030 -950 20040 -880
rect 20100 -950 20110 -880
rect 20030 -960 20110 -950
rect 20370 -880 20450 -870
rect 20370 -950 20380 -880
rect 20440 -950 20450 -880
rect 20370 -960 20450 -950
rect 20710 -880 20790 -870
rect 20710 -950 20720 -880
rect 20780 -950 20790 -880
rect 20710 -960 20790 -950
rect 21050 -880 21130 -870
rect 21050 -950 21060 -880
rect 21120 -950 21130 -880
rect 21050 -960 21130 -950
rect 21390 -880 21470 -870
rect 21390 -950 21400 -880
rect 21460 -950 21470 -880
rect 21390 -960 21470 -950
rect 21730 -880 21810 -870
rect 21730 -950 21740 -880
rect 21800 -950 21810 -880
rect 21730 -960 21810 -950
rect 22070 -880 22150 -870
rect 22070 -950 22080 -880
rect 22140 -950 22150 -880
rect 22070 -960 22150 -950
rect 22410 -880 22490 -870
rect 22410 -950 22420 -880
rect 22480 -950 22490 -880
rect 22410 -960 22490 -950
rect 22750 -880 22830 -870
rect 22750 -950 22760 -880
rect 22820 -950 22830 -880
rect 22750 -960 22830 -950
rect 23090 -880 23170 -870
rect 23090 -950 23100 -880
rect 23160 -950 23170 -880
rect 23090 -960 23170 -950
rect 23430 -880 23510 -870
rect 23430 -950 23440 -880
rect 23500 -950 23510 -880
rect 23430 -960 23510 -950
rect 23770 -880 23850 -870
rect 23770 -950 23780 -880
rect 23840 -950 23850 -880
rect 23770 -960 23850 -950
rect 24110 -880 24190 -870
rect 24110 -950 24120 -880
rect 24180 -950 24190 -880
rect 24110 -960 24190 -950
rect 24450 -880 24530 -870
rect 24450 -950 24460 -880
rect 24520 -950 24530 -880
rect 24450 -960 24530 -950
rect 24790 -880 24870 -870
rect 24790 -950 24800 -880
rect 24860 -950 24870 -880
rect 24790 -960 24870 -950
rect 25130 -880 25210 -870
rect 25130 -950 25140 -880
rect 25200 -950 25210 -880
rect 25130 -960 25210 -950
rect 25470 -880 25550 -870
rect 25470 -950 25480 -880
rect 25540 -950 25550 -880
rect 25470 -960 25550 -950
rect 25810 -880 25890 -870
rect 25810 -950 25820 -880
rect 25880 -950 25890 -880
rect 25810 -960 25890 -950
rect 26150 -880 26230 -870
rect 26150 -950 26160 -880
rect 26220 -950 26230 -880
rect 26150 -960 26230 -950
rect 26490 -880 26570 -870
rect 26490 -950 26500 -880
rect 26560 -950 26570 -880
rect 26490 -960 26570 -950
rect 26830 -880 26910 -870
rect 26830 -950 26840 -880
rect 26900 -950 26910 -880
rect 26830 -960 26910 -950
rect 27170 -880 27250 -870
rect 27170 -950 27180 -880
rect 27240 -950 27250 -880
rect 27170 -960 27250 -950
rect 27510 -880 27590 -870
rect 27510 -950 27520 -880
rect 27580 -950 27590 -880
rect 27510 -960 27590 -950
rect 27850 -880 27930 -870
rect 27850 -950 27860 -880
rect 27920 -950 27930 -880
rect 27850 -960 27930 -950
rect 28190 -880 28270 -870
rect 28190 -950 28200 -880
rect 28260 -950 28270 -880
rect 28190 -960 28270 -950
rect 28530 -880 28610 -870
rect 28530 -950 28540 -880
rect 28600 -950 28610 -880
rect 28530 -960 28610 -950
rect 28870 -880 28950 -870
rect 28870 -950 28880 -880
rect 28940 -950 28950 -880
rect 28870 -960 28950 -950
rect 29210 -880 29290 -870
rect 29210 -950 29220 -880
rect 29280 -950 29290 -880
rect 29210 -960 29290 -950
rect 29550 -880 29630 -870
rect 29550 -950 29560 -880
rect 29620 -950 29630 -880
rect 29550 -960 29630 -950
rect 29890 -880 29970 -870
rect 29890 -950 29900 -880
rect 29960 -950 29970 -880
rect 29890 -960 29970 -950
rect 30230 -880 30310 -870
rect 30230 -950 30240 -880
rect 30300 -950 30310 -880
rect 30230 -960 30310 -950
rect 30570 -880 30650 -870
rect 30570 -950 30580 -880
rect 30640 -950 30650 -880
rect 30570 -960 30650 -950
rect 30910 -880 30990 -870
rect 30910 -950 30920 -880
rect 30980 -950 30990 -880
rect 30910 -960 30990 -950
rect 31250 -880 31330 -870
rect 31250 -950 31260 -880
rect 31320 -950 31330 -880
rect 31250 -960 31330 -950
rect 31590 -880 31670 -870
rect 31590 -950 31600 -880
rect 31660 -950 31670 -880
rect 31590 -960 31670 -950
rect 31930 -880 32010 -870
rect 31930 -950 31940 -880
rect 32000 -950 32010 -880
rect 31930 -960 32010 -950
rect 32270 -880 32350 -870
rect 32270 -950 32280 -880
rect 32340 -950 32350 -880
rect 32270 -960 32350 -950
rect 32610 -880 32690 -870
rect 32610 -950 32620 -880
rect 32680 -950 32690 -880
rect 32610 -960 32690 -950
rect 32950 -880 33030 -870
rect 32950 -950 32960 -880
rect 33020 -950 33030 -880
rect 32950 -960 33030 -950
rect 33290 -880 33370 -870
rect 33290 -950 33300 -880
rect 33360 -950 33370 -880
rect 33290 -960 33370 -950
rect 33630 -880 33710 -870
rect 33630 -950 33640 -880
rect 33700 -950 33710 -880
rect 33630 -960 33710 -950
rect 33970 -880 34050 -870
rect 33970 -950 33980 -880
rect 34040 -950 34050 -880
rect 33970 -960 34050 -950
rect 34310 -880 34390 -870
rect 34310 -950 34320 -880
rect 34380 -950 34390 -880
rect 34310 -960 34390 -950
rect 34650 -880 34730 -870
rect 34650 -950 34660 -880
rect 34720 -950 34730 -880
rect 34650 -960 34730 -950
rect 34990 -880 35070 -870
rect 34990 -950 35000 -880
rect 35060 -950 35070 -880
rect 34990 -960 35070 -950
rect 35330 -880 35410 -870
rect 35330 -950 35340 -880
rect 35400 -950 35410 -880
rect 35330 -960 35410 -950
rect 35670 -880 35750 -870
rect 35670 -950 35680 -880
rect 35740 -950 35750 -880
rect 35670 -960 35750 -950
rect 36010 -880 36090 -870
rect 36010 -950 36020 -880
rect 36080 -950 36090 -880
rect 36010 -960 36090 -950
rect 36350 -880 36430 -870
rect 36350 -950 36360 -880
rect 36420 -950 36430 -880
rect 36350 -960 36430 -950
rect 36690 -880 36770 -870
rect 36690 -950 36700 -880
rect 36760 -950 36770 -880
rect 36690 -960 36770 -950
rect 37030 -880 37110 -870
rect 37030 -950 37040 -880
rect 37100 -950 37110 -880
rect 37030 -960 37110 -950
rect 37370 -880 37450 -870
rect 37370 -950 37380 -880
rect 37440 -950 37450 -880
rect 37370 -960 37450 -950
rect 37710 -880 37790 -870
rect 37710 -950 37720 -880
rect 37780 -950 37790 -880
rect 37710 -960 37790 -950
rect 38050 -880 38130 -870
rect 38050 -950 38060 -880
rect 38120 -950 38130 -880
rect 38050 -960 38130 -950
rect 38390 -880 38470 -870
rect 38390 -950 38400 -880
rect 38460 -950 38470 -880
rect 38390 -960 38470 -950
rect 38730 -880 38810 -870
rect 38730 -950 38740 -880
rect 38800 -950 38810 -880
rect 38730 -960 38810 -950
rect 39070 -880 39150 -870
rect 39070 -950 39080 -880
rect 39140 -950 39150 -880
rect 39070 -960 39150 -950
rect 39410 -880 39490 -870
rect 39410 -950 39420 -880
rect 39480 -950 39490 -880
rect 39410 -960 39490 -950
rect 39750 -880 39830 -870
rect 39750 -950 39760 -880
rect 39820 -950 39830 -880
rect 39750 -960 39830 -950
rect 40090 -880 40170 -870
rect 40090 -950 40100 -880
rect 40160 -950 40170 -880
rect 40090 -960 40170 -950
rect 40430 -880 40510 -870
rect 40430 -950 40440 -880
rect 40500 -950 40510 -880
rect 40430 -960 40510 -950
rect 40770 -880 40850 -870
rect 40770 -950 40780 -880
rect 40840 -950 40850 -880
rect 40770 -960 40850 -950
rect 41110 -880 41190 -870
rect 41110 -950 41120 -880
rect 41180 -950 41190 -880
rect 41110 -960 41190 -950
rect 41450 -880 41530 -870
rect 41450 -950 41460 -880
rect 41520 -950 41530 -880
rect 41450 -960 41530 -950
rect 41790 -880 41870 -870
rect 41790 -950 41800 -880
rect 41860 -950 41870 -880
rect 41790 -960 41870 -950
rect 42130 -880 42210 -870
rect 42130 -950 42140 -880
rect 42200 -950 42210 -880
rect 42130 -960 42210 -950
rect 42470 -880 42550 -870
rect 42470 -950 42480 -880
rect 42540 -950 42550 -880
rect 42470 -960 42550 -950
rect 42810 -880 42890 -870
rect 42810 -950 42820 -880
rect 42880 -950 42890 -880
rect 42810 -960 42890 -950
rect 43150 -880 43230 -870
rect 43150 -950 43160 -880
rect 43220 -950 43230 -880
rect 43150 -960 43230 -950
rect 43490 -880 43570 -870
rect 43490 -950 43500 -880
rect 43560 -950 43570 -880
rect 43490 -960 43570 -950
rect 43830 -880 43910 -870
rect 43830 -950 43840 -880
rect 43900 -950 43910 -880
rect 43830 -960 43910 -950
rect 44170 -880 44250 -870
rect 44170 -950 44180 -880
rect 44240 -950 44250 -880
rect 44170 -960 44250 -950
rect 44510 -880 44590 -870
rect 44510 -950 44520 -880
rect 44580 -950 44590 -880
rect 44510 -960 44590 -950
rect 44850 -880 44930 -870
rect 44850 -950 44860 -880
rect 44920 -950 44930 -880
rect 44850 -960 44930 -950
rect 45190 -880 45270 -870
rect 45190 -950 45200 -880
rect 45260 -950 45270 -880
rect 45190 -960 45270 -950
rect 45530 -880 45610 -870
rect 45530 -950 45540 -880
rect 45600 -950 45610 -880
rect 45530 -960 45610 -950
rect 45870 -880 45950 -870
rect 45870 -950 45880 -880
rect 45940 -950 45950 -880
rect 45870 -960 45950 -950
rect 46210 -880 46290 -870
rect 46210 -950 46220 -880
rect 46280 -950 46290 -880
rect 46210 -960 46290 -950
rect 46550 -880 46630 -870
rect 46550 -950 46560 -880
rect 46620 -950 46630 -880
rect 46550 -960 46630 -950
rect 46890 -880 46970 -870
rect 46890 -950 46900 -880
rect 46960 -950 46970 -880
rect 46890 -960 46970 -950
rect 47230 -880 47310 -870
rect 47230 -950 47240 -880
rect 47300 -950 47310 -880
rect 47230 -960 47310 -950
rect 47570 -880 47650 -870
rect 47570 -950 47580 -880
rect 47640 -950 47650 -880
rect 47570 -960 47650 -950
rect 47910 -880 47990 -870
rect 47910 -950 47920 -880
rect 47980 -950 47990 -880
rect 47910 -960 47990 -950
rect 48250 -880 48330 -870
rect 48250 -950 48260 -880
rect 48320 -950 48330 -880
rect 48250 -960 48330 -950
rect 48590 -880 48670 -870
rect 48590 -950 48600 -880
rect 48660 -950 48670 -880
rect 48590 -960 48670 -950
rect 48930 -880 49010 -870
rect 48930 -950 48940 -880
rect 49000 -950 49010 -880
rect 48930 -960 49010 -950
rect 49270 -880 49350 -870
rect 49270 -950 49280 -880
rect 49340 -950 49350 -880
rect 49270 -960 49350 -950
rect 49610 -880 49690 -870
rect 49610 -950 49620 -880
rect 49680 -950 49690 -880
rect 49610 -960 49690 -950
rect 49950 -880 50030 -870
rect 49950 -950 49960 -880
rect 50020 -950 50030 -880
rect 49950 -960 50030 -950
rect 50290 -880 50370 -870
rect 50290 -950 50300 -880
rect 50360 -950 50370 -880
rect 50290 -960 50370 -950
rect 50630 -880 50710 -870
rect 50630 -950 50640 -880
rect 50700 -950 50710 -880
rect 50630 -960 50710 -950
rect 50970 -880 51050 -870
rect 50970 -950 50980 -880
rect 51040 -950 51050 -880
rect 50970 -960 51050 -950
rect 51310 -880 51390 -870
rect 51310 -950 51320 -880
rect 51380 -950 51390 -880
rect 51310 -960 51390 -950
rect 51650 -880 51730 -870
rect 51650 -950 51660 -880
rect 51720 -950 51730 -880
rect 51650 -960 51730 -950
rect 51990 -880 52070 -870
rect 51990 -950 52000 -880
rect 52060 -950 52070 -880
rect 51990 -960 52070 -950
rect 52330 -880 52410 -870
rect 52330 -950 52340 -880
rect 52400 -950 52410 -880
rect 52330 -960 52410 -950
rect 52670 -880 52750 -870
rect 52670 -950 52680 -880
rect 52740 -950 52750 -880
rect 52670 -960 52750 -950
rect 53010 -880 53090 -870
rect 53010 -950 53020 -880
rect 53080 -950 53090 -880
rect 53010 -960 53090 -950
rect 53350 -880 53430 -870
rect 53350 -950 53360 -880
rect 53420 -950 53430 -880
rect 53350 -960 53430 -950
rect 53690 -880 53770 -870
rect 53690 -950 53700 -880
rect 53760 -950 53770 -880
rect 53690 -960 53770 -950
rect 54030 -880 54110 -870
rect 54030 -950 54040 -880
rect 54100 -950 54110 -880
rect 54030 -960 54110 -950
rect 54370 -880 54450 -870
rect 54370 -950 54380 -880
rect 54440 -950 54450 -880
rect 54370 -960 54450 -950
rect 54710 -880 54790 -870
rect 54710 -950 54720 -880
rect 54780 -950 54790 -880
rect 54710 -960 54790 -950
rect 55050 -880 55130 -870
rect 55050 -950 55060 -880
rect 55120 -950 55130 -880
rect 55050 -960 55130 -950
rect 55390 -880 55470 -870
rect 55390 -950 55400 -880
rect 55460 -950 55470 -880
rect 55390 -960 55470 -950
rect 55730 -880 55810 -870
rect 55730 -950 55740 -880
rect 55800 -950 55810 -880
rect 55730 -960 55810 -950
rect 56070 -880 56150 -870
rect 56070 -950 56080 -880
rect 56140 -950 56150 -880
rect 56070 -960 56150 -950
rect 56410 -880 56490 -870
rect 56410 -950 56420 -880
rect 56480 -950 56490 -880
rect 56410 -960 56490 -950
rect 56750 -880 56830 -870
rect 56750 -950 56760 -880
rect 56820 -950 56830 -880
rect 56750 -960 56830 -950
rect 57090 -880 57170 -870
rect 57090 -950 57100 -880
rect 57160 -950 57170 -880
rect 57090 -960 57170 -950
rect 57430 -880 57510 -870
rect 57430 -950 57440 -880
rect 57500 -950 57510 -880
rect 57430 -960 57510 -950
rect 57770 -880 57850 -870
rect 57770 -950 57780 -880
rect 57840 -950 57850 -880
rect 57770 -960 57850 -950
rect 58110 -880 58190 -870
rect 58110 -950 58120 -880
rect 58180 -950 58190 -880
rect 58110 -960 58190 -950
rect 58450 -880 58530 -870
rect 58450 -950 58460 -880
rect 58520 -950 58530 -880
rect 58450 -960 58530 -950
rect 58790 -880 58870 -870
rect 58790 -950 58800 -880
rect 58860 -950 58870 -880
rect 58790 -960 58870 -950
rect 59130 -880 59210 -870
rect 59130 -950 59140 -880
rect 59200 -950 59210 -880
rect 59130 -960 59210 -950
rect 59470 -880 59550 -870
rect 59470 -950 59480 -880
rect 59540 -950 59550 -880
rect 59470 -960 59550 -950
rect 59810 -880 59890 -870
rect 59810 -950 59820 -880
rect 59880 -950 59890 -880
rect 59810 -960 59890 -950
rect 60150 -880 60230 -870
rect 60150 -950 60160 -880
rect 60220 -950 60230 -880
rect 60150 -960 60230 -950
rect 60490 -880 60570 -870
rect 60490 -950 60500 -880
rect 60560 -950 60570 -880
rect 60490 -960 60570 -950
rect 60830 -880 60910 -870
rect 60830 -950 60840 -880
rect 60900 -950 60910 -880
rect 60830 -960 60910 -950
rect 61170 -880 61250 -870
rect 61170 -950 61180 -880
rect 61240 -950 61250 -880
rect 61170 -960 61250 -950
rect 61510 -880 61590 -870
rect 61510 -950 61520 -880
rect 61580 -950 61590 -880
rect 61510 -960 61590 -950
rect 61850 -880 61930 -870
rect 61850 -950 61860 -880
rect 61920 -950 61930 -880
rect 61850 -960 61930 -950
rect 62190 -880 62270 -870
rect 62190 -950 62200 -880
rect 62260 -950 62270 -880
rect 62190 -960 62270 -950
rect 62530 -880 62610 -870
rect 62530 -950 62540 -880
rect 62600 -950 62610 -880
rect 62530 -960 62610 -950
rect 62870 -880 62950 -870
rect 62870 -950 62880 -880
rect 62940 -950 62950 -880
rect 62870 -960 62950 -950
rect 63210 -880 63290 -870
rect 63210 -950 63220 -880
rect 63280 -950 63290 -880
rect 63210 -960 63290 -950
rect 63550 -880 63630 -870
rect 63550 -950 63560 -880
rect 63620 -950 63630 -880
rect 63550 -960 63630 -950
rect 63890 -880 63970 -870
rect 63890 -950 63900 -880
rect 63960 -950 63970 -880
rect 63890 -960 63970 -950
rect 64230 -880 64310 -870
rect 64230 -950 64240 -880
rect 64300 -950 64310 -880
rect 64230 -960 64310 -950
rect 64570 -880 64650 -870
rect 64570 -950 64580 -880
rect 64640 -950 64650 -880
rect 64570 -960 64650 -950
rect 64910 -880 64990 -870
rect 64910 -950 64920 -880
rect 64980 -950 64990 -880
rect 64910 -960 64990 -950
rect 65250 -880 65330 -870
rect 65250 -950 65260 -880
rect 65320 -950 65330 -880
rect 65250 -960 65330 -950
rect 65590 -880 65670 -870
rect 65590 -950 65600 -880
rect 65660 -950 65670 -880
rect 65590 -960 65670 -950
rect 65930 -880 66010 -870
rect 65930 -950 65940 -880
rect 66000 -950 66010 -880
rect 65930 -960 66010 -950
rect 66270 -880 66350 -870
rect 66270 -950 66280 -880
rect 66340 -950 66350 -880
rect 66270 -960 66350 -950
rect 66610 -880 66690 -870
rect 66610 -950 66620 -880
rect 66680 -950 66690 -880
rect 66610 -960 66690 -950
rect 66950 -880 67030 -870
rect 66950 -950 66960 -880
rect 67020 -950 67030 -880
rect 66950 -960 67030 -950
rect 67290 -880 67370 -870
rect 67290 -950 67300 -880
rect 67360 -950 67370 -880
rect 67290 -960 67370 -950
rect 67630 -880 67710 -870
rect 67630 -950 67640 -880
rect 67700 -950 67710 -880
rect 67630 -960 67710 -950
rect 67970 -880 68050 -870
rect 67970 -950 67980 -880
rect 68040 -950 68050 -880
rect 67970 -960 68050 -950
rect 68310 -880 68390 -870
rect 68310 -950 68320 -880
rect 68380 -950 68390 -880
rect 68310 -960 68390 -950
rect 68650 -880 68730 -870
rect 68650 -950 68660 -880
rect 68720 -950 68730 -880
rect 68650 -960 68730 -950
rect 68990 -880 69070 -870
rect 68990 -950 69000 -880
rect 69060 -950 69070 -880
rect 68990 -960 69070 -950
rect 69330 -880 69410 -870
rect 69330 -950 69340 -880
rect 69400 -950 69410 -880
rect 69330 -960 69410 -950
rect 69670 -880 69750 -870
rect 69670 -950 69680 -880
rect 69740 -950 69750 -880
rect 69670 -960 69750 -950
rect 70010 -880 70090 -870
rect 70010 -950 70020 -880
rect 70080 -950 70090 -880
rect 70010 -960 70090 -950
rect 70350 -880 70430 -870
rect 70350 -950 70360 -880
rect 70420 -950 70430 -880
rect 70350 -960 70430 -950
rect 70690 -880 70770 -870
rect 70690 -950 70700 -880
rect 70760 -950 70770 -880
rect 70690 -960 70770 -950
rect 71030 -880 71110 -870
rect 71030 -950 71040 -880
rect 71100 -950 71110 -880
rect 71030 -960 71110 -950
rect 71370 -880 71450 -870
rect 71370 -950 71380 -880
rect 71440 -950 71450 -880
rect 71370 -960 71450 -950
rect 71710 -880 71790 -870
rect 71710 -950 71720 -880
rect 71780 -950 71790 -880
rect 71710 -960 71790 -950
rect 72050 -880 72130 -870
rect 72050 -950 72060 -880
rect 72120 -950 72130 -880
rect 72050 -960 72130 -950
rect 72390 -880 72470 -870
rect 72390 -950 72400 -880
rect 72460 -950 72470 -880
rect 72390 -960 72470 -950
rect 72730 -880 72810 -870
rect 72730 -950 72740 -880
rect 72800 -950 72810 -880
rect 72730 -960 72810 -950
rect 73070 -880 73150 -870
rect 73070 -950 73080 -880
rect 73140 -950 73150 -880
rect 73070 -960 73150 -950
rect 73410 -880 73490 -870
rect 73410 -950 73420 -880
rect 73480 -950 73490 -880
rect 73410 -960 73490 -950
rect 73750 -880 73830 -870
rect 73750 -950 73760 -880
rect 73820 -950 73830 -880
rect 73750 -960 73830 -950
rect 74090 -880 74170 -870
rect 74090 -950 74100 -880
rect 74160 -950 74170 -880
rect 74090 -960 74170 -950
rect 74430 -880 74510 -870
rect 74430 -950 74440 -880
rect 74500 -950 74510 -880
rect 74430 -960 74510 -950
rect 74770 -880 74850 -870
rect 74770 -950 74780 -880
rect 74840 -950 74850 -880
rect 74770 -960 74850 -950
rect 75110 -880 75190 -870
rect 75110 -950 75120 -880
rect 75180 -950 75190 -880
rect 75110 -960 75190 -950
rect 75450 -880 75530 -870
rect 75450 -950 75460 -880
rect 75520 -950 75530 -880
rect 75450 -960 75530 -950
rect 75790 -880 75870 -870
rect 75790 -950 75800 -880
rect 75860 -950 75870 -880
rect 75790 -960 75870 -950
rect 76130 -880 76210 -870
rect 76130 -950 76140 -880
rect 76200 -950 76210 -880
rect 76130 -960 76210 -950
rect 76470 -880 76550 -870
rect 76470 -950 76480 -880
rect 76540 -950 76550 -880
rect 76470 -960 76550 -950
rect 76810 -880 76890 -870
rect 76810 -950 76820 -880
rect 76880 -950 76890 -880
rect 76810 -960 76890 -950
rect 77150 -880 77230 -870
rect 77150 -950 77160 -880
rect 77220 -950 77230 -880
rect 77150 -960 77230 -950
rect 77490 -880 77570 -870
rect 77490 -950 77500 -880
rect 77560 -950 77570 -880
rect 77490 -960 77570 -950
rect 77830 -880 77910 -870
rect 77830 -950 77840 -880
rect 77900 -950 77910 -880
rect 77830 -960 77910 -950
rect 78170 -880 78250 -870
rect 78170 -950 78180 -880
rect 78240 -950 78250 -880
rect 78170 -960 78250 -950
rect 78510 -880 78590 -870
rect 78510 -950 78520 -880
rect 78580 -950 78590 -880
rect 78510 -960 78590 -950
rect 78850 -880 78930 -870
rect 78850 -950 78860 -880
rect 78920 -950 78930 -880
rect 78850 -960 78930 -950
rect 79190 -880 79270 -870
rect 79190 -950 79200 -880
rect 79260 -950 79270 -880
rect 79190 -960 79270 -950
rect 79530 -880 79610 -870
rect 79530 -950 79540 -880
rect 79600 -950 79610 -880
rect 79530 -960 79610 -950
rect 79870 -880 79950 -870
rect 79870 -950 79880 -880
rect 79940 -950 79950 -880
rect 79870 -960 79950 -950
rect 80210 -880 80290 -870
rect 80210 -950 80220 -880
rect 80280 -950 80290 -880
rect 80210 -960 80290 -950
rect 80550 -880 80630 -870
rect 80550 -950 80560 -880
rect 80620 -950 80630 -880
rect 80550 -960 80630 -950
rect 80890 -880 80970 -870
rect 80890 -950 80900 -880
rect 80960 -950 80970 -880
rect 80890 -960 80970 -950
rect 81230 -880 81310 -870
rect 81230 -950 81240 -880
rect 81300 -950 81310 -880
rect 81230 -960 81310 -950
rect 81570 -880 81650 -870
rect 81570 -950 81580 -880
rect 81640 -950 81650 -880
rect 81570 -960 81650 -950
rect 81910 -880 81990 -870
rect 81910 -950 81920 -880
rect 81980 -950 81990 -880
rect 81910 -960 81990 -950
rect 82250 -880 82330 -870
rect 82250 -950 82260 -880
rect 82320 -950 82330 -880
rect 82250 -960 82330 -950
rect 82590 -880 82670 -870
rect 82590 -950 82600 -880
rect 82660 -950 82670 -880
rect 82590 -960 82670 -950
rect 82930 -880 83010 -870
rect 82930 -950 82940 -880
rect 83000 -950 83010 -880
rect 82930 -960 83010 -950
rect 83270 -880 83350 -870
rect 83270 -950 83280 -880
rect 83340 -950 83350 -880
rect 83270 -960 83350 -950
rect 83610 -880 83690 -870
rect 83610 -950 83620 -880
rect 83680 -950 83690 -880
rect 83610 -960 83690 -950
rect 83950 -880 84030 -870
rect 83950 -950 83960 -880
rect 84020 -950 84030 -880
rect 83950 -960 84030 -950
rect 84290 -880 84370 -870
rect 84290 -950 84300 -880
rect 84360 -950 84370 -880
rect 84290 -960 84370 -950
rect 84630 -880 84710 -870
rect 84630 -950 84640 -880
rect 84700 -950 84710 -880
rect 84630 -960 84710 -950
rect 84970 -880 85050 -870
rect 84970 -950 84980 -880
rect 85040 -950 85050 -880
rect 84970 -960 85050 -950
rect 85310 -880 85390 -870
rect 85310 -950 85320 -880
rect 85380 -950 85390 -880
rect 85310 -960 85390 -950
rect 85650 -880 85730 -870
rect 85650 -950 85660 -880
rect 85720 -950 85730 -880
rect 85650 -960 85730 -950
rect 85990 -880 86070 -870
rect 85990 -950 86000 -880
rect 86060 -950 86070 -880
rect 85990 -960 86070 -950
rect 86330 -880 86410 -870
rect 86330 -950 86340 -880
rect 86400 -950 86410 -880
rect 86330 -960 86410 -950
rect 86670 -880 86750 -870
rect 86670 -950 86680 -880
rect 86740 -950 86750 -880
rect 86670 -960 86750 -950
rect 87010 -880 87090 -870
rect 87010 -950 87020 -880
rect 87080 -950 87090 -880
rect 87010 -960 87090 -950
rect 130 -1100 230 -1080
rect 470 -1100 570 -1080
rect 810 -1100 910 -1080
rect 1150 -1100 1250 -1080
rect 1490 -1100 1590 -1080
rect 1830 -1100 1930 -1080
rect 2170 -1100 2270 -1080
rect 2510 -1100 2610 -1080
rect 2850 -1100 2950 -1080
rect 3190 -1100 3290 -1080
rect 3530 -1100 3630 -1080
rect 3870 -1100 3970 -1080
rect 4210 -1100 4310 -1080
rect 4550 -1100 4650 -1080
rect 4890 -1100 4990 -1080
rect 5230 -1100 5330 -1080
rect 5570 -1100 5670 -1080
rect 5910 -1100 6010 -1080
rect 6250 -1100 6350 -1080
rect 6590 -1100 6690 -1080
rect 6930 -1100 7030 -1080
rect 7270 -1100 7370 -1080
rect 7610 -1100 7710 -1080
rect 7950 -1100 8050 -1080
rect 8290 -1100 8390 -1080
rect 8630 -1100 8730 -1080
rect 8970 -1100 9070 -1080
rect 9310 -1100 9410 -1080
rect 9650 -1100 9750 -1080
rect 9990 -1100 10090 -1080
rect 10330 -1100 10430 -1080
rect 10670 -1100 10770 -1080
rect 11010 -1100 11110 -1080
rect 11350 -1100 11450 -1080
rect 11690 -1100 11790 -1080
rect 12030 -1100 12130 -1080
rect 12370 -1100 12470 -1080
rect 12710 -1100 12810 -1080
rect 13050 -1100 13150 -1080
rect 13390 -1100 13490 -1080
rect 13730 -1100 13830 -1080
rect 14070 -1100 14170 -1080
rect 14410 -1100 14510 -1080
rect 14750 -1100 14850 -1080
rect 15090 -1100 15190 -1080
rect 15430 -1100 15530 -1080
rect 15770 -1100 15870 -1080
rect 16110 -1100 16210 -1080
rect 16450 -1100 16550 -1080
rect 16790 -1100 16890 -1080
rect 17130 -1100 17230 -1080
rect 17470 -1100 17570 -1080
rect 17810 -1100 17910 -1080
rect 18150 -1100 18250 -1080
rect 18490 -1100 18590 -1080
rect 18830 -1100 18930 -1080
rect 19170 -1100 19270 -1080
rect 19510 -1100 19610 -1080
rect 19850 -1100 19950 -1080
rect 20190 -1100 20290 -1080
rect 20530 -1100 20630 -1080
rect 20870 -1100 20970 -1080
rect 21210 -1100 21310 -1080
rect 21550 -1100 21650 -1080
rect 21890 -1100 21990 -1080
rect 22230 -1100 22330 -1080
rect 22570 -1100 22670 -1080
rect 22910 -1100 23010 -1080
rect 23250 -1100 23350 -1080
rect 23590 -1100 23690 -1080
rect 23930 -1100 24030 -1080
rect 24270 -1100 24370 -1080
rect 24610 -1100 24710 -1080
rect 24950 -1100 25050 -1080
rect 25290 -1100 25390 -1080
rect 25630 -1100 25730 -1080
rect 25970 -1100 26070 -1080
rect 26310 -1100 26410 -1080
rect 26650 -1100 26750 -1080
rect 26990 -1100 27090 -1080
rect 27330 -1100 27430 -1080
rect 27670 -1100 27770 -1080
rect 28010 -1100 28110 -1080
rect 28350 -1100 28450 -1080
rect 28690 -1100 28790 -1080
rect 29030 -1100 29130 -1080
rect 29370 -1100 29470 -1080
rect 29710 -1100 29810 -1080
rect 30050 -1100 30150 -1080
rect 30390 -1100 30490 -1080
rect 30730 -1100 30830 -1080
rect 31070 -1100 31170 -1080
rect 31410 -1100 31510 -1080
rect 31750 -1100 31850 -1080
rect 32090 -1100 32190 -1080
rect 32430 -1100 32530 -1080
rect 32770 -1100 32870 -1080
rect 33110 -1100 33210 -1080
rect 33450 -1100 33550 -1080
rect 33790 -1100 33890 -1080
rect 34130 -1100 34230 -1080
rect 34470 -1100 34570 -1080
rect 34810 -1100 34910 -1080
rect 35150 -1100 35250 -1080
rect 35490 -1100 35590 -1080
rect 35830 -1100 35930 -1080
rect 36170 -1100 36270 -1080
rect 36510 -1100 36610 -1080
rect 36850 -1100 36950 -1080
rect 37190 -1100 37290 -1080
rect 37530 -1100 37630 -1080
rect 37870 -1100 37970 -1080
rect 38210 -1100 38310 -1080
rect 38550 -1100 38650 -1080
rect 38890 -1100 38990 -1080
rect 39230 -1100 39330 -1080
rect 39570 -1100 39670 -1080
rect 39910 -1100 40010 -1080
rect 40250 -1100 40350 -1080
rect 40590 -1100 40690 -1080
rect 40930 -1100 41030 -1080
rect 41270 -1100 41370 -1080
rect 41610 -1100 41710 -1080
rect 41950 -1100 42050 -1080
rect 42290 -1100 42390 -1080
rect 42630 -1100 42730 -1080
rect 42970 -1100 43070 -1080
rect 43310 -1100 43410 -1080
rect 43650 -1100 43750 -1080
rect 43990 -1100 44090 -1080
rect 44330 -1100 44430 -1080
rect 44670 -1100 44770 -1080
rect 45010 -1100 45110 -1080
rect 45350 -1100 45450 -1080
rect 45690 -1100 45790 -1080
rect 46030 -1100 46130 -1080
rect 46370 -1100 46470 -1080
rect 46710 -1100 46810 -1080
rect 47050 -1100 47150 -1080
rect 47390 -1100 47490 -1080
rect 47730 -1100 47830 -1080
rect 48070 -1100 48170 -1080
rect 48410 -1100 48510 -1080
rect 48750 -1100 48850 -1080
rect 49090 -1100 49190 -1080
rect 49430 -1100 49530 -1080
rect 49770 -1100 49870 -1080
rect 50110 -1100 50210 -1080
rect 50450 -1100 50550 -1080
rect 50790 -1100 50890 -1080
rect 51130 -1100 51230 -1080
rect 51470 -1100 51570 -1080
rect 51810 -1100 51910 -1080
rect 52150 -1100 52250 -1080
rect 52490 -1100 52590 -1080
rect 52830 -1100 52930 -1080
rect 53170 -1100 53270 -1080
rect 53510 -1100 53610 -1080
rect 53850 -1100 53950 -1080
rect 54190 -1100 54290 -1080
rect 54530 -1100 54630 -1080
rect 54870 -1100 54970 -1080
rect 55210 -1100 55310 -1080
rect 55550 -1100 55650 -1080
rect 55890 -1100 55990 -1080
rect 56230 -1100 56330 -1080
rect 56570 -1100 56670 -1080
rect 56910 -1100 57010 -1080
rect 57250 -1100 57350 -1080
rect 57590 -1100 57690 -1080
rect 57930 -1100 58030 -1080
rect 58270 -1100 58370 -1080
rect 58610 -1100 58710 -1080
rect 58950 -1100 59050 -1080
rect 59290 -1100 59390 -1080
rect 59630 -1100 59730 -1080
rect 59970 -1100 60070 -1080
rect 60310 -1100 60410 -1080
rect 60650 -1100 60750 -1080
rect 60990 -1100 61090 -1080
rect 61330 -1100 61430 -1080
rect 61670 -1100 61770 -1080
rect 62010 -1100 62110 -1080
rect 62350 -1100 62450 -1080
rect 62690 -1100 62790 -1080
rect 63030 -1100 63130 -1080
rect 63370 -1100 63470 -1080
rect 63710 -1100 63810 -1080
rect 64050 -1100 64150 -1080
rect 64390 -1100 64490 -1080
rect 64730 -1100 64830 -1080
rect 65070 -1100 65170 -1080
rect 65410 -1100 65510 -1080
rect 65750 -1100 65850 -1080
rect 66090 -1100 66190 -1080
rect 66430 -1100 66530 -1080
rect 66770 -1100 66870 -1080
rect 67110 -1100 67210 -1080
rect 67450 -1100 67550 -1080
rect 67790 -1100 67890 -1080
rect 68130 -1100 68230 -1080
rect 68470 -1100 68570 -1080
rect 68810 -1100 68910 -1080
rect 69150 -1100 69250 -1080
rect 69490 -1100 69590 -1080
rect 69830 -1100 69930 -1080
rect 70170 -1100 70270 -1080
rect 70510 -1100 70610 -1080
rect 70850 -1100 70950 -1080
rect 71190 -1100 71290 -1080
rect 71530 -1100 71630 -1080
rect 71870 -1100 71970 -1080
rect 72210 -1100 72310 -1080
rect 72550 -1100 72650 -1080
rect 72890 -1100 72990 -1080
rect 73230 -1100 73330 -1080
rect 73570 -1100 73670 -1080
rect 73910 -1100 74010 -1080
rect 74250 -1100 74350 -1080
rect 74590 -1100 74690 -1080
rect 74930 -1100 75030 -1080
rect 75270 -1100 75370 -1080
rect 75610 -1100 75710 -1080
rect 75950 -1100 76050 -1080
rect 76290 -1100 76390 -1080
rect 76630 -1100 76730 -1080
rect 76970 -1100 77070 -1080
rect 77310 -1100 77410 -1080
rect 77650 -1100 77750 -1080
rect 77990 -1100 78090 -1080
rect 78330 -1100 78430 -1080
rect 78670 -1100 78770 -1080
rect 79010 -1100 79110 -1080
rect 79350 -1100 79450 -1080
rect 79690 -1100 79790 -1080
rect 80030 -1100 80130 -1080
rect 80370 -1100 80470 -1080
rect 80710 -1100 80810 -1080
rect 81050 -1100 81150 -1080
rect 81390 -1100 81490 -1080
rect 81730 -1100 81830 -1080
rect 82070 -1100 82170 -1080
rect 82410 -1100 82510 -1080
rect 82750 -1100 82850 -1080
rect 83090 -1100 83190 -1080
rect 83430 -1100 83530 -1080
rect 83770 -1100 83870 -1080
rect 84110 -1100 84210 -1080
rect 84450 -1100 84550 -1080
rect 84790 -1100 84890 -1080
rect 85130 -1100 85230 -1080
rect 85470 -1100 85570 -1080
rect 85810 -1100 85910 -1080
rect 86150 -1100 86250 -1080
rect 86490 -1100 86590 -1080
rect 86830 -1100 86930 -1080
rect 87170 -1100 87270 -1080
rect 110 -1160 150 -1100
rect 210 -1160 490 -1100
rect 550 -1160 830 -1100
rect 890 -1160 1170 -1100
rect 1230 -1160 1510 -1100
rect 1570 -1160 1850 -1100
rect 1910 -1160 2190 -1100
rect 2250 -1160 2530 -1100
rect 2590 -1160 2870 -1100
rect 2930 -1160 3210 -1100
rect 3270 -1160 3550 -1100
rect 3610 -1160 3890 -1100
rect 3950 -1160 4230 -1100
rect 4290 -1160 4570 -1100
rect 4630 -1160 4910 -1100
rect 4970 -1160 5250 -1100
rect 5310 -1160 5590 -1100
rect 5650 -1160 5930 -1100
rect 5990 -1160 6270 -1100
rect 6330 -1160 6610 -1100
rect 6670 -1160 6950 -1100
rect 7010 -1160 7290 -1100
rect 7350 -1160 7630 -1100
rect 7690 -1160 7970 -1100
rect 8030 -1160 8310 -1100
rect 8370 -1160 8650 -1100
rect 8710 -1160 8990 -1100
rect 9050 -1160 9330 -1100
rect 9390 -1160 9670 -1100
rect 9730 -1160 10010 -1100
rect 10070 -1160 10350 -1100
rect 10410 -1160 10690 -1100
rect 10750 -1160 11030 -1100
rect 11090 -1160 11370 -1100
rect 11430 -1160 11710 -1100
rect 11770 -1160 12050 -1100
rect 12110 -1160 12390 -1100
rect 12450 -1160 12730 -1100
rect 12790 -1160 13070 -1100
rect 13130 -1160 13410 -1100
rect 13470 -1160 13750 -1100
rect 13810 -1160 14090 -1100
rect 14150 -1160 14430 -1100
rect 14490 -1160 14770 -1100
rect 14830 -1160 15110 -1100
rect 15170 -1160 15450 -1100
rect 15510 -1160 15790 -1100
rect 15850 -1160 16130 -1100
rect 16190 -1160 16470 -1100
rect 16530 -1160 16810 -1100
rect 16870 -1160 17150 -1100
rect 17210 -1160 17490 -1100
rect 17550 -1160 17830 -1100
rect 17890 -1160 18170 -1100
rect 18230 -1160 18510 -1100
rect 18570 -1160 18850 -1100
rect 18910 -1160 19190 -1100
rect 19250 -1160 19530 -1100
rect 19590 -1160 19870 -1100
rect 19930 -1160 20210 -1100
rect 20270 -1160 20550 -1100
rect 20610 -1160 20890 -1100
rect 20950 -1160 21230 -1100
rect 21290 -1160 21570 -1100
rect 21630 -1160 21910 -1100
rect 21970 -1160 22250 -1100
rect 22310 -1160 22590 -1100
rect 22650 -1160 22930 -1100
rect 22990 -1160 23270 -1100
rect 23330 -1160 23610 -1100
rect 23670 -1160 23950 -1100
rect 24010 -1160 24290 -1100
rect 24350 -1160 24630 -1100
rect 24690 -1160 24970 -1100
rect 25030 -1160 25310 -1100
rect 25370 -1160 25650 -1100
rect 25710 -1160 25990 -1100
rect 26050 -1160 26330 -1100
rect 26390 -1160 26670 -1100
rect 26730 -1160 27010 -1100
rect 27070 -1160 27350 -1100
rect 27410 -1160 27690 -1100
rect 27750 -1160 28030 -1100
rect 28090 -1160 28370 -1100
rect 28430 -1160 28710 -1100
rect 28770 -1160 29050 -1100
rect 29110 -1160 29390 -1100
rect 29450 -1160 29730 -1100
rect 29790 -1160 30070 -1100
rect 30130 -1160 30410 -1100
rect 30470 -1160 30750 -1100
rect 30810 -1160 31090 -1100
rect 31150 -1160 31430 -1100
rect 31490 -1160 31770 -1100
rect 31830 -1160 32110 -1100
rect 32170 -1160 32450 -1100
rect 32510 -1160 32790 -1100
rect 32850 -1160 33130 -1100
rect 33190 -1160 33470 -1100
rect 33530 -1160 33810 -1100
rect 33870 -1160 34150 -1100
rect 34210 -1160 34490 -1100
rect 34550 -1160 34830 -1100
rect 34890 -1160 35170 -1100
rect 35230 -1160 35510 -1100
rect 35570 -1160 35850 -1100
rect 35910 -1160 36190 -1100
rect 36250 -1160 36530 -1100
rect 36590 -1160 36870 -1100
rect 36930 -1160 37210 -1100
rect 37270 -1160 37550 -1100
rect 37610 -1160 37890 -1100
rect 37950 -1160 38230 -1100
rect 38290 -1160 38570 -1100
rect 38630 -1160 38910 -1100
rect 38970 -1160 39250 -1100
rect 39310 -1160 39590 -1100
rect 39650 -1160 39930 -1100
rect 39990 -1160 40270 -1100
rect 40330 -1160 40610 -1100
rect 40670 -1160 40950 -1100
rect 41010 -1160 41290 -1100
rect 41350 -1160 41630 -1100
rect 41690 -1160 41970 -1100
rect 42030 -1160 42310 -1100
rect 42370 -1160 42650 -1100
rect 42710 -1160 42990 -1100
rect 43050 -1160 43330 -1100
rect 43390 -1160 43670 -1100
rect 43730 -1160 44010 -1100
rect 44070 -1160 44350 -1100
rect 44410 -1160 44690 -1100
rect 44750 -1160 45030 -1100
rect 45090 -1160 45370 -1100
rect 45430 -1160 45710 -1100
rect 45770 -1160 46050 -1100
rect 46110 -1160 46390 -1100
rect 46450 -1160 46730 -1100
rect 46790 -1160 47070 -1100
rect 47130 -1160 47410 -1100
rect 47470 -1160 47750 -1100
rect 47810 -1160 48090 -1100
rect 48150 -1160 48430 -1100
rect 48490 -1160 48770 -1100
rect 48830 -1160 49110 -1100
rect 49170 -1160 49450 -1100
rect 49510 -1160 49790 -1100
rect 49850 -1160 50130 -1100
rect 50190 -1160 50470 -1100
rect 50530 -1160 50810 -1100
rect 50870 -1160 51150 -1100
rect 51210 -1160 51490 -1100
rect 51550 -1160 51830 -1100
rect 51890 -1160 52170 -1100
rect 52230 -1160 52510 -1100
rect 52570 -1160 52850 -1100
rect 52910 -1160 53190 -1100
rect 53250 -1160 53530 -1100
rect 53590 -1160 53870 -1100
rect 53930 -1160 54210 -1100
rect 54270 -1160 54550 -1100
rect 54610 -1160 54890 -1100
rect 54950 -1160 55230 -1100
rect 55290 -1160 55570 -1100
rect 55630 -1160 55910 -1100
rect 55970 -1160 56250 -1100
rect 56310 -1160 56590 -1100
rect 56650 -1160 56930 -1100
rect 56990 -1160 57270 -1100
rect 57330 -1160 57610 -1100
rect 57670 -1160 57950 -1100
rect 58010 -1160 58290 -1100
rect 58350 -1160 58630 -1100
rect 58690 -1160 58970 -1100
rect 59030 -1160 59310 -1100
rect 59370 -1160 59650 -1100
rect 59710 -1160 59990 -1100
rect 60050 -1160 60330 -1100
rect 60390 -1160 60670 -1100
rect 60730 -1160 61010 -1100
rect 61070 -1160 61350 -1100
rect 61410 -1160 61690 -1100
rect 61750 -1160 62030 -1100
rect 62090 -1160 62370 -1100
rect 62430 -1160 62710 -1100
rect 62770 -1160 63050 -1100
rect 63110 -1160 63390 -1100
rect 63450 -1160 63730 -1100
rect 63790 -1160 64070 -1100
rect 64130 -1160 64410 -1100
rect 64470 -1160 64750 -1100
rect 64810 -1160 65090 -1100
rect 65150 -1160 65430 -1100
rect 65490 -1160 65770 -1100
rect 65830 -1160 66110 -1100
rect 66170 -1160 66450 -1100
rect 66510 -1160 66790 -1100
rect 66850 -1160 67130 -1100
rect 67190 -1160 67470 -1100
rect 67530 -1160 67810 -1100
rect 67870 -1160 68150 -1100
rect 68210 -1160 68490 -1100
rect 68550 -1160 68830 -1100
rect 68890 -1160 69170 -1100
rect 69230 -1160 69510 -1100
rect 69570 -1160 69850 -1100
rect 69910 -1160 70190 -1100
rect 70250 -1160 70530 -1100
rect 70590 -1160 70870 -1100
rect 70930 -1160 71210 -1100
rect 71270 -1160 71550 -1100
rect 71610 -1160 71890 -1100
rect 71950 -1160 72230 -1100
rect 72290 -1160 72570 -1100
rect 72630 -1160 72910 -1100
rect 72970 -1160 73250 -1100
rect 73310 -1160 73590 -1100
rect 73650 -1160 73930 -1100
rect 73990 -1160 74270 -1100
rect 74330 -1160 74610 -1100
rect 74670 -1160 74950 -1100
rect 75010 -1160 75290 -1100
rect 75350 -1160 75630 -1100
rect 75690 -1160 75970 -1100
rect 76030 -1160 76310 -1100
rect 76370 -1160 76650 -1100
rect 76710 -1160 76990 -1100
rect 77050 -1160 77330 -1100
rect 77390 -1160 77670 -1100
rect 77730 -1160 78010 -1100
rect 78070 -1160 78350 -1100
rect 78410 -1160 78690 -1100
rect 78750 -1160 79030 -1100
rect 79090 -1160 79370 -1100
rect 79430 -1160 79710 -1100
rect 79770 -1160 80050 -1100
rect 80110 -1160 80390 -1100
rect 80450 -1160 80730 -1100
rect 80790 -1160 81070 -1100
rect 81130 -1160 81410 -1100
rect 81470 -1160 81750 -1100
rect 81810 -1160 82090 -1100
rect 82150 -1160 82430 -1100
rect 82490 -1160 82770 -1100
rect 82830 -1160 83110 -1100
rect 83170 -1160 83450 -1100
rect 83510 -1160 83790 -1100
rect 83850 -1160 84130 -1100
rect 84190 -1160 84470 -1100
rect 84530 -1160 84810 -1100
rect 84870 -1160 85150 -1100
rect 85210 -1160 85490 -1100
rect 85550 -1160 85830 -1100
rect 85890 -1160 86170 -1100
rect 86230 -1160 86510 -1100
rect 86570 -1160 86850 -1100
rect 86910 -1160 87190 -1100
rect 87250 -1160 87270 -1100
rect 130 -1180 230 -1160
rect 470 -1180 570 -1160
rect 810 -1180 910 -1160
rect 1150 -1180 1250 -1160
rect 1490 -1180 1590 -1160
rect 1830 -1180 1930 -1160
rect 2170 -1180 2270 -1160
rect 2510 -1180 2610 -1160
rect 2850 -1180 2950 -1160
rect 3190 -1180 3290 -1160
rect 3530 -1180 3630 -1160
rect 3870 -1180 3970 -1160
rect 4210 -1180 4310 -1160
rect 4550 -1180 4650 -1160
rect 4890 -1180 4990 -1160
rect 5230 -1180 5330 -1160
rect 5570 -1180 5670 -1160
rect 5910 -1180 6010 -1160
rect 6250 -1180 6350 -1160
rect 6590 -1180 6690 -1160
rect 6930 -1180 7030 -1160
rect 7270 -1180 7370 -1160
rect 7610 -1180 7710 -1160
rect 7950 -1180 8050 -1160
rect 8290 -1180 8390 -1160
rect 8630 -1180 8730 -1160
rect 8970 -1180 9070 -1160
rect 9310 -1180 9410 -1160
rect 9650 -1180 9750 -1160
rect 9990 -1180 10090 -1160
rect 10330 -1180 10430 -1160
rect 10670 -1180 10770 -1160
rect 11010 -1180 11110 -1160
rect 11350 -1180 11450 -1160
rect 11690 -1180 11790 -1160
rect 12030 -1180 12130 -1160
rect 12370 -1180 12470 -1160
rect 12710 -1180 12810 -1160
rect 13050 -1180 13150 -1160
rect 13390 -1180 13490 -1160
rect 13730 -1180 13830 -1160
rect 14070 -1180 14170 -1160
rect 14410 -1180 14510 -1160
rect 14750 -1180 14850 -1160
rect 15090 -1180 15190 -1160
rect 15430 -1180 15530 -1160
rect 15770 -1180 15870 -1160
rect 16110 -1180 16210 -1160
rect 16450 -1180 16550 -1160
rect 16790 -1180 16890 -1160
rect 17130 -1180 17230 -1160
rect 17470 -1180 17570 -1160
rect 17810 -1180 17910 -1160
rect 18150 -1180 18250 -1160
rect 18490 -1180 18590 -1160
rect 18830 -1180 18930 -1160
rect 19170 -1180 19270 -1160
rect 19510 -1180 19610 -1160
rect 19850 -1180 19950 -1160
rect 20190 -1180 20290 -1160
rect 20530 -1180 20630 -1160
rect 20870 -1180 20970 -1160
rect 21210 -1180 21310 -1160
rect 21550 -1180 21650 -1160
rect 21890 -1180 21990 -1160
rect 22230 -1180 22330 -1160
rect 22570 -1180 22670 -1160
rect 22910 -1180 23010 -1160
rect 23250 -1180 23350 -1160
rect 23590 -1180 23690 -1160
rect 23930 -1180 24030 -1160
rect 24270 -1180 24370 -1160
rect 24610 -1180 24710 -1160
rect 24950 -1180 25050 -1160
rect 25290 -1180 25390 -1160
rect 25630 -1180 25730 -1160
rect 25970 -1180 26070 -1160
rect 26310 -1180 26410 -1160
rect 26650 -1180 26750 -1160
rect 26990 -1180 27090 -1160
rect 27330 -1180 27430 -1160
rect 27670 -1180 27770 -1160
rect 28010 -1180 28110 -1160
rect 28350 -1180 28450 -1160
rect 28690 -1180 28790 -1160
rect 29030 -1180 29130 -1160
rect 29370 -1180 29470 -1160
rect 29710 -1180 29810 -1160
rect 30050 -1180 30150 -1160
rect 30390 -1180 30490 -1160
rect 30730 -1180 30830 -1160
rect 31070 -1180 31170 -1160
rect 31410 -1180 31510 -1160
rect 31750 -1180 31850 -1160
rect 32090 -1180 32190 -1160
rect 32430 -1180 32530 -1160
rect 32770 -1180 32870 -1160
rect 33110 -1180 33210 -1160
rect 33450 -1180 33550 -1160
rect 33790 -1180 33890 -1160
rect 34130 -1180 34230 -1160
rect 34470 -1180 34570 -1160
rect 34810 -1180 34910 -1160
rect 35150 -1180 35250 -1160
rect 35490 -1180 35590 -1160
rect 35830 -1180 35930 -1160
rect 36170 -1180 36270 -1160
rect 36510 -1180 36610 -1160
rect 36850 -1180 36950 -1160
rect 37190 -1180 37290 -1160
rect 37530 -1180 37630 -1160
rect 37870 -1180 37970 -1160
rect 38210 -1180 38310 -1160
rect 38550 -1180 38650 -1160
rect 38890 -1180 38990 -1160
rect 39230 -1180 39330 -1160
rect 39570 -1180 39670 -1160
rect 39910 -1180 40010 -1160
rect 40250 -1180 40350 -1160
rect 40590 -1180 40690 -1160
rect 40930 -1180 41030 -1160
rect 41270 -1180 41370 -1160
rect 41610 -1180 41710 -1160
rect 41950 -1180 42050 -1160
rect 42290 -1180 42390 -1160
rect 42630 -1180 42730 -1160
rect 42970 -1180 43070 -1160
rect 43310 -1180 43410 -1160
rect 43650 -1180 43750 -1160
rect 43990 -1180 44090 -1160
rect 44330 -1180 44430 -1160
rect 44670 -1180 44770 -1160
rect 45010 -1180 45110 -1160
rect 45350 -1180 45450 -1160
rect 45690 -1180 45790 -1160
rect 46030 -1180 46130 -1160
rect 46370 -1180 46470 -1160
rect 46710 -1180 46810 -1160
rect 47050 -1180 47150 -1160
rect 47390 -1180 47490 -1160
rect 47730 -1180 47830 -1160
rect 48070 -1180 48170 -1160
rect 48410 -1180 48510 -1160
rect 48750 -1180 48850 -1160
rect 49090 -1180 49190 -1160
rect 49430 -1180 49530 -1160
rect 49770 -1180 49870 -1160
rect 50110 -1180 50210 -1160
rect 50450 -1180 50550 -1160
rect 50790 -1180 50890 -1160
rect 51130 -1180 51230 -1160
rect 51470 -1180 51570 -1160
rect 51810 -1180 51910 -1160
rect 52150 -1180 52250 -1160
rect 52490 -1180 52590 -1160
rect 52830 -1180 52930 -1160
rect 53170 -1180 53270 -1160
rect 53510 -1180 53610 -1160
rect 53850 -1180 53950 -1160
rect 54190 -1180 54290 -1160
rect 54530 -1180 54630 -1160
rect 54870 -1180 54970 -1160
rect 55210 -1180 55310 -1160
rect 55550 -1180 55650 -1160
rect 55890 -1180 55990 -1160
rect 56230 -1180 56330 -1160
rect 56570 -1180 56670 -1160
rect 56910 -1180 57010 -1160
rect 57250 -1180 57350 -1160
rect 57590 -1180 57690 -1160
rect 57930 -1180 58030 -1160
rect 58270 -1180 58370 -1160
rect 58610 -1180 58710 -1160
rect 58950 -1180 59050 -1160
rect 59290 -1180 59390 -1160
rect 59630 -1180 59730 -1160
rect 59970 -1180 60070 -1160
rect 60310 -1180 60410 -1160
rect 60650 -1180 60750 -1160
rect 60990 -1180 61090 -1160
rect 61330 -1180 61430 -1160
rect 61670 -1180 61770 -1160
rect 62010 -1180 62110 -1160
rect 62350 -1180 62450 -1160
rect 62690 -1180 62790 -1160
rect 63030 -1180 63130 -1160
rect 63370 -1180 63470 -1160
rect 63710 -1180 63810 -1160
rect 64050 -1180 64150 -1160
rect 64390 -1180 64490 -1160
rect 64730 -1180 64830 -1160
rect 65070 -1180 65170 -1160
rect 65410 -1180 65510 -1160
rect 65750 -1180 65850 -1160
rect 66090 -1180 66190 -1160
rect 66430 -1180 66530 -1160
rect 66770 -1180 66870 -1160
rect 67110 -1180 67210 -1160
rect 67450 -1180 67550 -1160
rect 67790 -1180 67890 -1160
rect 68130 -1180 68230 -1160
rect 68470 -1180 68570 -1160
rect 68810 -1180 68910 -1160
rect 69150 -1180 69250 -1160
rect 69490 -1180 69590 -1160
rect 69830 -1180 69930 -1160
rect 70170 -1180 70270 -1160
rect 70510 -1180 70610 -1160
rect 70850 -1180 70950 -1160
rect 71190 -1180 71290 -1160
rect 71530 -1180 71630 -1160
rect 71870 -1180 71970 -1160
rect 72210 -1180 72310 -1160
rect 72550 -1180 72650 -1160
rect 72890 -1180 72990 -1160
rect 73230 -1180 73330 -1160
rect 73570 -1180 73670 -1160
rect 73910 -1180 74010 -1160
rect 74250 -1180 74350 -1160
rect 74590 -1180 74690 -1160
rect 74930 -1180 75030 -1160
rect 75270 -1180 75370 -1160
rect 75610 -1180 75710 -1160
rect 75950 -1180 76050 -1160
rect 76290 -1180 76390 -1160
rect 76630 -1180 76730 -1160
rect 76970 -1180 77070 -1160
rect 77310 -1180 77410 -1160
rect 77650 -1180 77750 -1160
rect 77990 -1180 78090 -1160
rect 78330 -1180 78430 -1160
rect 78670 -1180 78770 -1160
rect 79010 -1180 79110 -1160
rect 79350 -1180 79450 -1160
rect 79690 -1180 79790 -1160
rect 80030 -1180 80130 -1160
rect 80370 -1180 80470 -1160
rect 80710 -1180 80810 -1160
rect 81050 -1180 81150 -1160
rect 81390 -1180 81490 -1160
rect 81730 -1180 81830 -1160
rect 82070 -1180 82170 -1160
rect 82410 -1180 82510 -1160
rect 82750 -1180 82850 -1160
rect 83090 -1180 83190 -1160
rect 83430 -1180 83530 -1160
rect 83770 -1180 83870 -1160
rect 84110 -1180 84210 -1160
rect 84450 -1180 84550 -1160
rect 84790 -1180 84890 -1160
rect 85130 -1180 85230 -1160
rect 85470 -1180 85570 -1160
rect 85810 -1180 85910 -1160
rect 86150 -1180 86250 -1160
rect 86490 -1180 86590 -1160
rect 86830 -1180 86930 -1160
rect 87170 -1180 87270 -1160
rect 130 -1300 230 -1280
rect 470 -1300 570 -1280
rect 810 -1300 910 -1280
rect 1150 -1300 1250 -1280
rect 1490 -1300 1590 -1280
rect 1830 -1300 1930 -1280
rect 2170 -1300 2270 -1280
rect 2510 -1300 2610 -1280
rect 2850 -1300 2950 -1280
rect 3190 -1300 3290 -1280
rect 3530 -1300 3630 -1280
rect 3870 -1300 3970 -1280
rect 4210 -1300 4310 -1280
rect 4550 -1300 4650 -1280
rect 4890 -1300 4990 -1280
rect 5230 -1300 5330 -1280
rect 5570 -1300 5670 -1280
rect 5910 -1300 6010 -1280
rect 6250 -1300 6350 -1280
rect 6590 -1300 6690 -1280
rect 6930 -1300 7030 -1280
rect 7270 -1300 7370 -1280
rect 7610 -1300 7710 -1280
rect 7950 -1300 8050 -1280
rect 8290 -1300 8390 -1280
rect 8630 -1300 8730 -1280
rect 8970 -1300 9070 -1280
rect 9310 -1300 9410 -1280
rect 9650 -1300 9750 -1280
rect 9990 -1300 10090 -1280
rect 10330 -1300 10430 -1280
rect 10670 -1300 10770 -1280
rect 11010 -1300 11110 -1280
rect 11350 -1300 11450 -1280
rect 11690 -1300 11790 -1280
rect 12030 -1300 12130 -1280
rect 12370 -1300 12470 -1280
rect 12710 -1300 12810 -1280
rect 13050 -1300 13150 -1280
rect 13390 -1300 13490 -1280
rect 13730 -1300 13830 -1280
rect 14070 -1300 14170 -1280
rect 14410 -1300 14510 -1280
rect 14750 -1300 14850 -1280
rect 15090 -1300 15190 -1280
rect 15430 -1300 15530 -1280
rect 15770 -1300 15870 -1280
rect 16110 -1300 16210 -1280
rect 16450 -1300 16550 -1280
rect 16790 -1300 16890 -1280
rect 17130 -1300 17230 -1280
rect 17470 -1300 17570 -1280
rect 17810 -1300 17910 -1280
rect 18150 -1300 18250 -1280
rect 18490 -1300 18590 -1280
rect 18830 -1300 18930 -1280
rect 19170 -1300 19270 -1280
rect 19510 -1300 19610 -1280
rect 19850 -1300 19950 -1280
rect 20190 -1300 20290 -1280
rect 20530 -1300 20630 -1280
rect 20870 -1300 20970 -1280
rect 21210 -1300 21310 -1280
rect 21550 -1300 21650 -1280
rect 21890 -1300 21990 -1280
rect 22230 -1300 22330 -1280
rect 22570 -1300 22670 -1280
rect 22910 -1300 23010 -1280
rect 23250 -1300 23350 -1280
rect 23590 -1300 23690 -1280
rect 23930 -1300 24030 -1280
rect 24270 -1300 24370 -1280
rect 24610 -1300 24710 -1280
rect 24950 -1300 25050 -1280
rect 25290 -1300 25390 -1280
rect 25630 -1300 25730 -1280
rect 25970 -1300 26070 -1280
rect 26310 -1300 26410 -1280
rect 26650 -1300 26750 -1280
rect 26990 -1300 27090 -1280
rect 27330 -1300 27430 -1280
rect 27670 -1300 27770 -1280
rect 28010 -1300 28110 -1280
rect 28350 -1300 28450 -1280
rect 28690 -1300 28790 -1280
rect 29030 -1300 29130 -1280
rect 29370 -1300 29470 -1280
rect 29710 -1300 29810 -1280
rect 30050 -1300 30150 -1280
rect 30390 -1300 30490 -1280
rect 30730 -1300 30830 -1280
rect 31070 -1300 31170 -1280
rect 31410 -1300 31510 -1280
rect 31750 -1300 31850 -1280
rect 32090 -1300 32190 -1280
rect 32430 -1300 32530 -1280
rect 32770 -1300 32870 -1280
rect 33110 -1300 33210 -1280
rect 33450 -1300 33550 -1280
rect 33790 -1300 33890 -1280
rect 34130 -1300 34230 -1280
rect 34470 -1300 34570 -1280
rect 34810 -1300 34910 -1280
rect 35150 -1300 35250 -1280
rect 35490 -1300 35590 -1280
rect 35830 -1300 35930 -1280
rect 36170 -1300 36270 -1280
rect 36510 -1300 36610 -1280
rect 36850 -1300 36950 -1280
rect 37190 -1300 37290 -1280
rect 37530 -1300 37630 -1280
rect 37870 -1300 37970 -1280
rect 38210 -1300 38310 -1280
rect 38550 -1300 38650 -1280
rect 38890 -1300 38990 -1280
rect 39230 -1300 39330 -1280
rect 39570 -1300 39670 -1280
rect 39910 -1300 40010 -1280
rect 40250 -1300 40350 -1280
rect 40590 -1300 40690 -1280
rect 40930 -1300 41030 -1280
rect 41270 -1300 41370 -1280
rect 41610 -1300 41710 -1280
rect 41950 -1300 42050 -1280
rect 42290 -1300 42390 -1280
rect 42630 -1300 42730 -1280
rect 42970 -1300 43070 -1280
rect 43310 -1300 43410 -1280
rect 43650 -1300 43750 -1280
rect 43990 -1300 44090 -1280
rect 44330 -1300 44430 -1280
rect 44670 -1300 44770 -1280
rect 45010 -1300 45110 -1280
rect 45350 -1300 45450 -1280
rect 45690 -1300 45790 -1280
rect 46030 -1300 46130 -1280
rect 46370 -1300 46470 -1280
rect 46710 -1300 46810 -1280
rect 47050 -1300 47150 -1280
rect 47390 -1300 47490 -1280
rect 47730 -1300 47830 -1280
rect 48070 -1300 48170 -1280
rect 48410 -1300 48510 -1280
rect 48750 -1300 48850 -1280
rect 49090 -1300 49190 -1280
rect 49430 -1300 49530 -1280
rect 49770 -1300 49870 -1280
rect 50110 -1300 50210 -1280
rect 50450 -1300 50550 -1280
rect 50790 -1300 50890 -1280
rect 51130 -1300 51230 -1280
rect 51470 -1300 51570 -1280
rect 51810 -1300 51910 -1280
rect 52150 -1300 52250 -1280
rect 52490 -1300 52590 -1280
rect 52830 -1300 52930 -1280
rect 53170 -1300 53270 -1280
rect 53510 -1300 53610 -1280
rect 53850 -1300 53950 -1280
rect 54190 -1300 54290 -1280
rect 54530 -1300 54630 -1280
rect 54870 -1300 54970 -1280
rect 55210 -1300 55310 -1280
rect 55550 -1300 55650 -1280
rect 55890 -1300 55990 -1280
rect 56230 -1300 56330 -1280
rect 56570 -1300 56670 -1280
rect 56910 -1300 57010 -1280
rect 57250 -1300 57350 -1280
rect 57590 -1300 57690 -1280
rect 57930 -1300 58030 -1280
rect 58270 -1300 58370 -1280
rect 58610 -1300 58710 -1280
rect 58950 -1300 59050 -1280
rect 59290 -1300 59390 -1280
rect 59630 -1300 59730 -1280
rect 59970 -1300 60070 -1280
rect 60310 -1300 60410 -1280
rect 60650 -1300 60750 -1280
rect 60990 -1300 61090 -1280
rect 61330 -1300 61430 -1280
rect 61670 -1300 61770 -1280
rect 62010 -1300 62110 -1280
rect 62350 -1300 62450 -1280
rect 62690 -1300 62790 -1280
rect 63030 -1300 63130 -1280
rect 63370 -1300 63470 -1280
rect 63710 -1300 63810 -1280
rect 64050 -1300 64150 -1280
rect 64390 -1300 64490 -1280
rect 64730 -1300 64830 -1280
rect 65070 -1300 65170 -1280
rect 65410 -1300 65510 -1280
rect 65750 -1300 65850 -1280
rect 66090 -1300 66190 -1280
rect 66430 -1300 66530 -1280
rect 66770 -1300 66870 -1280
rect 67110 -1300 67210 -1280
rect 67450 -1300 67550 -1280
rect 67790 -1300 67890 -1280
rect 68130 -1300 68230 -1280
rect 68470 -1300 68570 -1280
rect 68810 -1300 68910 -1280
rect 69150 -1300 69250 -1280
rect 69490 -1300 69590 -1280
rect 69830 -1300 69930 -1280
rect 70170 -1300 70270 -1280
rect 70510 -1300 70610 -1280
rect 70850 -1300 70950 -1280
rect 71190 -1300 71290 -1280
rect 71530 -1300 71630 -1280
rect 71870 -1300 71970 -1280
rect 72210 -1300 72310 -1280
rect 72550 -1300 72650 -1280
rect 72890 -1300 72990 -1280
rect 73230 -1300 73330 -1280
rect 73570 -1300 73670 -1280
rect 73910 -1300 74010 -1280
rect 74250 -1300 74350 -1280
rect 74590 -1300 74690 -1280
rect 74930 -1300 75030 -1280
rect 75270 -1300 75370 -1280
rect 75610 -1300 75710 -1280
rect 75950 -1300 76050 -1280
rect 76290 -1300 76390 -1280
rect 76630 -1300 76730 -1280
rect 76970 -1300 77070 -1280
rect 77310 -1300 77410 -1280
rect 77650 -1300 77750 -1280
rect 77990 -1300 78090 -1280
rect 78330 -1300 78430 -1280
rect 78670 -1300 78770 -1280
rect 79010 -1300 79110 -1280
rect 79350 -1300 79450 -1280
rect 79690 -1300 79790 -1280
rect 80030 -1300 80130 -1280
rect 80370 -1300 80470 -1280
rect 80710 -1300 80810 -1280
rect 81050 -1300 81150 -1280
rect 81390 -1300 81490 -1280
rect 81730 -1300 81830 -1280
rect 82070 -1300 82170 -1280
rect 82410 -1300 82510 -1280
rect 82750 -1300 82850 -1280
rect 83090 -1300 83190 -1280
rect 83430 -1300 83530 -1280
rect 83770 -1300 83870 -1280
rect 84110 -1300 84210 -1280
rect 84450 -1300 84550 -1280
rect 84790 -1300 84890 -1280
rect 85130 -1300 85230 -1280
rect 85470 -1300 85570 -1280
rect 85810 -1300 85910 -1280
rect 86150 -1300 86250 -1280
rect 86490 -1300 86590 -1280
rect 86830 -1300 86930 -1280
rect 87170 -1300 87270 -1280
rect 110 -1360 150 -1300
rect 210 -1360 490 -1300
rect 550 -1360 830 -1300
rect 890 -1360 1170 -1300
rect 1230 -1360 1510 -1300
rect 1570 -1360 1850 -1300
rect 1910 -1360 2190 -1300
rect 2250 -1360 2530 -1300
rect 2590 -1360 2870 -1300
rect 2930 -1360 3210 -1300
rect 3270 -1360 3550 -1300
rect 3610 -1360 3890 -1300
rect 3950 -1360 4230 -1300
rect 4290 -1360 4570 -1300
rect 4630 -1360 4910 -1300
rect 4970 -1360 5250 -1300
rect 5310 -1360 5590 -1300
rect 5650 -1360 5930 -1300
rect 5990 -1360 6270 -1300
rect 6330 -1360 6610 -1300
rect 6670 -1360 6950 -1300
rect 7010 -1360 7290 -1300
rect 7350 -1360 7630 -1300
rect 7690 -1360 7970 -1300
rect 8030 -1360 8310 -1300
rect 8370 -1360 8650 -1300
rect 8710 -1360 8990 -1300
rect 9050 -1360 9330 -1300
rect 9390 -1360 9670 -1300
rect 9730 -1360 10010 -1300
rect 10070 -1360 10350 -1300
rect 10410 -1360 10690 -1300
rect 10750 -1360 11030 -1300
rect 11090 -1360 11370 -1300
rect 11430 -1360 11710 -1300
rect 11770 -1360 12050 -1300
rect 12110 -1360 12390 -1300
rect 12450 -1360 12730 -1300
rect 12790 -1360 13070 -1300
rect 13130 -1360 13410 -1300
rect 13470 -1360 13750 -1300
rect 13810 -1360 14090 -1300
rect 14150 -1360 14430 -1300
rect 14490 -1360 14770 -1300
rect 14830 -1360 15110 -1300
rect 15170 -1360 15450 -1300
rect 15510 -1360 15790 -1300
rect 15850 -1360 16130 -1300
rect 16190 -1360 16470 -1300
rect 16530 -1360 16810 -1300
rect 16870 -1360 17150 -1300
rect 17210 -1360 17490 -1300
rect 17550 -1360 17830 -1300
rect 17890 -1360 18170 -1300
rect 18230 -1360 18510 -1300
rect 18570 -1360 18850 -1300
rect 18910 -1360 19190 -1300
rect 19250 -1360 19530 -1300
rect 19590 -1360 19870 -1300
rect 19930 -1360 20210 -1300
rect 20270 -1360 20550 -1300
rect 20610 -1360 20890 -1300
rect 20950 -1360 21230 -1300
rect 21290 -1360 21570 -1300
rect 21630 -1360 21910 -1300
rect 21970 -1360 22250 -1300
rect 22310 -1360 22590 -1300
rect 22650 -1360 22930 -1300
rect 22990 -1360 23270 -1300
rect 23330 -1360 23610 -1300
rect 23670 -1360 23950 -1300
rect 24010 -1360 24290 -1300
rect 24350 -1360 24630 -1300
rect 24690 -1360 24970 -1300
rect 25030 -1360 25310 -1300
rect 25370 -1360 25650 -1300
rect 25710 -1360 25990 -1300
rect 26050 -1360 26330 -1300
rect 26390 -1360 26670 -1300
rect 26730 -1360 27010 -1300
rect 27070 -1360 27350 -1300
rect 27410 -1360 27690 -1300
rect 27750 -1360 28030 -1300
rect 28090 -1360 28370 -1300
rect 28430 -1360 28710 -1300
rect 28770 -1360 29050 -1300
rect 29110 -1360 29390 -1300
rect 29450 -1360 29730 -1300
rect 29790 -1360 30070 -1300
rect 30130 -1360 30410 -1300
rect 30470 -1360 30750 -1300
rect 30810 -1360 31090 -1300
rect 31150 -1360 31430 -1300
rect 31490 -1360 31770 -1300
rect 31830 -1360 32110 -1300
rect 32170 -1360 32450 -1300
rect 32510 -1360 32790 -1300
rect 32850 -1360 33130 -1300
rect 33190 -1360 33470 -1300
rect 33530 -1360 33810 -1300
rect 33870 -1360 34150 -1300
rect 34210 -1360 34490 -1300
rect 34550 -1360 34830 -1300
rect 34890 -1360 35170 -1300
rect 35230 -1360 35510 -1300
rect 35570 -1360 35850 -1300
rect 35910 -1360 36190 -1300
rect 36250 -1360 36530 -1300
rect 36590 -1360 36870 -1300
rect 36930 -1360 37210 -1300
rect 37270 -1360 37550 -1300
rect 37610 -1360 37890 -1300
rect 37950 -1360 38230 -1300
rect 38290 -1360 38570 -1300
rect 38630 -1360 38910 -1300
rect 38970 -1360 39250 -1300
rect 39310 -1360 39590 -1300
rect 39650 -1360 39930 -1300
rect 39990 -1360 40270 -1300
rect 40330 -1360 40610 -1300
rect 40670 -1360 40950 -1300
rect 41010 -1360 41290 -1300
rect 41350 -1360 41630 -1300
rect 41690 -1360 41970 -1300
rect 42030 -1360 42310 -1300
rect 42370 -1360 42650 -1300
rect 42710 -1360 42990 -1300
rect 43050 -1360 43330 -1300
rect 43390 -1360 43670 -1300
rect 43730 -1360 44010 -1300
rect 44070 -1360 44350 -1300
rect 44410 -1360 44690 -1300
rect 44750 -1360 45030 -1300
rect 45090 -1360 45370 -1300
rect 45430 -1360 45710 -1300
rect 45770 -1360 46050 -1300
rect 46110 -1360 46390 -1300
rect 46450 -1360 46730 -1300
rect 46790 -1360 47070 -1300
rect 47130 -1360 47410 -1300
rect 47470 -1360 47750 -1300
rect 47810 -1360 48090 -1300
rect 48150 -1360 48430 -1300
rect 48490 -1360 48770 -1300
rect 48830 -1360 49110 -1300
rect 49170 -1360 49450 -1300
rect 49510 -1360 49790 -1300
rect 49850 -1360 50130 -1300
rect 50190 -1360 50470 -1300
rect 50530 -1360 50810 -1300
rect 50870 -1360 51150 -1300
rect 51210 -1360 51490 -1300
rect 51550 -1360 51830 -1300
rect 51890 -1360 52170 -1300
rect 52230 -1360 52510 -1300
rect 52570 -1360 52850 -1300
rect 52910 -1360 53190 -1300
rect 53250 -1360 53530 -1300
rect 53590 -1360 53870 -1300
rect 53930 -1360 54210 -1300
rect 54270 -1360 54550 -1300
rect 54610 -1360 54890 -1300
rect 54950 -1360 55230 -1300
rect 55290 -1360 55570 -1300
rect 55630 -1360 55910 -1300
rect 55970 -1360 56250 -1300
rect 56310 -1360 56590 -1300
rect 56650 -1360 56930 -1300
rect 56990 -1360 57270 -1300
rect 57330 -1360 57610 -1300
rect 57670 -1360 57950 -1300
rect 58010 -1360 58290 -1300
rect 58350 -1360 58630 -1300
rect 58690 -1360 58970 -1300
rect 59030 -1360 59310 -1300
rect 59370 -1360 59650 -1300
rect 59710 -1360 59990 -1300
rect 60050 -1360 60330 -1300
rect 60390 -1360 60670 -1300
rect 60730 -1360 61010 -1300
rect 61070 -1360 61350 -1300
rect 61410 -1360 61690 -1300
rect 61750 -1360 62030 -1300
rect 62090 -1360 62370 -1300
rect 62430 -1360 62710 -1300
rect 62770 -1360 63050 -1300
rect 63110 -1360 63390 -1300
rect 63450 -1360 63730 -1300
rect 63790 -1360 64070 -1300
rect 64130 -1360 64410 -1300
rect 64470 -1360 64750 -1300
rect 64810 -1360 65090 -1300
rect 65150 -1360 65430 -1300
rect 65490 -1360 65770 -1300
rect 65830 -1360 66110 -1300
rect 66170 -1360 66450 -1300
rect 66510 -1360 66790 -1300
rect 66850 -1360 67130 -1300
rect 67190 -1360 67470 -1300
rect 67530 -1360 67810 -1300
rect 67870 -1360 68150 -1300
rect 68210 -1360 68490 -1300
rect 68550 -1360 68830 -1300
rect 68890 -1360 69170 -1300
rect 69230 -1360 69510 -1300
rect 69570 -1360 69850 -1300
rect 69910 -1360 70190 -1300
rect 70250 -1360 70530 -1300
rect 70590 -1360 70870 -1300
rect 70930 -1360 71210 -1300
rect 71270 -1360 71550 -1300
rect 71610 -1360 71890 -1300
rect 71950 -1360 72230 -1300
rect 72290 -1360 72570 -1300
rect 72630 -1360 72910 -1300
rect 72970 -1360 73250 -1300
rect 73310 -1360 73590 -1300
rect 73650 -1360 73930 -1300
rect 73990 -1360 74270 -1300
rect 74330 -1360 74610 -1300
rect 74670 -1360 74950 -1300
rect 75010 -1360 75290 -1300
rect 75350 -1360 75630 -1300
rect 75690 -1360 75970 -1300
rect 76030 -1360 76310 -1300
rect 76370 -1360 76650 -1300
rect 76710 -1360 76990 -1300
rect 77050 -1360 77330 -1300
rect 77390 -1360 77670 -1300
rect 77730 -1360 78010 -1300
rect 78070 -1360 78350 -1300
rect 78410 -1360 78690 -1300
rect 78750 -1360 79030 -1300
rect 79090 -1360 79370 -1300
rect 79430 -1360 79710 -1300
rect 79770 -1360 80050 -1300
rect 80110 -1360 80390 -1300
rect 80450 -1360 80730 -1300
rect 80790 -1360 81070 -1300
rect 81130 -1360 81410 -1300
rect 81470 -1360 81750 -1300
rect 81810 -1360 82090 -1300
rect 82150 -1360 82430 -1300
rect 82490 -1360 82770 -1300
rect 82830 -1360 83110 -1300
rect 83170 -1360 83450 -1300
rect 83510 -1360 83790 -1300
rect 83850 -1360 84130 -1300
rect 84190 -1360 84470 -1300
rect 84530 -1360 84810 -1300
rect 84870 -1360 85150 -1300
rect 85210 -1360 85490 -1300
rect 85550 -1360 85830 -1300
rect 85890 -1360 86170 -1300
rect 86230 -1360 86510 -1300
rect 86570 -1360 86850 -1300
rect 86910 -1360 87190 -1300
rect 87250 -1360 87270 -1300
rect 130 -1380 230 -1360
rect 470 -1380 570 -1360
rect 810 -1380 910 -1360
rect 1150 -1380 1250 -1360
rect 1490 -1380 1590 -1360
rect 1830 -1380 1930 -1360
rect 2170 -1380 2270 -1360
rect 2510 -1380 2610 -1360
rect 2850 -1380 2950 -1360
rect 3190 -1380 3290 -1360
rect 3530 -1380 3630 -1360
rect 3870 -1380 3970 -1360
rect 4210 -1380 4310 -1360
rect 4550 -1380 4650 -1360
rect 4890 -1380 4990 -1360
rect 5230 -1380 5330 -1360
rect 5570 -1380 5670 -1360
rect 5910 -1380 6010 -1360
rect 6250 -1380 6350 -1360
rect 6590 -1380 6690 -1360
rect 6930 -1380 7030 -1360
rect 7270 -1380 7370 -1360
rect 7610 -1380 7710 -1360
rect 7950 -1380 8050 -1360
rect 8290 -1380 8390 -1360
rect 8630 -1380 8730 -1360
rect 8970 -1380 9070 -1360
rect 9310 -1380 9410 -1360
rect 9650 -1380 9750 -1360
rect 9990 -1380 10090 -1360
rect 10330 -1380 10430 -1360
rect 10670 -1380 10770 -1360
rect 11010 -1380 11110 -1360
rect 11350 -1380 11450 -1360
rect 11690 -1380 11790 -1360
rect 12030 -1380 12130 -1360
rect 12370 -1380 12470 -1360
rect 12710 -1380 12810 -1360
rect 13050 -1380 13150 -1360
rect 13390 -1380 13490 -1360
rect 13730 -1380 13830 -1360
rect 14070 -1380 14170 -1360
rect 14410 -1380 14510 -1360
rect 14750 -1380 14850 -1360
rect 15090 -1380 15190 -1360
rect 15430 -1380 15530 -1360
rect 15770 -1380 15870 -1360
rect 16110 -1380 16210 -1360
rect 16450 -1380 16550 -1360
rect 16790 -1380 16890 -1360
rect 17130 -1380 17230 -1360
rect 17470 -1380 17570 -1360
rect 17810 -1380 17910 -1360
rect 18150 -1380 18250 -1360
rect 18490 -1380 18590 -1360
rect 18830 -1380 18930 -1360
rect 19170 -1380 19270 -1360
rect 19510 -1380 19610 -1360
rect 19850 -1380 19950 -1360
rect 20190 -1380 20290 -1360
rect 20530 -1380 20630 -1360
rect 20870 -1380 20970 -1360
rect 21210 -1380 21310 -1360
rect 21550 -1380 21650 -1360
rect 21890 -1380 21990 -1360
rect 22230 -1380 22330 -1360
rect 22570 -1380 22670 -1360
rect 22910 -1380 23010 -1360
rect 23250 -1380 23350 -1360
rect 23590 -1380 23690 -1360
rect 23930 -1380 24030 -1360
rect 24270 -1380 24370 -1360
rect 24610 -1380 24710 -1360
rect 24950 -1380 25050 -1360
rect 25290 -1380 25390 -1360
rect 25630 -1380 25730 -1360
rect 25970 -1380 26070 -1360
rect 26310 -1380 26410 -1360
rect 26650 -1380 26750 -1360
rect 26990 -1380 27090 -1360
rect 27330 -1380 27430 -1360
rect 27670 -1380 27770 -1360
rect 28010 -1380 28110 -1360
rect 28350 -1380 28450 -1360
rect 28690 -1380 28790 -1360
rect 29030 -1380 29130 -1360
rect 29370 -1380 29470 -1360
rect 29710 -1380 29810 -1360
rect 30050 -1380 30150 -1360
rect 30390 -1380 30490 -1360
rect 30730 -1380 30830 -1360
rect 31070 -1380 31170 -1360
rect 31410 -1380 31510 -1360
rect 31750 -1380 31850 -1360
rect 32090 -1380 32190 -1360
rect 32430 -1380 32530 -1360
rect 32770 -1380 32870 -1360
rect 33110 -1380 33210 -1360
rect 33450 -1380 33550 -1360
rect 33790 -1380 33890 -1360
rect 34130 -1380 34230 -1360
rect 34470 -1380 34570 -1360
rect 34810 -1380 34910 -1360
rect 35150 -1380 35250 -1360
rect 35490 -1380 35590 -1360
rect 35830 -1380 35930 -1360
rect 36170 -1380 36270 -1360
rect 36510 -1380 36610 -1360
rect 36850 -1380 36950 -1360
rect 37190 -1380 37290 -1360
rect 37530 -1380 37630 -1360
rect 37870 -1380 37970 -1360
rect 38210 -1380 38310 -1360
rect 38550 -1380 38650 -1360
rect 38890 -1380 38990 -1360
rect 39230 -1380 39330 -1360
rect 39570 -1380 39670 -1360
rect 39910 -1380 40010 -1360
rect 40250 -1380 40350 -1360
rect 40590 -1380 40690 -1360
rect 40930 -1380 41030 -1360
rect 41270 -1380 41370 -1360
rect 41610 -1380 41710 -1360
rect 41950 -1380 42050 -1360
rect 42290 -1380 42390 -1360
rect 42630 -1380 42730 -1360
rect 42970 -1380 43070 -1360
rect 43310 -1380 43410 -1360
rect 43650 -1380 43750 -1360
rect 43990 -1380 44090 -1360
rect 44330 -1380 44430 -1360
rect 44670 -1380 44770 -1360
rect 45010 -1380 45110 -1360
rect 45350 -1380 45450 -1360
rect 45690 -1380 45790 -1360
rect 46030 -1380 46130 -1360
rect 46370 -1380 46470 -1360
rect 46710 -1380 46810 -1360
rect 47050 -1380 47150 -1360
rect 47390 -1380 47490 -1360
rect 47730 -1380 47830 -1360
rect 48070 -1380 48170 -1360
rect 48410 -1380 48510 -1360
rect 48750 -1380 48850 -1360
rect 49090 -1380 49190 -1360
rect 49430 -1380 49530 -1360
rect 49770 -1380 49870 -1360
rect 50110 -1380 50210 -1360
rect 50450 -1380 50550 -1360
rect 50790 -1380 50890 -1360
rect 51130 -1380 51230 -1360
rect 51470 -1380 51570 -1360
rect 51810 -1380 51910 -1360
rect 52150 -1380 52250 -1360
rect 52490 -1380 52590 -1360
rect 52830 -1380 52930 -1360
rect 53170 -1380 53270 -1360
rect 53510 -1380 53610 -1360
rect 53850 -1380 53950 -1360
rect 54190 -1380 54290 -1360
rect 54530 -1380 54630 -1360
rect 54870 -1380 54970 -1360
rect 55210 -1380 55310 -1360
rect 55550 -1380 55650 -1360
rect 55890 -1380 55990 -1360
rect 56230 -1380 56330 -1360
rect 56570 -1380 56670 -1360
rect 56910 -1380 57010 -1360
rect 57250 -1380 57350 -1360
rect 57590 -1380 57690 -1360
rect 57930 -1380 58030 -1360
rect 58270 -1380 58370 -1360
rect 58610 -1380 58710 -1360
rect 58950 -1380 59050 -1360
rect 59290 -1380 59390 -1360
rect 59630 -1380 59730 -1360
rect 59970 -1380 60070 -1360
rect 60310 -1380 60410 -1360
rect 60650 -1380 60750 -1360
rect 60990 -1380 61090 -1360
rect 61330 -1380 61430 -1360
rect 61670 -1380 61770 -1360
rect 62010 -1380 62110 -1360
rect 62350 -1380 62450 -1360
rect 62690 -1380 62790 -1360
rect 63030 -1380 63130 -1360
rect 63370 -1380 63470 -1360
rect 63710 -1380 63810 -1360
rect 64050 -1380 64150 -1360
rect 64390 -1380 64490 -1360
rect 64730 -1380 64830 -1360
rect 65070 -1380 65170 -1360
rect 65410 -1380 65510 -1360
rect 65750 -1380 65850 -1360
rect 66090 -1380 66190 -1360
rect 66430 -1380 66530 -1360
rect 66770 -1380 66870 -1360
rect 67110 -1380 67210 -1360
rect 67450 -1380 67550 -1360
rect 67790 -1380 67890 -1360
rect 68130 -1380 68230 -1360
rect 68470 -1380 68570 -1360
rect 68810 -1380 68910 -1360
rect 69150 -1380 69250 -1360
rect 69490 -1380 69590 -1360
rect 69830 -1380 69930 -1360
rect 70170 -1380 70270 -1360
rect 70510 -1380 70610 -1360
rect 70850 -1380 70950 -1360
rect 71190 -1380 71290 -1360
rect 71530 -1380 71630 -1360
rect 71870 -1380 71970 -1360
rect 72210 -1380 72310 -1360
rect 72550 -1380 72650 -1360
rect 72890 -1380 72990 -1360
rect 73230 -1380 73330 -1360
rect 73570 -1380 73670 -1360
rect 73910 -1380 74010 -1360
rect 74250 -1380 74350 -1360
rect 74590 -1380 74690 -1360
rect 74930 -1380 75030 -1360
rect 75270 -1380 75370 -1360
rect 75610 -1380 75710 -1360
rect 75950 -1380 76050 -1360
rect 76290 -1380 76390 -1360
rect 76630 -1380 76730 -1360
rect 76970 -1380 77070 -1360
rect 77310 -1380 77410 -1360
rect 77650 -1380 77750 -1360
rect 77990 -1380 78090 -1360
rect 78330 -1380 78430 -1360
rect 78670 -1380 78770 -1360
rect 79010 -1380 79110 -1360
rect 79350 -1380 79450 -1360
rect 79690 -1380 79790 -1360
rect 80030 -1380 80130 -1360
rect 80370 -1380 80470 -1360
rect 80710 -1380 80810 -1360
rect 81050 -1380 81150 -1360
rect 81390 -1380 81490 -1360
rect 81730 -1380 81830 -1360
rect 82070 -1380 82170 -1360
rect 82410 -1380 82510 -1360
rect 82750 -1380 82850 -1360
rect 83090 -1380 83190 -1360
rect 83430 -1380 83530 -1360
rect 83770 -1380 83870 -1360
rect 84110 -1380 84210 -1360
rect 84450 -1380 84550 -1360
rect 84790 -1380 84890 -1360
rect 85130 -1380 85230 -1360
rect 85470 -1380 85570 -1360
rect 85810 -1380 85910 -1360
rect 86150 -1380 86250 -1360
rect 86490 -1380 86590 -1360
rect 86830 -1380 86930 -1360
rect 87170 -1380 87270 -1360
rect 770 -1470 970 -1440
rect 770 -1540 830 -1470
rect 910 -1540 970 -1470
rect 770 -1570 970 -1540
rect 4940 -1470 5140 -1440
rect 4940 -1540 5000 -1470
rect 5080 -1540 5140 -1470
rect 4940 -1570 5140 -1540
rect 8970 -1470 9170 -1440
rect 8970 -1540 9030 -1470
rect 9110 -1540 9170 -1470
rect 8970 -1570 9170 -1540
rect 13000 -1470 13200 -1440
rect 13000 -1540 13060 -1470
rect 13140 -1540 13200 -1470
rect 13000 -1570 13200 -1540
rect 17040 -1470 17240 -1440
rect 17040 -1540 17100 -1470
rect 17180 -1540 17240 -1470
rect 17040 -1570 17240 -1540
rect 21140 -1470 21340 -1440
rect 21140 -1540 21200 -1470
rect 21280 -1540 21340 -1470
rect 21140 -1570 21340 -1540
rect 25250 -1470 25450 -1440
rect 25250 -1540 25310 -1470
rect 25390 -1540 25450 -1470
rect 25250 -1570 25450 -1540
rect 29350 -1470 29550 -1440
rect 29350 -1540 29410 -1470
rect 29490 -1540 29550 -1470
rect 29350 -1570 29550 -1540
rect 33380 -1470 33580 -1440
rect 33380 -1540 33440 -1470
rect 33520 -1540 33580 -1470
rect 33380 -1570 33580 -1540
rect 37490 -1470 37690 -1440
rect 37490 -1540 37550 -1470
rect 37630 -1540 37690 -1470
rect 37490 -1570 37690 -1540
rect 41590 -1470 41790 -1440
rect 41590 -1540 41650 -1470
rect 41730 -1540 41790 -1470
rect 41590 -1570 41790 -1540
rect 47040 -1470 47240 -1440
rect 47040 -1540 47100 -1470
rect 47180 -1540 47240 -1470
rect 47040 -1570 47240 -1540
rect 51120 -1470 51320 -1440
rect 51120 -1540 51180 -1470
rect 51260 -1540 51320 -1470
rect 51120 -1570 51320 -1540
rect 55230 -1470 55430 -1440
rect 55230 -1540 55290 -1470
rect 55370 -1540 55430 -1470
rect 55230 -1570 55430 -1540
rect 59260 -1470 59460 -1440
rect 59260 -1540 59320 -1470
rect 59400 -1540 59460 -1470
rect 59260 -1570 59460 -1540
rect 63360 -1470 63560 -1440
rect 63360 -1540 63420 -1470
rect 63500 -1540 63560 -1470
rect 63360 -1570 63560 -1540
rect 67470 -1470 67670 -1440
rect 67470 -1540 67530 -1470
rect 67610 -1540 67670 -1470
rect 67470 -1570 67670 -1540
rect 71500 -1470 71700 -1440
rect 71500 -1540 71560 -1470
rect 71640 -1540 71700 -1470
rect 71500 -1570 71700 -1540
rect 75750 -1470 75950 -1440
rect 75750 -1540 75810 -1470
rect 75890 -1540 75950 -1470
rect 75750 -1570 75950 -1540
rect 79710 -1470 79910 -1440
rect 79710 -1540 79770 -1470
rect 79850 -1540 79910 -1470
rect 79710 -1570 79910 -1540
rect 83890 -1470 84090 -1440
rect 83890 -1540 83950 -1470
rect 84030 -1540 84090 -1470
rect 83890 -1570 84090 -1540
rect 86450 -1474 86648 -1444
rect 86450 -1544 86508 -1474
rect 86588 -1544 86648 -1474
rect 86450 -1572 86648 -1544
<< via2 >>
rect 1300 650 1390 710
rect 6390 630 6490 690
rect 790 520 870 590
rect 2170 520 2250 590
rect 3550 520 3630 590
rect 5210 520 5290 590
rect 8040 520 8120 590
rect 10800 520 10880 590
rect 13430 520 13510 590
rect 16470 520 16550 590
rect 20540 520 20620 590
rect 24680 520 24760 590
rect 28760 520 28840 590
rect 32910 520 32990 590
rect 36780 520 36860 590
rect 40920 520 41000 590
rect 44910 520 44990 590
rect 48990 520 49070 590
rect 53080 520 53160 590
rect 57240 520 57320 590
rect 30 350 90 410
rect 450 350 510 410
rect 1130 350 1190 410
rect 1520 350 1580 410
rect 2880 350 2940 410
rect 4240 350 4300 410
rect 4540 350 4600 410
rect 5900 350 5960 410
rect 7260 350 7320 410
rect 8620 350 8680 410
rect 9980 350 10040 410
rect 11340 350 11400 410
rect 12700 350 12760 410
rect 14060 350 14120 410
rect 15420 350 15480 410
rect 15720 350 15780 410
rect 17080 350 17140 410
rect 18440 350 18500 410
rect 19800 350 19860 410
rect 21160 350 21220 410
rect 22520 350 22580 410
rect 23880 350 23940 410
rect 25240 350 25300 410
rect 26600 350 26660 410
rect 27960 350 28020 410
rect 29320 350 29380 410
rect 30680 350 30740 410
rect 32040 350 32100 410
rect 33400 350 33460 410
rect 34760 350 34820 410
rect 36120 350 36180 410
rect 37480 350 37540 410
rect 38840 350 38900 410
rect 40200 350 40260 410
rect 41560 350 41620 410
rect 42920 350 42980 410
rect 44280 350 44340 410
rect 45640 350 45700 410
rect 47000 350 47060 410
rect 48360 350 48420 410
rect 49720 350 49780 410
rect 51080 350 51140 410
rect 52440 350 52500 410
rect 53800 350 53860 410
rect 55160 350 55220 410
rect 56520 350 56580 410
rect 57880 350 57940 410
rect 59240 350 59300 410
rect 620 130 680 200
rect 960 130 1020 200
rect 1690 130 1750 200
rect 2030 130 2090 200
rect 2370 130 2430 200
rect 2710 130 2770 200
rect 3050 130 3110 200
rect 3390 130 3450 200
rect 3730 130 3790 200
rect 4070 130 4130 200
rect 4710 130 4770 200
rect 5050 130 5110 200
rect 5390 130 5450 200
rect 5730 130 5790 200
rect 6070 130 6130 200
rect 6410 130 6470 200
rect 6750 130 6810 200
rect 7090 130 7150 200
rect 7430 130 7490 200
rect 7770 130 7830 200
rect 8110 130 8170 200
rect 8450 130 8510 200
rect 8790 130 8850 200
rect 9130 130 9190 200
rect 9470 130 9530 200
rect 9810 130 9870 200
rect 10150 130 10210 200
rect 10490 130 10550 200
rect 10830 130 10890 200
rect 11170 130 11230 200
rect 11510 130 11570 200
rect 11850 130 11910 200
rect 12190 130 12250 200
rect 12530 130 12590 200
rect 12870 130 12930 200
rect 13210 130 13270 200
rect 13550 130 13610 200
rect 13890 130 13950 200
rect 14230 130 14290 200
rect 14570 130 14630 200
rect 14910 130 14970 200
rect 15250 130 15310 200
rect 15890 130 15950 200
rect 16230 130 16290 200
rect 16570 130 16630 200
rect 16910 130 16970 200
rect 17250 130 17310 200
rect 17590 130 17650 200
rect 17930 130 17990 200
rect 18270 130 18330 200
rect 18610 130 18670 200
rect 18950 130 19010 200
rect 19290 130 19350 200
rect 19630 130 19690 200
rect 19970 130 20030 200
rect 20310 130 20370 200
rect 20650 130 20710 200
rect 20990 130 21050 200
rect 21330 130 21390 200
rect 21670 130 21730 200
rect 22010 130 22070 200
rect 22350 130 22410 200
rect 22690 130 22750 200
rect 23030 130 23090 200
rect 23370 130 23430 200
rect 23710 130 23770 200
rect 24050 130 24110 200
rect 24390 130 24450 200
rect 24730 130 24790 200
rect 25070 130 25130 200
rect 25410 130 25470 200
rect 25750 130 25810 200
rect 26090 130 26150 200
rect 26430 130 26490 200
rect 26770 130 26830 200
rect 27110 130 27170 200
rect 27450 130 27510 200
rect 27790 130 27850 200
rect 28130 130 28190 200
rect 28470 130 28530 200
rect 28810 130 28870 200
rect 29150 130 29210 200
rect 29490 130 29550 200
rect 29830 130 29890 200
rect 30170 130 30230 200
rect 30510 130 30570 200
rect 30850 130 30910 200
rect 31190 130 31250 200
rect 31530 130 31590 200
rect 31870 130 31930 200
rect 32210 130 32270 200
rect 32550 130 32610 200
rect 32890 130 32950 200
rect 33230 130 33290 200
rect 33570 130 33630 200
rect 33910 130 33970 200
rect 34250 130 34310 200
rect 34590 130 34650 200
rect 34930 130 34990 200
rect 35270 130 35330 200
rect 35610 130 35670 200
rect 35950 130 36010 200
rect 36290 130 36350 200
rect 36630 130 36690 200
rect 36970 130 37030 200
rect 37310 130 37370 200
rect 37650 130 37710 200
rect 37990 130 38050 200
rect 38330 130 38390 200
rect 38670 130 38730 200
rect 39010 130 39070 200
rect 39350 130 39410 200
rect 39690 130 39750 200
rect 40030 130 40090 200
rect 40370 130 40430 200
rect 40710 130 40770 200
rect 41050 130 41110 200
rect 41390 130 41450 200
rect 41730 130 41790 200
rect 42070 130 42130 200
rect 42410 130 42470 200
rect 42750 130 42810 200
rect 43090 130 43150 200
rect 43430 130 43490 200
rect 43770 130 43830 200
rect 44110 130 44170 200
rect 44450 130 44510 200
rect 44790 130 44850 200
rect 45130 130 45190 200
rect 45470 130 45530 200
rect 45810 130 45870 200
rect 46150 130 46210 200
rect 46490 130 46550 200
rect 46830 130 46890 200
rect 47170 130 47230 200
rect 47510 130 47570 200
rect 47850 130 47910 200
rect 48190 130 48250 200
rect 48530 130 48590 200
rect 48870 130 48930 200
rect 49210 130 49270 200
rect 49550 130 49610 200
rect 49890 130 49950 200
rect 50230 130 50290 200
rect 50570 130 50630 200
rect 50910 130 50970 200
rect 51250 130 51310 200
rect 51590 130 51650 200
rect 51930 130 51990 200
rect 52270 130 52330 200
rect 52610 130 52670 200
rect 52950 130 53010 200
rect 53290 130 53350 200
rect 53630 130 53690 200
rect 53970 130 54030 200
rect 54310 130 54370 200
rect 54650 130 54710 200
rect 54990 130 55050 200
rect 55330 130 55390 200
rect 55670 130 55730 200
rect 56010 130 56070 200
rect 56350 130 56410 200
rect 56690 130 56750 200
rect 57030 130 57090 200
rect 57370 130 57430 200
rect 57710 130 57770 200
rect 58050 130 58110 200
rect 58390 130 58450 200
rect 58730 130 58790 200
rect 59070 130 59130 200
rect 450 20 510 80
rect 1130 20 1190 80
rect 1520 20 1580 80
rect 2880 20 2940 80
rect 4880 20 4940 80
rect 6240 20 6300 80
rect 7260 20 7320 80
rect 8620 20 8680 80
rect 9980 20 10040 80
rect 11000 20 11060 80
rect 16400 20 16460 80
rect 17760 20 17820 80
rect 18780 20 18840 80
rect 20140 20 20200 80
rect 21500 20 21560 80
rect 22520 20 22580 80
rect 23880 20 23940 80
rect 24560 20 24620 80
rect 28300 20 28360 80
rect 29660 20 29720 80
rect 30680 20 30740 80
rect 32040 20 32100 80
rect 33400 20 33460 80
rect 34420 20 34480 80
rect 35780 20 35840 80
rect 36460 20 36520 80
rect 42580 20 42640 80
rect 44620 20 44680 80
rect 48360 20 48420 80
rect 49720 20 49780 80
rect 50740 20 50800 80
rect 52100 20 52160 80
rect 53460 20 53520 80
rect 55500 20 55560 80
rect 30 -120 90 -60
rect 1300 -130 1400 -50
rect 4380 -130 4480 -50
rect 15560 -130 15660 -50
rect 2120 -390 2350 -260
rect 5138 -398 5368 -268
rect 7624 -398 7854 -268
rect 9044 -398 9274 -268
rect 13668 -394 13898 -264
rect 16868 -394 17098 -264
rect 20424 -394 20654 -264
rect 25758 -394 25988 -264
rect 28602 -394 28832 -264
rect 32514 -394 32744 -264
rect 34670 -394 34900 -264
rect 37492 -394 37722 -264
rect 40692 -394 40922 -264
rect 45668 -394 45898 -264
rect 48868 -394 49098 -264
rect 51002 -394 51232 -264
rect 54558 -394 54788 -264
rect 57402 -394 57632 -264
rect 61314 -394 61544 -264
rect 64158 -394 64388 -264
rect 67714 -394 67944 -264
rect 70558 -394 70788 -264
rect 74468 -394 74698 -264
rect 78380 -394 78610 -264
rect 82292 -394 82522 -264
rect 86202 -394 86432 -264
rect 15930 -520 16000 -460
rect 31230 -520 31300 -460
rect 59110 -520 59180 -460
rect 150 -730 210 -670
rect 1510 -730 1570 -670
rect 2870 -730 2930 -670
rect 4570 -730 4630 -670
rect 5930 -730 5990 -670
rect 6950 -730 7010 -670
rect 8310 -730 8370 -670
rect 9670 -730 9730 -670
rect 10690 -730 10750 -670
rect 11710 -730 11770 -670
rect 13070 -730 13130 -670
rect 14430 -730 14490 -670
rect 16130 -730 16190 -670
rect 17490 -730 17550 -670
rect 18510 -730 18570 -670
rect 19870 -730 19930 -670
rect 21230 -730 21290 -670
rect 22250 -730 22310 -670
rect 23610 -730 23670 -670
rect 24970 -730 25030 -670
rect 26330 -730 26390 -670
rect 28030 -730 28090 -670
rect 29390 -730 29450 -670
rect 30410 -730 30470 -670
rect 31770 -730 31830 -670
rect 33130 -730 33190 -670
rect 34150 -730 34210 -670
rect 35510 -730 35570 -670
rect 36870 -730 36930 -670
rect 38230 -730 38290 -670
rect 39930 -730 39990 -670
rect 41290 -730 41350 -670
rect 42310 -730 42370 -670
rect 43670 -730 43730 -670
rect 45030 -730 45090 -670
rect 46390 -730 46450 -670
rect 48090 -730 48150 -670
rect 49450 -730 49510 -670
rect 50470 -730 50530 -670
rect 51830 -730 51890 -670
rect 53190 -730 53250 -670
rect 54210 -730 54270 -670
rect 55230 -730 55290 -670
rect 56590 -730 56650 -670
rect 57950 -730 58010 -670
rect 59650 -730 59710 -670
rect 61010 -730 61070 -670
rect 62030 -730 62090 -670
rect 63390 -730 63450 -670
rect 64750 -730 64810 -670
rect 65770 -730 65830 -670
rect 67130 -730 67190 -670
rect 68490 -730 68550 -670
rect 69850 -730 69910 -670
rect 71550 -730 71610 -670
rect 72910 -730 72970 -670
rect 73930 -730 73990 -670
rect 75290 -730 75350 -670
rect 76650 -730 76710 -670
rect 77670 -730 77730 -670
rect 79030 -730 79090 -670
rect 80390 -730 80450 -670
rect 81750 -730 81810 -670
rect 83450 -730 83510 -670
rect 84810 -730 84870 -670
rect 85830 -730 85890 -670
rect 87190 -730 87250 -670
rect 320 -950 380 -880
rect 660 -950 720 -880
rect 1000 -950 1060 -880
rect 1340 -950 1400 -880
rect 1680 -950 1740 -880
rect 2020 -950 2080 -880
rect 2360 -950 2420 -880
rect 2700 -950 2760 -880
rect 3040 -950 3100 -880
rect 3380 -950 3440 -880
rect 3720 -950 3780 -880
rect 4060 -950 4120 -880
rect 4400 -950 4460 -880
rect 4740 -950 4800 -880
rect 5080 -950 5140 -880
rect 5420 -950 5480 -880
rect 5760 -950 5820 -880
rect 6100 -950 6160 -880
rect 6440 -950 6500 -880
rect 6780 -950 6840 -880
rect 7120 -950 7180 -880
rect 7460 -950 7520 -880
rect 7800 -950 7860 -880
rect 8140 -950 8200 -880
rect 8480 -950 8540 -880
rect 8820 -950 8880 -880
rect 9160 -950 9220 -880
rect 9500 -950 9560 -880
rect 9840 -950 9900 -880
rect 10180 -950 10240 -880
rect 10520 -950 10580 -880
rect 10860 -950 10920 -880
rect 11200 -950 11260 -880
rect 11540 -950 11600 -880
rect 11880 -950 11940 -880
rect 12220 -950 12280 -880
rect 12560 -950 12620 -880
rect 12900 -950 12960 -880
rect 13240 -950 13300 -880
rect 13580 -950 13640 -880
rect 13920 -950 13980 -880
rect 14260 -950 14320 -880
rect 14600 -950 14660 -880
rect 14940 -950 15000 -880
rect 15280 -950 15340 -880
rect 15620 -950 15680 -880
rect 15960 -950 16020 -880
rect 16300 -950 16360 -880
rect 16640 -950 16700 -880
rect 16980 -950 17040 -880
rect 17320 -950 17380 -880
rect 17660 -950 17720 -880
rect 18000 -950 18060 -880
rect 18340 -950 18400 -880
rect 18680 -950 18740 -880
rect 19020 -950 19080 -880
rect 19360 -950 19420 -880
rect 19700 -950 19760 -880
rect 20040 -950 20100 -880
rect 20380 -950 20440 -880
rect 20720 -950 20780 -880
rect 21060 -950 21120 -880
rect 21400 -950 21460 -880
rect 21740 -950 21800 -880
rect 22080 -950 22140 -880
rect 22420 -950 22480 -880
rect 22760 -950 22820 -880
rect 23100 -950 23160 -880
rect 23440 -950 23500 -880
rect 23780 -950 23840 -880
rect 24120 -950 24180 -880
rect 24460 -950 24520 -880
rect 24800 -950 24860 -880
rect 25140 -950 25200 -880
rect 25480 -950 25540 -880
rect 25820 -950 25880 -880
rect 26160 -950 26220 -880
rect 26500 -950 26560 -880
rect 26840 -950 26900 -880
rect 27180 -950 27240 -880
rect 27520 -950 27580 -880
rect 27860 -950 27920 -880
rect 28200 -950 28260 -880
rect 28540 -950 28600 -880
rect 28880 -950 28940 -880
rect 29220 -950 29280 -880
rect 29560 -950 29620 -880
rect 29900 -950 29960 -880
rect 30240 -950 30300 -880
rect 30580 -950 30640 -880
rect 30920 -950 30980 -880
rect 31260 -950 31320 -880
rect 31600 -950 31660 -880
rect 31940 -950 32000 -880
rect 32280 -950 32340 -880
rect 32620 -950 32680 -880
rect 32960 -950 33020 -880
rect 33300 -950 33360 -880
rect 33640 -950 33700 -880
rect 33980 -950 34040 -880
rect 34320 -950 34380 -880
rect 34660 -950 34720 -880
rect 35000 -950 35060 -880
rect 35340 -950 35400 -880
rect 35680 -950 35740 -880
rect 36020 -950 36080 -880
rect 36360 -950 36420 -880
rect 36700 -950 36760 -880
rect 37040 -950 37100 -880
rect 37380 -950 37440 -880
rect 37720 -950 37780 -880
rect 38060 -950 38120 -880
rect 38400 -950 38460 -880
rect 38740 -950 38800 -880
rect 39080 -950 39140 -880
rect 39420 -950 39480 -880
rect 39760 -950 39820 -880
rect 40100 -950 40160 -880
rect 40440 -950 40500 -880
rect 40780 -950 40840 -880
rect 41120 -950 41180 -880
rect 41460 -950 41520 -880
rect 41800 -950 41860 -880
rect 42140 -950 42200 -880
rect 42480 -950 42540 -880
rect 42820 -950 42880 -880
rect 43160 -950 43220 -880
rect 43500 -950 43560 -880
rect 43840 -950 43900 -880
rect 44180 -950 44240 -880
rect 44520 -950 44580 -880
rect 44860 -950 44920 -880
rect 45200 -950 45260 -880
rect 45540 -950 45600 -880
rect 45880 -950 45940 -880
rect 46220 -950 46280 -880
rect 46560 -950 46620 -880
rect 46900 -950 46960 -880
rect 47240 -950 47300 -880
rect 47580 -950 47640 -880
rect 47920 -950 47980 -880
rect 48260 -950 48320 -880
rect 48600 -950 48660 -880
rect 48940 -950 49000 -880
rect 49280 -950 49340 -880
rect 49620 -950 49680 -880
rect 49960 -950 50020 -880
rect 50300 -950 50360 -880
rect 50640 -950 50700 -880
rect 50980 -950 51040 -880
rect 51320 -950 51380 -880
rect 51660 -950 51720 -880
rect 52000 -950 52060 -880
rect 52340 -950 52400 -880
rect 52680 -950 52740 -880
rect 53020 -950 53080 -880
rect 53360 -950 53420 -880
rect 53700 -950 53760 -880
rect 54040 -950 54100 -880
rect 54380 -950 54440 -880
rect 54720 -950 54780 -880
rect 55060 -950 55120 -880
rect 55400 -950 55460 -880
rect 55740 -950 55800 -880
rect 56080 -950 56140 -880
rect 56420 -950 56480 -880
rect 56760 -950 56820 -880
rect 57100 -950 57160 -880
rect 57440 -950 57500 -880
rect 57780 -950 57840 -880
rect 58120 -950 58180 -880
rect 58460 -950 58520 -880
rect 58800 -950 58860 -880
rect 59140 -950 59200 -880
rect 59480 -950 59540 -880
rect 59820 -950 59880 -880
rect 60160 -950 60220 -880
rect 60500 -950 60560 -880
rect 60840 -950 60900 -880
rect 61180 -950 61240 -880
rect 61520 -950 61580 -880
rect 61860 -950 61920 -880
rect 62200 -950 62260 -880
rect 62540 -950 62600 -880
rect 62880 -950 62940 -880
rect 63220 -950 63280 -880
rect 63560 -950 63620 -880
rect 63900 -950 63960 -880
rect 64240 -950 64300 -880
rect 64580 -950 64640 -880
rect 64920 -950 64980 -880
rect 65260 -950 65320 -880
rect 65600 -950 65660 -880
rect 65940 -950 66000 -880
rect 66280 -950 66340 -880
rect 66620 -950 66680 -880
rect 66960 -950 67020 -880
rect 67300 -950 67360 -880
rect 67640 -950 67700 -880
rect 67980 -950 68040 -880
rect 68320 -950 68380 -880
rect 68660 -950 68720 -880
rect 69000 -950 69060 -880
rect 69340 -950 69400 -880
rect 69680 -950 69740 -880
rect 70020 -950 70080 -880
rect 70360 -950 70420 -880
rect 70700 -950 70760 -880
rect 71040 -950 71100 -880
rect 71380 -950 71440 -880
rect 71720 -950 71780 -880
rect 72060 -950 72120 -880
rect 72400 -950 72460 -880
rect 72740 -950 72800 -880
rect 73080 -950 73140 -880
rect 73420 -950 73480 -880
rect 73760 -950 73820 -880
rect 74100 -950 74160 -880
rect 74440 -950 74500 -880
rect 74780 -950 74840 -880
rect 75120 -950 75180 -880
rect 75460 -950 75520 -880
rect 75800 -950 75860 -880
rect 76140 -950 76200 -880
rect 76480 -950 76540 -880
rect 76820 -950 76880 -880
rect 77160 -950 77220 -880
rect 77500 -950 77560 -880
rect 77840 -950 77900 -880
rect 78180 -950 78240 -880
rect 78520 -950 78580 -880
rect 78860 -950 78920 -880
rect 79200 -950 79260 -880
rect 79540 -950 79600 -880
rect 79880 -950 79940 -880
rect 80220 -950 80280 -880
rect 80560 -950 80620 -880
rect 80900 -950 80960 -880
rect 81240 -950 81300 -880
rect 81580 -950 81640 -880
rect 81920 -950 81980 -880
rect 82260 -950 82320 -880
rect 82600 -950 82660 -880
rect 82940 -950 83000 -880
rect 83280 -950 83340 -880
rect 83620 -950 83680 -880
rect 83960 -950 84020 -880
rect 84300 -950 84360 -880
rect 84640 -950 84700 -880
rect 84980 -950 85040 -880
rect 85320 -950 85380 -880
rect 85660 -950 85720 -880
rect 86000 -950 86060 -880
rect 86340 -950 86400 -880
rect 86680 -950 86740 -880
rect 87020 -950 87080 -880
rect 150 -1160 210 -1100
rect 1510 -1160 1570 -1100
rect 2870 -1160 2930 -1100
rect 4230 -1160 4290 -1100
rect 5590 -1160 5650 -1100
rect 6950 -1160 7010 -1100
rect 8310 -1160 8370 -1100
rect 9670 -1160 9730 -1100
rect 11030 -1160 11090 -1100
rect 12390 -1160 12450 -1100
rect 13750 -1160 13810 -1100
rect 15110 -1160 15170 -1100
rect 16470 -1160 16530 -1100
rect 17830 -1160 17890 -1100
rect 19190 -1160 19250 -1100
rect 20550 -1160 20610 -1100
rect 21910 -1160 21970 -1100
rect 23270 -1160 23330 -1100
rect 24630 -1160 24690 -1100
rect 25990 -1160 26050 -1100
rect 27350 -1160 27410 -1100
rect 28710 -1160 28770 -1100
rect 30070 -1160 30130 -1100
rect 31430 -1160 31490 -1100
rect 32790 -1160 32850 -1100
rect 34150 -1160 34210 -1100
rect 35510 -1160 35570 -1100
rect 36870 -1160 36930 -1100
rect 38230 -1160 38290 -1100
rect 39590 -1160 39650 -1100
rect 40950 -1160 41010 -1100
rect 42310 -1160 42370 -1100
rect 43670 -1160 43730 -1100
rect 45030 -1160 45090 -1100
rect 46390 -1160 46450 -1100
rect 47750 -1160 47810 -1100
rect 49110 -1160 49170 -1100
rect 50470 -1160 50530 -1100
rect 51830 -1160 51890 -1100
rect 53190 -1160 53250 -1100
rect 54550 -1160 54610 -1100
rect 55910 -1160 55970 -1100
rect 57270 -1160 57330 -1100
rect 58630 -1160 58690 -1100
rect 59990 -1160 60050 -1100
rect 61350 -1160 61410 -1100
rect 62710 -1160 62770 -1100
rect 64070 -1160 64130 -1100
rect 65430 -1160 65490 -1100
rect 66790 -1160 66850 -1100
rect 68150 -1160 68210 -1100
rect 69510 -1160 69570 -1100
rect 70870 -1160 70930 -1100
rect 72230 -1160 72290 -1100
rect 73590 -1160 73650 -1100
rect 74950 -1160 75010 -1100
rect 76310 -1160 76370 -1100
rect 77670 -1160 77730 -1100
rect 79030 -1160 79090 -1100
rect 80390 -1160 80450 -1100
rect 81750 -1160 81810 -1100
rect 83110 -1160 83170 -1100
rect 84470 -1160 84530 -1100
rect 85830 -1160 85890 -1100
rect 150 -1360 210 -1300
rect 1510 -1360 1570 -1300
rect 2870 -1360 2930 -1300
rect 4230 -1360 4290 -1300
rect 5590 -1360 5650 -1300
rect 6950 -1360 7010 -1300
rect 8310 -1360 8370 -1300
rect 9670 -1360 9730 -1300
rect 11030 -1360 11090 -1300
rect 12390 -1360 12450 -1300
rect 13750 -1360 13810 -1300
rect 15110 -1360 15170 -1300
rect 16470 -1360 16530 -1300
rect 17830 -1360 17890 -1300
rect 19190 -1360 19250 -1300
rect 20550 -1360 20610 -1300
rect 21910 -1360 21970 -1300
rect 23270 -1360 23330 -1300
rect 24630 -1360 24690 -1300
rect 25990 -1360 26050 -1300
rect 27350 -1360 27410 -1300
rect 28710 -1360 28770 -1300
rect 30070 -1360 30130 -1300
rect 31430 -1360 31490 -1300
rect 32790 -1360 32850 -1300
rect 34150 -1360 34210 -1300
rect 35510 -1360 35570 -1300
rect 36870 -1360 36930 -1300
rect 38230 -1360 38290 -1300
rect 39590 -1360 39650 -1300
rect 40950 -1360 41010 -1300
rect 42310 -1360 42370 -1300
rect 43670 -1360 43730 -1300
rect 45030 -1360 45090 -1300
rect 46390 -1360 46450 -1300
rect 47750 -1360 47810 -1300
rect 49110 -1360 49170 -1300
rect 50470 -1360 50530 -1300
rect 51830 -1360 51890 -1300
rect 53190 -1360 53250 -1300
rect 54550 -1360 54610 -1300
rect 55910 -1360 55970 -1300
rect 57270 -1360 57330 -1300
rect 58630 -1360 58690 -1300
rect 59990 -1360 60050 -1300
rect 61350 -1360 61410 -1300
rect 62710 -1360 62770 -1300
rect 64070 -1360 64130 -1300
rect 65430 -1360 65490 -1300
rect 66790 -1360 66850 -1300
rect 68150 -1360 68210 -1300
rect 69510 -1360 69570 -1300
rect 70870 -1360 70930 -1300
rect 72230 -1360 72290 -1300
rect 73590 -1360 73650 -1300
rect 74950 -1360 75010 -1300
rect 76310 -1360 76370 -1300
rect 77670 -1360 77730 -1300
rect 79030 -1360 79090 -1300
rect 80390 -1360 80450 -1300
rect 81750 -1360 81810 -1300
rect 83110 -1360 83170 -1300
rect 84470 -1360 84530 -1300
rect 85830 -1360 85890 -1300
rect 830 -1540 910 -1470
rect 5000 -1540 5080 -1470
rect 9030 -1540 9110 -1470
rect 13060 -1540 13140 -1470
rect 17100 -1540 17180 -1470
rect 21200 -1540 21280 -1470
rect 25310 -1540 25390 -1470
rect 29410 -1540 29490 -1470
rect 33440 -1540 33520 -1470
rect 37550 -1540 37630 -1470
rect 41650 -1540 41730 -1470
rect 47100 -1540 47180 -1470
rect 51180 -1540 51260 -1470
rect 55290 -1540 55370 -1470
rect 59320 -1540 59400 -1470
rect 63420 -1540 63500 -1470
rect 67530 -1540 67610 -1470
rect 71560 -1540 71640 -1470
rect 75810 -1540 75890 -1470
rect 79770 -1540 79850 -1470
rect 83950 -1540 84030 -1470
rect 86508 -1544 86588 -1474
<< metal3 >>
rect 1280 710 1410 730
rect 1280 650 1300 710
rect 1390 650 1410 710
rect -20 620 140 630
rect -20 530 0 620
rect 120 530 140 620
rect 730 590 930 620
rect -20 520 140 530
rect 400 570 560 580
rect 10 410 110 520
rect 400 480 420 570
rect 540 480 560 570
rect 730 520 790 590
rect 870 520 930 590
rect 730 490 930 520
rect 1080 570 1200 580
rect 400 470 560 480
rect 1080 480 1090 570
rect 1190 480 1200 570
rect 1080 470 1200 480
rect 10 350 30 410
rect 90 350 110 410
rect 10 330 110 350
rect 430 410 530 470
rect 430 350 450 410
rect 510 350 530 410
rect 430 330 530 350
rect 1110 430 1200 470
rect 1110 410 1210 430
rect 1110 350 1130 410
rect 1190 350 1210 410
rect 1110 330 1210 350
rect 590 210 710 220
rect 590 120 610 210
rect 690 120 710 210
rect 590 110 710 120
rect 930 210 1050 220
rect 930 120 950 210
rect 1030 120 1050 210
rect 930 110 1050 120
rect 1280 210 1410 650
rect 6370 690 6510 710
rect 6370 630 6390 690
rect 6490 630 6510 690
rect 2110 590 2310 620
rect 1470 570 1630 580
rect 1470 480 1490 570
rect 1610 480 1630 570
rect 2110 520 2170 590
rect 2250 520 2310 590
rect 3490 590 3690 620
rect 2110 490 2310 520
rect 2830 570 2990 580
rect 1470 470 1630 480
rect 2830 480 2850 570
rect 2970 480 2990 570
rect 3490 520 3550 590
rect 3630 520 3690 590
rect 5150 590 5350 620
rect 6370 610 6510 630
rect 3490 490 3690 520
rect 4190 570 4350 580
rect 2830 470 2990 480
rect 4190 480 4210 570
rect 4330 480 4350 570
rect 4190 470 4350 480
rect 4490 570 4650 580
rect 4490 480 4510 570
rect 4630 480 4650 570
rect 5150 520 5210 590
rect 5290 520 5350 590
rect 5150 490 5350 520
rect 5850 570 6010 580
rect 4490 470 4650 480
rect 5850 480 5870 570
rect 5990 480 6010 570
rect 5850 470 6010 480
rect 1500 410 1600 470
rect 1500 350 1520 410
rect 1580 350 1600 410
rect 1500 330 1600 350
rect 2860 410 2960 470
rect 2860 350 2880 410
rect 2940 350 2960 410
rect 2860 330 2960 350
rect 4220 410 4320 470
rect 4220 350 4240 410
rect 4300 350 4320 410
rect 4220 330 4320 350
rect 4520 410 4620 470
rect 4520 350 4540 410
rect 4600 350 4620 410
rect 4520 330 4620 350
rect 5880 410 5980 470
rect 5880 350 5900 410
rect 5960 350 5980 410
rect 5880 330 5980 350
rect 1280 120 1290 210
rect 1400 120 1410 210
rect 430 80 530 100
rect 430 20 450 80
rect 510 20 530 80
rect 10 -60 110 -40
rect 10 -120 30 -60
rect 90 -120 110 -60
rect 10 -140 110 -120
rect 30 -250 90 -140
rect -40 -270 270 -250
rect 430 -260 530 20
rect 1110 80 1210 100
rect 1110 20 1130 80
rect 1190 20 1210 80
rect 1110 -260 1210 20
rect 1280 -50 1410 120
rect 1660 210 1780 220
rect 1660 120 1680 210
rect 1760 120 1780 210
rect 1660 110 1780 120
rect 2000 210 2120 220
rect 2000 120 2020 210
rect 2100 120 2120 210
rect 2000 110 2120 120
rect 2340 210 2460 220
rect 2340 120 2360 210
rect 2440 120 2460 210
rect 2340 110 2460 120
rect 2680 210 2800 220
rect 2680 120 2700 210
rect 2780 120 2800 210
rect 2680 110 2800 120
rect 3020 210 3140 220
rect 3020 120 3040 210
rect 3120 120 3140 210
rect 3020 110 3140 120
rect 3360 210 3480 220
rect 3360 120 3380 210
rect 3460 120 3480 210
rect 3360 110 3480 120
rect 3700 210 3820 220
rect 3700 120 3720 210
rect 3800 120 3820 210
rect 3700 110 3820 120
rect 4040 210 4160 220
rect 4040 120 4060 210
rect 4140 120 4160 210
rect 4040 110 4160 120
rect 4360 210 4490 230
rect 6390 220 6490 610
rect 7980 590 8180 620
rect 7210 570 7370 580
rect 7210 480 7230 570
rect 7350 480 7370 570
rect 7980 520 8040 590
rect 8120 520 8180 590
rect 10740 590 10940 620
rect 7980 490 8180 520
rect 8570 570 8730 580
rect 7210 470 7370 480
rect 8570 480 8590 570
rect 8710 480 8730 570
rect 8570 470 8730 480
rect 9930 570 10090 580
rect 9930 480 9950 570
rect 10070 480 10090 570
rect 10740 520 10800 590
rect 10880 520 10940 590
rect 13370 590 13570 620
rect 10740 490 10940 520
rect 11290 570 11450 580
rect 9930 470 10090 480
rect 11290 480 11310 570
rect 11430 480 11450 570
rect 11290 470 11450 480
rect 12650 570 12810 580
rect 12650 480 12670 570
rect 12790 480 12810 570
rect 13370 520 13430 590
rect 13510 520 13570 590
rect 16410 590 16610 620
rect 13370 490 13570 520
rect 14010 570 14170 580
rect 12650 470 12810 480
rect 14010 480 14030 570
rect 14150 480 14170 570
rect 14010 470 14170 480
rect 15370 570 15530 580
rect 15370 480 15390 570
rect 15510 480 15530 570
rect 15370 470 15530 480
rect 15670 570 15830 580
rect 15670 480 15690 570
rect 15810 480 15830 570
rect 16410 520 16470 590
rect 16550 520 16610 590
rect 20480 590 20680 620
rect 16410 490 16610 520
rect 17030 570 17190 580
rect 15670 470 15830 480
rect 17030 480 17050 570
rect 17170 480 17190 570
rect 17030 470 17190 480
rect 18390 570 18550 580
rect 18390 480 18410 570
rect 18530 480 18550 570
rect 18390 470 18550 480
rect 19750 570 19910 580
rect 19750 480 19770 570
rect 19890 480 19910 570
rect 20480 520 20540 590
rect 20620 520 20680 590
rect 24620 590 24820 620
rect 20480 490 20680 520
rect 21110 570 21270 580
rect 19750 470 19910 480
rect 21110 480 21130 570
rect 21250 480 21270 570
rect 21110 470 21270 480
rect 22470 570 22630 580
rect 22470 480 22490 570
rect 22610 480 22630 570
rect 22470 470 22630 480
rect 23830 570 23990 580
rect 23830 480 23850 570
rect 23970 480 23990 570
rect 24620 520 24680 590
rect 24760 520 24820 590
rect 28700 590 28900 620
rect 24620 490 24820 520
rect 25190 570 25350 580
rect 23830 470 23990 480
rect 25190 480 25210 570
rect 25330 480 25350 570
rect 25190 470 25350 480
rect 26550 570 26710 580
rect 26550 480 26570 570
rect 26690 480 26710 570
rect 26550 470 26710 480
rect 27910 570 28070 580
rect 27910 480 27930 570
rect 28050 480 28070 570
rect 28700 520 28760 590
rect 28840 520 28900 590
rect 32850 590 33050 620
rect 28700 490 28900 520
rect 29270 570 29430 580
rect 27910 470 28070 480
rect 29270 480 29290 570
rect 29410 480 29430 570
rect 29270 470 29430 480
rect 30630 570 30790 580
rect 30630 480 30650 570
rect 30770 480 30790 570
rect 30630 470 30790 480
rect 31990 570 32150 580
rect 31990 480 32010 570
rect 32130 480 32150 570
rect 32850 520 32910 590
rect 32990 520 33050 590
rect 36720 590 36920 620
rect 32850 490 33050 520
rect 33350 570 33510 580
rect 31990 470 32150 480
rect 33350 480 33370 570
rect 33490 480 33510 570
rect 33350 470 33510 480
rect 34710 570 34870 580
rect 34710 480 34730 570
rect 34850 480 34870 570
rect 34710 470 34870 480
rect 36070 570 36230 580
rect 36070 480 36090 570
rect 36210 480 36230 570
rect 36720 520 36780 590
rect 36860 520 36920 590
rect 40860 590 41060 620
rect 36720 490 36920 520
rect 37430 570 37590 580
rect 36070 470 36230 480
rect 37430 480 37450 570
rect 37570 480 37590 570
rect 37430 470 37590 480
rect 38790 570 38950 580
rect 38790 480 38810 570
rect 38930 480 38950 570
rect 38790 470 38950 480
rect 40150 570 40310 580
rect 40150 480 40170 570
rect 40290 480 40310 570
rect 40860 520 40920 590
rect 41000 520 41060 590
rect 44850 590 45050 620
rect 40860 490 41060 520
rect 41510 570 41670 580
rect 40150 470 40310 480
rect 41510 480 41530 570
rect 41650 480 41670 570
rect 41510 470 41670 480
rect 42870 570 43030 580
rect 42870 480 42890 570
rect 43010 480 43030 570
rect 42870 470 43030 480
rect 44230 570 44390 580
rect 44230 480 44250 570
rect 44370 480 44390 570
rect 44850 520 44910 590
rect 44990 520 45050 590
rect 48930 590 49130 620
rect 44850 490 45050 520
rect 45590 570 45750 580
rect 44230 470 44390 480
rect 45590 480 45610 570
rect 45730 480 45750 570
rect 45590 470 45750 480
rect 46950 570 47110 580
rect 46950 480 46970 570
rect 47090 480 47110 570
rect 46950 470 47110 480
rect 48310 570 48470 580
rect 48310 480 48330 570
rect 48450 480 48470 570
rect 48930 520 48990 590
rect 49070 520 49130 590
rect 53020 590 53220 620
rect 48930 490 49130 520
rect 49670 570 49830 580
rect 48310 470 48470 480
rect 49670 480 49690 570
rect 49810 480 49830 570
rect 49670 470 49830 480
rect 51030 570 51190 580
rect 51030 480 51050 570
rect 51170 480 51190 570
rect 51030 470 51190 480
rect 52390 570 52550 580
rect 52390 480 52410 570
rect 52530 480 52550 570
rect 53020 520 53080 590
rect 53160 520 53220 590
rect 57180 590 57380 620
rect 53020 490 53220 520
rect 53750 570 53910 580
rect 52390 470 52550 480
rect 53750 480 53770 570
rect 53890 480 53910 570
rect 53750 470 53910 480
rect 55110 570 55270 580
rect 55110 480 55130 570
rect 55250 480 55270 570
rect 55110 470 55270 480
rect 56470 570 56630 580
rect 56470 480 56490 570
rect 56610 480 56630 570
rect 57180 520 57240 590
rect 57320 520 57380 590
rect 57180 490 57380 520
rect 57830 570 57990 580
rect 56470 470 56630 480
rect 57830 480 57850 570
rect 57970 480 57990 570
rect 57830 470 57990 480
rect 59190 570 59340 580
rect 59190 480 59210 570
rect 59330 480 59340 570
rect 59190 470 59340 480
rect 7240 410 7340 470
rect 7240 350 7260 410
rect 7320 350 7340 410
rect 7240 330 7340 350
rect 8600 410 8700 470
rect 8600 350 8620 410
rect 8680 350 8700 410
rect 8600 330 8700 350
rect 9960 410 10060 470
rect 9960 350 9980 410
rect 10040 350 10060 410
rect 9960 330 10060 350
rect 11320 410 11420 470
rect 11320 350 11340 410
rect 11400 350 11420 410
rect 11320 330 11420 350
rect 12680 410 12780 470
rect 12680 350 12700 410
rect 12760 350 12780 410
rect 12680 330 12780 350
rect 14040 410 14140 470
rect 14040 350 14060 410
rect 14120 350 14140 410
rect 14040 330 14140 350
rect 15400 410 15500 470
rect 15400 350 15420 410
rect 15480 350 15500 410
rect 15400 330 15500 350
rect 15700 410 15800 470
rect 15700 350 15720 410
rect 15780 350 15800 410
rect 15700 330 15800 350
rect 17060 410 17160 470
rect 17060 350 17080 410
rect 17140 350 17160 410
rect 17060 330 17160 350
rect 18420 410 18520 470
rect 18420 350 18440 410
rect 18500 350 18520 410
rect 18420 330 18520 350
rect 19780 410 19880 470
rect 19780 350 19800 410
rect 19860 350 19880 410
rect 19780 330 19880 350
rect 21140 410 21240 470
rect 21140 350 21160 410
rect 21220 350 21240 410
rect 21140 330 21240 350
rect 22500 410 22600 470
rect 22500 350 22520 410
rect 22580 350 22600 410
rect 22500 330 22600 350
rect 23860 410 23960 470
rect 23860 350 23880 410
rect 23940 350 23960 410
rect 23860 330 23960 350
rect 25220 410 25320 470
rect 25220 350 25240 410
rect 25300 350 25320 410
rect 25220 330 25320 350
rect 26580 410 26680 470
rect 26580 350 26600 410
rect 26660 350 26680 410
rect 26580 330 26680 350
rect 27940 410 28040 470
rect 27940 350 27960 410
rect 28020 350 28040 410
rect 27940 330 28040 350
rect 29300 410 29400 470
rect 29300 350 29320 410
rect 29380 350 29400 410
rect 29300 330 29400 350
rect 30660 410 30760 470
rect 30660 350 30680 410
rect 30740 350 30760 410
rect 30660 330 30760 350
rect 32020 410 32120 470
rect 32020 350 32040 410
rect 32100 350 32120 410
rect 32020 330 32120 350
rect 33380 410 33480 470
rect 33380 350 33400 410
rect 33460 350 33480 410
rect 33380 330 33480 350
rect 34740 410 34840 470
rect 34740 350 34760 410
rect 34820 350 34840 410
rect 34740 330 34840 350
rect 36100 410 36200 470
rect 36100 350 36120 410
rect 36180 350 36200 410
rect 36100 330 36200 350
rect 37460 410 37560 470
rect 37460 350 37480 410
rect 37540 350 37560 410
rect 37460 330 37560 350
rect 38820 410 38920 470
rect 38820 350 38840 410
rect 38900 350 38920 410
rect 38820 330 38920 350
rect 40180 410 40280 470
rect 40180 350 40200 410
rect 40260 350 40280 410
rect 40180 330 40280 350
rect 41540 410 41640 470
rect 41540 350 41560 410
rect 41620 350 41640 410
rect 41540 330 41640 350
rect 42900 410 43000 470
rect 42900 350 42920 410
rect 42980 350 43000 410
rect 42900 330 43000 350
rect 44260 410 44360 470
rect 44260 350 44280 410
rect 44340 350 44360 410
rect 44260 330 44360 350
rect 45620 410 45720 470
rect 45620 350 45640 410
rect 45700 350 45720 410
rect 45620 330 45720 350
rect 46980 410 47080 470
rect 46980 350 47000 410
rect 47060 350 47080 410
rect 46980 330 47080 350
rect 48340 410 48440 470
rect 48340 350 48360 410
rect 48420 350 48440 410
rect 48340 330 48440 350
rect 49700 410 49800 470
rect 49700 350 49720 410
rect 49780 350 49800 410
rect 49700 330 49800 350
rect 51060 410 51160 470
rect 51060 350 51080 410
rect 51140 350 51160 410
rect 51060 330 51160 350
rect 52420 410 52520 470
rect 52420 350 52440 410
rect 52500 350 52520 410
rect 52420 330 52520 350
rect 53780 410 53880 470
rect 53780 350 53800 410
rect 53860 350 53880 410
rect 53780 330 53880 350
rect 55140 410 55240 470
rect 55140 350 55160 410
rect 55220 350 55240 410
rect 55140 330 55240 350
rect 56500 410 56600 470
rect 56500 350 56520 410
rect 56580 350 56600 410
rect 56500 330 56600 350
rect 57860 410 57960 470
rect 57860 350 57880 410
rect 57940 350 57960 410
rect 57860 330 57960 350
rect 59220 410 59320 470
rect 59220 350 59240 410
rect 59300 350 59320 410
rect 59220 330 59320 350
rect 4360 120 4370 210
rect 4480 120 4490 210
rect 1280 -130 1300 -50
rect 1400 -130 1410 -50
rect 1280 -160 1410 -130
rect 1500 80 1600 100
rect 1500 20 1520 80
rect 1580 20 1600 80
rect 1500 -260 1600 20
rect 2860 80 2960 100
rect 2860 20 2880 80
rect 2940 20 2960 80
rect 2860 0 2960 20
rect 2070 -260 2400 -240
rect 2880 -260 2940 0
rect 4360 -50 4490 120
rect 4680 210 4800 220
rect 4680 120 4700 210
rect 4780 120 4800 210
rect 4680 110 4800 120
rect 5020 210 5140 220
rect 5020 120 5040 210
rect 5120 120 5140 210
rect 5020 110 5140 120
rect 5360 210 5480 220
rect 5360 120 5380 210
rect 5460 120 5480 210
rect 5360 110 5480 120
rect 5700 210 5820 220
rect 5700 120 5720 210
rect 5800 120 5820 210
rect 5700 110 5820 120
rect 6040 210 6160 220
rect 6040 120 6060 210
rect 6140 120 6160 210
rect 6040 110 6160 120
rect 6380 210 6500 220
rect 6380 120 6400 210
rect 6480 120 6500 210
rect 6380 110 6500 120
rect 6720 210 6840 220
rect 6720 120 6740 210
rect 6820 120 6840 210
rect 6720 110 6840 120
rect 7060 210 7180 220
rect 7060 120 7080 210
rect 7160 120 7180 210
rect 7060 110 7180 120
rect 7400 210 7520 220
rect 7400 120 7420 210
rect 7500 120 7520 210
rect 7400 110 7520 120
rect 7740 210 7860 220
rect 7740 120 7760 210
rect 7840 120 7860 210
rect 7740 110 7860 120
rect 8080 210 8200 220
rect 8080 120 8100 210
rect 8180 120 8200 210
rect 8080 110 8200 120
rect 8420 210 8540 220
rect 8420 120 8440 210
rect 8520 120 8540 210
rect 8420 110 8540 120
rect 8760 210 8880 220
rect 8760 120 8780 210
rect 8860 120 8880 210
rect 8760 110 8880 120
rect 9100 210 9220 220
rect 9100 120 9120 210
rect 9200 120 9220 210
rect 9100 110 9220 120
rect 9440 210 9560 220
rect 9440 120 9460 210
rect 9540 120 9560 210
rect 9440 110 9560 120
rect 9780 210 9900 220
rect 9780 120 9800 210
rect 9880 120 9900 210
rect 9780 110 9900 120
rect 10120 210 10240 220
rect 10120 120 10140 210
rect 10220 120 10240 210
rect 10120 110 10240 120
rect 10460 210 10580 220
rect 10460 120 10480 210
rect 10560 120 10580 210
rect 10460 110 10580 120
rect 10800 210 10920 220
rect 10800 120 10820 210
rect 10900 120 10920 210
rect 10800 110 10920 120
rect 11140 210 11260 220
rect 11140 120 11160 210
rect 11240 120 11260 210
rect 11140 110 11260 120
rect 11480 210 11600 220
rect 11480 120 11500 210
rect 11580 120 11600 210
rect 11480 110 11600 120
rect 11820 210 11940 220
rect 11820 120 11840 210
rect 11920 120 11940 210
rect 11820 110 11940 120
rect 12160 210 12280 220
rect 12160 120 12180 210
rect 12260 120 12280 210
rect 12160 110 12280 120
rect 12500 210 12620 220
rect 12500 120 12520 210
rect 12600 120 12620 210
rect 12500 110 12620 120
rect 12840 210 12960 220
rect 12840 120 12860 210
rect 12940 120 12960 210
rect 12840 110 12960 120
rect 13180 210 13300 220
rect 13180 120 13200 210
rect 13280 120 13300 210
rect 13180 110 13300 120
rect 13520 210 13640 220
rect 13520 120 13540 210
rect 13620 120 13640 210
rect 13520 110 13640 120
rect 13860 210 13980 220
rect 13860 120 13880 210
rect 13960 120 13980 210
rect 13860 110 13980 120
rect 14200 210 14320 220
rect 14200 120 14220 210
rect 14300 120 14320 210
rect 14200 110 14320 120
rect 14540 210 14660 220
rect 14540 120 14560 210
rect 14640 120 14660 210
rect 14540 110 14660 120
rect 14880 210 15000 220
rect 14880 120 14900 210
rect 14980 120 15000 210
rect 14880 110 15000 120
rect 15220 210 15340 220
rect 15220 120 15240 210
rect 15320 120 15340 210
rect 15220 110 15340 120
rect 15540 210 15670 230
rect 15540 120 15550 210
rect 15660 120 15670 210
rect 4860 80 4960 100
rect 4860 20 4880 80
rect 4940 20 4960 80
rect 4860 0 4960 20
rect 6220 80 6320 100
rect 6220 20 6240 80
rect 6300 20 6320 80
rect 6220 0 6320 20
rect 7240 80 7340 100
rect 7240 20 7260 80
rect 7320 20 7340 80
rect 7240 0 7340 20
rect 8600 80 8700 100
rect 8600 20 8620 80
rect 8680 20 8700 80
rect 8600 0 8700 20
rect 9960 80 10060 100
rect 9960 20 9980 80
rect 10040 20 10060 80
rect 9960 0 10060 20
rect 10980 80 11080 100
rect 10980 20 11000 80
rect 11060 20 11080 80
rect 10980 0 11080 20
rect 4360 -130 4380 -50
rect 4480 -130 4490 -50
rect 4360 -140 4490 -130
rect 4880 -250 4940 0
rect 4570 -260 4630 -250
rect -40 -370 0 -270
rect 100 -370 130 -270
rect 230 -370 270 -270
rect -40 -400 270 -370
rect 390 -280 570 -260
rect 390 -380 430 -280
rect 530 -380 570 -280
rect 390 -400 570 -380
rect 1070 -280 1250 -260
rect 1070 -380 1110 -280
rect 1210 -380 1250 -280
rect 1070 -400 1250 -380
rect 1450 -270 1630 -260
rect 1450 -370 1490 -270
rect 1590 -370 1630 -270
rect 1450 -390 1630 -370
rect 2070 -390 2120 -260
rect 2350 -390 2400 -260
rect 130 -670 230 -400
rect 130 -730 150 -670
rect 210 -730 230 -670
rect 130 -750 230 -730
rect 1490 -670 1590 -390
rect 2070 -410 2400 -390
rect 2820 -280 3000 -260
rect 2820 -380 2860 -280
rect 2960 -380 3000 -280
rect 2820 -400 3000 -380
rect 4510 -280 4690 -260
rect 4510 -380 4550 -280
rect 4650 -380 4690 -280
rect 4510 -400 4690 -380
rect 4820 -270 5000 -250
rect 4820 -370 4860 -270
rect 4960 -370 5000 -270
rect 4820 -390 5000 -370
rect 5088 -268 5418 -248
rect 6240 -250 6300 0
rect 4870 -400 4930 -390
rect 5088 -398 5138 -268
rect 5368 -398 5418 -268
rect 5870 -270 6050 -250
rect 5870 -370 5910 -270
rect 6010 -370 6050 -270
rect 5870 -390 6050 -370
rect 6180 -270 6360 -250
rect 6180 -370 6220 -270
rect 6320 -370 6360 -270
rect 6180 -390 6360 -370
rect 6890 -270 7070 -250
rect 7260 -260 7320 0
rect 6890 -370 6930 -270
rect 7030 -370 7070 -270
rect 6890 -390 7070 -370
rect 7200 -280 7380 -260
rect 7200 -380 7240 -280
rect 7340 -380 7380 -280
rect 2870 -650 2930 -400
rect 4560 -410 4640 -400
rect 4570 -650 4630 -410
rect 5088 -418 5418 -398
rect 5930 -650 5990 -390
rect 6950 -650 7010 -390
rect 7200 -400 7380 -380
rect 7574 -268 7904 -248
rect 8620 -250 8680 0
rect 8310 -260 8370 -250
rect 7574 -398 7624 -268
rect 7854 -398 7904 -268
rect 7574 -418 7904 -398
rect 8250 -280 8430 -260
rect 8250 -380 8290 -280
rect 8390 -380 8430 -280
rect 8250 -400 8430 -380
rect 8560 -270 8740 -250
rect 8560 -370 8600 -270
rect 8700 -370 8740 -270
rect 8560 -390 8740 -370
rect 8994 -268 9324 -248
rect 9980 -250 10040 0
rect 8610 -400 8670 -390
rect 8994 -398 9044 -268
rect 9274 -398 9324 -268
rect 9610 -270 9790 -250
rect 9610 -370 9650 -270
rect 9750 -370 9790 -270
rect 9610 -390 9790 -370
rect 9920 -270 10100 -250
rect 9920 -370 9960 -270
rect 10060 -370 10100 -270
rect 9920 -390 10100 -370
rect 10630 -270 10810 -250
rect 11000 -260 11060 0
rect 15540 -50 15670 120
rect 15860 210 15980 220
rect 15860 120 15880 210
rect 15960 120 15980 210
rect 15860 110 15980 120
rect 16200 210 16320 220
rect 16200 120 16220 210
rect 16300 120 16320 210
rect 16200 110 16320 120
rect 16540 210 16660 220
rect 16540 120 16560 210
rect 16640 120 16660 210
rect 16540 110 16660 120
rect 16880 210 17000 220
rect 16880 120 16900 210
rect 16980 120 17000 210
rect 16880 110 17000 120
rect 17220 210 17340 220
rect 17220 120 17240 210
rect 17320 120 17340 210
rect 17220 110 17340 120
rect 17560 210 17680 220
rect 17560 120 17580 210
rect 17660 120 17680 210
rect 17560 110 17680 120
rect 17900 210 18020 220
rect 17900 120 17920 210
rect 18000 120 18020 210
rect 17900 110 18020 120
rect 18240 210 18360 220
rect 18240 120 18260 210
rect 18340 120 18360 210
rect 18240 110 18360 120
rect 18580 210 18700 220
rect 18580 120 18600 210
rect 18680 120 18700 210
rect 18580 110 18700 120
rect 18920 210 19040 220
rect 18920 120 18940 210
rect 19020 120 19040 210
rect 18920 110 19040 120
rect 19260 210 19380 220
rect 19260 120 19280 210
rect 19360 120 19380 210
rect 19260 110 19380 120
rect 19600 210 19720 220
rect 19600 120 19620 210
rect 19700 120 19720 210
rect 19600 110 19720 120
rect 19940 210 20060 220
rect 19940 120 19960 210
rect 20040 120 20060 210
rect 19940 110 20060 120
rect 20280 210 20400 220
rect 20280 120 20300 210
rect 20380 120 20400 210
rect 20280 110 20400 120
rect 20620 210 20740 220
rect 20620 120 20640 210
rect 20720 120 20740 210
rect 20620 110 20740 120
rect 20960 210 21080 220
rect 20960 120 20980 210
rect 21060 120 21080 210
rect 20960 110 21080 120
rect 21300 210 21420 220
rect 21300 120 21320 210
rect 21400 120 21420 210
rect 21300 110 21420 120
rect 21640 210 21760 220
rect 21640 120 21660 210
rect 21740 120 21760 210
rect 21640 110 21760 120
rect 21980 210 22100 220
rect 21980 120 22000 210
rect 22080 120 22100 210
rect 21980 110 22100 120
rect 22320 210 22440 220
rect 22320 120 22340 210
rect 22420 120 22440 210
rect 22320 110 22440 120
rect 22660 210 22780 220
rect 22660 120 22680 210
rect 22760 120 22780 210
rect 22660 110 22780 120
rect 23000 210 23120 220
rect 23000 120 23020 210
rect 23100 120 23120 210
rect 23000 110 23120 120
rect 23340 210 23460 220
rect 23340 120 23360 210
rect 23440 120 23460 210
rect 23340 110 23460 120
rect 23680 210 23800 220
rect 23680 120 23700 210
rect 23780 120 23800 210
rect 23680 110 23800 120
rect 24020 210 24140 220
rect 24020 120 24040 210
rect 24120 120 24140 210
rect 24020 110 24140 120
rect 24360 210 24480 220
rect 24360 120 24380 210
rect 24460 120 24480 210
rect 24360 110 24480 120
rect 24700 210 24820 220
rect 24700 120 24720 210
rect 24800 120 24820 210
rect 24700 110 24820 120
rect 25040 210 25160 220
rect 25040 120 25060 210
rect 25140 120 25160 210
rect 25040 110 25160 120
rect 25380 210 25500 220
rect 25380 120 25400 210
rect 25480 120 25500 210
rect 25380 110 25500 120
rect 25720 210 25840 220
rect 25720 120 25740 210
rect 25820 120 25840 210
rect 25720 110 25840 120
rect 26060 210 26180 220
rect 26060 120 26080 210
rect 26160 120 26180 210
rect 26060 110 26180 120
rect 26400 210 26520 220
rect 26400 120 26420 210
rect 26500 120 26520 210
rect 26400 110 26520 120
rect 26740 210 26860 220
rect 26740 120 26760 210
rect 26840 120 26860 210
rect 26740 110 26860 120
rect 27080 210 27200 220
rect 27080 120 27100 210
rect 27180 120 27200 210
rect 27080 110 27200 120
rect 27420 210 27540 220
rect 27420 120 27440 210
rect 27520 120 27540 210
rect 27420 110 27540 120
rect 27760 210 27880 220
rect 27760 120 27780 210
rect 27860 120 27880 210
rect 27760 110 27880 120
rect 28100 210 28220 220
rect 28100 120 28120 210
rect 28200 120 28220 210
rect 28100 110 28220 120
rect 28440 210 28560 220
rect 28440 120 28460 210
rect 28540 120 28560 210
rect 28440 110 28560 120
rect 28780 210 28900 220
rect 28780 120 28800 210
rect 28880 120 28900 210
rect 28780 110 28900 120
rect 29120 210 29240 220
rect 29120 120 29140 210
rect 29220 120 29240 210
rect 29120 110 29240 120
rect 29460 210 29580 220
rect 29460 120 29480 210
rect 29560 120 29580 210
rect 29460 110 29580 120
rect 29800 210 29920 220
rect 29800 120 29820 210
rect 29900 120 29920 210
rect 29800 110 29920 120
rect 30140 210 30260 220
rect 30140 120 30160 210
rect 30240 120 30260 210
rect 30140 110 30260 120
rect 30480 210 30600 220
rect 30480 120 30500 210
rect 30580 120 30600 210
rect 30480 110 30600 120
rect 30820 210 30940 220
rect 30820 120 30840 210
rect 30920 120 30940 210
rect 30820 110 30940 120
rect 31160 210 31280 220
rect 31160 120 31180 210
rect 31260 120 31280 210
rect 31160 110 31280 120
rect 31500 210 31620 220
rect 31500 120 31520 210
rect 31600 120 31620 210
rect 31500 110 31620 120
rect 31840 210 31960 220
rect 31840 120 31860 210
rect 31940 120 31960 210
rect 31840 110 31960 120
rect 32180 210 32300 220
rect 32180 120 32200 210
rect 32280 120 32300 210
rect 32180 110 32300 120
rect 32520 210 32640 220
rect 32520 120 32540 210
rect 32620 120 32640 210
rect 32520 110 32640 120
rect 32860 210 32980 220
rect 32860 120 32880 210
rect 32960 120 32980 210
rect 32860 110 32980 120
rect 33200 210 33320 220
rect 33200 120 33220 210
rect 33300 120 33320 210
rect 33200 110 33320 120
rect 33540 210 33660 220
rect 33540 120 33560 210
rect 33640 120 33660 210
rect 33540 110 33660 120
rect 33880 210 34000 220
rect 33880 120 33900 210
rect 33980 120 34000 210
rect 33880 110 34000 120
rect 34220 210 34340 220
rect 34220 120 34240 210
rect 34320 120 34340 210
rect 34220 110 34340 120
rect 34560 210 34680 220
rect 34560 120 34580 210
rect 34660 120 34680 210
rect 34560 110 34680 120
rect 34900 210 35020 220
rect 34900 120 34920 210
rect 35000 120 35020 210
rect 34900 110 35020 120
rect 35240 210 35360 220
rect 35240 120 35260 210
rect 35340 120 35360 210
rect 35240 110 35360 120
rect 35580 210 35700 220
rect 35580 120 35600 210
rect 35680 120 35700 210
rect 35580 110 35700 120
rect 35920 210 36040 220
rect 35920 120 35940 210
rect 36020 120 36040 210
rect 35920 110 36040 120
rect 36260 210 36380 220
rect 36260 120 36280 210
rect 36360 120 36380 210
rect 36260 110 36380 120
rect 36600 210 36720 220
rect 36600 120 36620 210
rect 36700 120 36720 210
rect 36600 110 36720 120
rect 36940 210 37060 220
rect 36940 120 36960 210
rect 37040 120 37060 210
rect 36940 110 37060 120
rect 37280 210 37400 220
rect 37280 120 37300 210
rect 37380 120 37400 210
rect 37280 110 37400 120
rect 37620 210 37740 220
rect 37620 120 37640 210
rect 37720 120 37740 210
rect 37620 110 37740 120
rect 37960 210 38080 220
rect 37960 120 37980 210
rect 38060 120 38080 210
rect 37960 110 38080 120
rect 38300 210 38420 220
rect 38300 120 38320 210
rect 38400 120 38420 210
rect 38300 110 38420 120
rect 38640 210 38760 220
rect 38640 120 38660 210
rect 38740 120 38760 210
rect 38640 110 38760 120
rect 38980 210 39100 220
rect 38980 120 39000 210
rect 39080 120 39100 210
rect 38980 110 39100 120
rect 39320 210 39440 220
rect 39320 120 39340 210
rect 39420 120 39440 210
rect 39320 110 39440 120
rect 39660 210 39780 220
rect 39660 120 39680 210
rect 39760 120 39780 210
rect 39660 110 39780 120
rect 40000 210 40120 220
rect 40000 120 40020 210
rect 40100 120 40120 210
rect 40000 110 40120 120
rect 40340 210 40460 220
rect 40340 120 40360 210
rect 40440 120 40460 210
rect 40340 110 40460 120
rect 40680 210 40800 220
rect 40680 120 40700 210
rect 40780 120 40800 210
rect 40680 110 40800 120
rect 41020 210 41140 220
rect 41020 120 41040 210
rect 41120 120 41140 210
rect 41020 110 41140 120
rect 41360 210 41480 220
rect 41360 120 41380 210
rect 41460 120 41480 210
rect 41360 110 41480 120
rect 41700 210 41820 220
rect 41700 120 41720 210
rect 41800 120 41820 210
rect 41700 110 41820 120
rect 42040 210 42160 220
rect 42040 120 42060 210
rect 42140 120 42160 210
rect 42040 110 42160 120
rect 42380 210 42500 220
rect 42380 120 42400 210
rect 42480 120 42500 210
rect 42380 110 42500 120
rect 42720 210 42840 220
rect 42720 120 42740 210
rect 42820 120 42840 210
rect 42720 110 42840 120
rect 43060 210 43180 220
rect 43060 120 43080 210
rect 43160 120 43180 210
rect 43060 110 43180 120
rect 43400 210 43520 220
rect 43400 120 43420 210
rect 43500 120 43520 210
rect 43400 110 43520 120
rect 43740 210 43860 220
rect 43740 120 43760 210
rect 43840 120 43860 210
rect 43740 110 43860 120
rect 44080 210 44200 220
rect 44080 120 44100 210
rect 44180 120 44200 210
rect 44080 110 44200 120
rect 44420 210 44540 220
rect 44420 120 44440 210
rect 44520 120 44540 210
rect 44420 110 44540 120
rect 44760 210 44880 220
rect 44760 120 44780 210
rect 44860 120 44880 210
rect 44760 110 44880 120
rect 45100 210 45220 220
rect 45100 120 45120 210
rect 45200 120 45220 210
rect 45100 110 45220 120
rect 45440 210 45560 220
rect 45440 120 45460 210
rect 45540 120 45560 210
rect 45440 110 45560 120
rect 45780 210 45900 220
rect 45780 120 45800 210
rect 45880 120 45900 210
rect 45780 110 45900 120
rect 46120 210 46240 220
rect 46120 120 46140 210
rect 46220 120 46240 210
rect 46120 110 46240 120
rect 46460 210 46580 220
rect 46460 120 46480 210
rect 46560 120 46580 210
rect 46460 110 46580 120
rect 46800 210 46920 220
rect 46800 120 46820 210
rect 46900 120 46920 210
rect 46800 110 46920 120
rect 47140 210 47260 220
rect 47140 120 47160 210
rect 47240 120 47260 210
rect 47140 110 47260 120
rect 47480 210 47600 220
rect 47480 120 47500 210
rect 47580 120 47600 210
rect 47480 110 47600 120
rect 47820 210 47940 220
rect 47820 120 47840 210
rect 47920 120 47940 210
rect 47820 110 47940 120
rect 48160 210 48280 220
rect 48160 120 48180 210
rect 48260 120 48280 210
rect 48160 110 48280 120
rect 48500 210 48620 220
rect 48500 120 48520 210
rect 48600 120 48620 210
rect 48500 110 48620 120
rect 48840 210 48960 220
rect 48840 120 48860 210
rect 48940 120 48960 210
rect 48840 110 48960 120
rect 49180 210 49300 220
rect 49180 120 49200 210
rect 49280 120 49300 210
rect 49180 110 49300 120
rect 49520 210 49640 220
rect 49520 120 49540 210
rect 49620 120 49640 210
rect 49520 110 49640 120
rect 49860 210 49980 220
rect 49860 120 49880 210
rect 49960 120 49980 210
rect 49860 110 49980 120
rect 50200 210 50320 220
rect 50200 120 50220 210
rect 50300 120 50320 210
rect 50200 110 50320 120
rect 50540 210 50660 220
rect 50540 120 50560 210
rect 50640 120 50660 210
rect 50540 110 50660 120
rect 50880 210 51000 220
rect 50880 120 50900 210
rect 50980 120 51000 210
rect 50880 110 51000 120
rect 51220 210 51340 220
rect 51220 120 51240 210
rect 51320 120 51340 210
rect 51220 110 51340 120
rect 51560 210 51680 220
rect 51560 120 51580 210
rect 51660 120 51680 210
rect 51560 110 51680 120
rect 51900 210 52020 220
rect 51900 120 51920 210
rect 52000 120 52020 210
rect 51900 110 52020 120
rect 52240 210 52360 220
rect 52240 120 52260 210
rect 52340 120 52360 210
rect 52240 110 52360 120
rect 52580 210 52700 220
rect 52580 120 52600 210
rect 52680 120 52700 210
rect 52580 110 52700 120
rect 52920 210 53040 220
rect 52920 120 52940 210
rect 53020 120 53040 210
rect 52920 110 53040 120
rect 53260 210 53380 220
rect 53260 120 53280 210
rect 53360 120 53380 210
rect 53260 110 53380 120
rect 53600 210 53720 220
rect 53600 120 53620 210
rect 53700 120 53720 210
rect 53600 110 53720 120
rect 53940 210 54060 220
rect 53940 120 53960 210
rect 54040 120 54060 210
rect 53940 110 54060 120
rect 54280 210 54400 220
rect 54280 120 54300 210
rect 54380 120 54400 210
rect 54280 110 54400 120
rect 54620 210 54740 220
rect 54620 120 54640 210
rect 54720 120 54740 210
rect 54620 110 54740 120
rect 54960 210 55080 220
rect 54960 120 54980 210
rect 55060 120 55080 210
rect 54960 110 55080 120
rect 55300 210 55420 220
rect 55300 120 55320 210
rect 55400 120 55420 210
rect 55300 110 55420 120
rect 55640 210 55760 220
rect 55640 120 55660 210
rect 55740 120 55760 210
rect 55640 110 55760 120
rect 55980 210 56100 220
rect 55980 120 56000 210
rect 56080 120 56100 210
rect 55980 110 56100 120
rect 56320 210 56440 220
rect 56320 120 56340 210
rect 56420 120 56440 210
rect 56320 110 56440 120
rect 56660 210 56780 220
rect 56660 120 56680 210
rect 56760 120 56780 210
rect 56660 110 56780 120
rect 57000 210 57120 220
rect 57000 120 57020 210
rect 57100 120 57120 210
rect 57000 110 57120 120
rect 57340 210 57460 220
rect 57340 120 57360 210
rect 57440 120 57460 210
rect 57340 110 57460 120
rect 57680 210 57800 220
rect 57680 120 57700 210
rect 57780 120 57800 210
rect 57680 110 57800 120
rect 58020 210 58140 220
rect 58020 120 58040 210
rect 58120 120 58140 210
rect 58020 110 58140 120
rect 58360 210 58480 220
rect 58360 120 58380 210
rect 58460 120 58480 210
rect 58360 110 58480 120
rect 58700 210 58820 220
rect 58700 120 58720 210
rect 58800 120 58820 210
rect 58700 110 58820 120
rect 59040 210 59160 220
rect 59040 120 59060 210
rect 59140 120 59160 210
rect 59040 110 59160 120
rect 15540 -130 15560 -50
rect 15660 -130 15670 -50
rect 15540 -140 15670 -130
rect 10630 -370 10670 -270
rect 10770 -370 10810 -270
rect 10630 -390 10810 -370
rect 10940 -280 11120 -260
rect 10940 -380 10980 -280
rect 11080 -380 11120 -280
rect 8300 -410 8380 -400
rect 8310 -650 8370 -410
rect 8994 -418 9324 -398
rect 9670 -650 9730 -390
rect 10690 -650 10750 -390
rect 10940 -400 11120 -380
rect 11690 -270 11830 -250
rect 11990 -260 12090 -220
rect 12670 -260 12770 -220
rect 13060 -260 13160 -220
rect 11790 -370 11830 -270
rect 11690 -390 11830 -370
rect 11950 -280 12130 -260
rect 11950 -380 11990 -280
rect 12090 -380 12130 -280
rect 1490 -730 1510 -670
rect 1570 -730 1590 -670
rect 1490 -750 1590 -730
rect 2850 -670 2950 -650
rect 2850 -730 2870 -670
rect 2930 -730 2950 -670
rect 2850 -750 2950 -730
rect 4550 -670 4650 -650
rect 4550 -730 4570 -670
rect 4630 -730 4650 -670
rect 4550 -750 4650 -730
rect 5910 -670 6010 -650
rect 5910 -730 5930 -670
rect 5990 -730 6010 -670
rect 5910 -750 6010 -730
rect 6930 -670 7030 -650
rect 6930 -730 6950 -670
rect 7010 -730 7030 -670
rect 6930 -750 7030 -730
rect 8290 -670 8390 -650
rect 8290 -730 8310 -670
rect 8370 -730 8390 -670
rect 8290 -750 8390 -730
rect 9650 -670 9750 -650
rect 9650 -730 9670 -670
rect 9730 -730 9750 -670
rect 9650 -750 9750 -730
rect 10670 -670 10770 -650
rect 10670 -730 10690 -670
rect 10750 -730 10770 -670
rect 10670 -750 10770 -730
rect 11690 -670 11790 -390
rect 11950 -400 12130 -380
rect 12630 -280 12810 -260
rect 12630 -380 12670 -280
rect 12770 -380 12810 -280
rect 12630 -400 12810 -380
rect 13010 -270 13190 -260
rect 13010 -370 13050 -270
rect 13150 -370 13190 -270
rect 13010 -390 13190 -370
rect 13618 -264 13948 -244
rect 14440 -260 14500 -220
rect 11690 -730 11710 -670
rect 11770 -730 11790 -670
rect 11690 -750 11790 -730
rect 13050 -670 13150 -390
rect 13618 -394 13668 -264
rect 13898 -394 13948 -264
rect 13618 -414 13948 -394
rect 14380 -280 14560 -260
rect 14380 -380 14420 -280
rect 14520 -380 14560 -280
rect 14380 -400 14560 -380
rect 14430 -650 14490 -400
rect 15870 -450 15970 110
rect 16380 80 16480 100
rect 16380 20 16400 80
rect 16460 20 16480 80
rect 16380 0 16480 20
rect 17740 80 17840 100
rect 17740 20 17760 80
rect 17820 20 17840 80
rect 17740 0 17840 20
rect 18760 80 18860 100
rect 18760 20 18780 80
rect 18840 20 18860 80
rect 18760 0 18860 20
rect 20120 80 20220 100
rect 20120 20 20140 80
rect 20200 20 20220 80
rect 20120 0 20220 20
rect 21480 80 21580 100
rect 21480 20 21500 80
rect 21560 20 21580 80
rect 21480 0 21580 20
rect 22500 80 22600 100
rect 22500 20 22520 80
rect 22580 20 22600 80
rect 22500 0 22600 20
rect 23860 80 23960 100
rect 23860 20 23880 80
rect 23940 20 23960 80
rect 23860 0 23960 20
rect 24540 80 24640 100
rect 24540 20 24560 80
rect 24620 20 24640 80
rect 24540 0 24640 20
rect 28280 80 28380 100
rect 28280 20 28300 80
rect 28360 20 28380 80
rect 28280 0 28380 20
rect 29640 80 29740 100
rect 29640 20 29660 80
rect 29720 20 29740 80
rect 29640 0 29740 20
rect 30660 80 30760 100
rect 30660 20 30680 80
rect 30740 20 30760 80
rect 30660 0 30760 20
rect 16400 -250 16460 0
rect 16130 -260 16190 -250
rect 16070 -280 16250 -260
rect 16070 -380 16110 -280
rect 16210 -380 16250 -280
rect 16070 -400 16250 -380
rect 16340 -270 16520 -250
rect 16340 -370 16380 -270
rect 16480 -370 16520 -270
rect 16340 -390 16520 -370
rect 16818 -264 17148 -244
rect 17760 -250 17820 0
rect 16390 -400 16450 -390
rect 16818 -394 16868 -264
rect 17098 -394 17148 -264
rect 17430 -270 17610 -250
rect 17430 -370 17470 -270
rect 17570 -370 17610 -270
rect 17430 -390 17610 -370
rect 17700 -270 17880 -250
rect 17700 -370 17740 -270
rect 17840 -370 17880 -270
rect 17700 -390 17880 -370
rect 18450 -270 18630 -250
rect 18780 -260 18840 0
rect 20140 -250 20200 0
rect 19870 -260 19930 -250
rect 18450 -370 18490 -270
rect 18590 -370 18630 -270
rect 18450 -390 18630 -370
rect 18720 -280 18900 -260
rect 18720 -380 18760 -280
rect 18860 -380 18900 -280
rect 16120 -410 16200 -400
rect 15850 -460 16010 -450
rect 15850 -520 15930 -460
rect 16000 -520 16010 -460
rect 15850 -610 16010 -520
rect 16130 -650 16190 -410
rect 16818 -414 17148 -394
rect 17490 -650 17550 -390
rect 18510 -650 18570 -390
rect 18720 -400 18900 -380
rect 19810 -280 19990 -260
rect 19810 -380 19850 -280
rect 19950 -380 19990 -280
rect 19810 -400 19990 -380
rect 20080 -270 20260 -250
rect 20080 -370 20120 -270
rect 20220 -370 20260 -270
rect 20080 -390 20260 -370
rect 20374 -264 20704 -244
rect 21500 -250 21560 0
rect 20130 -400 20190 -390
rect 20374 -394 20424 -264
rect 20654 -394 20704 -264
rect 21170 -270 21350 -250
rect 21170 -370 21210 -270
rect 21310 -370 21350 -270
rect 21170 -390 21350 -370
rect 21440 -270 21620 -250
rect 21440 -370 21480 -270
rect 21580 -370 21620 -270
rect 21440 -390 21620 -370
rect 22190 -270 22370 -250
rect 22520 -260 22580 0
rect 23880 -220 23940 0
rect 24560 -220 24620 0
rect 22190 -370 22230 -270
rect 22330 -370 22370 -270
rect 22190 -390 22370 -370
rect 22460 -280 22640 -260
rect 22460 -380 22500 -280
rect 22600 -380 22640 -280
rect 19860 -410 19940 -400
rect 19870 -650 19930 -410
rect 20374 -414 20704 -394
rect 21230 -650 21290 -390
rect 22250 -650 22310 -390
rect 22460 -400 22640 -380
rect 23590 -270 23730 -250
rect 23860 -260 23960 -220
rect 24530 -260 24630 -220
rect 24960 -260 25060 -220
rect 23690 -370 23730 -270
rect 23590 -390 23730 -370
rect 23820 -280 24000 -260
rect 23820 -380 23860 -280
rect 23960 -380 24000 -280
rect 13050 -730 13070 -670
rect 13130 -730 13150 -670
rect 13050 -750 13150 -730
rect 14410 -670 14510 -650
rect 14410 -730 14430 -670
rect 14490 -730 14510 -670
rect 14410 -750 14510 -730
rect 16110 -670 16210 -650
rect 16110 -730 16130 -670
rect 16190 -730 16210 -670
rect 16110 -750 16210 -730
rect 17470 -670 17570 -650
rect 17470 -730 17490 -670
rect 17550 -730 17570 -670
rect 17470 -750 17570 -730
rect 18490 -670 18590 -650
rect 18490 -730 18510 -670
rect 18570 -730 18590 -670
rect 18490 -750 18590 -730
rect 19850 -670 19950 -650
rect 19850 -730 19870 -670
rect 19930 -730 19950 -670
rect 19850 -750 19950 -730
rect 21210 -670 21310 -650
rect 21210 -730 21230 -670
rect 21290 -730 21310 -670
rect 21210 -750 21310 -730
rect 22230 -670 22330 -650
rect 22230 -730 22250 -670
rect 22310 -730 22330 -670
rect 22230 -750 22330 -730
rect 23590 -670 23690 -390
rect 23820 -400 24000 -380
rect 24490 -280 24670 -260
rect 24490 -380 24530 -280
rect 24630 -380 24670 -280
rect 24490 -400 24670 -380
rect 24910 -270 25090 -260
rect 24910 -370 24950 -270
rect 25050 -370 25090 -270
rect 24910 -390 25090 -370
rect 25708 -264 26038 -244
rect 26340 -260 26400 -220
rect 28300 -250 28360 0
rect 28030 -260 28090 -250
rect 23590 -730 23610 -670
rect 23670 -730 23690 -670
rect 23590 -750 23690 -730
rect 24950 -670 25050 -390
rect 25708 -394 25758 -264
rect 25988 -394 26038 -264
rect 25708 -414 26038 -394
rect 26280 -280 26460 -260
rect 26280 -380 26320 -280
rect 26420 -380 26460 -280
rect 26280 -400 26460 -380
rect 27970 -280 28150 -260
rect 27970 -380 28010 -280
rect 28110 -380 28150 -280
rect 27970 -400 28150 -380
rect 28240 -270 28420 -250
rect 28240 -370 28280 -270
rect 28380 -370 28420 -270
rect 28240 -390 28420 -370
rect 28552 -264 28882 -244
rect 29660 -250 29720 0
rect 28290 -400 28350 -390
rect 28552 -394 28602 -264
rect 28832 -394 28882 -264
rect 29330 -270 29510 -250
rect 29330 -370 29370 -270
rect 29470 -370 29510 -270
rect 29330 -390 29510 -370
rect 29600 -270 29780 -250
rect 29600 -370 29640 -270
rect 29740 -370 29780 -270
rect 29600 -390 29780 -370
rect 30350 -270 30530 -250
rect 30680 -260 30740 0
rect 30350 -370 30390 -270
rect 30490 -370 30530 -270
rect 30350 -390 30530 -370
rect 30620 -280 30800 -260
rect 30620 -380 30660 -280
rect 30760 -380 30800 -280
rect 26330 -650 26390 -400
rect 28020 -410 28100 -400
rect 28030 -650 28090 -410
rect 28552 -414 28882 -394
rect 29390 -650 29450 -390
rect 30410 -650 30470 -390
rect 30620 -400 30800 -380
rect 31170 -450 31270 110
rect 32020 80 32120 100
rect 32020 20 32040 80
rect 32100 20 32120 80
rect 32020 0 32120 20
rect 33380 80 33480 100
rect 33380 20 33400 80
rect 33460 20 33480 80
rect 33380 0 33480 20
rect 34400 80 34500 100
rect 34400 20 34420 80
rect 34480 20 34500 80
rect 34400 0 34500 20
rect 35760 80 35860 100
rect 35760 20 35780 80
rect 35840 20 35860 80
rect 35760 0 35860 20
rect 36440 80 36540 100
rect 36440 20 36460 80
rect 36520 20 36540 80
rect 36440 0 36540 20
rect 42560 80 42660 100
rect 42560 20 42580 80
rect 42640 20 42660 80
rect 42560 0 42660 20
rect 44600 80 44700 100
rect 44600 20 44620 80
rect 44680 20 44700 80
rect 44600 0 44700 20
rect 48340 80 48440 100
rect 48340 20 48360 80
rect 48420 20 48440 80
rect 48340 0 48440 20
rect 49700 80 49800 100
rect 49700 20 49720 80
rect 49780 20 49800 80
rect 49700 0 49800 20
rect 50720 80 50820 100
rect 50720 20 50740 80
rect 50800 20 50820 80
rect 50720 0 50820 20
rect 52080 80 52180 100
rect 52080 20 52100 80
rect 52160 20 52180 80
rect 52080 0 52180 20
rect 53440 80 53540 100
rect 53440 20 53460 80
rect 53520 20 53540 80
rect 53440 0 53540 20
rect 55480 80 55580 100
rect 55480 20 55500 80
rect 55560 20 55580 80
rect 55480 0 55580 20
rect 32040 -250 32100 0
rect 31770 -260 31830 -250
rect 31710 -280 31890 -260
rect 31710 -380 31750 -280
rect 31850 -380 31890 -280
rect 31710 -400 31890 -380
rect 31980 -270 32160 -250
rect 31980 -370 32020 -270
rect 32120 -370 32160 -270
rect 31980 -390 32160 -370
rect 32464 -264 32794 -244
rect 33400 -250 33460 0
rect 32030 -400 32090 -390
rect 32464 -394 32514 -264
rect 32744 -394 32794 -264
rect 33070 -270 33250 -250
rect 33070 -370 33110 -270
rect 33210 -370 33250 -270
rect 33070 -390 33250 -370
rect 33340 -270 33520 -250
rect 33340 -370 33380 -270
rect 33480 -370 33520 -270
rect 33340 -390 33520 -370
rect 34090 -270 34270 -250
rect 34420 -260 34480 0
rect 35780 -220 35840 0
rect 36460 -220 36520 0
rect 34090 -370 34130 -270
rect 34230 -370 34270 -270
rect 34090 -390 34270 -370
rect 34360 -280 34540 -260
rect 34360 -380 34400 -280
rect 34500 -380 34540 -280
rect 31760 -410 31840 -400
rect 31150 -460 31310 -450
rect 31150 -520 31230 -460
rect 31300 -520 31310 -460
rect 31150 -610 31310 -520
rect 31770 -650 31830 -410
rect 32464 -414 32794 -394
rect 33130 -650 33190 -390
rect 34150 -650 34210 -390
rect 34360 -400 34540 -380
rect 34620 -264 34950 -244
rect 34620 -394 34670 -264
rect 34900 -394 34950 -264
rect 34620 -414 34950 -394
rect 35490 -270 35630 -250
rect 35760 -260 35860 -220
rect 36430 -260 36530 -220
rect 36860 -260 36960 -220
rect 35590 -370 35630 -270
rect 35490 -390 35630 -370
rect 35720 -280 35900 -260
rect 35720 -380 35760 -280
rect 35860 -380 35900 -280
rect 24950 -730 24970 -670
rect 25030 -730 25050 -670
rect 24950 -750 25050 -730
rect 26310 -670 26410 -650
rect 26310 -730 26330 -670
rect 26390 -730 26410 -670
rect 26310 -750 26410 -730
rect 28010 -670 28110 -650
rect 28010 -730 28030 -670
rect 28090 -730 28110 -670
rect 28010 -750 28110 -730
rect 29370 -670 29470 -650
rect 29370 -730 29390 -670
rect 29450 -730 29470 -670
rect 29370 -750 29470 -730
rect 30390 -670 30490 -650
rect 30390 -730 30410 -670
rect 30470 -730 30490 -670
rect 30390 -750 30490 -730
rect 31750 -670 31850 -650
rect 31750 -730 31770 -670
rect 31830 -730 31850 -670
rect 31750 -750 31850 -730
rect 33110 -670 33210 -650
rect 33110 -730 33130 -670
rect 33190 -730 33210 -670
rect 33110 -750 33210 -730
rect 34130 -670 34230 -650
rect 34130 -730 34150 -670
rect 34210 -730 34230 -670
rect 34130 -750 34230 -730
rect 35490 -670 35590 -390
rect 35720 -400 35900 -380
rect 36390 -280 36570 -260
rect 36390 -380 36430 -280
rect 36530 -380 36570 -280
rect 36390 -400 36570 -380
rect 36810 -270 36990 -260
rect 36810 -370 36850 -270
rect 36950 -370 36990 -270
rect 36810 -390 36990 -370
rect 37442 -264 37772 -244
rect 38240 -260 38300 -220
rect 39930 -260 39990 -250
rect 35490 -730 35510 -670
rect 35570 -730 35590 -670
rect 35490 -750 35590 -730
rect 36850 -670 36950 -390
rect 37442 -394 37492 -264
rect 37722 -394 37772 -264
rect 37442 -414 37772 -394
rect 38180 -280 38360 -260
rect 38180 -380 38220 -280
rect 38320 -380 38360 -280
rect 38180 -400 38360 -380
rect 39870 -280 40050 -260
rect 39870 -380 39910 -280
rect 40010 -380 40050 -280
rect 39870 -400 40050 -380
rect 40642 -264 40972 -244
rect 40642 -394 40692 -264
rect 40922 -394 40972 -264
rect 41230 -270 41410 -250
rect 41230 -370 41270 -270
rect 41370 -370 41410 -270
rect 41230 -390 41410 -370
rect 42250 -270 42430 -250
rect 42580 -260 42640 0
rect 44620 -220 44680 0
rect 43630 -260 43790 -250
rect 44600 -260 44700 -220
rect 42250 -370 42290 -270
rect 42390 -370 42430 -270
rect 42250 -390 42430 -370
rect 42520 -280 42700 -260
rect 42520 -380 42560 -280
rect 42660 -380 42700 -280
rect 38230 -650 38290 -400
rect 39920 -410 40000 -400
rect 39930 -650 39990 -410
rect 40642 -414 40972 -394
rect 41290 -650 41350 -390
rect 42310 -650 42370 -390
rect 42520 -400 42700 -380
rect 43610 -270 43790 -260
rect 43610 -380 43650 -270
rect 43750 -380 43790 -270
rect 43610 -400 43790 -380
rect 44560 -280 44740 -260
rect 44560 -380 44600 -280
rect 44700 -380 44740 -280
rect 44560 -400 44740 -380
rect 44970 -270 45150 -260
rect 44970 -370 45010 -270
rect 45110 -370 45150 -270
rect 44970 -390 45150 -370
rect 45618 -264 45948 -244
rect 48360 -250 48420 0
rect 48090 -260 48150 -250
rect 36850 -730 36870 -670
rect 36930 -730 36950 -670
rect 36850 -750 36950 -730
rect 38210 -670 38310 -650
rect 38210 -730 38230 -670
rect 38290 -730 38310 -670
rect 38210 -750 38310 -730
rect 39910 -670 40010 -650
rect 39910 -730 39930 -670
rect 39990 -730 40010 -670
rect 39910 -750 40010 -730
rect 41270 -670 41370 -650
rect 41270 -730 41290 -670
rect 41350 -730 41370 -670
rect 41270 -750 41370 -730
rect 42290 -670 42390 -650
rect 42290 -730 42310 -670
rect 42370 -730 42390 -670
rect 42290 -750 42390 -730
rect 43650 -670 43750 -400
rect 43650 -730 43670 -670
rect 43730 -730 43750 -670
rect 43650 -750 43750 -730
rect 45010 -670 45110 -390
rect 45618 -394 45668 -264
rect 45898 -394 45948 -264
rect 45618 -414 45948 -394
rect 46340 -280 46520 -260
rect 46340 -380 46380 -280
rect 46480 -380 46520 -280
rect 46340 -400 46520 -380
rect 48030 -280 48210 -260
rect 48030 -380 48070 -280
rect 48170 -380 48210 -280
rect 48030 -400 48210 -380
rect 48300 -270 48480 -250
rect 48300 -370 48340 -270
rect 48440 -370 48480 -270
rect 48300 -390 48480 -370
rect 48818 -264 49148 -244
rect 49720 -250 49780 0
rect 48350 -400 48410 -390
rect 48818 -394 48868 -264
rect 49098 -394 49148 -264
rect 49390 -270 49570 -250
rect 49390 -370 49430 -270
rect 49530 -370 49570 -270
rect 49390 -390 49570 -370
rect 49660 -270 49840 -250
rect 49660 -370 49700 -270
rect 49800 -370 49840 -270
rect 49660 -390 49840 -370
rect 50410 -270 50590 -250
rect 50740 -260 50800 0
rect 50410 -370 50450 -270
rect 50550 -370 50590 -270
rect 50410 -390 50590 -370
rect 50680 -280 50860 -260
rect 50680 -380 50720 -280
rect 50820 -380 50860 -280
rect 46390 -650 46450 -400
rect 48080 -410 48160 -400
rect 48090 -650 48150 -410
rect 48818 -414 49148 -394
rect 49450 -650 49510 -390
rect 50470 -650 50530 -390
rect 50680 -400 50860 -380
rect 50952 -264 51282 -244
rect 52100 -250 52160 0
rect 53460 -250 53520 0
rect 55500 -220 55560 0
rect 51830 -260 51890 -250
rect 50952 -394 51002 -264
rect 51232 -394 51282 -264
rect 50952 -414 51282 -394
rect 51770 -280 51950 -260
rect 51770 -380 51810 -280
rect 51910 -380 51950 -280
rect 51770 -400 51950 -380
rect 52040 -270 52220 -250
rect 52040 -370 52080 -270
rect 52180 -370 52220 -270
rect 52040 -390 52220 -370
rect 53130 -270 53310 -250
rect 53130 -370 53170 -270
rect 53270 -370 53310 -270
rect 53130 -390 53310 -370
rect 53400 -270 53580 -250
rect 53400 -370 53440 -270
rect 53540 -370 53580 -270
rect 53400 -390 53580 -370
rect 54150 -270 54330 -250
rect 54150 -370 54190 -270
rect 54290 -370 54330 -270
rect 54150 -390 54330 -370
rect 54508 -264 54838 -244
rect 52090 -400 52150 -390
rect 51820 -410 51900 -400
rect 51830 -650 51890 -410
rect 53190 -650 53250 -390
rect 54210 -650 54270 -390
rect 54508 -394 54558 -264
rect 54788 -394 54838 -264
rect 54508 -414 54838 -394
rect 55210 -270 55350 -250
rect 55480 -260 55580 -220
rect 56580 -260 56680 -220
rect 55310 -370 55350 -270
rect 55210 -390 55350 -370
rect 55440 -280 55620 -260
rect 55440 -380 55480 -280
rect 55580 -380 55620 -280
rect 45010 -730 45030 -670
rect 45090 -730 45110 -670
rect 45010 -750 45110 -730
rect 46370 -670 46470 -650
rect 46370 -730 46390 -670
rect 46450 -730 46470 -670
rect 46370 -750 46470 -730
rect 48070 -670 48170 -650
rect 48070 -730 48090 -670
rect 48150 -730 48170 -670
rect 48070 -750 48170 -730
rect 49430 -670 49530 -650
rect 49430 -730 49450 -670
rect 49510 -730 49530 -670
rect 49430 -750 49530 -730
rect 50450 -670 50550 -650
rect 50450 -730 50470 -670
rect 50530 -730 50550 -670
rect 50450 -750 50550 -730
rect 51810 -670 51910 -650
rect 51810 -730 51830 -670
rect 51890 -730 51910 -670
rect 51810 -750 51910 -730
rect 53170 -670 53270 -650
rect 53170 -730 53190 -670
rect 53250 -730 53270 -670
rect 53170 -750 53270 -730
rect 54190 -670 54290 -650
rect 54190 -730 54210 -670
rect 54270 -730 54290 -670
rect 54190 -750 54290 -730
rect 55210 -670 55310 -390
rect 55440 -400 55620 -380
rect 56530 -270 56710 -260
rect 56530 -370 56570 -270
rect 56670 -370 56710 -270
rect 56530 -390 56710 -370
rect 57352 -264 57682 -244
rect 57960 -260 58020 -220
rect 55210 -730 55230 -670
rect 55290 -730 55310 -670
rect 55210 -750 55310 -730
rect 56570 -670 56670 -390
rect 57352 -394 57402 -264
rect 57632 -394 57682 -264
rect 57352 -414 57682 -394
rect 57900 -280 58080 -260
rect 57900 -380 57940 -280
rect 58040 -380 58080 -280
rect 57900 -400 58080 -380
rect 57950 -650 58010 -400
rect 59060 -450 59140 110
rect 59650 -260 59710 -250
rect 59590 -280 59770 -260
rect 59590 -380 59630 -280
rect 59730 -380 59770 -280
rect 59590 -400 59770 -380
rect 60950 -270 61130 -250
rect 60950 -370 60990 -270
rect 61090 -370 61130 -270
rect 60950 -390 61130 -370
rect 61264 -264 61594 -244
rect 59640 -410 59720 -400
rect 59030 -460 59190 -450
rect 59030 -520 59110 -460
rect 59180 -520 59190 -460
rect 59030 -610 59190 -520
rect 59650 -650 59710 -410
rect 61010 -650 61070 -390
rect 61264 -394 61314 -264
rect 61544 -394 61594 -264
rect 61970 -270 62150 -250
rect 63390 -260 63450 -250
rect 61970 -370 62010 -270
rect 62110 -370 62150 -270
rect 61970 -390 62150 -370
rect 63330 -280 63510 -260
rect 63330 -380 63370 -280
rect 63470 -380 63510 -280
rect 61264 -414 61594 -394
rect 62030 -650 62090 -390
rect 63330 -400 63510 -380
rect 64108 -264 64438 -244
rect 64108 -394 64158 -264
rect 64388 -394 64438 -264
rect 64690 -270 64870 -250
rect 64690 -370 64730 -270
rect 64830 -370 64870 -270
rect 64690 -390 64870 -370
rect 65710 -270 65890 -250
rect 65710 -370 65750 -270
rect 65850 -370 65890 -270
rect 65710 -390 65890 -370
rect 67110 -270 67250 -250
rect 67210 -370 67250 -270
rect 67110 -390 67250 -370
rect 67664 -264 67994 -244
rect 68480 -260 68580 -220
rect 69860 -260 69920 -220
rect 63380 -410 63460 -400
rect 63390 -650 63450 -410
rect 64108 -414 64438 -394
rect 64750 -650 64810 -390
rect 65770 -650 65830 -390
rect 56570 -730 56590 -670
rect 56650 -730 56670 -670
rect 56570 -750 56670 -730
rect 57930 -670 58030 -650
rect 57930 -730 57950 -670
rect 58010 -730 58030 -670
rect 57930 -750 58030 -730
rect 59630 -670 59730 -650
rect 59630 -730 59650 -670
rect 59710 -730 59730 -670
rect 59630 -750 59730 -730
rect 60990 -670 61090 -650
rect 60990 -730 61010 -670
rect 61070 -730 61090 -670
rect 60990 -750 61090 -730
rect 62010 -670 62110 -650
rect 62010 -730 62030 -670
rect 62090 -730 62110 -670
rect 62010 -750 62110 -730
rect 63370 -670 63470 -650
rect 63370 -730 63390 -670
rect 63450 -730 63470 -670
rect 63370 -750 63470 -730
rect 64730 -670 64830 -650
rect 64730 -730 64750 -670
rect 64810 -730 64830 -670
rect 64730 -750 64830 -730
rect 65750 -670 65850 -650
rect 65750 -730 65770 -670
rect 65830 -730 65850 -670
rect 65750 -750 65850 -730
rect 67110 -670 67210 -390
rect 67664 -394 67714 -264
rect 67944 -394 67994 -264
rect 68430 -270 68610 -260
rect 68430 -370 68470 -270
rect 68570 -370 68610 -270
rect 68430 -390 68610 -370
rect 69800 -280 69980 -260
rect 69800 -380 69840 -280
rect 69940 -380 69980 -280
rect 67664 -414 67994 -394
rect 67110 -730 67130 -670
rect 67190 -730 67210 -670
rect 67110 -750 67210 -730
rect 68470 -670 68570 -390
rect 69800 -400 69980 -380
rect 70508 -264 70838 -244
rect 71550 -260 71610 -250
rect 70508 -394 70558 -264
rect 70788 -394 70838 -264
rect 69850 -650 69910 -400
rect 70508 -414 70838 -394
rect 71490 -280 71670 -260
rect 71490 -380 71530 -280
rect 71630 -380 71670 -280
rect 71490 -400 71670 -380
rect 72850 -270 73030 -250
rect 72850 -370 72890 -270
rect 72990 -370 73030 -270
rect 72850 -390 73030 -370
rect 73870 -270 74050 -250
rect 73870 -370 73910 -270
rect 74010 -370 74050 -270
rect 73870 -390 74050 -370
rect 74418 -264 74748 -244
rect 75290 -260 75350 -250
rect 71540 -410 71620 -400
rect 71550 -650 71610 -410
rect 72910 -650 72970 -390
rect 73930 -650 73990 -390
rect 74418 -394 74468 -264
rect 74698 -394 74748 -264
rect 74418 -414 74748 -394
rect 75230 -280 75410 -260
rect 75230 -380 75270 -280
rect 75370 -380 75410 -280
rect 75230 -400 75410 -380
rect 76590 -270 76770 -250
rect 76590 -370 76630 -270
rect 76730 -370 76770 -270
rect 76590 -390 76770 -370
rect 77610 -270 77790 -250
rect 77610 -370 77650 -270
rect 77750 -370 77790 -270
rect 77610 -390 77790 -370
rect 78330 -264 78660 -244
rect 75280 -410 75360 -400
rect 75290 -650 75350 -410
rect 76650 -650 76710 -390
rect 77670 -650 77730 -390
rect 78330 -394 78380 -264
rect 78610 -394 78660 -264
rect 78330 -414 78660 -394
rect 79010 -270 79150 -250
rect 80380 -260 80480 -220
rect 81760 -260 81820 -220
rect 79110 -370 79150 -270
rect 79010 -390 79150 -370
rect 80330 -270 80510 -260
rect 80330 -370 80370 -270
rect 80470 -370 80510 -270
rect 80330 -390 80510 -370
rect 81700 -280 81880 -260
rect 81700 -380 81740 -280
rect 81840 -380 81880 -280
rect 68470 -730 68490 -670
rect 68550 -730 68570 -670
rect 68470 -750 68570 -730
rect 69830 -670 69930 -650
rect 69830 -730 69850 -670
rect 69910 -730 69930 -670
rect 69830 -750 69930 -730
rect 71530 -670 71630 -650
rect 71530 -730 71550 -670
rect 71610 -730 71630 -670
rect 71530 -750 71630 -730
rect 72890 -670 72990 -650
rect 72890 -730 72910 -670
rect 72970 -730 72990 -670
rect 72890 -750 72990 -730
rect 73910 -670 74010 -650
rect 73910 -730 73930 -670
rect 73990 -730 74010 -670
rect 73910 -750 74010 -730
rect 75270 -670 75370 -650
rect 75270 -730 75290 -670
rect 75350 -730 75370 -670
rect 75270 -750 75370 -730
rect 76630 -670 76730 -650
rect 76630 -730 76650 -670
rect 76710 -730 76730 -670
rect 76630 -750 76730 -730
rect 77650 -670 77750 -650
rect 77650 -730 77670 -670
rect 77730 -730 77750 -670
rect 77650 -750 77750 -730
rect 79010 -670 79110 -390
rect 79010 -730 79030 -670
rect 79090 -730 79110 -670
rect 79010 -750 79110 -730
rect 80370 -670 80470 -390
rect 81700 -400 81880 -380
rect 82242 -264 82572 -244
rect 83450 -260 83510 -250
rect 82242 -394 82292 -264
rect 82522 -394 82572 -264
rect 81750 -650 81810 -400
rect 82242 -414 82572 -394
rect 83390 -280 83570 -260
rect 83390 -380 83430 -280
rect 83530 -380 83570 -280
rect 83390 -400 83570 -380
rect 84750 -270 84930 -250
rect 84750 -370 84790 -270
rect 84890 -370 84930 -270
rect 84750 -390 84930 -370
rect 85770 -270 85950 -250
rect 85770 -370 85810 -270
rect 85910 -370 85950 -270
rect 85770 -390 85950 -370
rect 86152 -264 86482 -244
rect 87190 -260 87250 -250
rect 83440 -410 83520 -400
rect 83450 -650 83510 -410
rect 84810 -650 84870 -390
rect 85830 -650 85890 -390
rect 86152 -394 86202 -264
rect 86432 -394 86482 -264
rect 86152 -414 86482 -394
rect 87130 -280 87310 -260
rect 87130 -380 87170 -280
rect 87270 -380 87310 -280
rect 87130 -400 87310 -380
rect 87180 -410 87260 -400
rect 87190 -650 87250 -410
rect 80370 -730 80390 -670
rect 80450 -730 80470 -670
rect 80370 -750 80470 -730
rect 81730 -670 81830 -650
rect 81730 -730 81750 -670
rect 81810 -730 81830 -670
rect 81730 -750 81830 -730
rect 83430 -670 83530 -650
rect 83430 -730 83450 -670
rect 83510 -730 83530 -670
rect 83430 -750 83530 -730
rect 84790 -670 84890 -650
rect 84790 -730 84810 -670
rect 84870 -730 84890 -670
rect 84790 -750 84890 -730
rect 85810 -670 85910 -650
rect 85810 -730 85830 -670
rect 85890 -730 85910 -670
rect 85810 -750 85910 -730
rect 87170 -670 87270 -650
rect 87170 -730 87190 -670
rect 87250 -730 87270 -670
rect 87170 -750 87270 -730
rect 290 -870 410 -860
rect 290 -960 310 -870
rect 390 -960 410 -870
rect 290 -970 410 -960
rect 630 -870 750 -860
rect 630 -960 650 -870
rect 730 -960 750 -870
rect 630 -970 750 -960
rect 970 -870 1090 -860
rect 970 -960 990 -870
rect 1070 -960 1090 -870
rect 970 -970 1090 -960
rect 1310 -870 1430 -860
rect 1310 -960 1330 -870
rect 1410 -960 1430 -870
rect 1310 -970 1430 -960
rect 1650 -870 1770 -860
rect 1650 -960 1670 -870
rect 1750 -960 1770 -870
rect 1650 -970 1770 -960
rect 1990 -870 2110 -860
rect 1990 -960 2010 -870
rect 2090 -960 2110 -870
rect 1990 -970 2110 -960
rect 2330 -870 2450 -860
rect 2330 -960 2350 -870
rect 2430 -960 2450 -870
rect 2330 -970 2450 -960
rect 2670 -870 2790 -860
rect 2670 -960 2690 -870
rect 2770 -960 2790 -870
rect 2670 -970 2790 -960
rect 3010 -870 3130 -860
rect 3010 -960 3030 -870
rect 3110 -960 3130 -870
rect 3010 -970 3130 -960
rect 3350 -870 3470 -860
rect 3350 -960 3370 -870
rect 3450 -960 3470 -870
rect 3350 -970 3470 -960
rect 3690 -870 3810 -860
rect 3690 -960 3710 -870
rect 3790 -960 3810 -870
rect 3690 -970 3810 -960
rect 4030 -870 4150 -860
rect 4030 -960 4050 -870
rect 4130 -960 4150 -870
rect 4030 -970 4150 -960
rect 4370 -870 4490 -860
rect 4370 -960 4390 -870
rect 4470 -960 4490 -870
rect 4370 -970 4490 -960
rect 4710 -870 4830 -860
rect 4710 -960 4730 -870
rect 4810 -960 4830 -870
rect 4710 -970 4830 -960
rect 5050 -870 5170 -860
rect 5050 -960 5070 -870
rect 5150 -960 5170 -870
rect 5050 -970 5170 -960
rect 5390 -870 5510 -860
rect 5390 -960 5410 -870
rect 5490 -960 5510 -870
rect 5390 -970 5510 -960
rect 5730 -870 5850 -860
rect 5730 -960 5750 -870
rect 5830 -960 5850 -870
rect 5730 -970 5850 -960
rect 6070 -870 6190 -860
rect 6070 -960 6090 -870
rect 6170 -960 6190 -870
rect 6070 -970 6190 -960
rect 6410 -870 6530 -860
rect 6410 -960 6430 -870
rect 6510 -960 6530 -870
rect 6410 -970 6530 -960
rect 6750 -870 6870 -860
rect 6750 -960 6770 -870
rect 6850 -960 6870 -870
rect 6750 -970 6870 -960
rect 7090 -870 7210 -860
rect 7090 -960 7110 -870
rect 7190 -960 7210 -870
rect 7090 -970 7210 -960
rect 7430 -870 7550 -860
rect 7430 -960 7450 -870
rect 7530 -960 7550 -870
rect 7430 -970 7550 -960
rect 7770 -870 7890 -860
rect 7770 -960 7790 -870
rect 7870 -960 7890 -870
rect 7770 -970 7890 -960
rect 8110 -870 8230 -860
rect 8110 -960 8130 -870
rect 8210 -960 8230 -870
rect 8110 -970 8230 -960
rect 8450 -870 8570 -860
rect 8450 -960 8470 -870
rect 8550 -960 8570 -870
rect 8450 -970 8570 -960
rect 8790 -870 8910 -860
rect 8790 -960 8810 -870
rect 8890 -960 8910 -870
rect 8790 -970 8910 -960
rect 9130 -870 9250 -860
rect 9130 -960 9150 -870
rect 9230 -960 9250 -870
rect 9130 -970 9250 -960
rect 9470 -870 9590 -860
rect 9470 -960 9490 -870
rect 9570 -960 9590 -870
rect 9470 -970 9590 -960
rect 9810 -870 9930 -860
rect 9810 -960 9830 -870
rect 9910 -960 9930 -870
rect 9810 -970 9930 -960
rect 10150 -870 10270 -860
rect 10150 -960 10170 -870
rect 10250 -960 10270 -870
rect 10150 -970 10270 -960
rect 10490 -870 10610 -860
rect 10490 -960 10510 -870
rect 10590 -960 10610 -870
rect 10490 -970 10610 -960
rect 10830 -870 10950 -860
rect 10830 -960 10850 -870
rect 10930 -960 10950 -870
rect 10830 -970 10950 -960
rect 11170 -870 11290 -860
rect 11170 -960 11190 -870
rect 11270 -960 11290 -870
rect 11170 -970 11290 -960
rect 11510 -870 11630 -860
rect 11510 -960 11530 -870
rect 11610 -960 11630 -870
rect 11510 -970 11630 -960
rect 11850 -870 11970 -860
rect 11850 -960 11870 -870
rect 11950 -960 11970 -870
rect 11850 -970 11970 -960
rect 12190 -870 12310 -860
rect 12190 -960 12210 -870
rect 12290 -960 12310 -870
rect 12190 -970 12310 -960
rect 12530 -870 12650 -860
rect 12530 -960 12550 -870
rect 12630 -960 12650 -870
rect 12530 -970 12650 -960
rect 12870 -870 12990 -860
rect 12870 -960 12890 -870
rect 12970 -960 12990 -870
rect 12870 -970 12990 -960
rect 13210 -870 13330 -860
rect 13210 -960 13230 -870
rect 13310 -960 13330 -870
rect 13210 -970 13330 -960
rect 13550 -870 13670 -860
rect 13550 -960 13570 -870
rect 13650 -960 13670 -870
rect 13550 -970 13670 -960
rect 13890 -870 14010 -860
rect 13890 -960 13910 -870
rect 13990 -960 14010 -870
rect 13890 -970 14010 -960
rect 14230 -870 14350 -860
rect 14230 -960 14250 -870
rect 14330 -960 14350 -870
rect 14230 -970 14350 -960
rect 14570 -870 14690 -860
rect 14570 -960 14590 -870
rect 14670 -960 14690 -870
rect 14570 -970 14690 -960
rect 14910 -870 15030 -860
rect 14910 -960 14930 -870
rect 15010 -960 15030 -870
rect 14910 -970 15030 -960
rect 15250 -870 15370 -860
rect 15250 -960 15270 -870
rect 15350 -960 15370 -870
rect 15250 -970 15370 -960
rect 15590 -870 15710 -860
rect 15590 -960 15610 -870
rect 15690 -960 15710 -870
rect 15590 -970 15710 -960
rect 15930 -870 16050 -860
rect 15930 -960 15950 -870
rect 16030 -960 16050 -870
rect 15930 -970 16050 -960
rect 16270 -870 16390 -860
rect 16270 -960 16290 -870
rect 16370 -960 16390 -870
rect 16270 -970 16390 -960
rect 16610 -870 16730 -860
rect 16610 -960 16630 -870
rect 16710 -960 16730 -870
rect 16610 -970 16730 -960
rect 16950 -870 17070 -860
rect 16950 -960 16970 -870
rect 17050 -960 17070 -870
rect 16950 -970 17070 -960
rect 17290 -870 17410 -860
rect 17290 -960 17310 -870
rect 17390 -960 17410 -870
rect 17290 -970 17410 -960
rect 17630 -870 17750 -860
rect 17630 -960 17650 -870
rect 17730 -960 17750 -870
rect 17630 -970 17750 -960
rect 17970 -870 18090 -860
rect 17970 -960 17990 -870
rect 18070 -960 18090 -870
rect 17970 -970 18090 -960
rect 18310 -870 18430 -860
rect 18310 -960 18330 -870
rect 18410 -960 18430 -870
rect 18310 -970 18430 -960
rect 18650 -870 18770 -860
rect 18650 -960 18670 -870
rect 18750 -960 18770 -870
rect 18650 -970 18770 -960
rect 18990 -870 19110 -860
rect 18990 -960 19010 -870
rect 19090 -960 19110 -870
rect 18990 -970 19110 -960
rect 19330 -870 19450 -860
rect 19330 -960 19350 -870
rect 19430 -960 19450 -870
rect 19330 -970 19450 -960
rect 19670 -870 19790 -860
rect 19670 -960 19690 -870
rect 19770 -960 19790 -870
rect 19670 -970 19790 -960
rect 20010 -870 20130 -860
rect 20010 -960 20030 -870
rect 20110 -960 20130 -870
rect 20010 -970 20130 -960
rect 20350 -870 20470 -860
rect 20350 -960 20370 -870
rect 20450 -960 20470 -870
rect 20350 -970 20470 -960
rect 20690 -870 20810 -860
rect 20690 -960 20710 -870
rect 20790 -960 20810 -870
rect 20690 -970 20810 -960
rect 21030 -870 21150 -860
rect 21030 -960 21050 -870
rect 21130 -960 21150 -870
rect 21030 -970 21150 -960
rect 21370 -870 21490 -860
rect 21370 -960 21390 -870
rect 21470 -960 21490 -870
rect 21370 -970 21490 -960
rect 21710 -870 21830 -860
rect 21710 -960 21730 -870
rect 21810 -960 21830 -870
rect 21710 -970 21830 -960
rect 22050 -870 22170 -860
rect 22050 -960 22070 -870
rect 22150 -960 22170 -870
rect 22050 -970 22170 -960
rect 22390 -870 22510 -860
rect 22390 -960 22410 -870
rect 22490 -960 22510 -870
rect 22390 -970 22510 -960
rect 22730 -870 22850 -860
rect 22730 -960 22750 -870
rect 22830 -960 22850 -870
rect 22730 -970 22850 -960
rect 23070 -870 23190 -860
rect 23070 -960 23090 -870
rect 23170 -960 23190 -870
rect 23070 -970 23190 -960
rect 23410 -870 23530 -860
rect 23410 -960 23430 -870
rect 23510 -960 23530 -870
rect 23410 -970 23530 -960
rect 23750 -870 23870 -860
rect 23750 -960 23770 -870
rect 23850 -960 23870 -870
rect 23750 -970 23870 -960
rect 24090 -870 24210 -860
rect 24090 -960 24110 -870
rect 24190 -960 24210 -870
rect 24090 -970 24210 -960
rect 24430 -870 24550 -860
rect 24430 -960 24450 -870
rect 24530 -960 24550 -870
rect 24430 -970 24550 -960
rect 24770 -870 24890 -860
rect 24770 -960 24790 -870
rect 24870 -960 24890 -870
rect 24770 -970 24890 -960
rect 25110 -870 25230 -860
rect 25110 -960 25130 -870
rect 25210 -960 25230 -870
rect 25110 -970 25230 -960
rect 25450 -870 25570 -860
rect 25450 -960 25470 -870
rect 25550 -960 25570 -870
rect 25450 -970 25570 -960
rect 25790 -870 25910 -860
rect 25790 -960 25810 -870
rect 25890 -960 25910 -870
rect 25790 -970 25910 -960
rect 26130 -870 26250 -860
rect 26130 -960 26150 -870
rect 26230 -960 26250 -870
rect 26130 -970 26250 -960
rect 26470 -870 26590 -860
rect 26470 -960 26490 -870
rect 26570 -960 26590 -870
rect 26470 -970 26590 -960
rect 26810 -870 26930 -860
rect 26810 -960 26830 -870
rect 26910 -960 26930 -870
rect 26810 -970 26930 -960
rect 27150 -870 27270 -860
rect 27150 -960 27170 -870
rect 27250 -960 27270 -870
rect 27150 -970 27270 -960
rect 27490 -870 27610 -860
rect 27490 -960 27510 -870
rect 27590 -960 27610 -870
rect 27490 -970 27610 -960
rect 27830 -870 27950 -860
rect 27830 -960 27850 -870
rect 27930 -960 27950 -870
rect 27830 -970 27950 -960
rect 28170 -870 28290 -860
rect 28170 -960 28190 -870
rect 28270 -960 28290 -870
rect 28170 -970 28290 -960
rect 28510 -870 28630 -860
rect 28510 -960 28530 -870
rect 28610 -960 28630 -870
rect 28510 -970 28630 -960
rect 28850 -870 28970 -860
rect 28850 -960 28870 -870
rect 28950 -960 28970 -870
rect 28850 -970 28970 -960
rect 29190 -870 29310 -860
rect 29190 -960 29210 -870
rect 29290 -960 29310 -870
rect 29190 -970 29310 -960
rect 29530 -870 29650 -860
rect 29530 -960 29550 -870
rect 29630 -960 29650 -870
rect 29530 -970 29650 -960
rect 29870 -870 29990 -860
rect 29870 -960 29890 -870
rect 29970 -960 29990 -870
rect 29870 -970 29990 -960
rect 30210 -870 30330 -860
rect 30210 -960 30230 -870
rect 30310 -960 30330 -870
rect 30210 -970 30330 -960
rect 30550 -870 30670 -860
rect 30550 -960 30570 -870
rect 30650 -960 30670 -870
rect 30550 -970 30670 -960
rect 30890 -870 31010 -860
rect 30890 -960 30910 -870
rect 30990 -960 31010 -870
rect 30890 -970 31010 -960
rect 31230 -870 31350 -860
rect 31230 -960 31250 -870
rect 31330 -960 31350 -870
rect 31230 -970 31350 -960
rect 31570 -870 31690 -860
rect 31570 -960 31590 -870
rect 31670 -960 31690 -870
rect 31570 -970 31690 -960
rect 31910 -870 32030 -860
rect 31910 -960 31930 -870
rect 32010 -960 32030 -870
rect 31910 -970 32030 -960
rect 32250 -870 32370 -860
rect 32250 -960 32270 -870
rect 32350 -960 32370 -870
rect 32250 -970 32370 -960
rect 32590 -870 32710 -860
rect 32590 -960 32610 -870
rect 32690 -960 32710 -870
rect 32590 -970 32710 -960
rect 32930 -870 33050 -860
rect 32930 -960 32950 -870
rect 33030 -960 33050 -870
rect 32930 -970 33050 -960
rect 33270 -870 33390 -860
rect 33270 -960 33290 -870
rect 33370 -960 33390 -870
rect 33270 -970 33390 -960
rect 33610 -870 33730 -860
rect 33610 -960 33630 -870
rect 33710 -960 33730 -870
rect 33610 -970 33730 -960
rect 33950 -870 34070 -860
rect 33950 -960 33970 -870
rect 34050 -960 34070 -870
rect 33950 -970 34070 -960
rect 34290 -870 34410 -860
rect 34290 -960 34310 -870
rect 34390 -960 34410 -870
rect 34290 -970 34410 -960
rect 34630 -870 34750 -860
rect 34630 -960 34650 -870
rect 34730 -960 34750 -870
rect 34630 -970 34750 -960
rect 34970 -870 35090 -860
rect 34970 -960 34990 -870
rect 35070 -960 35090 -870
rect 34970 -970 35090 -960
rect 35310 -870 35430 -860
rect 35310 -960 35330 -870
rect 35410 -960 35430 -870
rect 35310 -970 35430 -960
rect 35650 -870 35770 -860
rect 35650 -960 35670 -870
rect 35750 -960 35770 -870
rect 35650 -970 35770 -960
rect 35990 -870 36110 -860
rect 35990 -960 36010 -870
rect 36090 -960 36110 -870
rect 35990 -970 36110 -960
rect 36330 -870 36450 -860
rect 36330 -960 36350 -870
rect 36430 -960 36450 -870
rect 36330 -970 36450 -960
rect 36670 -870 36790 -860
rect 36670 -960 36690 -870
rect 36770 -960 36790 -870
rect 36670 -970 36790 -960
rect 37010 -870 37130 -860
rect 37010 -960 37030 -870
rect 37110 -960 37130 -870
rect 37010 -970 37130 -960
rect 37350 -870 37470 -860
rect 37350 -960 37370 -870
rect 37450 -960 37470 -870
rect 37350 -970 37470 -960
rect 37690 -870 37810 -860
rect 37690 -960 37710 -870
rect 37790 -960 37810 -870
rect 37690 -970 37810 -960
rect 38030 -870 38150 -860
rect 38030 -960 38050 -870
rect 38130 -960 38150 -870
rect 38030 -970 38150 -960
rect 38370 -870 38490 -860
rect 38370 -960 38390 -870
rect 38470 -960 38490 -870
rect 38370 -970 38490 -960
rect 38710 -870 38830 -860
rect 38710 -960 38730 -870
rect 38810 -960 38830 -870
rect 38710 -970 38830 -960
rect 39050 -870 39170 -860
rect 39050 -960 39070 -870
rect 39150 -960 39170 -870
rect 39050 -970 39170 -960
rect 39390 -870 39510 -860
rect 39390 -960 39410 -870
rect 39490 -960 39510 -870
rect 39390 -970 39510 -960
rect 39730 -870 39850 -860
rect 39730 -960 39750 -870
rect 39830 -960 39850 -870
rect 39730 -970 39850 -960
rect 40070 -870 40190 -860
rect 40070 -960 40090 -870
rect 40170 -960 40190 -870
rect 40070 -970 40190 -960
rect 40410 -870 40530 -860
rect 40410 -960 40430 -870
rect 40510 -960 40530 -870
rect 40410 -970 40530 -960
rect 40750 -870 40870 -860
rect 40750 -960 40770 -870
rect 40850 -960 40870 -870
rect 40750 -970 40870 -960
rect 41090 -870 41210 -860
rect 41090 -960 41110 -870
rect 41190 -960 41210 -870
rect 41090 -970 41210 -960
rect 41430 -870 41550 -860
rect 41430 -960 41450 -870
rect 41530 -960 41550 -870
rect 41430 -970 41550 -960
rect 41770 -870 41890 -860
rect 41770 -960 41790 -870
rect 41870 -960 41890 -870
rect 41770 -970 41890 -960
rect 42110 -870 42230 -860
rect 42110 -960 42130 -870
rect 42210 -960 42230 -870
rect 42110 -970 42230 -960
rect 42450 -870 42570 -860
rect 42450 -960 42470 -870
rect 42550 -960 42570 -870
rect 42450 -970 42570 -960
rect 42790 -870 42910 -860
rect 42790 -960 42810 -870
rect 42890 -960 42910 -870
rect 42790 -970 42910 -960
rect 43130 -870 43250 -860
rect 43130 -960 43150 -870
rect 43230 -960 43250 -870
rect 43130 -970 43250 -960
rect 43470 -870 43590 -860
rect 43470 -960 43490 -870
rect 43570 -960 43590 -870
rect 43470 -970 43590 -960
rect 43810 -870 43930 -860
rect 43810 -960 43830 -870
rect 43910 -960 43930 -870
rect 43810 -970 43930 -960
rect 44150 -870 44270 -860
rect 44150 -960 44170 -870
rect 44250 -960 44270 -870
rect 44150 -970 44270 -960
rect 44490 -870 44610 -860
rect 44490 -960 44510 -870
rect 44590 -960 44610 -870
rect 44490 -970 44610 -960
rect 44830 -870 44950 -860
rect 44830 -960 44850 -870
rect 44930 -960 44950 -870
rect 44830 -970 44950 -960
rect 45170 -870 45290 -860
rect 45170 -960 45190 -870
rect 45270 -960 45290 -870
rect 45170 -970 45290 -960
rect 45510 -870 45630 -860
rect 45510 -960 45530 -870
rect 45610 -960 45630 -870
rect 45510 -970 45630 -960
rect 45850 -870 45970 -860
rect 45850 -960 45870 -870
rect 45950 -960 45970 -870
rect 45850 -970 45970 -960
rect 46190 -870 46310 -860
rect 46190 -960 46210 -870
rect 46290 -960 46310 -870
rect 46190 -970 46310 -960
rect 46530 -870 46650 -860
rect 46530 -960 46550 -870
rect 46630 -960 46650 -870
rect 46530 -970 46650 -960
rect 46870 -870 46990 -860
rect 46870 -960 46890 -870
rect 46970 -960 46990 -870
rect 46870 -970 46990 -960
rect 47210 -870 47330 -860
rect 47210 -960 47230 -870
rect 47310 -960 47330 -870
rect 47210 -970 47330 -960
rect 47550 -870 47670 -860
rect 47550 -960 47570 -870
rect 47650 -960 47670 -870
rect 47550 -970 47670 -960
rect 47890 -870 48010 -860
rect 47890 -960 47910 -870
rect 47990 -960 48010 -870
rect 47890 -970 48010 -960
rect 48230 -870 48350 -860
rect 48230 -960 48250 -870
rect 48330 -960 48350 -870
rect 48230 -970 48350 -960
rect 48570 -870 48690 -860
rect 48570 -960 48590 -870
rect 48670 -960 48690 -870
rect 48570 -970 48690 -960
rect 48910 -870 49030 -860
rect 48910 -960 48930 -870
rect 49010 -960 49030 -870
rect 48910 -970 49030 -960
rect 49250 -870 49370 -860
rect 49250 -960 49270 -870
rect 49350 -960 49370 -870
rect 49250 -970 49370 -960
rect 49590 -870 49710 -860
rect 49590 -960 49610 -870
rect 49690 -960 49710 -870
rect 49590 -970 49710 -960
rect 49930 -870 50050 -860
rect 49930 -960 49950 -870
rect 50030 -960 50050 -870
rect 49930 -970 50050 -960
rect 50270 -870 50390 -860
rect 50270 -960 50290 -870
rect 50370 -960 50390 -870
rect 50270 -970 50390 -960
rect 50610 -870 50730 -860
rect 50610 -960 50630 -870
rect 50710 -960 50730 -870
rect 50610 -970 50730 -960
rect 50950 -870 51070 -860
rect 50950 -960 50970 -870
rect 51050 -960 51070 -870
rect 50950 -970 51070 -960
rect 51290 -870 51410 -860
rect 51290 -960 51310 -870
rect 51390 -960 51410 -870
rect 51290 -970 51410 -960
rect 51630 -870 51750 -860
rect 51630 -960 51650 -870
rect 51730 -960 51750 -870
rect 51630 -970 51750 -960
rect 51970 -870 52090 -860
rect 51970 -960 51990 -870
rect 52070 -960 52090 -870
rect 51970 -970 52090 -960
rect 52310 -870 52430 -860
rect 52310 -960 52330 -870
rect 52410 -960 52430 -870
rect 52310 -970 52430 -960
rect 52650 -870 52770 -860
rect 52650 -960 52670 -870
rect 52750 -960 52770 -870
rect 52650 -970 52770 -960
rect 52990 -870 53110 -860
rect 52990 -960 53010 -870
rect 53090 -960 53110 -870
rect 52990 -970 53110 -960
rect 53330 -870 53450 -860
rect 53330 -960 53350 -870
rect 53430 -960 53450 -870
rect 53330 -970 53450 -960
rect 53670 -870 53790 -860
rect 53670 -960 53690 -870
rect 53770 -960 53790 -870
rect 53670 -970 53790 -960
rect 54010 -870 54130 -860
rect 54010 -960 54030 -870
rect 54110 -960 54130 -870
rect 54010 -970 54130 -960
rect 54350 -870 54470 -860
rect 54350 -960 54370 -870
rect 54450 -960 54470 -870
rect 54350 -970 54470 -960
rect 54690 -870 54810 -860
rect 54690 -960 54710 -870
rect 54790 -960 54810 -870
rect 54690 -970 54810 -960
rect 55030 -870 55150 -860
rect 55030 -960 55050 -870
rect 55130 -960 55150 -870
rect 55030 -970 55150 -960
rect 55370 -870 55490 -860
rect 55370 -960 55390 -870
rect 55470 -960 55490 -870
rect 55370 -970 55490 -960
rect 55710 -870 55830 -860
rect 55710 -960 55730 -870
rect 55810 -960 55830 -870
rect 55710 -970 55830 -960
rect 56050 -870 56170 -860
rect 56050 -960 56070 -870
rect 56150 -960 56170 -870
rect 56050 -970 56170 -960
rect 56390 -870 56510 -860
rect 56390 -960 56410 -870
rect 56490 -960 56510 -870
rect 56390 -970 56510 -960
rect 56730 -870 56850 -860
rect 56730 -960 56750 -870
rect 56830 -960 56850 -870
rect 56730 -970 56850 -960
rect 57070 -870 57190 -860
rect 57070 -960 57090 -870
rect 57170 -960 57190 -870
rect 57070 -970 57190 -960
rect 57410 -870 57530 -860
rect 57410 -960 57430 -870
rect 57510 -960 57530 -870
rect 57410 -970 57530 -960
rect 57750 -870 57870 -860
rect 57750 -960 57770 -870
rect 57850 -960 57870 -870
rect 57750 -970 57870 -960
rect 58090 -870 58210 -860
rect 58090 -960 58110 -870
rect 58190 -960 58210 -870
rect 58090 -970 58210 -960
rect 58430 -870 58550 -860
rect 58430 -960 58450 -870
rect 58530 -960 58550 -870
rect 58430 -970 58550 -960
rect 58770 -870 58890 -860
rect 58770 -960 58790 -870
rect 58870 -960 58890 -870
rect 58770 -970 58890 -960
rect 59110 -870 59230 -860
rect 59110 -960 59130 -870
rect 59210 -960 59230 -870
rect 59110 -970 59230 -960
rect 59450 -870 59570 -860
rect 59450 -960 59470 -870
rect 59550 -960 59570 -870
rect 59450 -970 59570 -960
rect 59790 -870 59910 -860
rect 59790 -960 59810 -870
rect 59890 -960 59910 -870
rect 59790 -970 59910 -960
rect 60130 -870 60250 -860
rect 60130 -960 60150 -870
rect 60230 -960 60250 -870
rect 60130 -970 60250 -960
rect 60470 -870 60590 -860
rect 60470 -960 60490 -870
rect 60570 -960 60590 -870
rect 60470 -970 60590 -960
rect 60810 -870 60930 -860
rect 60810 -960 60830 -870
rect 60910 -960 60930 -870
rect 60810 -970 60930 -960
rect 61150 -870 61270 -860
rect 61150 -960 61170 -870
rect 61250 -960 61270 -870
rect 61150 -970 61270 -960
rect 61490 -870 61610 -860
rect 61490 -960 61510 -870
rect 61590 -960 61610 -870
rect 61490 -970 61610 -960
rect 61830 -870 61950 -860
rect 61830 -960 61850 -870
rect 61930 -960 61950 -870
rect 61830 -970 61950 -960
rect 62170 -870 62290 -860
rect 62170 -960 62190 -870
rect 62270 -960 62290 -870
rect 62170 -970 62290 -960
rect 62510 -870 62630 -860
rect 62510 -960 62530 -870
rect 62610 -960 62630 -870
rect 62510 -970 62630 -960
rect 62850 -870 62970 -860
rect 62850 -960 62870 -870
rect 62950 -960 62970 -870
rect 62850 -970 62970 -960
rect 63190 -870 63310 -860
rect 63190 -960 63210 -870
rect 63290 -960 63310 -870
rect 63190 -970 63310 -960
rect 63530 -870 63650 -860
rect 63530 -960 63550 -870
rect 63630 -960 63650 -870
rect 63530 -970 63650 -960
rect 63870 -870 63990 -860
rect 63870 -960 63890 -870
rect 63970 -960 63990 -870
rect 63870 -970 63990 -960
rect 64210 -870 64330 -860
rect 64210 -960 64230 -870
rect 64310 -960 64330 -870
rect 64210 -970 64330 -960
rect 64550 -870 64670 -860
rect 64550 -960 64570 -870
rect 64650 -960 64670 -870
rect 64550 -970 64670 -960
rect 64890 -870 65010 -860
rect 64890 -960 64910 -870
rect 64990 -960 65010 -870
rect 64890 -970 65010 -960
rect 65230 -870 65350 -860
rect 65230 -960 65250 -870
rect 65330 -960 65350 -870
rect 65230 -970 65350 -960
rect 65570 -870 65690 -860
rect 65570 -960 65590 -870
rect 65670 -960 65690 -870
rect 65570 -970 65690 -960
rect 65910 -870 66030 -860
rect 65910 -960 65930 -870
rect 66010 -960 66030 -870
rect 65910 -970 66030 -960
rect 66250 -870 66370 -860
rect 66250 -960 66270 -870
rect 66350 -960 66370 -870
rect 66250 -970 66370 -960
rect 66590 -870 66710 -860
rect 66590 -960 66610 -870
rect 66690 -960 66710 -870
rect 66590 -970 66710 -960
rect 66930 -870 67050 -860
rect 66930 -960 66950 -870
rect 67030 -960 67050 -870
rect 66930 -970 67050 -960
rect 67270 -870 67390 -860
rect 67270 -960 67290 -870
rect 67370 -960 67390 -870
rect 67270 -970 67390 -960
rect 67610 -870 67730 -860
rect 67610 -960 67630 -870
rect 67710 -960 67730 -870
rect 67610 -970 67730 -960
rect 67950 -870 68070 -860
rect 67950 -960 67970 -870
rect 68050 -960 68070 -870
rect 67950 -970 68070 -960
rect 68290 -870 68410 -860
rect 68290 -960 68310 -870
rect 68390 -960 68410 -870
rect 68290 -970 68410 -960
rect 68630 -870 68750 -860
rect 68630 -960 68650 -870
rect 68730 -960 68750 -870
rect 68630 -970 68750 -960
rect 68970 -870 69090 -860
rect 68970 -960 68990 -870
rect 69070 -960 69090 -870
rect 68970 -970 69090 -960
rect 69310 -870 69430 -860
rect 69310 -960 69330 -870
rect 69410 -960 69430 -870
rect 69310 -970 69430 -960
rect 69650 -870 69770 -860
rect 69650 -960 69670 -870
rect 69750 -960 69770 -870
rect 69650 -970 69770 -960
rect 69990 -870 70110 -860
rect 69990 -960 70010 -870
rect 70090 -960 70110 -870
rect 69990 -970 70110 -960
rect 70330 -870 70450 -860
rect 70330 -960 70350 -870
rect 70430 -960 70450 -870
rect 70330 -970 70450 -960
rect 70670 -870 70790 -860
rect 70670 -960 70690 -870
rect 70770 -960 70790 -870
rect 70670 -970 70790 -960
rect 71010 -870 71130 -860
rect 71010 -960 71030 -870
rect 71110 -960 71130 -870
rect 71010 -970 71130 -960
rect 71350 -870 71470 -860
rect 71350 -960 71370 -870
rect 71450 -960 71470 -870
rect 71350 -970 71470 -960
rect 71690 -870 71810 -860
rect 71690 -960 71710 -870
rect 71790 -960 71810 -870
rect 71690 -970 71810 -960
rect 72030 -870 72150 -860
rect 72030 -960 72050 -870
rect 72130 -960 72150 -870
rect 72030 -970 72150 -960
rect 72370 -870 72490 -860
rect 72370 -960 72390 -870
rect 72470 -960 72490 -870
rect 72370 -970 72490 -960
rect 72710 -870 72830 -860
rect 72710 -960 72730 -870
rect 72810 -960 72830 -870
rect 72710 -970 72830 -960
rect 73050 -870 73170 -860
rect 73050 -960 73070 -870
rect 73150 -960 73170 -870
rect 73050 -970 73170 -960
rect 73390 -870 73510 -860
rect 73390 -960 73410 -870
rect 73490 -960 73510 -870
rect 73390 -970 73510 -960
rect 73730 -870 73850 -860
rect 73730 -960 73750 -870
rect 73830 -960 73850 -870
rect 73730 -970 73850 -960
rect 74070 -870 74190 -860
rect 74070 -960 74090 -870
rect 74170 -960 74190 -870
rect 74070 -970 74190 -960
rect 74410 -870 74530 -860
rect 74410 -960 74430 -870
rect 74510 -960 74530 -870
rect 74410 -970 74530 -960
rect 74750 -870 74870 -860
rect 74750 -960 74770 -870
rect 74850 -960 74870 -870
rect 74750 -970 74870 -960
rect 75090 -870 75210 -860
rect 75090 -960 75110 -870
rect 75190 -960 75210 -870
rect 75090 -970 75210 -960
rect 75430 -870 75550 -860
rect 75430 -960 75450 -870
rect 75530 -960 75550 -870
rect 75430 -970 75550 -960
rect 75770 -870 75890 -860
rect 75770 -960 75790 -870
rect 75870 -960 75890 -870
rect 75770 -970 75890 -960
rect 76110 -870 76230 -860
rect 76110 -960 76130 -870
rect 76210 -960 76230 -870
rect 76110 -970 76230 -960
rect 76450 -870 76570 -860
rect 76450 -960 76470 -870
rect 76550 -960 76570 -870
rect 76450 -970 76570 -960
rect 76790 -870 76910 -860
rect 76790 -960 76810 -870
rect 76890 -960 76910 -870
rect 76790 -970 76910 -960
rect 77130 -870 77250 -860
rect 77130 -960 77150 -870
rect 77230 -960 77250 -870
rect 77130 -970 77250 -960
rect 77470 -870 77590 -860
rect 77470 -960 77490 -870
rect 77570 -960 77590 -870
rect 77470 -970 77590 -960
rect 77810 -870 77930 -860
rect 77810 -960 77830 -870
rect 77910 -960 77930 -870
rect 77810 -970 77930 -960
rect 78150 -870 78270 -860
rect 78150 -960 78170 -870
rect 78250 -960 78270 -870
rect 78150 -970 78270 -960
rect 78490 -870 78610 -860
rect 78490 -960 78510 -870
rect 78590 -960 78610 -870
rect 78490 -970 78610 -960
rect 78830 -870 78950 -860
rect 78830 -960 78850 -870
rect 78930 -960 78950 -870
rect 78830 -970 78950 -960
rect 79170 -870 79290 -860
rect 79170 -960 79190 -870
rect 79270 -960 79290 -870
rect 79170 -970 79290 -960
rect 79510 -870 79630 -860
rect 79510 -960 79530 -870
rect 79610 -960 79630 -870
rect 79510 -970 79630 -960
rect 79850 -870 79970 -860
rect 79850 -960 79870 -870
rect 79950 -960 79970 -870
rect 79850 -970 79970 -960
rect 80190 -870 80310 -860
rect 80190 -960 80210 -870
rect 80290 -960 80310 -870
rect 80190 -970 80310 -960
rect 80530 -870 80650 -860
rect 80530 -960 80550 -870
rect 80630 -960 80650 -870
rect 80530 -970 80650 -960
rect 80870 -870 80990 -860
rect 80870 -960 80890 -870
rect 80970 -960 80990 -870
rect 80870 -970 80990 -960
rect 81210 -870 81330 -860
rect 81210 -960 81230 -870
rect 81310 -960 81330 -870
rect 81210 -970 81330 -960
rect 81550 -870 81670 -860
rect 81550 -960 81570 -870
rect 81650 -960 81670 -870
rect 81550 -970 81670 -960
rect 81890 -870 82010 -860
rect 81890 -960 81910 -870
rect 81990 -960 82010 -870
rect 81890 -970 82010 -960
rect 82230 -870 82350 -860
rect 82230 -960 82250 -870
rect 82330 -960 82350 -870
rect 82230 -970 82350 -960
rect 82570 -870 82690 -860
rect 82570 -960 82590 -870
rect 82670 -960 82690 -870
rect 82570 -970 82690 -960
rect 82910 -870 83030 -860
rect 82910 -960 82930 -870
rect 83010 -960 83030 -870
rect 82910 -970 83030 -960
rect 83250 -870 83370 -860
rect 83250 -960 83270 -870
rect 83350 -960 83370 -870
rect 83250 -970 83370 -960
rect 83590 -870 83710 -860
rect 83590 -960 83610 -870
rect 83690 -960 83710 -870
rect 83590 -970 83710 -960
rect 83930 -870 84050 -860
rect 83930 -960 83950 -870
rect 84030 -960 84050 -870
rect 83930 -970 84050 -960
rect 84270 -870 84390 -860
rect 84270 -960 84290 -870
rect 84370 -960 84390 -870
rect 84270 -970 84390 -960
rect 84610 -870 84730 -860
rect 84610 -960 84630 -870
rect 84710 -960 84730 -870
rect 84610 -970 84730 -960
rect 84950 -870 85070 -860
rect 84950 -960 84970 -870
rect 85050 -960 85070 -870
rect 84950 -970 85070 -960
rect 85290 -870 85410 -860
rect 85290 -960 85310 -870
rect 85390 -960 85410 -870
rect 85290 -970 85410 -960
rect 85630 -870 85750 -860
rect 85630 -960 85650 -870
rect 85730 -960 85750 -870
rect 85630 -970 85750 -960
rect 85970 -870 86090 -860
rect 85970 -960 85990 -870
rect 86070 -960 86090 -870
rect 85970 -970 86090 -960
rect 86310 -870 86430 -860
rect 86310 -960 86330 -870
rect 86410 -960 86430 -870
rect 86310 -970 86430 -960
rect 86650 -870 86770 -860
rect 86650 -960 86670 -870
rect 86750 -960 86770 -870
rect 86650 -970 86770 -960
rect 86990 -870 87110 -860
rect 86990 -960 87010 -870
rect 87090 -960 87110 -870
rect 86990 -970 87110 -960
rect 130 -1100 230 -1080
rect 130 -1160 150 -1100
rect 210 -1160 230 -1100
rect 130 -1300 230 -1160
rect 130 -1360 150 -1300
rect 210 -1360 230 -1300
rect 130 -1420 230 -1360
rect 1490 -1100 1590 -1080
rect 1490 -1160 1510 -1100
rect 1570 -1160 1590 -1100
rect 1490 -1300 1590 -1160
rect 1490 -1360 1510 -1300
rect 1570 -1360 1590 -1300
rect 1490 -1420 1590 -1360
rect 2850 -1100 2950 -1080
rect 2850 -1160 2870 -1100
rect 2930 -1160 2950 -1100
rect 2850 -1300 2950 -1160
rect 2850 -1360 2870 -1300
rect 2930 -1360 2950 -1300
rect 2850 -1420 2950 -1360
rect 4210 -1100 4310 -1080
rect 4210 -1160 4230 -1100
rect 4290 -1160 4310 -1100
rect 4210 -1300 4310 -1160
rect 4210 -1360 4230 -1300
rect 4290 -1360 4310 -1300
rect 4210 -1420 4310 -1360
rect 5570 -1100 5670 -1080
rect 5570 -1160 5590 -1100
rect 5650 -1160 5670 -1100
rect 5570 -1300 5670 -1160
rect 5570 -1360 5590 -1300
rect 5650 -1360 5670 -1300
rect 5570 -1420 5670 -1360
rect 6930 -1100 7030 -1080
rect 6930 -1160 6950 -1100
rect 7010 -1160 7030 -1100
rect 6930 -1300 7030 -1160
rect 6930 -1360 6950 -1300
rect 7010 -1360 7030 -1300
rect 6930 -1420 7030 -1360
rect 8290 -1100 8390 -1080
rect 8290 -1160 8310 -1100
rect 8370 -1160 8390 -1100
rect 8290 -1300 8390 -1160
rect 8290 -1360 8310 -1300
rect 8370 -1360 8390 -1300
rect 8290 -1420 8390 -1360
rect 9650 -1100 9750 -1080
rect 9650 -1160 9670 -1100
rect 9730 -1160 9750 -1100
rect 9650 -1300 9750 -1160
rect 9650 -1360 9670 -1300
rect 9730 -1360 9750 -1300
rect 9650 -1420 9750 -1360
rect 11010 -1100 11110 -1080
rect 11010 -1160 11030 -1100
rect 11090 -1160 11110 -1100
rect 11010 -1300 11110 -1160
rect 11010 -1360 11030 -1300
rect 11090 -1360 11110 -1300
rect 11010 -1420 11110 -1360
rect 12370 -1100 12470 -1080
rect 12370 -1160 12390 -1100
rect 12450 -1160 12470 -1100
rect 12370 -1300 12470 -1160
rect 12370 -1360 12390 -1300
rect 12450 -1360 12470 -1300
rect 12370 -1420 12470 -1360
rect 13730 -1100 13830 -1080
rect 13730 -1160 13750 -1100
rect 13810 -1160 13830 -1100
rect 13730 -1300 13830 -1160
rect 13730 -1360 13750 -1300
rect 13810 -1360 13830 -1300
rect 13730 -1420 13830 -1360
rect 15090 -1100 15190 -1080
rect 15090 -1160 15110 -1100
rect 15170 -1160 15190 -1100
rect 15090 -1300 15190 -1160
rect 15090 -1360 15110 -1300
rect 15170 -1360 15190 -1300
rect 15090 -1420 15190 -1360
rect 16450 -1100 16550 -1080
rect 16450 -1160 16470 -1100
rect 16530 -1160 16550 -1100
rect 16450 -1300 16550 -1160
rect 16450 -1360 16470 -1300
rect 16530 -1360 16550 -1300
rect 16450 -1420 16550 -1360
rect 17810 -1100 17910 -1080
rect 17810 -1160 17830 -1100
rect 17890 -1160 17910 -1100
rect 17810 -1300 17910 -1160
rect 17810 -1360 17830 -1300
rect 17890 -1360 17910 -1300
rect 17810 -1420 17910 -1360
rect 19170 -1100 19270 -1080
rect 19170 -1160 19190 -1100
rect 19250 -1160 19270 -1100
rect 19170 -1300 19270 -1160
rect 19170 -1360 19190 -1300
rect 19250 -1360 19270 -1300
rect 19170 -1420 19270 -1360
rect 20530 -1100 20630 -1080
rect 20530 -1160 20550 -1100
rect 20610 -1160 20630 -1100
rect 20530 -1300 20630 -1160
rect 20530 -1360 20550 -1300
rect 20610 -1360 20630 -1300
rect 20530 -1420 20630 -1360
rect 21890 -1100 21990 -1080
rect 21890 -1160 21910 -1100
rect 21970 -1160 21990 -1100
rect 21890 -1300 21990 -1160
rect 21890 -1360 21910 -1300
rect 21970 -1360 21990 -1300
rect 21890 -1420 21990 -1360
rect 23250 -1100 23350 -1080
rect 23250 -1160 23270 -1100
rect 23330 -1160 23350 -1100
rect 23250 -1300 23350 -1160
rect 23250 -1360 23270 -1300
rect 23330 -1360 23350 -1300
rect 23250 -1420 23350 -1360
rect 24610 -1100 24710 -1080
rect 24610 -1160 24630 -1100
rect 24690 -1160 24710 -1100
rect 24610 -1300 24710 -1160
rect 24610 -1360 24630 -1300
rect 24690 -1360 24710 -1300
rect 24610 -1420 24710 -1360
rect 25970 -1100 26070 -1080
rect 25970 -1160 25990 -1100
rect 26050 -1160 26070 -1100
rect 25970 -1300 26070 -1160
rect 25970 -1360 25990 -1300
rect 26050 -1360 26070 -1300
rect 25970 -1420 26070 -1360
rect 27330 -1100 27430 -1080
rect 27330 -1160 27350 -1100
rect 27410 -1160 27430 -1100
rect 27330 -1300 27430 -1160
rect 27330 -1360 27350 -1300
rect 27410 -1360 27430 -1300
rect 27330 -1420 27430 -1360
rect 28690 -1100 28790 -1080
rect 28690 -1160 28710 -1100
rect 28770 -1160 28790 -1100
rect 28690 -1300 28790 -1160
rect 28690 -1360 28710 -1300
rect 28770 -1360 28790 -1300
rect 28690 -1420 28790 -1360
rect 30050 -1100 30150 -1080
rect 30050 -1160 30070 -1100
rect 30130 -1160 30150 -1100
rect 30050 -1300 30150 -1160
rect 30050 -1360 30070 -1300
rect 30130 -1360 30150 -1300
rect 30050 -1420 30150 -1360
rect 31410 -1100 31510 -1080
rect 31410 -1160 31430 -1100
rect 31490 -1160 31510 -1100
rect 31410 -1300 31510 -1160
rect 31410 -1360 31430 -1300
rect 31490 -1360 31510 -1300
rect 31410 -1420 31510 -1360
rect 32770 -1100 32870 -1080
rect 32770 -1160 32790 -1100
rect 32850 -1160 32870 -1100
rect 32770 -1300 32870 -1160
rect 32770 -1360 32790 -1300
rect 32850 -1360 32870 -1300
rect 32770 -1420 32870 -1360
rect 34130 -1100 34230 -1080
rect 34130 -1160 34150 -1100
rect 34210 -1160 34230 -1100
rect 34130 -1300 34230 -1160
rect 34130 -1360 34150 -1300
rect 34210 -1360 34230 -1300
rect 34130 -1420 34230 -1360
rect 35490 -1100 35590 -1080
rect 35490 -1160 35510 -1100
rect 35570 -1160 35590 -1100
rect 35490 -1300 35590 -1160
rect 35490 -1360 35510 -1300
rect 35570 -1360 35590 -1300
rect 35490 -1420 35590 -1360
rect 36850 -1100 36950 -1080
rect 36850 -1160 36870 -1100
rect 36930 -1160 36950 -1100
rect 36850 -1300 36950 -1160
rect 36850 -1360 36870 -1300
rect 36930 -1360 36950 -1300
rect 36850 -1420 36950 -1360
rect 38210 -1100 38310 -1080
rect 38210 -1160 38230 -1100
rect 38290 -1160 38310 -1100
rect 38210 -1300 38310 -1160
rect 38210 -1360 38230 -1300
rect 38290 -1360 38310 -1300
rect 38210 -1420 38310 -1360
rect 39570 -1100 39670 -1080
rect 39570 -1160 39590 -1100
rect 39650 -1160 39670 -1100
rect 39570 -1300 39670 -1160
rect 39570 -1360 39590 -1300
rect 39650 -1360 39670 -1300
rect 39570 -1420 39670 -1360
rect 40930 -1100 41030 -1080
rect 40930 -1160 40950 -1100
rect 41010 -1160 41030 -1100
rect 40930 -1300 41030 -1160
rect 40930 -1360 40950 -1300
rect 41010 -1360 41030 -1300
rect 40930 -1420 41030 -1360
rect 42290 -1100 42390 -1080
rect 42290 -1160 42310 -1100
rect 42370 -1160 42390 -1100
rect 42290 -1300 42390 -1160
rect 42290 -1360 42310 -1300
rect 42370 -1360 42390 -1300
rect 42290 -1420 42390 -1360
rect 43650 -1100 43750 -1080
rect 43650 -1160 43670 -1100
rect 43730 -1160 43750 -1100
rect 43650 -1300 43750 -1160
rect 43650 -1360 43670 -1300
rect 43730 -1360 43750 -1300
rect 43650 -1420 43750 -1360
rect 45010 -1100 45110 -1080
rect 45010 -1160 45030 -1100
rect 45090 -1160 45110 -1100
rect 45010 -1300 45110 -1160
rect 45010 -1360 45030 -1300
rect 45090 -1360 45110 -1300
rect 45010 -1420 45110 -1360
rect 46370 -1100 46470 -1080
rect 46370 -1160 46390 -1100
rect 46450 -1160 46470 -1100
rect 46370 -1300 46470 -1160
rect 46370 -1360 46390 -1300
rect 46450 -1360 46470 -1300
rect 46370 -1420 46470 -1360
rect 47730 -1100 47830 -1080
rect 47730 -1160 47750 -1100
rect 47810 -1160 47830 -1100
rect 47730 -1300 47830 -1160
rect 47730 -1360 47750 -1300
rect 47810 -1360 47830 -1300
rect 47730 -1420 47830 -1360
rect 49090 -1100 49190 -1080
rect 49090 -1160 49110 -1100
rect 49170 -1160 49190 -1100
rect 49090 -1300 49190 -1160
rect 49090 -1360 49110 -1300
rect 49170 -1360 49190 -1300
rect 49090 -1420 49190 -1360
rect 50450 -1100 50550 -1080
rect 50450 -1160 50470 -1100
rect 50530 -1160 50550 -1100
rect 50450 -1300 50550 -1160
rect 50450 -1360 50470 -1300
rect 50530 -1360 50550 -1300
rect 50450 -1420 50550 -1360
rect 51810 -1100 51910 -1080
rect 51810 -1160 51830 -1100
rect 51890 -1160 51910 -1100
rect 51810 -1300 51910 -1160
rect 51810 -1360 51830 -1300
rect 51890 -1360 51910 -1300
rect 51810 -1420 51910 -1360
rect 53170 -1100 53270 -1080
rect 53170 -1160 53190 -1100
rect 53250 -1160 53270 -1100
rect 53170 -1300 53270 -1160
rect 53170 -1360 53190 -1300
rect 53250 -1360 53270 -1300
rect 53170 -1420 53270 -1360
rect 54530 -1100 54630 -1080
rect 54530 -1160 54550 -1100
rect 54610 -1160 54630 -1100
rect 54530 -1300 54630 -1160
rect 54530 -1360 54550 -1300
rect 54610 -1360 54630 -1300
rect 54530 -1420 54630 -1360
rect 55890 -1100 55990 -1080
rect 55890 -1160 55910 -1100
rect 55970 -1160 55990 -1100
rect 55890 -1300 55990 -1160
rect 55890 -1360 55910 -1300
rect 55970 -1360 55990 -1300
rect 55890 -1420 55990 -1360
rect 57250 -1100 57350 -1080
rect 57250 -1160 57270 -1100
rect 57330 -1160 57350 -1100
rect 57250 -1300 57350 -1160
rect 57250 -1360 57270 -1300
rect 57330 -1360 57350 -1300
rect 57250 -1420 57350 -1360
rect 58610 -1100 58710 -1080
rect 58610 -1160 58630 -1100
rect 58690 -1160 58710 -1100
rect 58610 -1300 58710 -1160
rect 58610 -1360 58630 -1300
rect 58690 -1360 58710 -1300
rect 58610 -1420 58710 -1360
rect 59970 -1100 60070 -1080
rect 59970 -1160 59990 -1100
rect 60050 -1160 60070 -1100
rect 59970 -1300 60070 -1160
rect 59970 -1360 59990 -1300
rect 60050 -1360 60070 -1300
rect 59970 -1420 60070 -1360
rect 61330 -1100 61430 -1080
rect 61330 -1160 61350 -1100
rect 61410 -1160 61430 -1100
rect 61330 -1300 61430 -1160
rect 61330 -1360 61350 -1300
rect 61410 -1360 61430 -1300
rect 61330 -1420 61430 -1360
rect 62690 -1100 62790 -1080
rect 62690 -1160 62710 -1100
rect 62770 -1160 62790 -1100
rect 62690 -1300 62790 -1160
rect 62690 -1360 62710 -1300
rect 62770 -1360 62790 -1300
rect 62690 -1420 62790 -1360
rect 64050 -1100 64150 -1080
rect 64050 -1160 64070 -1100
rect 64130 -1160 64150 -1100
rect 64050 -1300 64150 -1160
rect 64050 -1360 64070 -1300
rect 64130 -1360 64150 -1300
rect 64050 -1420 64150 -1360
rect 65410 -1100 65510 -1080
rect 65410 -1160 65430 -1100
rect 65490 -1160 65510 -1100
rect 65410 -1300 65510 -1160
rect 65410 -1360 65430 -1300
rect 65490 -1360 65510 -1300
rect 65410 -1420 65510 -1360
rect 66770 -1100 66870 -1080
rect 66770 -1160 66790 -1100
rect 66850 -1160 66870 -1100
rect 66770 -1300 66870 -1160
rect 66770 -1360 66790 -1300
rect 66850 -1360 66870 -1300
rect 66770 -1420 66870 -1360
rect 68130 -1100 68230 -1080
rect 68130 -1160 68150 -1100
rect 68210 -1160 68230 -1100
rect 68130 -1300 68230 -1160
rect 68130 -1360 68150 -1300
rect 68210 -1360 68230 -1300
rect 68130 -1420 68230 -1360
rect 69490 -1100 69590 -1080
rect 69490 -1160 69510 -1100
rect 69570 -1160 69590 -1100
rect 69490 -1300 69590 -1160
rect 69490 -1360 69510 -1300
rect 69570 -1360 69590 -1300
rect 69490 -1420 69590 -1360
rect 70850 -1100 70950 -1080
rect 70850 -1160 70870 -1100
rect 70930 -1160 70950 -1100
rect 70850 -1300 70950 -1160
rect 70850 -1360 70870 -1300
rect 70930 -1360 70950 -1300
rect 70850 -1420 70950 -1360
rect 72210 -1100 72310 -1080
rect 72210 -1160 72230 -1100
rect 72290 -1160 72310 -1100
rect 72210 -1300 72310 -1160
rect 72210 -1360 72230 -1300
rect 72290 -1360 72310 -1300
rect 72210 -1420 72310 -1360
rect 73570 -1100 73670 -1080
rect 73570 -1160 73590 -1100
rect 73650 -1160 73670 -1100
rect 73570 -1300 73670 -1160
rect 73570 -1360 73590 -1300
rect 73650 -1360 73670 -1300
rect 73570 -1420 73670 -1360
rect 74930 -1100 75030 -1080
rect 74930 -1160 74950 -1100
rect 75010 -1160 75030 -1100
rect 74930 -1300 75030 -1160
rect 74930 -1360 74950 -1300
rect 75010 -1360 75030 -1300
rect 74930 -1420 75030 -1360
rect 76290 -1100 76390 -1080
rect 76290 -1160 76310 -1100
rect 76370 -1160 76390 -1100
rect 76290 -1300 76390 -1160
rect 76290 -1360 76310 -1300
rect 76370 -1360 76390 -1300
rect 76290 -1420 76390 -1360
rect 77650 -1100 77750 -1080
rect 77650 -1160 77670 -1100
rect 77730 -1160 77750 -1100
rect 77650 -1300 77750 -1160
rect 77650 -1360 77670 -1300
rect 77730 -1360 77750 -1300
rect 77650 -1420 77750 -1360
rect 79010 -1100 79110 -1080
rect 79010 -1160 79030 -1100
rect 79090 -1160 79110 -1100
rect 79010 -1300 79110 -1160
rect 79010 -1360 79030 -1300
rect 79090 -1360 79110 -1300
rect 79010 -1420 79110 -1360
rect 80370 -1100 80470 -1080
rect 80370 -1160 80390 -1100
rect 80450 -1160 80470 -1100
rect 80370 -1300 80470 -1160
rect 80370 -1360 80390 -1300
rect 80450 -1360 80470 -1300
rect 80370 -1420 80470 -1360
rect 81730 -1100 81830 -1080
rect 81730 -1160 81750 -1100
rect 81810 -1160 81830 -1100
rect 81730 -1300 81830 -1160
rect 81730 -1360 81750 -1300
rect 81810 -1360 81830 -1300
rect 81730 -1420 81830 -1360
rect 83090 -1100 83190 -1080
rect 83090 -1160 83110 -1100
rect 83170 -1160 83190 -1100
rect 83090 -1300 83190 -1160
rect 83090 -1360 83110 -1300
rect 83170 -1360 83190 -1300
rect 83090 -1420 83190 -1360
rect 84450 -1100 84550 -1080
rect 84450 -1160 84470 -1100
rect 84530 -1160 84550 -1100
rect 84450 -1300 84550 -1160
rect 84450 -1360 84470 -1300
rect 84530 -1360 84550 -1300
rect 84450 -1420 84550 -1360
rect 85810 -1100 85910 -1080
rect 85810 -1160 85830 -1100
rect 85890 -1160 85910 -1100
rect 85810 -1300 85910 -1160
rect 85810 -1360 85830 -1300
rect 85890 -1360 85910 -1300
rect 85810 -1420 85910 -1360
rect 100 -1430 260 -1420
rect 100 -1520 120 -1430
rect 240 -1520 260 -1430
rect 1460 -1430 1620 -1420
rect 100 -1530 260 -1520
rect 770 -1470 970 -1440
rect 770 -1540 830 -1470
rect 910 -1540 970 -1470
rect 1460 -1520 1480 -1430
rect 1600 -1520 1620 -1430
rect 1460 -1530 1620 -1520
rect 2820 -1430 2980 -1420
rect 2820 -1520 2840 -1430
rect 2960 -1520 2980 -1430
rect 2820 -1530 2980 -1520
rect 4180 -1430 4340 -1420
rect 4180 -1520 4200 -1430
rect 4320 -1520 4340 -1430
rect 5540 -1430 5700 -1420
rect 4180 -1530 4340 -1520
rect 4940 -1470 5140 -1440
rect 770 -1570 970 -1540
rect 4940 -1540 5000 -1470
rect 5080 -1540 5140 -1470
rect 5540 -1520 5560 -1430
rect 5680 -1520 5700 -1430
rect 5540 -1530 5700 -1520
rect 6900 -1430 7060 -1420
rect 6900 -1520 6920 -1430
rect 7040 -1520 7060 -1430
rect 6900 -1530 7060 -1520
rect 8260 -1430 8420 -1420
rect 8260 -1520 8280 -1430
rect 8400 -1520 8420 -1430
rect 9620 -1430 9780 -1420
rect 8260 -1530 8420 -1520
rect 8970 -1470 9170 -1440
rect 4940 -1570 5140 -1540
rect 8970 -1540 9030 -1470
rect 9110 -1540 9170 -1470
rect 9620 -1520 9640 -1430
rect 9760 -1520 9780 -1430
rect 9620 -1530 9780 -1520
rect 10980 -1430 11140 -1420
rect 10980 -1520 11000 -1430
rect 11120 -1520 11140 -1430
rect 10980 -1530 11140 -1520
rect 12340 -1430 12500 -1420
rect 12340 -1520 12360 -1430
rect 12480 -1520 12500 -1430
rect 13700 -1430 13860 -1420
rect 12340 -1530 12500 -1520
rect 13000 -1470 13200 -1440
rect 8970 -1570 9170 -1540
rect 13000 -1540 13060 -1470
rect 13140 -1540 13200 -1470
rect 13700 -1520 13720 -1430
rect 13840 -1520 13860 -1430
rect 13700 -1530 13860 -1520
rect 15060 -1430 15220 -1420
rect 15060 -1520 15080 -1430
rect 15200 -1520 15220 -1430
rect 15060 -1530 15220 -1520
rect 16420 -1430 16580 -1420
rect 16420 -1520 16440 -1430
rect 16560 -1520 16580 -1430
rect 17780 -1430 17940 -1420
rect 16420 -1530 16580 -1520
rect 17040 -1470 17240 -1440
rect 13000 -1570 13200 -1540
rect 17040 -1540 17100 -1470
rect 17180 -1540 17240 -1470
rect 17780 -1520 17800 -1430
rect 17920 -1520 17940 -1430
rect 17780 -1530 17940 -1520
rect 19140 -1430 19300 -1420
rect 19140 -1520 19160 -1430
rect 19280 -1520 19300 -1430
rect 19140 -1530 19300 -1520
rect 20500 -1430 20660 -1420
rect 20500 -1520 20520 -1430
rect 20640 -1520 20660 -1430
rect 21860 -1430 22020 -1420
rect 20500 -1530 20660 -1520
rect 21140 -1470 21340 -1440
rect 17040 -1570 17240 -1540
rect 21140 -1540 21200 -1470
rect 21280 -1540 21340 -1470
rect 21860 -1520 21880 -1430
rect 22000 -1520 22020 -1430
rect 21860 -1530 22020 -1520
rect 23220 -1430 23380 -1420
rect 23220 -1520 23240 -1430
rect 23360 -1520 23380 -1430
rect 23220 -1530 23380 -1520
rect 24580 -1430 24740 -1420
rect 24580 -1520 24600 -1430
rect 24720 -1520 24740 -1430
rect 25940 -1430 26100 -1420
rect 24580 -1530 24740 -1520
rect 25250 -1470 25450 -1440
rect 21140 -1570 21340 -1540
rect 25250 -1540 25310 -1470
rect 25390 -1540 25450 -1470
rect 25940 -1520 25960 -1430
rect 26080 -1520 26100 -1430
rect 25940 -1530 26100 -1520
rect 27300 -1430 27460 -1420
rect 27300 -1520 27320 -1430
rect 27440 -1520 27460 -1430
rect 27300 -1530 27460 -1520
rect 28660 -1430 28820 -1420
rect 28660 -1520 28680 -1430
rect 28800 -1520 28820 -1430
rect 30020 -1430 30180 -1420
rect 28660 -1530 28820 -1520
rect 29350 -1470 29550 -1440
rect 25250 -1570 25450 -1540
rect 29350 -1540 29410 -1470
rect 29490 -1540 29550 -1470
rect 30020 -1520 30040 -1430
rect 30160 -1520 30180 -1430
rect 30020 -1530 30180 -1520
rect 31380 -1430 31540 -1420
rect 31380 -1520 31400 -1430
rect 31520 -1520 31540 -1430
rect 31380 -1530 31540 -1520
rect 32740 -1430 32900 -1420
rect 32740 -1520 32760 -1430
rect 32880 -1520 32900 -1430
rect 34100 -1430 34260 -1420
rect 32740 -1530 32900 -1520
rect 33380 -1470 33580 -1440
rect 29350 -1570 29550 -1540
rect 33380 -1540 33440 -1470
rect 33520 -1540 33580 -1470
rect 34100 -1520 34120 -1430
rect 34240 -1520 34260 -1430
rect 34100 -1530 34260 -1520
rect 35460 -1430 35620 -1420
rect 35460 -1520 35480 -1430
rect 35600 -1520 35620 -1430
rect 35460 -1530 35620 -1520
rect 36820 -1430 36980 -1420
rect 36820 -1520 36840 -1430
rect 36960 -1520 36980 -1430
rect 38180 -1430 38340 -1420
rect 36820 -1530 36980 -1520
rect 37490 -1470 37690 -1440
rect 33380 -1570 33580 -1540
rect 37490 -1540 37550 -1470
rect 37630 -1540 37690 -1470
rect 38180 -1520 38200 -1430
rect 38320 -1520 38340 -1430
rect 38180 -1530 38340 -1520
rect 39540 -1430 39700 -1420
rect 39540 -1520 39560 -1430
rect 39680 -1520 39700 -1430
rect 39540 -1530 39700 -1520
rect 40900 -1430 41060 -1420
rect 40900 -1520 40920 -1430
rect 41040 -1520 41060 -1430
rect 42260 -1430 42420 -1420
rect 40900 -1530 41060 -1520
rect 41590 -1470 41790 -1440
rect 37490 -1570 37690 -1540
rect 41590 -1540 41650 -1470
rect 41730 -1540 41790 -1470
rect 42260 -1520 42280 -1430
rect 42400 -1520 42420 -1430
rect 42260 -1530 42420 -1520
rect 43630 -1430 43780 -1420
rect 43630 -1520 43640 -1430
rect 43760 -1520 43780 -1430
rect 43630 -1530 43780 -1520
rect 44980 -1430 45140 -1420
rect 44980 -1520 45000 -1430
rect 45120 -1520 45140 -1430
rect 44980 -1530 45140 -1520
rect 46340 -1430 46500 -1420
rect 46340 -1520 46360 -1430
rect 46480 -1520 46500 -1430
rect 47700 -1430 47860 -1420
rect 46340 -1530 46500 -1520
rect 47040 -1470 47240 -1440
rect 41590 -1570 41790 -1540
rect 47040 -1540 47100 -1470
rect 47180 -1540 47240 -1470
rect 47700 -1520 47720 -1430
rect 47840 -1520 47860 -1430
rect 47700 -1530 47860 -1520
rect 49060 -1430 49220 -1420
rect 49060 -1520 49080 -1430
rect 49200 -1520 49220 -1430
rect 49060 -1530 49220 -1520
rect 50420 -1430 50580 -1420
rect 50420 -1520 50440 -1430
rect 50560 -1520 50580 -1430
rect 51780 -1430 51940 -1420
rect 50420 -1530 50580 -1520
rect 51120 -1470 51320 -1440
rect 47040 -1570 47240 -1540
rect 51120 -1540 51180 -1470
rect 51260 -1540 51320 -1470
rect 51780 -1520 51800 -1430
rect 51920 -1520 51940 -1430
rect 51780 -1530 51940 -1520
rect 53140 -1430 53300 -1420
rect 53140 -1520 53160 -1430
rect 53280 -1520 53300 -1430
rect 53140 -1530 53300 -1520
rect 54500 -1430 54660 -1420
rect 54500 -1520 54520 -1430
rect 54640 -1520 54660 -1430
rect 55860 -1430 56020 -1420
rect 54500 -1530 54660 -1520
rect 55230 -1470 55430 -1440
rect 51120 -1570 51320 -1540
rect 55230 -1540 55290 -1470
rect 55370 -1540 55430 -1470
rect 55860 -1520 55880 -1430
rect 56000 -1520 56020 -1430
rect 55860 -1530 56020 -1520
rect 57220 -1430 57380 -1420
rect 57220 -1520 57240 -1430
rect 57360 -1520 57380 -1430
rect 57220 -1530 57380 -1520
rect 58580 -1430 58740 -1420
rect 58580 -1520 58600 -1430
rect 58720 -1520 58740 -1430
rect 59940 -1430 60100 -1420
rect 58580 -1530 58740 -1520
rect 59260 -1470 59460 -1440
rect 55230 -1570 55430 -1540
rect 59260 -1540 59320 -1470
rect 59400 -1540 59460 -1470
rect 59940 -1520 59960 -1430
rect 60080 -1520 60100 -1430
rect 59940 -1530 60100 -1520
rect 61300 -1430 61460 -1420
rect 61300 -1520 61320 -1430
rect 61440 -1520 61460 -1430
rect 61300 -1530 61460 -1520
rect 62660 -1430 62820 -1420
rect 62660 -1520 62680 -1430
rect 62800 -1520 62820 -1430
rect 64020 -1430 64180 -1420
rect 62660 -1530 62820 -1520
rect 63360 -1470 63560 -1440
rect 59260 -1570 59460 -1540
rect 63360 -1540 63420 -1470
rect 63500 -1540 63560 -1470
rect 64020 -1520 64040 -1430
rect 64160 -1520 64180 -1430
rect 64020 -1530 64180 -1520
rect 65380 -1430 65540 -1420
rect 65380 -1520 65400 -1430
rect 65520 -1520 65540 -1430
rect 65380 -1530 65540 -1520
rect 66740 -1430 66900 -1420
rect 66740 -1520 66760 -1430
rect 66880 -1520 66900 -1430
rect 68100 -1430 68260 -1420
rect 66740 -1530 66900 -1520
rect 67470 -1470 67670 -1440
rect 63360 -1570 63560 -1540
rect 67470 -1540 67530 -1470
rect 67610 -1540 67670 -1470
rect 68100 -1520 68120 -1430
rect 68240 -1520 68260 -1430
rect 68100 -1530 68260 -1520
rect 69460 -1430 69620 -1420
rect 69460 -1520 69480 -1430
rect 69600 -1520 69620 -1430
rect 69460 -1530 69620 -1520
rect 70820 -1430 70980 -1420
rect 70820 -1520 70840 -1430
rect 70960 -1520 70980 -1430
rect 72180 -1430 72340 -1420
rect 70820 -1530 70980 -1520
rect 71500 -1470 71700 -1440
rect 67470 -1570 67670 -1540
rect 71500 -1540 71560 -1470
rect 71640 -1540 71700 -1470
rect 72180 -1520 72200 -1430
rect 72320 -1520 72340 -1430
rect 72180 -1530 72340 -1520
rect 73540 -1430 73700 -1420
rect 73540 -1520 73560 -1430
rect 73680 -1520 73700 -1430
rect 73540 -1530 73700 -1520
rect 74900 -1430 75060 -1420
rect 74900 -1520 74920 -1430
rect 75040 -1520 75060 -1430
rect 76260 -1430 76420 -1420
rect 74900 -1530 75060 -1520
rect 75750 -1470 75950 -1440
rect 71500 -1570 71700 -1540
rect 75750 -1540 75810 -1470
rect 75890 -1540 75950 -1470
rect 76260 -1520 76280 -1430
rect 76400 -1520 76420 -1430
rect 76260 -1530 76420 -1520
rect 77620 -1430 77780 -1420
rect 77620 -1520 77640 -1430
rect 77760 -1520 77780 -1430
rect 77620 -1530 77780 -1520
rect 78980 -1430 79140 -1420
rect 78980 -1520 79000 -1430
rect 79120 -1520 79140 -1430
rect 80340 -1430 80500 -1420
rect 78980 -1530 79140 -1520
rect 79710 -1470 79910 -1440
rect 75750 -1570 75950 -1540
rect 79710 -1540 79770 -1470
rect 79850 -1540 79910 -1470
rect 80340 -1520 80360 -1430
rect 80480 -1520 80500 -1430
rect 80340 -1530 80500 -1520
rect 81700 -1430 81860 -1420
rect 81700 -1520 81720 -1430
rect 81840 -1520 81860 -1430
rect 81700 -1530 81860 -1520
rect 83060 -1430 83220 -1420
rect 83060 -1520 83080 -1430
rect 83200 -1520 83220 -1430
rect 84420 -1430 84580 -1420
rect 83060 -1530 83220 -1520
rect 83890 -1470 84090 -1440
rect 79710 -1570 79910 -1540
rect 83890 -1540 83950 -1470
rect 84030 -1540 84090 -1470
rect 84420 -1520 84440 -1430
rect 84560 -1520 84580 -1430
rect 84420 -1530 84580 -1520
rect 85780 -1430 85940 -1420
rect 85780 -1520 85800 -1430
rect 85920 -1520 85940 -1430
rect 85780 -1530 85940 -1520
rect 86450 -1474 86648 -1444
rect 83890 -1570 84090 -1540
rect 86450 -1544 86508 -1474
rect 86588 -1544 86648 -1474
rect 86450 -1572 86648 -1544
<< via3 >>
rect 0 530 120 620
rect 420 480 540 570
rect 790 520 870 590
rect 1090 480 1190 570
rect 610 200 690 210
rect 610 130 620 200
rect 620 130 680 200
rect 680 130 690 200
rect 610 120 690 130
rect 950 200 1030 210
rect 950 130 960 200
rect 960 130 1020 200
rect 1020 130 1030 200
rect 950 120 1030 130
rect 1490 480 1610 570
rect 2170 520 2250 590
rect 2850 480 2970 570
rect 3550 520 3630 590
rect 4210 480 4330 570
rect 4510 480 4630 570
rect 5210 520 5290 590
rect 5870 480 5990 570
rect 1290 120 1400 210
rect 1680 200 1760 210
rect 1680 130 1690 200
rect 1690 130 1750 200
rect 1750 130 1760 200
rect 1680 120 1760 130
rect 2020 200 2100 210
rect 2020 130 2030 200
rect 2030 130 2090 200
rect 2090 130 2100 200
rect 2020 120 2100 130
rect 2360 200 2440 210
rect 2360 130 2370 200
rect 2370 130 2430 200
rect 2430 130 2440 200
rect 2360 120 2440 130
rect 2700 200 2780 210
rect 2700 130 2710 200
rect 2710 130 2770 200
rect 2770 130 2780 200
rect 2700 120 2780 130
rect 3040 200 3120 210
rect 3040 130 3050 200
rect 3050 130 3110 200
rect 3110 130 3120 200
rect 3040 120 3120 130
rect 3380 200 3460 210
rect 3380 130 3390 200
rect 3390 130 3450 200
rect 3450 130 3460 200
rect 3380 120 3460 130
rect 3720 200 3800 210
rect 3720 130 3730 200
rect 3730 130 3790 200
rect 3790 130 3800 200
rect 3720 120 3800 130
rect 4060 200 4140 210
rect 4060 130 4070 200
rect 4070 130 4130 200
rect 4130 130 4140 200
rect 4060 120 4140 130
rect 7230 480 7350 570
rect 8040 520 8120 590
rect 8590 480 8710 570
rect 9950 480 10070 570
rect 10800 520 10880 590
rect 11310 480 11430 570
rect 12670 480 12790 570
rect 13430 520 13510 590
rect 14030 480 14150 570
rect 15390 480 15510 570
rect 15690 480 15810 570
rect 16470 520 16550 590
rect 17050 480 17170 570
rect 18410 480 18530 570
rect 19770 480 19890 570
rect 20540 520 20620 590
rect 21130 480 21250 570
rect 22490 480 22610 570
rect 23850 480 23970 570
rect 24680 520 24760 590
rect 25210 480 25330 570
rect 26570 480 26690 570
rect 27930 480 28050 570
rect 28760 520 28840 590
rect 29290 480 29410 570
rect 30650 480 30770 570
rect 32010 480 32130 570
rect 32910 520 32990 590
rect 33370 480 33490 570
rect 34730 480 34850 570
rect 36090 480 36210 570
rect 36780 520 36860 590
rect 37450 480 37570 570
rect 38810 480 38930 570
rect 40170 480 40290 570
rect 40920 520 41000 590
rect 41530 480 41650 570
rect 42890 480 43010 570
rect 44250 480 44370 570
rect 44910 520 44990 590
rect 45610 480 45730 570
rect 46970 480 47090 570
rect 48330 480 48450 570
rect 48990 520 49070 590
rect 49690 480 49810 570
rect 51050 480 51170 570
rect 52410 480 52530 570
rect 53080 520 53160 590
rect 53770 480 53890 570
rect 55130 480 55250 570
rect 56490 480 56610 570
rect 57240 520 57320 590
rect 57850 480 57970 570
rect 59210 480 59330 570
rect 4370 120 4480 210
rect 4700 200 4780 210
rect 4700 130 4710 200
rect 4710 130 4770 200
rect 4770 130 4780 200
rect 4700 120 4780 130
rect 5040 200 5120 210
rect 5040 130 5050 200
rect 5050 130 5110 200
rect 5110 130 5120 200
rect 5040 120 5120 130
rect 5380 200 5460 210
rect 5380 130 5390 200
rect 5390 130 5450 200
rect 5450 130 5460 200
rect 5380 120 5460 130
rect 5720 200 5800 210
rect 5720 130 5730 200
rect 5730 130 5790 200
rect 5790 130 5800 200
rect 5720 120 5800 130
rect 6060 200 6140 210
rect 6060 130 6070 200
rect 6070 130 6130 200
rect 6130 130 6140 200
rect 6060 120 6140 130
rect 6400 200 6480 210
rect 6400 130 6410 200
rect 6410 130 6470 200
rect 6470 130 6480 200
rect 6400 120 6480 130
rect 6740 200 6820 210
rect 6740 130 6750 200
rect 6750 130 6810 200
rect 6810 130 6820 200
rect 6740 120 6820 130
rect 7080 200 7160 210
rect 7080 130 7090 200
rect 7090 130 7150 200
rect 7150 130 7160 200
rect 7080 120 7160 130
rect 7420 200 7500 210
rect 7420 130 7430 200
rect 7430 130 7490 200
rect 7490 130 7500 200
rect 7420 120 7500 130
rect 7760 200 7840 210
rect 7760 130 7770 200
rect 7770 130 7830 200
rect 7830 130 7840 200
rect 7760 120 7840 130
rect 8100 200 8180 210
rect 8100 130 8110 200
rect 8110 130 8170 200
rect 8170 130 8180 200
rect 8100 120 8180 130
rect 8440 200 8520 210
rect 8440 130 8450 200
rect 8450 130 8510 200
rect 8510 130 8520 200
rect 8440 120 8520 130
rect 8780 200 8860 210
rect 8780 130 8790 200
rect 8790 130 8850 200
rect 8850 130 8860 200
rect 8780 120 8860 130
rect 9120 200 9200 210
rect 9120 130 9130 200
rect 9130 130 9190 200
rect 9190 130 9200 200
rect 9120 120 9200 130
rect 9460 200 9540 210
rect 9460 130 9470 200
rect 9470 130 9530 200
rect 9530 130 9540 200
rect 9460 120 9540 130
rect 9800 200 9880 210
rect 9800 130 9810 200
rect 9810 130 9870 200
rect 9870 130 9880 200
rect 9800 120 9880 130
rect 10140 200 10220 210
rect 10140 130 10150 200
rect 10150 130 10210 200
rect 10210 130 10220 200
rect 10140 120 10220 130
rect 10480 200 10560 210
rect 10480 130 10490 200
rect 10490 130 10550 200
rect 10550 130 10560 200
rect 10480 120 10560 130
rect 10820 200 10900 210
rect 10820 130 10830 200
rect 10830 130 10890 200
rect 10890 130 10900 200
rect 10820 120 10900 130
rect 11160 200 11240 210
rect 11160 130 11170 200
rect 11170 130 11230 200
rect 11230 130 11240 200
rect 11160 120 11240 130
rect 11500 200 11580 210
rect 11500 130 11510 200
rect 11510 130 11570 200
rect 11570 130 11580 200
rect 11500 120 11580 130
rect 11840 200 11920 210
rect 11840 130 11850 200
rect 11850 130 11910 200
rect 11910 130 11920 200
rect 11840 120 11920 130
rect 12180 200 12260 210
rect 12180 130 12190 200
rect 12190 130 12250 200
rect 12250 130 12260 200
rect 12180 120 12260 130
rect 12520 200 12600 210
rect 12520 130 12530 200
rect 12530 130 12590 200
rect 12590 130 12600 200
rect 12520 120 12600 130
rect 12860 200 12940 210
rect 12860 130 12870 200
rect 12870 130 12930 200
rect 12930 130 12940 200
rect 12860 120 12940 130
rect 13200 200 13280 210
rect 13200 130 13210 200
rect 13210 130 13270 200
rect 13270 130 13280 200
rect 13200 120 13280 130
rect 13540 200 13620 210
rect 13540 130 13550 200
rect 13550 130 13610 200
rect 13610 130 13620 200
rect 13540 120 13620 130
rect 13880 200 13960 210
rect 13880 130 13890 200
rect 13890 130 13950 200
rect 13950 130 13960 200
rect 13880 120 13960 130
rect 14220 200 14300 210
rect 14220 130 14230 200
rect 14230 130 14290 200
rect 14290 130 14300 200
rect 14220 120 14300 130
rect 14560 200 14640 210
rect 14560 130 14570 200
rect 14570 130 14630 200
rect 14630 130 14640 200
rect 14560 120 14640 130
rect 14900 200 14980 210
rect 14900 130 14910 200
rect 14910 130 14970 200
rect 14970 130 14980 200
rect 14900 120 14980 130
rect 15240 200 15320 210
rect 15240 130 15250 200
rect 15250 130 15310 200
rect 15310 130 15320 200
rect 15240 120 15320 130
rect 15550 120 15660 210
rect 0 -370 100 -270
rect 130 -370 230 -270
rect 430 -380 530 -280
rect 1110 -380 1210 -280
rect 1490 -370 1590 -270
rect 2120 -390 2350 -260
rect 2860 -380 2960 -280
rect 4550 -380 4650 -280
rect 4860 -370 4960 -270
rect 5138 -398 5368 -268
rect 5910 -370 6010 -270
rect 6220 -370 6320 -270
rect 6930 -370 7030 -270
rect 7240 -380 7340 -280
rect 7624 -398 7854 -268
rect 8290 -380 8390 -280
rect 8600 -370 8700 -270
rect 9044 -398 9274 -268
rect 9650 -370 9750 -270
rect 9960 -370 10060 -270
rect 15880 200 15960 210
rect 15880 130 15890 200
rect 15890 130 15950 200
rect 15950 130 15960 200
rect 15880 120 15960 130
rect 16220 200 16300 210
rect 16220 130 16230 200
rect 16230 130 16290 200
rect 16290 130 16300 200
rect 16220 120 16300 130
rect 16560 200 16640 210
rect 16560 130 16570 200
rect 16570 130 16630 200
rect 16630 130 16640 200
rect 16560 120 16640 130
rect 16900 200 16980 210
rect 16900 130 16910 200
rect 16910 130 16970 200
rect 16970 130 16980 200
rect 16900 120 16980 130
rect 17240 200 17320 210
rect 17240 130 17250 200
rect 17250 130 17310 200
rect 17310 130 17320 200
rect 17240 120 17320 130
rect 17580 200 17660 210
rect 17580 130 17590 200
rect 17590 130 17650 200
rect 17650 130 17660 200
rect 17580 120 17660 130
rect 17920 200 18000 210
rect 17920 130 17930 200
rect 17930 130 17990 200
rect 17990 130 18000 200
rect 17920 120 18000 130
rect 18260 200 18340 210
rect 18260 130 18270 200
rect 18270 130 18330 200
rect 18330 130 18340 200
rect 18260 120 18340 130
rect 18600 200 18680 210
rect 18600 130 18610 200
rect 18610 130 18670 200
rect 18670 130 18680 200
rect 18600 120 18680 130
rect 18940 200 19020 210
rect 18940 130 18950 200
rect 18950 130 19010 200
rect 19010 130 19020 200
rect 18940 120 19020 130
rect 19280 200 19360 210
rect 19280 130 19290 200
rect 19290 130 19350 200
rect 19350 130 19360 200
rect 19280 120 19360 130
rect 19620 200 19700 210
rect 19620 130 19630 200
rect 19630 130 19690 200
rect 19690 130 19700 200
rect 19620 120 19700 130
rect 19960 200 20040 210
rect 19960 130 19970 200
rect 19970 130 20030 200
rect 20030 130 20040 200
rect 19960 120 20040 130
rect 20300 200 20380 210
rect 20300 130 20310 200
rect 20310 130 20370 200
rect 20370 130 20380 200
rect 20300 120 20380 130
rect 20640 200 20720 210
rect 20640 130 20650 200
rect 20650 130 20710 200
rect 20710 130 20720 200
rect 20640 120 20720 130
rect 20980 200 21060 210
rect 20980 130 20990 200
rect 20990 130 21050 200
rect 21050 130 21060 200
rect 20980 120 21060 130
rect 21320 200 21400 210
rect 21320 130 21330 200
rect 21330 130 21390 200
rect 21390 130 21400 200
rect 21320 120 21400 130
rect 21660 200 21740 210
rect 21660 130 21670 200
rect 21670 130 21730 200
rect 21730 130 21740 200
rect 21660 120 21740 130
rect 22000 200 22080 210
rect 22000 130 22010 200
rect 22010 130 22070 200
rect 22070 130 22080 200
rect 22000 120 22080 130
rect 22340 200 22420 210
rect 22340 130 22350 200
rect 22350 130 22410 200
rect 22410 130 22420 200
rect 22340 120 22420 130
rect 22680 200 22760 210
rect 22680 130 22690 200
rect 22690 130 22750 200
rect 22750 130 22760 200
rect 22680 120 22760 130
rect 23020 200 23100 210
rect 23020 130 23030 200
rect 23030 130 23090 200
rect 23090 130 23100 200
rect 23020 120 23100 130
rect 23360 200 23440 210
rect 23360 130 23370 200
rect 23370 130 23430 200
rect 23430 130 23440 200
rect 23360 120 23440 130
rect 23700 200 23780 210
rect 23700 130 23710 200
rect 23710 130 23770 200
rect 23770 130 23780 200
rect 23700 120 23780 130
rect 24040 200 24120 210
rect 24040 130 24050 200
rect 24050 130 24110 200
rect 24110 130 24120 200
rect 24040 120 24120 130
rect 24380 200 24460 210
rect 24380 130 24390 200
rect 24390 130 24450 200
rect 24450 130 24460 200
rect 24380 120 24460 130
rect 24720 200 24800 210
rect 24720 130 24730 200
rect 24730 130 24790 200
rect 24790 130 24800 200
rect 24720 120 24800 130
rect 25060 200 25140 210
rect 25060 130 25070 200
rect 25070 130 25130 200
rect 25130 130 25140 200
rect 25060 120 25140 130
rect 25400 200 25480 210
rect 25400 130 25410 200
rect 25410 130 25470 200
rect 25470 130 25480 200
rect 25400 120 25480 130
rect 25740 200 25820 210
rect 25740 130 25750 200
rect 25750 130 25810 200
rect 25810 130 25820 200
rect 25740 120 25820 130
rect 26080 200 26160 210
rect 26080 130 26090 200
rect 26090 130 26150 200
rect 26150 130 26160 200
rect 26080 120 26160 130
rect 26420 200 26500 210
rect 26420 130 26430 200
rect 26430 130 26490 200
rect 26490 130 26500 200
rect 26420 120 26500 130
rect 26760 200 26840 210
rect 26760 130 26770 200
rect 26770 130 26830 200
rect 26830 130 26840 200
rect 26760 120 26840 130
rect 27100 200 27180 210
rect 27100 130 27110 200
rect 27110 130 27170 200
rect 27170 130 27180 200
rect 27100 120 27180 130
rect 27440 200 27520 210
rect 27440 130 27450 200
rect 27450 130 27510 200
rect 27510 130 27520 200
rect 27440 120 27520 130
rect 27780 200 27860 210
rect 27780 130 27790 200
rect 27790 130 27850 200
rect 27850 130 27860 200
rect 27780 120 27860 130
rect 28120 200 28200 210
rect 28120 130 28130 200
rect 28130 130 28190 200
rect 28190 130 28200 200
rect 28120 120 28200 130
rect 28460 200 28540 210
rect 28460 130 28470 200
rect 28470 130 28530 200
rect 28530 130 28540 200
rect 28460 120 28540 130
rect 28800 200 28880 210
rect 28800 130 28810 200
rect 28810 130 28870 200
rect 28870 130 28880 200
rect 28800 120 28880 130
rect 29140 200 29220 210
rect 29140 130 29150 200
rect 29150 130 29210 200
rect 29210 130 29220 200
rect 29140 120 29220 130
rect 29480 200 29560 210
rect 29480 130 29490 200
rect 29490 130 29550 200
rect 29550 130 29560 200
rect 29480 120 29560 130
rect 29820 200 29900 210
rect 29820 130 29830 200
rect 29830 130 29890 200
rect 29890 130 29900 200
rect 29820 120 29900 130
rect 30160 200 30240 210
rect 30160 130 30170 200
rect 30170 130 30230 200
rect 30230 130 30240 200
rect 30160 120 30240 130
rect 30500 200 30580 210
rect 30500 130 30510 200
rect 30510 130 30570 200
rect 30570 130 30580 200
rect 30500 120 30580 130
rect 30840 200 30920 210
rect 30840 130 30850 200
rect 30850 130 30910 200
rect 30910 130 30920 200
rect 30840 120 30920 130
rect 31180 200 31260 210
rect 31180 130 31190 200
rect 31190 130 31250 200
rect 31250 130 31260 200
rect 31180 120 31260 130
rect 31520 200 31600 210
rect 31520 130 31530 200
rect 31530 130 31590 200
rect 31590 130 31600 200
rect 31520 120 31600 130
rect 31860 200 31940 210
rect 31860 130 31870 200
rect 31870 130 31930 200
rect 31930 130 31940 200
rect 31860 120 31940 130
rect 32200 200 32280 210
rect 32200 130 32210 200
rect 32210 130 32270 200
rect 32270 130 32280 200
rect 32200 120 32280 130
rect 32540 200 32620 210
rect 32540 130 32550 200
rect 32550 130 32610 200
rect 32610 130 32620 200
rect 32540 120 32620 130
rect 32880 200 32960 210
rect 32880 130 32890 200
rect 32890 130 32950 200
rect 32950 130 32960 200
rect 32880 120 32960 130
rect 33220 200 33300 210
rect 33220 130 33230 200
rect 33230 130 33290 200
rect 33290 130 33300 200
rect 33220 120 33300 130
rect 33560 200 33640 210
rect 33560 130 33570 200
rect 33570 130 33630 200
rect 33630 130 33640 200
rect 33560 120 33640 130
rect 33900 200 33980 210
rect 33900 130 33910 200
rect 33910 130 33970 200
rect 33970 130 33980 200
rect 33900 120 33980 130
rect 34240 200 34320 210
rect 34240 130 34250 200
rect 34250 130 34310 200
rect 34310 130 34320 200
rect 34240 120 34320 130
rect 34580 200 34660 210
rect 34580 130 34590 200
rect 34590 130 34650 200
rect 34650 130 34660 200
rect 34580 120 34660 130
rect 34920 200 35000 210
rect 34920 130 34930 200
rect 34930 130 34990 200
rect 34990 130 35000 200
rect 34920 120 35000 130
rect 35260 200 35340 210
rect 35260 130 35270 200
rect 35270 130 35330 200
rect 35330 130 35340 200
rect 35260 120 35340 130
rect 35600 200 35680 210
rect 35600 130 35610 200
rect 35610 130 35670 200
rect 35670 130 35680 200
rect 35600 120 35680 130
rect 35940 200 36020 210
rect 35940 130 35950 200
rect 35950 130 36010 200
rect 36010 130 36020 200
rect 35940 120 36020 130
rect 36280 200 36360 210
rect 36280 130 36290 200
rect 36290 130 36350 200
rect 36350 130 36360 200
rect 36280 120 36360 130
rect 36620 200 36700 210
rect 36620 130 36630 200
rect 36630 130 36690 200
rect 36690 130 36700 200
rect 36620 120 36700 130
rect 36960 200 37040 210
rect 36960 130 36970 200
rect 36970 130 37030 200
rect 37030 130 37040 200
rect 36960 120 37040 130
rect 37300 200 37380 210
rect 37300 130 37310 200
rect 37310 130 37370 200
rect 37370 130 37380 200
rect 37300 120 37380 130
rect 37640 200 37720 210
rect 37640 130 37650 200
rect 37650 130 37710 200
rect 37710 130 37720 200
rect 37640 120 37720 130
rect 37980 200 38060 210
rect 37980 130 37990 200
rect 37990 130 38050 200
rect 38050 130 38060 200
rect 37980 120 38060 130
rect 38320 200 38400 210
rect 38320 130 38330 200
rect 38330 130 38390 200
rect 38390 130 38400 200
rect 38320 120 38400 130
rect 38660 200 38740 210
rect 38660 130 38670 200
rect 38670 130 38730 200
rect 38730 130 38740 200
rect 38660 120 38740 130
rect 39000 200 39080 210
rect 39000 130 39010 200
rect 39010 130 39070 200
rect 39070 130 39080 200
rect 39000 120 39080 130
rect 39340 200 39420 210
rect 39340 130 39350 200
rect 39350 130 39410 200
rect 39410 130 39420 200
rect 39340 120 39420 130
rect 39680 200 39760 210
rect 39680 130 39690 200
rect 39690 130 39750 200
rect 39750 130 39760 200
rect 39680 120 39760 130
rect 40020 200 40100 210
rect 40020 130 40030 200
rect 40030 130 40090 200
rect 40090 130 40100 200
rect 40020 120 40100 130
rect 40360 200 40440 210
rect 40360 130 40370 200
rect 40370 130 40430 200
rect 40430 130 40440 200
rect 40360 120 40440 130
rect 40700 200 40780 210
rect 40700 130 40710 200
rect 40710 130 40770 200
rect 40770 130 40780 200
rect 40700 120 40780 130
rect 41040 200 41120 210
rect 41040 130 41050 200
rect 41050 130 41110 200
rect 41110 130 41120 200
rect 41040 120 41120 130
rect 41380 200 41460 210
rect 41380 130 41390 200
rect 41390 130 41450 200
rect 41450 130 41460 200
rect 41380 120 41460 130
rect 41720 200 41800 210
rect 41720 130 41730 200
rect 41730 130 41790 200
rect 41790 130 41800 200
rect 41720 120 41800 130
rect 42060 200 42140 210
rect 42060 130 42070 200
rect 42070 130 42130 200
rect 42130 130 42140 200
rect 42060 120 42140 130
rect 42400 200 42480 210
rect 42400 130 42410 200
rect 42410 130 42470 200
rect 42470 130 42480 200
rect 42400 120 42480 130
rect 42740 200 42820 210
rect 42740 130 42750 200
rect 42750 130 42810 200
rect 42810 130 42820 200
rect 42740 120 42820 130
rect 43080 200 43160 210
rect 43080 130 43090 200
rect 43090 130 43150 200
rect 43150 130 43160 200
rect 43080 120 43160 130
rect 43420 200 43500 210
rect 43420 130 43430 200
rect 43430 130 43490 200
rect 43490 130 43500 200
rect 43420 120 43500 130
rect 43760 200 43840 210
rect 43760 130 43770 200
rect 43770 130 43830 200
rect 43830 130 43840 200
rect 43760 120 43840 130
rect 44100 200 44180 210
rect 44100 130 44110 200
rect 44110 130 44170 200
rect 44170 130 44180 200
rect 44100 120 44180 130
rect 44440 200 44520 210
rect 44440 130 44450 200
rect 44450 130 44510 200
rect 44510 130 44520 200
rect 44440 120 44520 130
rect 44780 200 44860 210
rect 44780 130 44790 200
rect 44790 130 44850 200
rect 44850 130 44860 200
rect 44780 120 44860 130
rect 45120 200 45200 210
rect 45120 130 45130 200
rect 45130 130 45190 200
rect 45190 130 45200 200
rect 45120 120 45200 130
rect 45460 200 45540 210
rect 45460 130 45470 200
rect 45470 130 45530 200
rect 45530 130 45540 200
rect 45460 120 45540 130
rect 45800 200 45880 210
rect 45800 130 45810 200
rect 45810 130 45870 200
rect 45870 130 45880 200
rect 45800 120 45880 130
rect 46140 200 46220 210
rect 46140 130 46150 200
rect 46150 130 46210 200
rect 46210 130 46220 200
rect 46140 120 46220 130
rect 46480 200 46560 210
rect 46480 130 46490 200
rect 46490 130 46550 200
rect 46550 130 46560 200
rect 46480 120 46560 130
rect 46820 200 46900 210
rect 46820 130 46830 200
rect 46830 130 46890 200
rect 46890 130 46900 200
rect 46820 120 46900 130
rect 47160 200 47240 210
rect 47160 130 47170 200
rect 47170 130 47230 200
rect 47230 130 47240 200
rect 47160 120 47240 130
rect 47500 200 47580 210
rect 47500 130 47510 200
rect 47510 130 47570 200
rect 47570 130 47580 200
rect 47500 120 47580 130
rect 47840 200 47920 210
rect 47840 130 47850 200
rect 47850 130 47910 200
rect 47910 130 47920 200
rect 47840 120 47920 130
rect 48180 200 48260 210
rect 48180 130 48190 200
rect 48190 130 48250 200
rect 48250 130 48260 200
rect 48180 120 48260 130
rect 48520 200 48600 210
rect 48520 130 48530 200
rect 48530 130 48590 200
rect 48590 130 48600 200
rect 48520 120 48600 130
rect 48860 200 48940 210
rect 48860 130 48870 200
rect 48870 130 48930 200
rect 48930 130 48940 200
rect 48860 120 48940 130
rect 49200 200 49280 210
rect 49200 130 49210 200
rect 49210 130 49270 200
rect 49270 130 49280 200
rect 49200 120 49280 130
rect 49540 200 49620 210
rect 49540 130 49550 200
rect 49550 130 49610 200
rect 49610 130 49620 200
rect 49540 120 49620 130
rect 49880 200 49960 210
rect 49880 130 49890 200
rect 49890 130 49950 200
rect 49950 130 49960 200
rect 49880 120 49960 130
rect 50220 200 50300 210
rect 50220 130 50230 200
rect 50230 130 50290 200
rect 50290 130 50300 200
rect 50220 120 50300 130
rect 50560 200 50640 210
rect 50560 130 50570 200
rect 50570 130 50630 200
rect 50630 130 50640 200
rect 50560 120 50640 130
rect 50900 200 50980 210
rect 50900 130 50910 200
rect 50910 130 50970 200
rect 50970 130 50980 200
rect 50900 120 50980 130
rect 51240 200 51320 210
rect 51240 130 51250 200
rect 51250 130 51310 200
rect 51310 130 51320 200
rect 51240 120 51320 130
rect 51580 200 51660 210
rect 51580 130 51590 200
rect 51590 130 51650 200
rect 51650 130 51660 200
rect 51580 120 51660 130
rect 51920 200 52000 210
rect 51920 130 51930 200
rect 51930 130 51990 200
rect 51990 130 52000 200
rect 51920 120 52000 130
rect 52260 200 52340 210
rect 52260 130 52270 200
rect 52270 130 52330 200
rect 52330 130 52340 200
rect 52260 120 52340 130
rect 52600 200 52680 210
rect 52600 130 52610 200
rect 52610 130 52670 200
rect 52670 130 52680 200
rect 52600 120 52680 130
rect 52940 200 53020 210
rect 52940 130 52950 200
rect 52950 130 53010 200
rect 53010 130 53020 200
rect 52940 120 53020 130
rect 53280 200 53360 210
rect 53280 130 53290 200
rect 53290 130 53350 200
rect 53350 130 53360 200
rect 53280 120 53360 130
rect 53620 200 53700 210
rect 53620 130 53630 200
rect 53630 130 53690 200
rect 53690 130 53700 200
rect 53620 120 53700 130
rect 53960 200 54040 210
rect 53960 130 53970 200
rect 53970 130 54030 200
rect 54030 130 54040 200
rect 53960 120 54040 130
rect 54300 200 54380 210
rect 54300 130 54310 200
rect 54310 130 54370 200
rect 54370 130 54380 200
rect 54300 120 54380 130
rect 54640 200 54720 210
rect 54640 130 54650 200
rect 54650 130 54710 200
rect 54710 130 54720 200
rect 54640 120 54720 130
rect 54980 200 55060 210
rect 54980 130 54990 200
rect 54990 130 55050 200
rect 55050 130 55060 200
rect 54980 120 55060 130
rect 55320 200 55400 210
rect 55320 130 55330 200
rect 55330 130 55390 200
rect 55390 130 55400 200
rect 55320 120 55400 130
rect 55660 200 55740 210
rect 55660 130 55670 200
rect 55670 130 55730 200
rect 55730 130 55740 200
rect 55660 120 55740 130
rect 56000 200 56080 210
rect 56000 130 56010 200
rect 56010 130 56070 200
rect 56070 130 56080 200
rect 56000 120 56080 130
rect 56340 200 56420 210
rect 56340 130 56350 200
rect 56350 130 56410 200
rect 56410 130 56420 200
rect 56340 120 56420 130
rect 56680 200 56760 210
rect 56680 130 56690 200
rect 56690 130 56750 200
rect 56750 130 56760 200
rect 56680 120 56760 130
rect 57020 200 57100 210
rect 57020 130 57030 200
rect 57030 130 57090 200
rect 57090 130 57100 200
rect 57020 120 57100 130
rect 57360 200 57440 210
rect 57360 130 57370 200
rect 57370 130 57430 200
rect 57430 130 57440 200
rect 57360 120 57440 130
rect 57700 200 57780 210
rect 57700 130 57710 200
rect 57710 130 57770 200
rect 57770 130 57780 200
rect 57700 120 57780 130
rect 58040 200 58120 210
rect 58040 130 58050 200
rect 58050 130 58110 200
rect 58110 130 58120 200
rect 58040 120 58120 130
rect 58380 200 58460 210
rect 58380 130 58390 200
rect 58390 130 58450 200
rect 58450 130 58460 200
rect 58380 120 58460 130
rect 58720 200 58800 210
rect 58720 130 58730 200
rect 58730 130 58790 200
rect 58790 130 58800 200
rect 58720 120 58800 130
rect 59060 200 59140 210
rect 59060 130 59070 200
rect 59070 130 59130 200
rect 59130 130 59140 200
rect 59060 120 59140 130
rect 10670 -370 10770 -270
rect 10980 -380 11080 -280
rect 11690 -370 11790 -270
rect 11990 -380 12090 -280
rect 12670 -380 12770 -280
rect 13050 -370 13150 -270
rect 13668 -394 13898 -264
rect 14420 -380 14520 -280
rect 16110 -380 16210 -280
rect 16380 -370 16480 -270
rect 16868 -394 17098 -264
rect 17470 -370 17570 -270
rect 17740 -370 17840 -270
rect 18490 -370 18590 -270
rect 18760 -380 18860 -280
rect 19850 -380 19950 -280
rect 20120 -370 20220 -270
rect 20424 -394 20654 -264
rect 21210 -370 21310 -270
rect 21480 -370 21580 -270
rect 22230 -370 22330 -270
rect 22500 -380 22600 -280
rect 23590 -370 23690 -270
rect 23860 -380 23960 -280
rect 24530 -380 24630 -280
rect 24950 -370 25050 -270
rect 25758 -394 25988 -264
rect 26320 -380 26420 -280
rect 28010 -380 28110 -280
rect 28280 -370 28380 -270
rect 28602 -394 28832 -264
rect 29370 -370 29470 -270
rect 29640 -370 29740 -270
rect 30390 -370 30490 -270
rect 30660 -380 30760 -280
rect 31750 -380 31850 -280
rect 32020 -370 32120 -270
rect 32514 -394 32744 -264
rect 33110 -370 33210 -270
rect 33380 -370 33480 -270
rect 34130 -370 34230 -270
rect 34400 -380 34500 -280
rect 34670 -394 34900 -264
rect 35490 -370 35590 -270
rect 35760 -380 35860 -280
rect 36430 -380 36530 -280
rect 36850 -370 36950 -270
rect 37492 -394 37722 -264
rect 38220 -380 38320 -280
rect 39910 -380 40010 -280
rect 40692 -394 40922 -264
rect 41270 -370 41370 -270
rect 42290 -370 42390 -270
rect 42560 -380 42660 -280
rect 43650 -380 43750 -270
rect 44600 -380 44700 -280
rect 45010 -370 45110 -270
rect 45668 -394 45898 -264
rect 46380 -380 46480 -280
rect 48070 -380 48170 -280
rect 48340 -370 48440 -270
rect 48868 -394 49098 -264
rect 49430 -370 49530 -270
rect 49700 -370 49800 -270
rect 50450 -370 50550 -270
rect 50720 -380 50820 -280
rect 51002 -394 51232 -264
rect 51810 -380 51910 -280
rect 52080 -370 52180 -270
rect 53170 -370 53270 -270
rect 53440 -370 53540 -270
rect 54190 -370 54290 -270
rect 54558 -394 54788 -264
rect 55210 -370 55310 -270
rect 55480 -380 55580 -280
rect 56570 -370 56670 -270
rect 57402 -394 57632 -264
rect 57940 -380 58040 -280
rect 59630 -380 59730 -280
rect 60990 -370 61090 -270
rect 61314 -394 61544 -264
rect 62010 -370 62110 -270
rect 63370 -380 63470 -280
rect 64158 -394 64388 -264
rect 64730 -370 64830 -270
rect 65750 -370 65850 -270
rect 67110 -370 67210 -270
rect 67714 -394 67944 -264
rect 68470 -370 68570 -270
rect 69840 -380 69940 -280
rect 70558 -394 70788 -264
rect 71530 -380 71630 -280
rect 72890 -370 72990 -270
rect 73910 -370 74010 -270
rect 74468 -394 74698 -264
rect 75270 -380 75370 -280
rect 76630 -370 76730 -270
rect 77650 -370 77750 -270
rect 78380 -394 78610 -264
rect 79010 -370 79110 -270
rect 80370 -370 80470 -270
rect 81740 -380 81840 -280
rect 82292 -394 82522 -264
rect 83430 -380 83530 -280
rect 84790 -370 84890 -270
rect 85810 -370 85910 -270
rect 86202 -394 86432 -264
rect 87170 -380 87270 -280
rect 310 -880 390 -870
rect 310 -950 320 -880
rect 320 -950 380 -880
rect 380 -950 390 -880
rect 310 -960 390 -950
rect 650 -880 730 -870
rect 650 -950 660 -880
rect 660 -950 720 -880
rect 720 -950 730 -880
rect 650 -960 730 -950
rect 990 -880 1070 -870
rect 990 -950 1000 -880
rect 1000 -950 1060 -880
rect 1060 -950 1070 -880
rect 990 -960 1070 -950
rect 1330 -880 1410 -870
rect 1330 -950 1340 -880
rect 1340 -950 1400 -880
rect 1400 -950 1410 -880
rect 1330 -960 1410 -950
rect 1670 -880 1750 -870
rect 1670 -950 1680 -880
rect 1680 -950 1740 -880
rect 1740 -950 1750 -880
rect 1670 -960 1750 -950
rect 2010 -880 2090 -870
rect 2010 -950 2020 -880
rect 2020 -950 2080 -880
rect 2080 -950 2090 -880
rect 2010 -960 2090 -950
rect 2350 -880 2430 -870
rect 2350 -950 2360 -880
rect 2360 -950 2420 -880
rect 2420 -950 2430 -880
rect 2350 -960 2430 -950
rect 2690 -880 2770 -870
rect 2690 -950 2700 -880
rect 2700 -950 2760 -880
rect 2760 -950 2770 -880
rect 2690 -960 2770 -950
rect 3030 -880 3110 -870
rect 3030 -950 3040 -880
rect 3040 -950 3100 -880
rect 3100 -950 3110 -880
rect 3030 -960 3110 -950
rect 3370 -880 3450 -870
rect 3370 -950 3380 -880
rect 3380 -950 3440 -880
rect 3440 -950 3450 -880
rect 3370 -960 3450 -950
rect 3710 -880 3790 -870
rect 3710 -950 3720 -880
rect 3720 -950 3780 -880
rect 3780 -950 3790 -880
rect 3710 -960 3790 -950
rect 4050 -880 4130 -870
rect 4050 -950 4060 -880
rect 4060 -950 4120 -880
rect 4120 -950 4130 -880
rect 4050 -960 4130 -950
rect 4390 -880 4470 -870
rect 4390 -950 4400 -880
rect 4400 -950 4460 -880
rect 4460 -950 4470 -880
rect 4390 -960 4470 -950
rect 4730 -880 4810 -870
rect 4730 -950 4740 -880
rect 4740 -950 4800 -880
rect 4800 -950 4810 -880
rect 4730 -960 4810 -950
rect 5070 -880 5150 -870
rect 5070 -950 5080 -880
rect 5080 -950 5140 -880
rect 5140 -950 5150 -880
rect 5070 -960 5150 -950
rect 5410 -880 5490 -870
rect 5410 -950 5420 -880
rect 5420 -950 5480 -880
rect 5480 -950 5490 -880
rect 5410 -960 5490 -950
rect 5750 -880 5830 -870
rect 5750 -950 5760 -880
rect 5760 -950 5820 -880
rect 5820 -950 5830 -880
rect 5750 -960 5830 -950
rect 6090 -880 6170 -870
rect 6090 -950 6100 -880
rect 6100 -950 6160 -880
rect 6160 -950 6170 -880
rect 6090 -960 6170 -950
rect 6430 -880 6510 -870
rect 6430 -950 6440 -880
rect 6440 -950 6500 -880
rect 6500 -950 6510 -880
rect 6430 -960 6510 -950
rect 6770 -880 6850 -870
rect 6770 -950 6780 -880
rect 6780 -950 6840 -880
rect 6840 -950 6850 -880
rect 6770 -960 6850 -950
rect 7110 -880 7190 -870
rect 7110 -950 7120 -880
rect 7120 -950 7180 -880
rect 7180 -950 7190 -880
rect 7110 -960 7190 -950
rect 7450 -880 7530 -870
rect 7450 -950 7460 -880
rect 7460 -950 7520 -880
rect 7520 -950 7530 -880
rect 7450 -960 7530 -950
rect 7790 -880 7870 -870
rect 7790 -950 7800 -880
rect 7800 -950 7860 -880
rect 7860 -950 7870 -880
rect 7790 -960 7870 -950
rect 8130 -880 8210 -870
rect 8130 -950 8140 -880
rect 8140 -950 8200 -880
rect 8200 -950 8210 -880
rect 8130 -960 8210 -950
rect 8470 -880 8550 -870
rect 8470 -950 8480 -880
rect 8480 -950 8540 -880
rect 8540 -950 8550 -880
rect 8470 -960 8550 -950
rect 8810 -880 8890 -870
rect 8810 -950 8820 -880
rect 8820 -950 8880 -880
rect 8880 -950 8890 -880
rect 8810 -960 8890 -950
rect 9150 -880 9230 -870
rect 9150 -950 9160 -880
rect 9160 -950 9220 -880
rect 9220 -950 9230 -880
rect 9150 -960 9230 -950
rect 9490 -880 9570 -870
rect 9490 -950 9500 -880
rect 9500 -950 9560 -880
rect 9560 -950 9570 -880
rect 9490 -960 9570 -950
rect 9830 -880 9910 -870
rect 9830 -950 9840 -880
rect 9840 -950 9900 -880
rect 9900 -950 9910 -880
rect 9830 -960 9910 -950
rect 10170 -880 10250 -870
rect 10170 -950 10180 -880
rect 10180 -950 10240 -880
rect 10240 -950 10250 -880
rect 10170 -960 10250 -950
rect 10510 -880 10590 -870
rect 10510 -950 10520 -880
rect 10520 -950 10580 -880
rect 10580 -950 10590 -880
rect 10510 -960 10590 -950
rect 10850 -880 10930 -870
rect 10850 -950 10860 -880
rect 10860 -950 10920 -880
rect 10920 -950 10930 -880
rect 10850 -960 10930 -950
rect 11190 -880 11270 -870
rect 11190 -950 11200 -880
rect 11200 -950 11260 -880
rect 11260 -950 11270 -880
rect 11190 -960 11270 -950
rect 11530 -880 11610 -870
rect 11530 -950 11540 -880
rect 11540 -950 11600 -880
rect 11600 -950 11610 -880
rect 11530 -960 11610 -950
rect 11870 -880 11950 -870
rect 11870 -950 11880 -880
rect 11880 -950 11940 -880
rect 11940 -950 11950 -880
rect 11870 -960 11950 -950
rect 12210 -880 12290 -870
rect 12210 -950 12220 -880
rect 12220 -950 12280 -880
rect 12280 -950 12290 -880
rect 12210 -960 12290 -950
rect 12550 -880 12630 -870
rect 12550 -950 12560 -880
rect 12560 -950 12620 -880
rect 12620 -950 12630 -880
rect 12550 -960 12630 -950
rect 12890 -880 12970 -870
rect 12890 -950 12900 -880
rect 12900 -950 12960 -880
rect 12960 -950 12970 -880
rect 12890 -960 12970 -950
rect 13230 -880 13310 -870
rect 13230 -950 13240 -880
rect 13240 -950 13300 -880
rect 13300 -950 13310 -880
rect 13230 -960 13310 -950
rect 13570 -880 13650 -870
rect 13570 -950 13580 -880
rect 13580 -950 13640 -880
rect 13640 -950 13650 -880
rect 13570 -960 13650 -950
rect 13910 -880 13990 -870
rect 13910 -950 13920 -880
rect 13920 -950 13980 -880
rect 13980 -950 13990 -880
rect 13910 -960 13990 -950
rect 14250 -880 14330 -870
rect 14250 -950 14260 -880
rect 14260 -950 14320 -880
rect 14320 -950 14330 -880
rect 14250 -960 14330 -950
rect 14590 -880 14670 -870
rect 14590 -950 14600 -880
rect 14600 -950 14660 -880
rect 14660 -950 14670 -880
rect 14590 -960 14670 -950
rect 14930 -880 15010 -870
rect 14930 -950 14940 -880
rect 14940 -950 15000 -880
rect 15000 -950 15010 -880
rect 14930 -960 15010 -950
rect 15270 -880 15350 -870
rect 15270 -950 15280 -880
rect 15280 -950 15340 -880
rect 15340 -950 15350 -880
rect 15270 -960 15350 -950
rect 15610 -880 15690 -870
rect 15610 -950 15620 -880
rect 15620 -950 15680 -880
rect 15680 -950 15690 -880
rect 15610 -960 15690 -950
rect 15950 -880 16030 -870
rect 15950 -950 15960 -880
rect 15960 -950 16020 -880
rect 16020 -950 16030 -880
rect 15950 -960 16030 -950
rect 16290 -880 16370 -870
rect 16290 -950 16300 -880
rect 16300 -950 16360 -880
rect 16360 -950 16370 -880
rect 16290 -960 16370 -950
rect 16630 -880 16710 -870
rect 16630 -950 16640 -880
rect 16640 -950 16700 -880
rect 16700 -950 16710 -880
rect 16630 -960 16710 -950
rect 16970 -880 17050 -870
rect 16970 -950 16980 -880
rect 16980 -950 17040 -880
rect 17040 -950 17050 -880
rect 16970 -960 17050 -950
rect 17310 -880 17390 -870
rect 17310 -950 17320 -880
rect 17320 -950 17380 -880
rect 17380 -950 17390 -880
rect 17310 -960 17390 -950
rect 17650 -880 17730 -870
rect 17650 -950 17660 -880
rect 17660 -950 17720 -880
rect 17720 -950 17730 -880
rect 17650 -960 17730 -950
rect 17990 -880 18070 -870
rect 17990 -950 18000 -880
rect 18000 -950 18060 -880
rect 18060 -950 18070 -880
rect 17990 -960 18070 -950
rect 18330 -880 18410 -870
rect 18330 -950 18340 -880
rect 18340 -950 18400 -880
rect 18400 -950 18410 -880
rect 18330 -960 18410 -950
rect 18670 -880 18750 -870
rect 18670 -950 18680 -880
rect 18680 -950 18740 -880
rect 18740 -950 18750 -880
rect 18670 -960 18750 -950
rect 19010 -880 19090 -870
rect 19010 -950 19020 -880
rect 19020 -950 19080 -880
rect 19080 -950 19090 -880
rect 19010 -960 19090 -950
rect 19350 -880 19430 -870
rect 19350 -950 19360 -880
rect 19360 -950 19420 -880
rect 19420 -950 19430 -880
rect 19350 -960 19430 -950
rect 19690 -880 19770 -870
rect 19690 -950 19700 -880
rect 19700 -950 19760 -880
rect 19760 -950 19770 -880
rect 19690 -960 19770 -950
rect 20030 -880 20110 -870
rect 20030 -950 20040 -880
rect 20040 -950 20100 -880
rect 20100 -950 20110 -880
rect 20030 -960 20110 -950
rect 20370 -880 20450 -870
rect 20370 -950 20380 -880
rect 20380 -950 20440 -880
rect 20440 -950 20450 -880
rect 20370 -960 20450 -950
rect 20710 -880 20790 -870
rect 20710 -950 20720 -880
rect 20720 -950 20780 -880
rect 20780 -950 20790 -880
rect 20710 -960 20790 -950
rect 21050 -880 21130 -870
rect 21050 -950 21060 -880
rect 21060 -950 21120 -880
rect 21120 -950 21130 -880
rect 21050 -960 21130 -950
rect 21390 -880 21470 -870
rect 21390 -950 21400 -880
rect 21400 -950 21460 -880
rect 21460 -950 21470 -880
rect 21390 -960 21470 -950
rect 21730 -880 21810 -870
rect 21730 -950 21740 -880
rect 21740 -950 21800 -880
rect 21800 -950 21810 -880
rect 21730 -960 21810 -950
rect 22070 -880 22150 -870
rect 22070 -950 22080 -880
rect 22080 -950 22140 -880
rect 22140 -950 22150 -880
rect 22070 -960 22150 -950
rect 22410 -880 22490 -870
rect 22410 -950 22420 -880
rect 22420 -950 22480 -880
rect 22480 -950 22490 -880
rect 22410 -960 22490 -950
rect 22750 -880 22830 -870
rect 22750 -950 22760 -880
rect 22760 -950 22820 -880
rect 22820 -950 22830 -880
rect 22750 -960 22830 -950
rect 23090 -880 23170 -870
rect 23090 -950 23100 -880
rect 23100 -950 23160 -880
rect 23160 -950 23170 -880
rect 23090 -960 23170 -950
rect 23430 -880 23510 -870
rect 23430 -950 23440 -880
rect 23440 -950 23500 -880
rect 23500 -950 23510 -880
rect 23430 -960 23510 -950
rect 23770 -880 23850 -870
rect 23770 -950 23780 -880
rect 23780 -950 23840 -880
rect 23840 -950 23850 -880
rect 23770 -960 23850 -950
rect 24110 -880 24190 -870
rect 24110 -950 24120 -880
rect 24120 -950 24180 -880
rect 24180 -950 24190 -880
rect 24110 -960 24190 -950
rect 24450 -880 24530 -870
rect 24450 -950 24460 -880
rect 24460 -950 24520 -880
rect 24520 -950 24530 -880
rect 24450 -960 24530 -950
rect 24790 -880 24870 -870
rect 24790 -950 24800 -880
rect 24800 -950 24860 -880
rect 24860 -950 24870 -880
rect 24790 -960 24870 -950
rect 25130 -880 25210 -870
rect 25130 -950 25140 -880
rect 25140 -950 25200 -880
rect 25200 -950 25210 -880
rect 25130 -960 25210 -950
rect 25470 -880 25550 -870
rect 25470 -950 25480 -880
rect 25480 -950 25540 -880
rect 25540 -950 25550 -880
rect 25470 -960 25550 -950
rect 25810 -880 25890 -870
rect 25810 -950 25820 -880
rect 25820 -950 25880 -880
rect 25880 -950 25890 -880
rect 25810 -960 25890 -950
rect 26150 -880 26230 -870
rect 26150 -950 26160 -880
rect 26160 -950 26220 -880
rect 26220 -950 26230 -880
rect 26150 -960 26230 -950
rect 26490 -880 26570 -870
rect 26490 -950 26500 -880
rect 26500 -950 26560 -880
rect 26560 -950 26570 -880
rect 26490 -960 26570 -950
rect 26830 -880 26910 -870
rect 26830 -950 26840 -880
rect 26840 -950 26900 -880
rect 26900 -950 26910 -880
rect 26830 -960 26910 -950
rect 27170 -880 27250 -870
rect 27170 -950 27180 -880
rect 27180 -950 27240 -880
rect 27240 -950 27250 -880
rect 27170 -960 27250 -950
rect 27510 -880 27590 -870
rect 27510 -950 27520 -880
rect 27520 -950 27580 -880
rect 27580 -950 27590 -880
rect 27510 -960 27590 -950
rect 27850 -880 27930 -870
rect 27850 -950 27860 -880
rect 27860 -950 27920 -880
rect 27920 -950 27930 -880
rect 27850 -960 27930 -950
rect 28190 -880 28270 -870
rect 28190 -950 28200 -880
rect 28200 -950 28260 -880
rect 28260 -950 28270 -880
rect 28190 -960 28270 -950
rect 28530 -880 28610 -870
rect 28530 -950 28540 -880
rect 28540 -950 28600 -880
rect 28600 -950 28610 -880
rect 28530 -960 28610 -950
rect 28870 -880 28950 -870
rect 28870 -950 28880 -880
rect 28880 -950 28940 -880
rect 28940 -950 28950 -880
rect 28870 -960 28950 -950
rect 29210 -880 29290 -870
rect 29210 -950 29220 -880
rect 29220 -950 29280 -880
rect 29280 -950 29290 -880
rect 29210 -960 29290 -950
rect 29550 -880 29630 -870
rect 29550 -950 29560 -880
rect 29560 -950 29620 -880
rect 29620 -950 29630 -880
rect 29550 -960 29630 -950
rect 29890 -880 29970 -870
rect 29890 -950 29900 -880
rect 29900 -950 29960 -880
rect 29960 -950 29970 -880
rect 29890 -960 29970 -950
rect 30230 -880 30310 -870
rect 30230 -950 30240 -880
rect 30240 -950 30300 -880
rect 30300 -950 30310 -880
rect 30230 -960 30310 -950
rect 30570 -880 30650 -870
rect 30570 -950 30580 -880
rect 30580 -950 30640 -880
rect 30640 -950 30650 -880
rect 30570 -960 30650 -950
rect 30910 -880 30990 -870
rect 30910 -950 30920 -880
rect 30920 -950 30980 -880
rect 30980 -950 30990 -880
rect 30910 -960 30990 -950
rect 31250 -880 31330 -870
rect 31250 -950 31260 -880
rect 31260 -950 31320 -880
rect 31320 -950 31330 -880
rect 31250 -960 31330 -950
rect 31590 -880 31670 -870
rect 31590 -950 31600 -880
rect 31600 -950 31660 -880
rect 31660 -950 31670 -880
rect 31590 -960 31670 -950
rect 31930 -880 32010 -870
rect 31930 -950 31940 -880
rect 31940 -950 32000 -880
rect 32000 -950 32010 -880
rect 31930 -960 32010 -950
rect 32270 -880 32350 -870
rect 32270 -950 32280 -880
rect 32280 -950 32340 -880
rect 32340 -950 32350 -880
rect 32270 -960 32350 -950
rect 32610 -880 32690 -870
rect 32610 -950 32620 -880
rect 32620 -950 32680 -880
rect 32680 -950 32690 -880
rect 32610 -960 32690 -950
rect 32950 -880 33030 -870
rect 32950 -950 32960 -880
rect 32960 -950 33020 -880
rect 33020 -950 33030 -880
rect 32950 -960 33030 -950
rect 33290 -880 33370 -870
rect 33290 -950 33300 -880
rect 33300 -950 33360 -880
rect 33360 -950 33370 -880
rect 33290 -960 33370 -950
rect 33630 -880 33710 -870
rect 33630 -950 33640 -880
rect 33640 -950 33700 -880
rect 33700 -950 33710 -880
rect 33630 -960 33710 -950
rect 33970 -880 34050 -870
rect 33970 -950 33980 -880
rect 33980 -950 34040 -880
rect 34040 -950 34050 -880
rect 33970 -960 34050 -950
rect 34310 -880 34390 -870
rect 34310 -950 34320 -880
rect 34320 -950 34380 -880
rect 34380 -950 34390 -880
rect 34310 -960 34390 -950
rect 34650 -880 34730 -870
rect 34650 -950 34660 -880
rect 34660 -950 34720 -880
rect 34720 -950 34730 -880
rect 34650 -960 34730 -950
rect 34990 -880 35070 -870
rect 34990 -950 35000 -880
rect 35000 -950 35060 -880
rect 35060 -950 35070 -880
rect 34990 -960 35070 -950
rect 35330 -880 35410 -870
rect 35330 -950 35340 -880
rect 35340 -950 35400 -880
rect 35400 -950 35410 -880
rect 35330 -960 35410 -950
rect 35670 -880 35750 -870
rect 35670 -950 35680 -880
rect 35680 -950 35740 -880
rect 35740 -950 35750 -880
rect 35670 -960 35750 -950
rect 36010 -880 36090 -870
rect 36010 -950 36020 -880
rect 36020 -950 36080 -880
rect 36080 -950 36090 -880
rect 36010 -960 36090 -950
rect 36350 -880 36430 -870
rect 36350 -950 36360 -880
rect 36360 -950 36420 -880
rect 36420 -950 36430 -880
rect 36350 -960 36430 -950
rect 36690 -880 36770 -870
rect 36690 -950 36700 -880
rect 36700 -950 36760 -880
rect 36760 -950 36770 -880
rect 36690 -960 36770 -950
rect 37030 -880 37110 -870
rect 37030 -950 37040 -880
rect 37040 -950 37100 -880
rect 37100 -950 37110 -880
rect 37030 -960 37110 -950
rect 37370 -880 37450 -870
rect 37370 -950 37380 -880
rect 37380 -950 37440 -880
rect 37440 -950 37450 -880
rect 37370 -960 37450 -950
rect 37710 -880 37790 -870
rect 37710 -950 37720 -880
rect 37720 -950 37780 -880
rect 37780 -950 37790 -880
rect 37710 -960 37790 -950
rect 38050 -880 38130 -870
rect 38050 -950 38060 -880
rect 38060 -950 38120 -880
rect 38120 -950 38130 -880
rect 38050 -960 38130 -950
rect 38390 -880 38470 -870
rect 38390 -950 38400 -880
rect 38400 -950 38460 -880
rect 38460 -950 38470 -880
rect 38390 -960 38470 -950
rect 38730 -880 38810 -870
rect 38730 -950 38740 -880
rect 38740 -950 38800 -880
rect 38800 -950 38810 -880
rect 38730 -960 38810 -950
rect 39070 -880 39150 -870
rect 39070 -950 39080 -880
rect 39080 -950 39140 -880
rect 39140 -950 39150 -880
rect 39070 -960 39150 -950
rect 39410 -880 39490 -870
rect 39410 -950 39420 -880
rect 39420 -950 39480 -880
rect 39480 -950 39490 -880
rect 39410 -960 39490 -950
rect 39750 -880 39830 -870
rect 39750 -950 39760 -880
rect 39760 -950 39820 -880
rect 39820 -950 39830 -880
rect 39750 -960 39830 -950
rect 40090 -880 40170 -870
rect 40090 -950 40100 -880
rect 40100 -950 40160 -880
rect 40160 -950 40170 -880
rect 40090 -960 40170 -950
rect 40430 -880 40510 -870
rect 40430 -950 40440 -880
rect 40440 -950 40500 -880
rect 40500 -950 40510 -880
rect 40430 -960 40510 -950
rect 40770 -880 40850 -870
rect 40770 -950 40780 -880
rect 40780 -950 40840 -880
rect 40840 -950 40850 -880
rect 40770 -960 40850 -950
rect 41110 -880 41190 -870
rect 41110 -950 41120 -880
rect 41120 -950 41180 -880
rect 41180 -950 41190 -880
rect 41110 -960 41190 -950
rect 41450 -880 41530 -870
rect 41450 -950 41460 -880
rect 41460 -950 41520 -880
rect 41520 -950 41530 -880
rect 41450 -960 41530 -950
rect 41790 -880 41870 -870
rect 41790 -950 41800 -880
rect 41800 -950 41860 -880
rect 41860 -950 41870 -880
rect 41790 -960 41870 -950
rect 42130 -880 42210 -870
rect 42130 -950 42140 -880
rect 42140 -950 42200 -880
rect 42200 -950 42210 -880
rect 42130 -960 42210 -950
rect 42470 -880 42550 -870
rect 42470 -950 42480 -880
rect 42480 -950 42540 -880
rect 42540 -950 42550 -880
rect 42470 -960 42550 -950
rect 42810 -880 42890 -870
rect 42810 -950 42820 -880
rect 42820 -950 42880 -880
rect 42880 -950 42890 -880
rect 42810 -960 42890 -950
rect 43150 -880 43230 -870
rect 43150 -950 43160 -880
rect 43160 -950 43220 -880
rect 43220 -950 43230 -880
rect 43150 -960 43230 -950
rect 43490 -880 43570 -870
rect 43490 -950 43500 -880
rect 43500 -950 43560 -880
rect 43560 -950 43570 -880
rect 43490 -960 43570 -950
rect 43830 -880 43910 -870
rect 43830 -950 43840 -880
rect 43840 -950 43900 -880
rect 43900 -950 43910 -880
rect 43830 -960 43910 -950
rect 44170 -880 44250 -870
rect 44170 -950 44180 -880
rect 44180 -950 44240 -880
rect 44240 -950 44250 -880
rect 44170 -960 44250 -950
rect 44510 -880 44590 -870
rect 44510 -950 44520 -880
rect 44520 -950 44580 -880
rect 44580 -950 44590 -880
rect 44510 -960 44590 -950
rect 44850 -880 44930 -870
rect 44850 -950 44860 -880
rect 44860 -950 44920 -880
rect 44920 -950 44930 -880
rect 44850 -960 44930 -950
rect 45190 -880 45270 -870
rect 45190 -950 45200 -880
rect 45200 -950 45260 -880
rect 45260 -950 45270 -880
rect 45190 -960 45270 -950
rect 45530 -880 45610 -870
rect 45530 -950 45540 -880
rect 45540 -950 45600 -880
rect 45600 -950 45610 -880
rect 45530 -960 45610 -950
rect 45870 -880 45950 -870
rect 45870 -950 45880 -880
rect 45880 -950 45940 -880
rect 45940 -950 45950 -880
rect 45870 -960 45950 -950
rect 46210 -880 46290 -870
rect 46210 -950 46220 -880
rect 46220 -950 46280 -880
rect 46280 -950 46290 -880
rect 46210 -960 46290 -950
rect 46550 -880 46630 -870
rect 46550 -950 46560 -880
rect 46560 -950 46620 -880
rect 46620 -950 46630 -880
rect 46550 -960 46630 -950
rect 46890 -880 46970 -870
rect 46890 -950 46900 -880
rect 46900 -950 46960 -880
rect 46960 -950 46970 -880
rect 46890 -960 46970 -950
rect 47230 -880 47310 -870
rect 47230 -950 47240 -880
rect 47240 -950 47300 -880
rect 47300 -950 47310 -880
rect 47230 -960 47310 -950
rect 47570 -880 47650 -870
rect 47570 -950 47580 -880
rect 47580 -950 47640 -880
rect 47640 -950 47650 -880
rect 47570 -960 47650 -950
rect 47910 -880 47990 -870
rect 47910 -950 47920 -880
rect 47920 -950 47980 -880
rect 47980 -950 47990 -880
rect 47910 -960 47990 -950
rect 48250 -880 48330 -870
rect 48250 -950 48260 -880
rect 48260 -950 48320 -880
rect 48320 -950 48330 -880
rect 48250 -960 48330 -950
rect 48590 -880 48670 -870
rect 48590 -950 48600 -880
rect 48600 -950 48660 -880
rect 48660 -950 48670 -880
rect 48590 -960 48670 -950
rect 48930 -880 49010 -870
rect 48930 -950 48940 -880
rect 48940 -950 49000 -880
rect 49000 -950 49010 -880
rect 48930 -960 49010 -950
rect 49270 -880 49350 -870
rect 49270 -950 49280 -880
rect 49280 -950 49340 -880
rect 49340 -950 49350 -880
rect 49270 -960 49350 -950
rect 49610 -880 49690 -870
rect 49610 -950 49620 -880
rect 49620 -950 49680 -880
rect 49680 -950 49690 -880
rect 49610 -960 49690 -950
rect 49950 -880 50030 -870
rect 49950 -950 49960 -880
rect 49960 -950 50020 -880
rect 50020 -950 50030 -880
rect 49950 -960 50030 -950
rect 50290 -880 50370 -870
rect 50290 -950 50300 -880
rect 50300 -950 50360 -880
rect 50360 -950 50370 -880
rect 50290 -960 50370 -950
rect 50630 -880 50710 -870
rect 50630 -950 50640 -880
rect 50640 -950 50700 -880
rect 50700 -950 50710 -880
rect 50630 -960 50710 -950
rect 50970 -880 51050 -870
rect 50970 -950 50980 -880
rect 50980 -950 51040 -880
rect 51040 -950 51050 -880
rect 50970 -960 51050 -950
rect 51310 -880 51390 -870
rect 51310 -950 51320 -880
rect 51320 -950 51380 -880
rect 51380 -950 51390 -880
rect 51310 -960 51390 -950
rect 51650 -880 51730 -870
rect 51650 -950 51660 -880
rect 51660 -950 51720 -880
rect 51720 -950 51730 -880
rect 51650 -960 51730 -950
rect 51990 -880 52070 -870
rect 51990 -950 52000 -880
rect 52000 -950 52060 -880
rect 52060 -950 52070 -880
rect 51990 -960 52070 -950
rect 52330 -880 52410 -870
rect 52330 -950 52340 -880
rect 52340 -950 52400 -880
rect 52400 -950 52410 -880
rect 52330 -960 52410 -950
rect 52670 -880 52750 -870
rect 52670 -950 52680 -880
rect 52680 -950 52740 -880
rect 52740 -950 52750 -880
rect 52670 -960 52750 -950
rect 53010 -880 53090 -870
rect 53010 -950 53020 -880
rect 53020 -950 53080 -880
rect 53080 -950 53090 -880
rect 53010 -960 53090 -950
rect 53350 -880 53430 -870
rect 53350 -950 53360 -880
rect 53360 -950 53420 -880
rect 53420 -950 53430 -880
rect 53350 -960 53430 -950
rect 53690 -880 53770 -870
rect 53690 -950 53700 -880
rect 53700 -950 53760 -880
rect 53760 -950 53770 -880
rect 53690 -960 53770 -950
rect 54030 -880 54110 -870
rect 54030 -950 54040 -880
rect 54040 -950 54100 -880
rect 54100 -950 54110 -880
rect 54030 -960 54110 -950
rect 54370 -880 54450 -870
rect 54370 -950 54380 -880
rect 54380 -950 54440 -880
rect 54440 -950 54450 -880
rect 54370 -960 54450 -950
rect 54710 -880 54790 -870
rect 54710 -950 54720 -880
rect 54720 -950 54780 -880
rect 54780 -950 54790 -880
rect 54710 -960 54790 -950
rect 55050 -880 55130 -870
rect 55050 -950 55060 -880
rect 55060 -950 55120 -880
rect 55120 -950 55130 -880
rect 55050 -960 55130 -950
rect 55390 -880 55470 -870
rect 55390 -950 55400 -880
rect 55400 -950 55460 -880
rect 55460 -950 55470 -880
rect 55390 -960 55470 -950
rect 55730 -880 55810 -870
rect 55730 -950 55740 -880
rect 55740 -950 55800 -880
rect 55800 -950 55810 -880
rect 55730 -960 55810 -950
rect 56070 -880 56150 -870
rect 56070 -950 56080 -880
rect 56080 -950 56140 -880
rect 56140 -950 56150 -880
rect 56070 -960 56150 -950
rect 56410 -880 56490 -870
rect 56410 -950 56420 -880
rect 56420 -950 56480 -880
rect 56480 -950 56490 -880
rect 56410 -960 56490 -950
rect 56750 -880 56830 -870
rect 56750 -950 56760 -880
rect 56760 -950 56820 -880
rect 56820 -950 56830 -880
rect 56750 -960 56830 -950
rect 57090 -880 57170 -870
rect 57090 -950 57100 -880
rect 57100 -950 57160 -880
rect 57160 -950 57170 -880
rect 57090 -960 57170 -950
rect 57430 -880 57510 -870
rect 57430 -950 57440 -880
rect 57440 -950 57500 -880
rect 57500 -950 57510 -880
rect 57430 -960 57510 -950
rect 57770 -880 57850 -870
rect 57770 -950 57780 -880
rect 57780 -950 57840 -880
rect 57840 -950 57850 -880
rect 57770 -960 57850 -950
rect 58110 -880 58190 -870
rect 58110 -950 58120 -880
rect 58120 -950 58180 -880
rect 58180 -950 58190 -880
rect 58110 -960 58190 -950
rect 58450 -880 58530 -870
rect 58450 -950 58460 -880
rect 58460 -950 58520 -880
rect 58520 -950 58530 -880
rect 58450 -960 58530 -950
rect 58790 -880 58870 -870
rect 58790 -950 58800 -880
rect 58800 -950 58860 -880
rect 58860 -950 58870 -880
rect 58790 -960 58870 -950
rect 59130 -880 59210 -870
rect 59130 -950 59140 -880
rect 59140 -950 59200 -880
rect 59200 -950 59210 -880
rect 59130 -960 59210 -950
rect 59470 -880 59550 -870
rect 59470 -950 59480 -880
rect 59480 -950 59540 -880
rect 59540 -950 59550 -880
rect 59470 -960 59550 -950
rect 59810 -880 59890 -870
rect 59810 -950 59820 -880
rect 59820 -950 59880 -880
rect 59880 -950 59890 -880
rect 59810 -960 59890 -950
rect 60150 -880 60230 -870
rect 60150 -950 60160 -880
rect 60160 -950 60220 -880
rect 60220 -950 60230 -880
rect 60150 -960 60230 -950
rect 60490 -880 60570 -870
rect 60490 -950 60500 -880
rect 60500 -950 60560 -880
rect 60560 -950 60570 -880
rect 60490 -960 60570 -950
rect 60830 -880 60910 -870
rect 60830 -950 60840 -880
rect 60840 -950 60900 -880
rect 60900 -950 60910 -880
rect 60830 -960 60910 -950
rect 61170 -880 61250 -870
rect 61170 -950 61180 -880
rect 61180 -950 61240 -880
rect 61240 -950 61250 -880
rect 61170 -960 61250 -950
rect 61510 -880 61590 -870
rect 61510 -950 61520 -880
rect 61520 -950 61580 -880
rect 61580 -950 61590 -880
rect 61510 -960 61590 -950
rect 61850 -880 61930 -870
rect 61850 -950 61860 -880
rect 61860 -950 61920 -880
rect 61920 -950 61930 -880
rect 61850 -960 61930 -950
rect 62190 -880 62270 -870
rect 62190 -950 62200 -880
rect 62200 -950 62260 -880
rect 62260 -950 62270 -880
rect 62190 -960 62270 -950
rect 62530 -880 62610 -870
rect 62530 -950 62540 -880
rect 62540 -950 62600 -880
rect 62600 -950 62610 -880
rect 62530 -960 62610 -950
rect 62870 -880 62950 -870
rect 62870 -950 62880 -880
rect 62880 -950 62940 -880
rect 62940 -950 62950 -880
rect 62870 -960 62950 -950
rect 63210 -880 63290 -870
rect 63210 -950 63220 -880
rect 63220 -950 63280 -880
rect 63280 -950 63290 -880
rect 63210 -960 63290 -950
rect 63550 -880 63630 -870
rect 63550 -950 63560 -880
rect 63560 -950 63620 -880
rect 63620 -950 63630 -880
rect 63550 -960 63630 -950
rect 63890 -880 63970 -870
rect 63890 -950 63900 -880
rect 63900 -950 63960 -880
rect 63960 -950 63970 -880
rect 63890 -960 63970 -950
rect 64230 -880 64310 -870
rect 64230 -950 64240 -880
rect 64240 -950 64300 -880
rect 64300 -950 64310 -880
rect 64230 -960 64310 -950
rect 64570 -880 64650 -870
rect 64570 -950 64580 -880
rect 64580 -950 64640 -880
rect 64640 -950 64650 -880
rect 64570 -960 64650 -950
rect 64910 -880 64990 -870
rect 64910 -950 64920 -880
rect 64920 -950 64980 -880
rect 64980 -950 64990 -880
rect 64910 -960 64990 -950
rect 65250 -880 65330 -870
rect 65250 -950 65260 -880
rect 65260 -950 65320 -880
rect 65320 -950 65330 -880
rect 65250 -960 65330 -950
rect 65590 -880 65670 -870
rect 65590 -950 65600 -880
rect 65600 -950 65660 -880
rect 65660 -950 65670 -880
rect 65590 -960 65670 -950
rect 65930 -880 66010 -870
rect 65930 -950 65940 -880
rect 65940 -950 66000 -880
rect 66000 -950 66010 -880
rect 65930 -960 66010 -950
rect 66270 -880 66350 -870
rect 66270 -950 66280 -880
rect 66280 -950 66340 -880
rect 66340 -950 66350 -880
rect 66270 -960 66350 -950
rect 66610 -880 66690 -870
rect 66610 -950 66620 -880
rect 66620 -950 66680 -880
rect 66680 -950 66690 -880
rect 66610 -960 66690 -950
rect 66950 -880 67030 -870
rect 66950 -950 66960 -880
rect 66960 -950 67020 -880
rect 67020 -950 67030 -880
rect 66950 -960 67030 -950
rect 67290 -880 67370 -870
rect 67290 -950 67300 -880
rect 67300 -950 67360 -880
rect 67360 -950 67370 -880
rect 67290 -960 67370 -950
rect 67630 -880 67710 -870
rect 67630 -950 67640 -880
rect 67640 -950 67700 -880
rect 67700 -950 67710 -880
rect 67630 -960 67710 -950
rect 67970 -880 68050 -870
rect 67970 -950 67980 -880
rect 67980 -950 68040 -880
rect 68040 -950 68050 -880
rect 67970 -960 68050 -950
rect 68310 -880 68390 -870
rect 68310 -950 68320 -880
rect 68320 -950 68380 -880
rect 68380 -950 68390 -880
rect 68310 -960 68390 -950
rect 68650 -880 68730 -870
rect 68650 -950 68660 -880
rect 68660 -950 68720 -880
rect 68720 -950 68730 -880
rect 68650 -960 68730 -950
rect 68990 -880 69070 -870
rect 68990 -950 69000 -880
rect 69000 -950 69060 -880
rect 69060 -950 69070 -880
rect 68990 -960 69070 -950
rect 69330 -880 69410 -870
rect 69330 -950 69340 -880
rect 69340 -950 69400 -880
rect 69400 -950 69410 -880
rect 69330 -960 69410 -950
rect 69670 -880 69750 -870
rect 69670 -950 69680 -880
rect 69680 -950 69740 -880
rect 69740 -950 69750 -880
rect 69670 -960 69750 -950
rect 70010 -880 70090 -870
rect 70010 -950 70020 -880
rect 70020 -950 70080 -880
rect 70080 -950 70090 -880
rect 70010 -960 70090 -950
rect 70350 -880 70430 -870
rect 70350 -950 70360 -880
rect 70360 -950 70420 -880
rect 70420 -950 70430 -880
rect 70350 -960 70430 -950
rect 70690 -880 70770 -870
rect 70690 -950 70700 -880
rect 70700 -950 70760 -880
rect 70760 -950 70770 -880
rect 70690 -960 70770 -950
rect 71030 -880 71110 -870
rect 71030 -950 71040 -880
rect 71040 -950 71100 -880
rect 71100 -950 71110 -880
rect 71030 -960 71110 -950
rect 71370 -880 71450 -870
rect 71370 -950 71380 -880
rect 71380 -950 71440 -880
rect 71440 -950 71450 -880
rect 71370 -960 71450 -950
rect 71710 -880 71790 -870
rect 71710 -950 71720 -880
rect 71720 -950 71780 -880
rect 71780 -950 71790 -880
rect 71710 -960 71790 -950
rect 72050 -880 72130 -870
rect 72050 -950 72060 -880
rect 72060 -950 72120 -880
rect 72120 -950 72130 -880
rect 72050 -960 72130 -950
rect 72390 -880 72470 -870
rect 72390 -950 72400 -880
rect 72400 -950 72460 -880
rect 72460 -950 72470 -880
rect 72390 -960 72470 -950
rect 72730 -880 72810 -870
rect 72730 -950 72740 -880
rect 72740 -950 72800 -880
rect 72800 -950 72810 -880
rect 72730 -960 72810 -950
rect 73070 -880 73150 -870
rect 73070 -950 73080 -880
rect 73080 -950 73140 -880
rect 73140 -950 73150 -880
rect 73070 -960 73150 -950
rect 73410 -880 73490 -870
rect 73410 -950 73420 -880
rect 73420 -950 73480 -880
rect 73480 -950 73490 -880
rect 73410 -960 73490 -950
rect 73750 -880 73830 -870
rect 73750 -950 73760 -880
rect 73760 -950 73820 -880
rect 73820 -950 73830 -880
rect 73750 -960 73830 -950
rect 74090 -880 74170 -870
rect 74090 -950 74100 -880
rect 74100 -950 74160 -880
rect 74160 -950 74170 -880
rect 74090 -960 74170 -950
rect 74430 -880 74510 -870
rect 74430 -950 74440 -880
rect 74440 -950 74500 -880
rect 74500 -950 74510 -880
rect 74430 -960 74510 -950
rect 74770 -880 74850 -870
rect 74770 -950 74780 -880
rect 74780 -950 74840 -880
rect 74840 -950 74850 -880
rect 74770 -960 74850 -950
rect 75110 -880 75190 -870
rect 75110 -950 75120 -880
rect 75120 -950 75180 -880
rect 75180 -950 75190 -880
rect 75110 -960 75190 -950
rect 75450 -880 75530 -870
rect 75450 -950 75460 -880
rect 75460 -950 75520 -880
rect 75520 -950 75530 -880
rect 75450 -960 75530 -950
rect 75790 -880 75870 -870
rect 75790 -950 75800 -880
rect 75800 -950 75860 -880
rect 75860 -950 75870 -880
rect 75790 -960 75870 -950
rect 76130 -880 76210 -870
rect 76130 -950 76140 -880
rect 76140 -950 76200 -880
rect 76200 -950 76210 -880
rect 76130 -960 76210 -950
rect 76470 -880 76550 -870
rect 76470 -950 76480 -880
rect 76480 -950 76540 -880
rect 76540 -950 76550 -880
rect 76470 -960 76550 -950
rect 76810 -880 76890 -870
rect 76810 -950 76820 -880
rect 76820 -950 76880 -880
rect 76880 -950 76890 -880
rect 76810 -960 76890 -950
rect 77150 -880 77230 -870
rect 77150 -950 77160 -880
rect 77160 -950 77220 -880
rect 77220 -950 77230 -880
rect 77150 -960 77230 -950
rect 77490 -880 77570 -870
rect 77490 -950 77500 -880
rect 77500 -950 77560 -880
rect 77560 -950 77570 -880
rect 77490 -960 77570 -950
rect 77830 -880 77910 -870
rect 77830 -950 77840 -880
rect 77840 -950 77900 -880
rect 77900 -950 77910 -880
rect 77830 -960 77910 -950
rect 78170 -880 78250 -870
rect 78170 -950 78180 -880
rect 78180 -950 78240 -880
rect 78240 -950 78250 -880
rect 78170 -960 78250 -950
rect 78510 -880 78590 -870
rect 78510 -950 78520 -880
rect 78520 -950 78580 -880
rect 78580 -950 78590 -880
rect 78510 -960 78590 -950
rect 78850 -880 78930 -870
rect 78850 -950 78860 -880
rect 78860 -950 78920 -880
rect 78920 -950 78930 -880
rect 78850 -960 78930 -950
rect 79190 -880 79270 -870
rect 79190 -950 79200 -880
rect 79200 -950 79260 -880
rect 79260 -950 79270 -880
rect 79190 -960 79270 -950
rect 79530 -880 79610 -870
rect 79530 -950 79540 -880
rect 79540 -950 79600 -880
rect 79600 -950 79610 -880
rect 79530 -960 79610 -950
rect 79870 -880 79950 -870
rect 79870 -950 79880 -880
rect 79880 -950 79940 -880
rect 79940 -950 79950 -880
rect 79870 -960 79950 -950
rect 80210 -880 80290 -870
rect 80210 -950 80220 -880
rect 80220 -950 80280 -880
rect 80280 -950 80290 -880
rect 80210 -960 80290 -950
rect 80550 -880 80630 -870
rect 80550 -950 80560 -880
rect 80560 -950 80620 -880
rect 80620 -950 80630 -880
rect 80550 -960 80630 -950
rect 80890 -880 80970 -870
rect 80890 -950 80900 -880
rect 80900 -950 80960 -880
rect 80960 -950 80970 -880
rect 80890 -960 80970 -950
rect 81230 -880 81310 -870
rect 81230 -950 81240 -880
rect 81240 -950 81300 -880
rect 81300 -950 81310 -880
rect 81230 -960 81310 -950
rect 81570 -880 81650 -870
rect 81570 -950 81580 -880
rect 81580 -950 81640 -880
rect 81640 -950 81650 -880
rect 81570 -960 81650 -950
rect 81910 -880 81990 -870
rect 81910 -950 81920 -880
rect 81920 -950 81980 -880
rect 81980 -950 81990 -880
rect 81910 -960 81990 -950
rect 82250 -880 82330 -870
rect 82250 -950 82260 -880
rect 82260 -950 82320 -880
rect 82320 -950 82330 -880
rect 82250 -960 82330 -950
rect 82590 -880 82670 -870
rect 82590 -950 82600 -880
rect 82600 -950 82660 -880
rect 82660 -950 82670 -880
rect 82590 -960 82670 -950
rect 82930 -880 83010 -870
rect 82930 -950 82940 -880
rect 82940 -950 83000 -880
rect 83000 -950 83010 -880
rect 82930 -960 83010 -950
rect 83270 -880 83350 -870
rect 83270 -950 83280 -880
rect 83280 -950 83340 -880
rect 83340 -950 83350 -880
rect 83270 -960 83350 -950
rect 83610 -880 83690 -870
rect 83610 -950 83620 -880
rect 83620 -950 83680 -880
rect 83680 -950 83690 -880
rect 83610 -960 83690 -950
rect 83950 -880 84030 -870
rect 83950 -950 83960 -880
rect 83960 -950 84020 -880
rect 84020 -950 84030 -880
rect 83950 -960 84030 -950
rect 84290 -880 84370 -870
rect 84290 -950 84300 -880
rect 84300 -950 84360 -880
rect 84360 -950 84370 -880
rect 84290 -960 84370 -950
rect 84630 -880 84710 -870
rect 84630 -950 84640 -880
rect 84640 -950 84700 -880
rect 84700 -950 84710 -880
rect 84630 -960 84710 -950
rect 84970 -880 85050 -870
rect 84970 -950 84980 -880
rect 84980 -950 85040 -880
rect 85040 -950 85050 -880
rect 84970 -960 85050 -950
rect 85310 -880 85390 -870
rect 85310 -950 85320 -880
rect 85320 -950 85380 -880
rect 85380 -950 85390 -880
rect 85310 -960 85390 -950
rect 85650 -880 85730 -870
rect 85650 -950 85660 -880
rect 85660 -950 85720 -880
rect 85720 -950 85730 -880
rect 85650 -960 85730 -950
rect 85990 -880 86070 -870
rect 85990 -950 86000 -880
rect 86000 -950 86060 -880
rect 86060 -950 86070 -880
rect 85990 -960 86070 -950
rect 86330 -880 86410 -870
rect 86330 -950 86340 -880
rect 86340 -950 86400 -880
rect 86400 -950 86410 -880
rect 86330 -960 86410 -950
rect 86670 -880 86750 -870
rect 86670 -950 86680 -880
rect 86680 -950 86740 -880
rect 86740 -950 86750 -880
rect 86670 -960 86750 -950
rect 87010 -880 87090 -870
rect 87010 -950 87020 -880
rect 87020 -950 87080 -880
rect 87080 -950 87090 -880
rect 87010 -960 87090 -950
rect 120 -1520 240 -1430
rect 830 -1540 910 -1470
rect 1480 -1520 1600 -1430
rect 2840 -1520 2960 -1430
rect 4200 -1520 4320 -1430
rect 5000 -1540 5080 -1470
rect 5560 -1520 5680 -1430
rect 6920 -1520 7040 -1430
rect 8280 -1520 8400 -1430
rect 9030 -1540 9110 -1470
rect 9640 -1520 9760 -1430
rect 11000 -1520 11120 -1430
rect 12360 -1520 12480 -1430
rect 13060 -1540 13140 -1470
rect 13720 -1520 13840 -1430
rect 15080 -1520 15200 -1430
rect 16440 -1520 16560 -1430
rect 17100 -1540 17180 -1470
rect 17800 -1520 17920 -1430
rect 19160 -1520 19280 -1430
rect 20520 -1520 20640 -1430
rect 21200 -1540 21280 -1470
rect 21880 -1520 22000 -1430
rect 23240 -1520 23360 -1430
rect 24600 -1520 24720 -1430
rect 25310 -1540 25390 -1470
rect 25960 -1520 26080 -1430
rect 27320 -1520 27440 -1430
rect 28680 -1520 28800 -1430
rect 29410 -1540 29490 -1470
rect 30040 -1520 30160 -1430
rect 31400 -1520 31520 -1430
rect 32760 -1520 32880 -1430
rect 33440 -1540 33520 -1470
rect 34120 -1520 34240 -1430
rect 35480 -1520 35600 -1430
rect 36840 -1520 36960 -1430
rect 37550 -1540 37630 -1470
rect 38200 -1520 38320 -1430
rect 39560 -1520 39680 -1430
rect 40920 -1520 41040 -1430
rect 41650 -1540 41730 -1470
rect 42280 -1520 42400 -1430
rect 43640 -1520 43760 -1430
rect 45000 -1520 45120 -1430
rect 46360 -1520 46480 -1430
rect 47100 -1540 47180 -1470
rect 47720 -1520 47840 -1430
rect 49080 -1520 49200 -1430
rect 50440 -1520 50560 -1430
rect 51180 -1540 51260 -1470
rect 51800 -1520 51920 -1430
rect 53160 -1520 53280 -1430
rect 54520 -1520 54640 -1430
rect 55290 -1540 55370 -1470
rect 55880 -1520 56000 -1430
rect 57240 -1520 57360 -1430
rect 58600 -1520 58720 -1430
rect 59320 -1540 59400 -1470
rect 59960 -1520 60080 -1430
rect 61320 -1520 61440 -1430
rect 62680 -1520 62800 -1430
rect 63420 -1540 63500 -1470
rect 64040 -1520 64160 -1430
rect 65400 -1520 65520 -1430
rect 66760 -1520 66880 -1430
rect 67530 -1540 67610 -1470
rect 68120 -1520 68240 -1430
rect 69480 -1520 69600 -1430
rect 70840 -1520 70960 -1430
rect 71560 -1540 71640 -1470
rect 72200 -1520 72320 -1430
rect 73560 -1520 73680 -1430
rect 74920 -1520 75040 -1430
rect 75810 -1540 75890 -1470
rect 76280 -1520 76400 -1430
rect 77640 -1520 77760 -1430
rect 79000 -1520 79120 -1430
rect 79770 -1540 79850 -1470
rect 80360 -1520 80480 -1430
rect 81720 -1520 81840 -1430
rect 83080 -1520 83200 -1430
rect 83950 -1540 84030 -1470
rect 84440 -1520 84560 -1430
rect 85800 -1520 85920 -1430
rect 86508 -1544 86588 -1474
<< metal4 >>
rect -520 670 -160 740
rect -520 660 -460 670
rect -564 410 -460 660
rect -520 400 -460 410
rect -200 660 -160 670
rect -200 620 360 660
rect -200 530 0 620
rect 120 580 360 620
rect 730 590 930 620
rect 730 580 790 590
rect 120 570 790 580
rect 120 530 420 570
rect -200 480 420 530
rect 540 520 790 570
rect 870 580 930 590
rect 2110 590 2310 620
rect 2110 580 2170 590
rect 870 570 1200 580
rect 870 520 1090 570
rect 540 480 1090 520
rect 1190 480 1200 570
rect -200 470 1200 480
rect 1470 570 2170 580
rect 1470 480 1490 570
rect 1610 520 2170 570
rect 2250 580 2310 590
rect 3490 590 3690 620
rect 3490 580 3550 590
rect 2250 570 3550 580
rect 2250 520 2850 570
rect 1610 480 2850 520
rect 2970 520 3550 570
rect 3630 580 3690 590
rect 5150 590 5350 620
rect 5150 580 5210 590
rect 3630 570 5210 580
rect 3630 520 4210 570
rect 2970 480 4210 520
rect 4330 480 4510 570
rect 4630 520 5210 570
rect 5290 580 5350 590
rect 7980 590 8180 620
rect 7980 580 8040 590
rect 5290 570 8040 580
rect 5290 520 5870 570
rect 4630 480 5870 520
rect 5990 480 7230 570
rect 7350 520 8040 570
rect 8120 580 8180 590
rect 10740 590 10940 620
rect 10740 580 10800 590
rect 8120 570 10800 580
rect 8120 520 8590 570
rect 7350 480 8590 520
rect 8710 480 9950 570
rect 10070 520 10800 570
rect 10880 580 10940 590
rect 13370 590 13570 620
rect 13370 580 13430 590
rect 10880 570 13430 580
rect 10880 520 11310 570
rect 10070 480 11310 520
rect 11430 480 12670 570
rect 12790 520 13430 570
rect 13510 580 13570 590
rect 16410 590 16610 620
rect 16410 580 16470 590
rect 13510 570 16470 580
rect 13510 520 14030 570
rect 12790 480 14030 520
rect 14150 480 15390 570
rect 15510 480 15690 570
rect 15810 520 16470 570
rect 16550 580 16610 590
rect 20480 590 20680 620
rect 20480 580 20540 590
rect 16550 570 20540 580
rect 16550 520 17050 570
rect 15810 480 17050 520
rect 17170 480 18410 570
rect 18530 480 19770 570
rect 19890 520 20540 570
rect 20620 580 20680 590
rect 24620 590 24820 620
rect 24620 580 24680 590
rect 20620 570 24680 580
rect 20620 520 21130 570
rect 19890 480 21130 520
rect 21250 480 22490 570
rect 22610 480 23850 570
rect 23970 520 24680 570
rect 24760 580 24820 590
rect 28700 590 28900 620
rect 28700 580 28760 590
rect 24760 570 28760 580
rect 24760 520 25210 570
rect 23970 480 25210 520
rect 25330 480 26570 570
rect 26690 480 27930 570
rect 28050 520 28760 570
rect 28840 580 28900 590
rect 32850 590 33050 620
rect 32850 580 32910 590
rect 28840 570 32910 580
rect 28840 520 29290 570
rect 28050 480 29290 520
rect 29410 480 30650 570
rect 30770 480 32010 570
rect 32130 520 32910 570
rect 32990 580 33050 590
rect 36720 590 36920 620
rect 36720 580 36780 590
rect 32990 570 36780 580
rect 32990 520 33370 570
rect 32130 480 33370 520
rect 33490 480 34730 570
rect 34850 480 36090 570
rect 36210 520 36780 570
rect 36860 580 36920 590
rect 40860 590 41060 620
rect 40860 580 40920 590
rect 36860 570 40920 580
rect 36860 520 37450 570
rect 36210 480 37450 520
rect 37570 480 38810 570
rect 38930 480 40170 570
rect 40290 520 40920 570
rect 41000 580 41060 590
rect 44850 590 45050 620
rect 44850 580 44910 590
rect 41000 570 44910 580
rect 41000 520 41530 570
rect 40290 480 41530 520
rect 41650 480 42890 570
rect 43010 480 44250 570
rect 44370 520 44910 570
rect 44990 580 45050 590
rect 48930 590 49130 620
rect 48930 580 48990 590
rect 44990 570 48990 580
rect 44990 520 45610 570
rect 44370 480 45610 520
rect 45730 480 46970 570
rect 47090 480 48330 570
rect 48450 520 48990 570
rect 49070 580 49130 590
rect 53020 590 53220 620
rect 53020 580 53080 590
rect 49070 570 53080 580
rect 49070 520 49690 570
rect 48450 480 49690 520
rect 49810 480 51050 570
rect 51170 480 52410 570
rect 52530 520 53080 570
rect 53160 580 53220 590
rect 57180 590 57380 620
rect 57180 580 57240 590
rect 53160 570 57240 580
rect 53160 520 53770 570
rect 52530 480 53770 520
rect 53890 480 55130 570
rect 55250 480 56490 570
rect 56610 520 57240 570
rect 57320 580 57380 590
rect 57320 570 59340 580
rect 57320 520 57850 570
rect 56610 480 57850 520
rect 57970 480 59210 570
rect 59330 480 59340 570
rect 1470 470 59340 480
rect -200 410 360 470
rect -200 400 -160 410
rect -520 280 -160 400
rect 590 210 1410 220
rect 590 120 610 210
rect 690 120 950 210
rect 1030 120 1290 210
rect 1400 120 1410 210
rect 590 110 1410 120
rect 1660 210 4490 220
rect 1660 120 1680 210
rect 1760 120 2020 210
rect 2100 120 2360 210
rect 2440 120 2700 210
rect 2780 120 3040 210
rect 3120 120 3380 210
rect 3460 120 3720 210
rect 3800 120 4060 210
rect 4140 120 4370 210
rect 4480 120 4490 210
rect 1660 110 4490 120
rect 4680 210 15670 220
rect 4680 120 4700 210
rect 4780 120 5040 210
rect 5120 120 5380 210
rect 5460 120 5720 210
rect 5800 120 6060 210
rect 6140 120 6400 210
rect 6480 120 6740 210
rect 6820 120 7080 210
rect 7160 120 7420 210
rect 7500 120 7760 210
rect 7840 120 8100 210
rect 8180 120 8440 210
rect 8520 120 8780 210
rect 8860 120 9120 210
rect 9200 120 9460 210
rect 9540 120 9800 210
rect 9880 120 10140 210
rect 10220 120 10480 210
rect 10560 120 10820 210
rect 10900 120 11160 210
rect 11240 120 11500 210
rect 11580 120 11840 210
rect 11920 120 12180 210
rect 12260 120 12520 210
rect 12600 120 12860 210
rect 12940 120 13200 210
rect 13280 120 13540 210
rect 13620 120 13880 210
rect 13960 120 14220 210
rect 14300 120 14560 210
rect 14640 120 14900 210
rect 14980 120 15240 210
rect 15320 120 15550 210
rect 15660 120 15670 210
rect 4680 110 15670 120
rect 15860 210 59200 220
rect 15860 120 15880 210
rect 15960 120 16220 210
rect 16300 120 16560 210
rect 16640 120 16900 210
rect 16980 120 17240 210
rect 17320 120 17580 210
rect 17660 120 17920 210
rect 18000 120 18260 210
rect 18340 120 18600 210
rect 18680 120 18940 210
rect 19020 120 19280 210
rect 19360 120 19620 210
rect 19700 120 19960 210
rect 20040 120 20300 210
rect 20380 120 20640 210
rect 20720 120 20980 210
rect 21060 120 21320 210
rect 21400 120 21660 210
rect 21740 120 22000 210
rect 22080 120 22340 210
rect 22420 120 22680 210
rect 22760 120 23020 210
rect 23100 120 23360 210
rect 23440 120 23700 210
rect 23780 120 24040 210
rect 24120 120 24380 210
rect 24460 120 24720 210
rect 24800 120 25060 210
rect 25140 120 25400 210
rect 25480 120 25740 210
rect 25820 120 26080 210
rect 26160 120 26420 210
rect 26500 120 26760 210
rect 26840 120 27100 210
rect 27180 120 27440 210
rect 27520 120 27780 210
rect 27860 120 28120 210
rect 28200 120 28460 210
rect 28540 120 28800 210
rect 28880 120 29140 210
rect 29220 120 29480 210
rect 29560 120 29820 210
rect 29900 120 30160 210
rect 30240 120 30500 210
rect 30580 120 30840 210
rect 30920 120 31180 210
rect 31260 120 31520 210
rect 31600 120 31860 210
rect 31940 120 32200 210
rect 32280 120 32540 210
rect 32620 120 32880 210
rect 32960 120 33220 210
rect 33300 120 33560 210
rect 33640 120 33900 210
rect 33980 120 34240 210
rect 34320 120 34580 210
rect 34660 120 34920 210
rect 35000 120 35260 210
rect 35340 120 35600 210
rect 35680 120 35940 210
rect 36020 120 36280 210
rect 36360 120 36620 210
rect 36700 120 36960 210
rect 37040 120 37300 210
rect 37380 120 37640 210
rect 37720 120 37980 210
rect 38060 120 38320 210
rect 38400 120 38660 210
rect 38740 120 39000 210
rect 39080 120 39340 210
rect 39420 120 39680 210
rect 39760 120 40020 210
rect 40100 120 40360 210
rect 40440 120 40700 210
rect 40780 120 41040 210
rect 41120 120 41380 210
rect 41460 120 41720 210
rect 41800 120 42060 210
rect 42140 120 42400 210
rect 42480 120 42740 210
rect 42820 120 43080 210
rect 43160 120 43420 210
rect 43500 120 43760 210
rect 43840 120 44100 210
rect 44180 120 44440 210
rect 44520 120 44780 210
rect 44860 120 45120 210
rect 45200 120 45460 210
rect 45540 120 45800 210
rect 45880 120 46140 210
rect 46220 120 46480 210
rect 46560 120 46820 210
rect 46900 120 47160 210
rect 47240 120 47500 210
rect 47580 120 47840 210
rect 47920 120 48180 210
rect 48260 120 48520 210
rect 48600 120 48860 210
rect 48940 120 49200 210
rect 49280 120 49540 210
rect 49620 120 49880 210
rect 49960 120 50220 210
rect 50300 120 50560 210
rect 50640 120 50900 210
rect 50980 120 51240 210
rect 51320 120 51580 210
rect 51660 120 51920 210
rect 52000 120 52260 210
rect 52340 120 52600 210
rect 52680 120 52940 210
rect 53020 120 53280 210
rect 53360 120 53620 210
rect 53700 120 53960 210
rect 54040 120 54300 210
rect 54380 120 54640 210
rect 54720 120 54980 210
rect 55060 120 55320 210
rect 55400 120 55660 210
rect 55740 120 56000 210
rect 56080 120 56340 210
rect 56420 120 56680 210
rect 56760 120 57020 210
rect 57100 120 57360 210
rect 57440 120 57700 210
rect 57780 120 58040 210
rect 58120 120 58380 210
rect 58460 120 58720 210
rect 58800 120 59060 210
rect 59140 120 59200 210
rect 15860 110 59200 120
rect -564 -220 350 -200
rect 79750 -220 80270 -210
rect -564 -260 87320 -220
rect -564 -270 2120 -260
rect -564 -370 0 -270
rect 100 -370 130 -270
rect 230 -280 1490 -270
rect 230 -370 430 -280
rect -564 -380 430 -370
rect 530 -380 1110 -280
rect 1210 -370 1490 -280
rect 1590 -370 2120 -270
rect 1210 -380 2120 -370
rect -564 -390 2120 -380
rect 2350 -264 87320 -260
rect 2350 -268 13668 -264
rect 2350 -270 5138 -268
rect 2350 -280 4860 -270
rect 2350 -380 2860 -280
rect 2960 -380 4550 -280
rect 4650 -370 4860 -280
rect 4960 -370 5138 -270
rect 4650 -380 5138 -370
rect 2350 -390 5138 -380
rect -564 -398 5138 -390
rect 5368 -270 7624 -268
rect 5368 -370 5910 -270
rect 6010 -370 6220 -270
rect 6320 -370 6930 -270
rect 7030 -280 7624 -270
rect 7030 -370 7240 -280
rect 5368 -380 7240 -370
rect 7340 -380 7624 -280
rect 5368 -398 7624 -380
rect 7854 -270 9044 -268
rect 7854 -280 8600 -270
rect 7854 -380 8290 -280
rect 8390 -370 8600 -280
rect 8700 -370 9044 -270
rect 8390 -380 9044 -370
rect 7854 -398 9044 -380
rect 9274 -270 13668 -268
rect 9274 -370 9650 -270
rect 9750 -370 9960 -270
rect 10060 -370 10670 -270
rect 10770 -280 11690 -270
rect 10770 -370 10980 -280
rect 9274 -380 10980 -370
rect 11080 -370 11690 -280
rect 11790 -280 13050 -270
rect 11790 -370 11990 -280
rect 11080 -380 11990 -370
rect 12090 -380 12670 -280
rect 12770 -370 13050 -280
rect 13150 -370 13668 -270
rect 12770 -380 13668 -370
rect 9274 -394 13668 -380
rect 13898 -270 16868 -264
rect 13898 -280 16380 -270
rect 13898 -380 14420 -280
rect 14520 -380 16110 -280
rect 16210 -370 16380 -280
rect 16480 -370 16868 -270
rect 16210 -380 16868 -370
rect 13898 -394 16868 -380
rect 17098 -270 20424 -264
rect 17098 -370 17470 -270
rect 17570 -370 17740 -270
rect 17840 -370 18490 -270
rect 18590 -280 20120 -270
rect 18590 -370 18760 -280
rect 17098 -380 18760 -370
rect 18860 -380 19850 -280
rect 19950 -370 20120 -280
rect 20220 -370 20424 -270
rect 19950 -380 20424 -370
rect 17098 -394 20424 -380
rect 20654 -270 25758 -264
rect 20654 -370 21210 -270
rect 21310 -370 21480 -270
rect 21580 -370 22230 -270
rect 22330 -280 23590 -270
rect 22330 -370 22500 -280
rect 20654 -380 22500 -370
rect 22600 -370 23590 -280
rect 23690 -280 24950 -270
rect 23690 -370 23860 -280
rect 22600 -380 23860 -370
rect 23960 -380 24530 -280
rect 24630 -370 24950 -280
rect 25050 -370 25758 -270
rect 24630 -380 25758 -370
rect 20654 -394 25758 -380
rect 25988 -270 28602 -264
rect 25988 -280 28280 -270
rect 25988 -380 26320 -280
rect 26420 -380 28010 -280
rect 28110 -370 28280 -280
rect 28380 -370 28602 -270
rect 28110 -380 28602 -370
rect 25988 -394 28602 -380
rect 28832 -270 32514 -264
rect 28832 -370 29370 -270
rect 29470 -370 29640 -270
rect 29740 -370 30390 -270
rect 30490 -280 32020 -270
rect 30490 -370 30660 -280
rect 28832 -380 30660 -370
rect 30760 -380 31750 -280
rect 31850 -370 32020 -280
rect 32120 -370 32514 -270
rect 31850 -380 32514 -370
rect 28832 -394 32514 -380
rect 32744 -270 34670 -264
rect 32744 -370 33110 -270
rect 33210 -370 33380 -270
rect 33480 -370 34130 -270
rect 34230 -280 34670 -270
rect 34230 -370 34400 -280
rect 32744 -380 34400 -370
rect 34500 -380 34670 -280
rect 32744 -394 34670 -380
rect 34900 -270 37492 -264
rect 34900 -370 35490 -270
rect 35590 -280 36850 -270
rect 35590 -370 35760 -280
rect 34900 -380 35760 -370
rect 35860 -380 36430 -280
rect 36530 -370 36850 -280
rect 36950 -370 37492 -270
rect 36530 -380 37492 -370
rect 34900 -394 37492 -380
rect 37722 -280 40692 -264
rect 37722 -380 38220 -280
rect 38320 -380 39910 -280
rect 40010 -380 40692 -280
rect 37722 -394 40692 -380
rect 40922 -270 45668 -264
rect 40922 -370 41270 -270
rect 41370 -370 42290 -270
rect 42390 -280 43650 -270
rect 42390 -370 42560 -280
rect 40922 -380 42560 -370
rect 42660 -380 43650 -280
rect 43750 -280 45010 -270
rect 43750 -380 44600 -280
rect 44700 -370 45010 -280
rect 45110 -370 45668 -270
rect 44700 -380 45668 -370
rect 40922 -394 45668 -380
rect 45898 -270 48868 -264
rect 45898 -280 48340 -270
rect 45898 -380 46380 -280
rect 46480 -380 48070 -280
rect 48170 -370 48340 -280
rect 48440 -370 48868 -270
rect 48170 -380 48868 -370
rect 45898 -394 48868 -380
rect 49098 -270 51002 -264
rect 49098 -370 49430 -270
rect 49530 -370 49700 -270
rect 49800 -370 50450 -270
rect 50550 -280 51002 -270
rect 50550 -370 50720 -280
rect 49098 -380 50720 -370
rect 50820 -380 51002 -280
rect 49098 -394 51002 -380
rect 51232 -270 54558 -264
rect 51232 -280 52080 -270
rect 51232 -380 51810 -280
rect 51910 -370 52080 -280
rect 52180 -370 53170 -270
rect 53270 -370 53440 -270
rect 53540 -370 54190 -270
rect 54290 -370 54558 -270
rect 51910 -380 54558 -370
rect 51232 -394 54558 -380
rect 54788 -270 57402 -264
rect 54788 -370 55210 -270
rect 55310 -280 56570 -270
rect 55310 -370 55480 -280
rect 54788 -380 55480 -370
rect 55580 -370 56570 -280
rect 56670 -370 57402 -270
rect 55580 -380 57402 -370
rect 54788 -394 57402 -380
rect 57632 -270 61314 -264
rect 57632 -280 60990 -270
rect 57632 -380 57940 -280
rect 58040 -380 59630 -280
rect 59730 -370 60990 -280
rect 61090 -370 61314 -270
rect 59730 -380 61314 -370
rect 57632 -394 61314 -380
rect 61544 -270 64158 -264
rect 61544 -370 62010 -270
rect 62110 -280 64158 -270
rect 62110 -370 63370 -280
rect 61544 -380 63370 -370
rect 63470 -380 64158 -280
rect 61544 -394 64158 -380
rect 64388 -270 67714 -264
rect 64388 -370 64730 -270
rect 64830 -370 65750 -270
rect 65850 -370 67110 -270
rect 67210 -370 67714 -270
rect 64388 -394 67714 -370
rect 67944 -270 70558 -264
rect 67944 -370 68470 -270
rect 68570 -280 70558 -270
rect 68570 -370 69840 -280
rect 67944 -380 69840 -370
rect 69940 -380 70558 -280
rect 67944 -394 70558 -380
rect 70788 -270 74468 -264
rect 70788 -280 72890 -270
rect 70788 -380 71530 -280
rect 71630 -370 72890 -280
rect 72990 -370 73910 -270
rect 74010 -370 74468 -270
rect 71630 -380 74468 -370
rect 70788 -394 74468 -380
rect 74698 -270 78380 -264
rect 74698 -280 76630 -270
rect 74698 -380 75270 -280
rect 75370 -370 76630 -280
rect 76730 -370 77650 -270
rect 77750 -370 78380 -270
rect 75370 -380 78380 -370
rect 74698 -394 78380 -380
rect 78610 -270 82292 -264
rect 78610 -370 79010 -270
rect 79110 -370 80370 -270
rect 80470 -280 82292 -270
rect 80470 -370 81740 -280
rect 78610 -380 81740 -370
rect 81840 -380 82292 -280
rect 78610 -394 82292 -380
rect 82522 -270 86202 -264
rect 82522 -280 84790 -270
rect 82522 -380 83430 -280
rect 83530 -370 84790 -280
rect 84890 -370 85810 -270
rect 85910 -370 86202 -270
rect 83530 -380 86202 -370
rect 82522 -394 86202 -380
rect 86432 -280 87320 -264
rect 86432 -380 87170 -280
rect 87270 -380 87320 -280
rect 86432 -394 87320 -380
rect 9274 -398 87320 -394
rect -564 -430 87320 -398
rect -564 -450 350 -430
rect 79750 -440 80270 -430
rect -940 -820 360 -790
rect -940 -860 550 -820
rect -940 -870 87300 -860
rect -940 -960 310 -870
rect 390 -960 650 -870
rect 730 -960 990 -870
rect 1070 -960 1330 -870
rect 1410 -960 1670 -870
rect 1750 -960 2010 -870
rect 2090 -960 2350 -870
rect 2430 -960 2690 -870
rect 2770 -960 3030 -870
rect 3110 -960 3370 -870
rect 3450 -960 3710 -870
rect 3790 -960 4050 -870
rect 4130 -960 4390 -870
rect 4470 -960 4730 -870
rect 4810 -960 5070 -870
rect 5150 -960 5410 -870
rect 5490 -960 5750 -870
rect 5830 -960 6090 -870
rect 6170 -960 6430 -870
rect 6510 -960 6770 -870
rect 6850 -960 7110 -870
rect 7190 -960 7450 -870
rect 7530 -960 7790 -870
rect 7870 -960 8130 -870
rect 8210 -960 8470 -870
rect 8550 -960 8810 -870
rect 8890 -960 9150 -870
rect 9230 -960 9490 -870
rect 9570 -960 9830 -870
rect 9910 -960 10170 -870
rect 10250 -960 10510 -870
rect 10590 -960 10850 -870
rect 10930 -960 11190 -870
rect 11270 -960 11530 -870
rect 11610 -960 11870 -870
rect 11950 -960 12210 -870
rect 12290 -960 12550 -870
rect 12630 -960 12890 -870
rect 12970 -960 13230 -870
rect 13310 -960 13570 -870
rect 13650 -960 13910 -870
rect 13990 -960 14250 -870
rect 14330 -960 14590 -870
rect 14670 -960 14930 -870
rect 15010 -960 15270 -870
rect 15350 -960 15610 -870
rect 15690 -960 15950 -870
rect 16030 -960 16290 -870
rect 16370 -960 16630 -870
rect 16710 -960 16970 -870
rect 17050 -960 17310 -870
rect 17390 -960 17650 -870
rect 17730 -960 17990 -870
rect 18070 -960 18330 -870
rect 18410 -960 18670 -870
rect 18750 -960 19010 -870
rect 19090 -960 19350 -870
rect 19430 -960 19690 -870
rect 19770 -960 20030 -870
rect 20110 -960 20370 -870
rect 20450 -960 20710 -870
rect 20790 -960 21050 -870
rect 21130 -960 21390 -870
rect 21470 -960 21730 -870
rect 21810 -960 22070 -870
rect 22150 -960 22410 -870
rect 22490 -960 22750 -870
rect 22830 -960 23090 -870
rect 23170 -960 23430 -870
rect 23510 -960 23770 -870
rect 23850 -960 24110 -870
rect 24190 -960 24450 -870
rect 24530 -960 24790 -870
rect 24870 -960 25130 -870
rect 25210 -960 25470 -870
rect 25550 -960 25810 -870
rect 25890 -960 26150 -870
rect 26230 -960 26490 -870
rect 26570 -960 26830 -870
rect 26910 -960 27170 -870
rect 27250 -960 27510 -870
rect 27590 -960 27850 -870
rect 27930 -960 28190 -870
rect 28270 -960 28530 -870
rect 28610 -960 28870 -870
rect 28950 -960 29210 -870
rect 29290 -960 29550 -870
rect 29630 -960 29890 -870
rect 29970 -960 30230 -870
rect 30310 -960 30570 -870
rect 30650 -960 30910 -870
rect 30990 -960 31250 -870
rect 31330 -960 31590 -870
rect 31670 -960 31930 -870
rect 32010 -960 32270 -870
rect 32350 -960 32610 -870
rect 32690 -960 32950 -870
rect 33030 -960 33290 -870
rect 33370 -960 33630 -870
rect 33710 -960 33970 -870
rect 34050 -960 34310 -870
rect 34390 -960 34650 -870
rect 34730 -960 34990 -870
rect 35070 -960 35330 -870
rect 35410 -960 35670 -870
rect 35750 -960 36010 -870
rect 36090 -960 36350 -870
rect 36430 -960 36690 -870
rect 36770 -960 37030 -870
rect 37110 -960 37370 -870
rect 37450 -960 37710 -870
rect 37790 -960 38050 -870
rect 38130 -960 38390 -870
rect 38470 -960 38730 -870
rect 38810 -960 39070 -870
rect 39150 -960 39410 -870
rect 39490 -960 39750 -870
rect 39830 -960 40090 -870
rect 40170 -960 40430 -870
rect 40510 -960 40770 -870
rect 40850 -960 41110 -870
rect 41190 -960 41450 -870
rect 41530 -960 41790 -870
rect 41870 -960 42130 -870
rect 42210 -960 42470 -870
rect 42550 -960 42810 -870
rect 42890 -960 43150 -870
rect 43230 -960 43490 -870
rect 43570 -960 43830 -870
rect 43910 -960 44170 -870
rect 44250 -960 44510 -870
rect 44590 -960 44850 -870
rect 44930 -960 45190 -870
rect 45270 -960 45530 -870
rect 45610 -960 45870 -870
rect 45950 -960 46210 -870
rect 46290 -960 46550 -870
rect 46630 -960 46890 -870
rect 46970 -960 47230 -870
rect 47310 -960 47570 -870
rect 47650 -960 47910 -870
rect 47990 -960 48250 -870
rect 48330 -960 48590 -870
rect 48670 -960 48930 -870
rect 49010 -960 49270 -870
rect 49350 -960 49610 -870
rect 49690 -960 49950 -870
rect 50030 -960 50290 -870
rect 50370 -960 50630 -870
rect 50710 -960 50970 -870
rect 51050 -960 51310 -870
rect 51390 -960 51650 -870
rect 51730 -960 51990 -870
rect 52070 -960 52330 -870
rect 52410 -960 52670 -870
rect 52750 -960 53010 -870
rect 53090 -960 53350 -870
rect 53430 -960 53690 -870
rect 53770 -960 54030 -870
rect 54110 -960 54370 -870
rect 54450 -960 54710 -870
rect 54790 -960 55050 -870
rect 55130 -960 55390 -870
rect 55470 -960 55730 -870
rect 55810 -960 56070 -870
rect 56150 -960 56410 -870
rect 56490 -960 56750 -870
rect 56830 -960 57090 -870
rect 57170 -960 57430 -870
rect 57510 -960 57770 -870
rect 57850 -960 58110 -870
rect 58190 -960 58450 -870
rect 58530 -960 58790 -870
rect 58870 -960 59130 -870
rect 59210 -960 59470 -870
rect 59550 -960 59810 -870
rect 59890 -960 60150 -870
rect 60230 -960 60490 -870
rect 60570 -960 60830 -870
rect 60910 -960 61170 -870
rect 61250 -960 61510 -870
rect 61590 -960 61850 -870
rect 61930 -960 62190 -870
rect 62270 -960 62530 -870
rect 62610 -960 62870 -870
rect 62950 -960 63210 -870
rect 63290 -960 63550 -870
rect 63630 -960 63890 -870
rect 63970 -960 64230 -870
rect 64310 -960 64570 -870
rect 64650 -960 64910 -870
rect 64990 -960 65250 -870
rect 65330 -960 65590 -870
rect 65670 -960 65930 -870
rect 66010 -960 66270 -870
rect 66350 -960 66610 -870
rect 66690 -960 66950 -870
rect 67030 -960 67290 -870
rect 67370 -960 67630 -870
rect 67710 -960 67970 -870
rect 68050 -960 68310 -870
rect 68390 -960 68650 -870
rect 68730 -960 68990 -870
rect 69070 -960 69330 -870
rect 69410 -960 69670 -870
rect 69750 -960 70010 -870
rect 70090 -960 70350 -870
rect 70430 -960 70690 -870
rect 70770 -960 71030 -870
rect 71110 -960 71370 -870
rect 71450 -960 71710 -870
rect 71790 -960 72050 -870
rect 72130 -960 72390 -870
rect 72470 -960 72730 -870
rect 72810 -960 73070 -870
rect 73150 -960 73410 -870
rect 73490 -960 73750 -870
rect 73830 -960 74090 -870
rect 74170 -960 74430 -870
rect 74510 -960 74770 -870
rect 74850 -960 75110 -870
rect 75190 -960 75450 -870
rect 75530 -960 75790 -870
rect 75870 -960 76130 -870
rect 76210 -960 76470 -870
rect 76550 -960 76810 -870
rect 76890 -960 77150 -870
rect 77230 -960 77490 -870
rect 77570 -960 77830 -870
rect 77910 -960 78170 -870
rect 78250 -960 78510 -870
rect 78590 -960 78850 -870
rect 78930 -960 79190 -870
rect 79270 -960 79530 -870
rect 79610 -960 79870 -870
rect 79950 -960 80210 -870
rect 80290 -960 80550 -870
rect 80630 -960 80890 -870
rect 80970 -960 81230 -870
rect 81310 -960 81570 -870
rect 81650 -960 81910 -870
rect 81990 -960 82250 -870
rect 82330 -960 82590 -870
rect 82670 -960 82930 -870
rect 83010 -960 83270 -870
rect 83350 -960 83610 -870
rect 83690 -960 83950 -870
rect 84030 -960 84290 -870
rect 84370 -960 84630 -870
rect 84710 -960 84970 -870
rect 85050 -960 85310 -870
rect 85390 -960 85650 -870
rect 85730 -960 85990 -870
rect 86070 -960 86330 -870
rect 86410 -960 86670 -870
rect 86750 -960 87010 -870
rect 87090 -960 87300 -870
rect -940 -970 87300 -960
rect -940 -1010 550 -970
rect -940 -1040 360 -1010
rect -490 -1340 -210 -1320
rect -490 -1400 -470 -1340
rect -560 -1550 -470 -1400
rect -490 -1610 -470 -1550
rect -210 -1420 390 -1400
rect -210 -1430 87320 -1420
rect -210 -1520 120 -1430
rect 240 -1470 1480 -1430
rect 240 -1520 830 -1470
rect -210 -1530 830 -1520
rect -210 -1550 390 -1530
rect 770 -1540 830 -1530
rect 910 -1520 1480 -1470
rect 1600 -1520 2840 -1430
rect 2960 -1520 4200 -1430
rect 4320 -1470 5560 -1430
rect 4320 -1520 5000 -1470
rect 910 -1530 5000 -1520
rect 910 -1540 970 -1530
rect 770 -1570 970 -1540
rect 4940 -1540 5000 -1530
rect 5080 -1520 5560 -1470
rect 5680 -1520 6920 -1430
rect 7040 -1520 8280 -1430
rect 8400 -1470 9640 -1430
rect 8400 -1520 9030 -1470
rect 5080 -1530 9030 -1520
rect 5080 -1540 5140 -1530
rect 4940 -1570 5140 -1540
rect 8970 -1540 9030 -1530
rect 9110 -1520 9640 -1470
rect 9760 -1520 11000 -1430
rect 11120 -1520 12360 -1430
rect 12480 -1470 13720 -1430
rect 12480 -1520 13060 -1470
rect 9110 -1530 13060 -1520
rect 9110 -1540 9170 -1530
rect 8970 -1570 9170 -1540
rect 13000 -1540 13060 -1530
rect 13140 -1520 13720 -1470
rect 13840 -1520 15080 -1430
rect 15200 -1520 16440 -1430
rect 16560 -1470 17800 -1430
rect 16560 -1520 17100 -1470
rect 13140 -1530 17100 -1520
rect 13140 -1540 13200 -1530
rect 13000 -1570 13200 -1540
rect 17040 -1540 17100 -1530
rect 17180 -1520 17800 -1470
rect 17920 -1520 19160 -1430
rect 19280 -1520 20520 -1430
rect 20640 -1470 21880 -1430
rect 20640 -1520 21200 -1470
rect 17180 -1530 21200 -1520
rect 17180 -1540 17240 -1530
rect 17040 -1570 17240 -1540
rect 21140 -1540 21200 -1530
rect 21280 -1520 21880 -1470
rect 22000 -1520 23240 -1430
rect 23360 -1520 24600 -1430
rect 24720 -1470 25960 -1430
rect 24720 -1520 25310 -1470
rect 21280 -1530 25310 -1520
rect 21280 -1540 21340 -1530
rect 21140 -1570 21340 -1540
rect 25250 -1540 25310 -1530
rect 25390 -1520 25960 -1470
rect 26080 -1520 27320 -1430
rect 27440 -1520 28680 -1430
rect 28800 -1470 30040 -1430
rect 28800 -1520 29410 -1470
rect 25390 -1530 29410 -1520
rect 25390 -1540 25450 -1530
rect 25250 -1570 25450 -1540
rect 29350 -1540 29410 -1530
rect 29490 -1520 30040 -1470
rect 30160 -1520 31400 -1430
rect 31520 -1520 32760 -1430
rect 32880 -1470 34120 -1430
rect 32880 -1520 33440 -1470
rect 29490 -1530 33440 -1520
rect 29490 -1540 29550 -1530
rect 29350 -1570 29550 -1540
rect 33380 -1540 33440 -1530
rect 33520 -1520 34120 -1470
rect 34240 -1520 35480 -1430
rect 35600 -1520 36840 -1430
rect 36960 -1470 38200 -1430
rect 36960 -1520 37550 -1470
rect 33520 -1530 37550 -1520
rect 33520 -1540 33580 -1530
rect 33380 -1570 33580 -1540
rect 37490 -1540 37550 -1530
rect 37630 -1520 38200 -1470
rect 38320 -1520 39560 -1430
rect 39680 -1520 40920 -1430
rect 41040 -1470 42280 -1430
rect 41040 -1520 41650 -1470
rect 37630 -1530 41650 -1520
rect 37630 -1540 37690 -1530
rect 37490 -1570 37690 -1540
rect 41590 -1540 41650 -1530
rect 41730 -1520 42280 -1470
rect 42400 -1520 43640 -1430
rect 43760 -1520 45000 -1430
rect 45120 -1520 46360 -1430
rect 46480 -1470 47720 -1430
rect 46480 -1520 47100 -1470
rect 41730 -1530 47100 -1520
rect 41730 -1540 41790 -1530
rect 41590 -1570 41790 -1540
rect 47040 -1540 47100 -1530
rect 47180 -1520 47720 -1470
rect 47840 -1520 49080 -1430
rect 49200 -1520 50440 -1430
rect 50560 -1470 51800 -1430
rect 50560 -1520 51180 -1470
rect 47180 -1530 51180 -1520
rect 47180 -1540 47240 -1530
rect 47040 -1570 47240 -1540
rect 51120 -1540 51180 -1530
rect 51260 -1520 51800 -1470
rect 51920 -1520 53160 -1430
rect 53280 -1520 54520 -1430
rect 54640 -1470 55880 -1430
rect 54640 -1520 55290 -1470
rect 51260 -1530 55290 -1520
rect 51260 -1540 51320 -1530
rect 51120 -1570 51320 -1540
rect 55230 -1540 55290 -1530
rect 55370 -1520 55880 -1470
rect 56000 -1520 57240 -1430
rect 57360 -1520 58600 -1430
rect 58720 -1470 59960 -1430
rect 58720 -1520 59320 -1470
rect 55370 -1530 59320 -1520
rect 55370 -1540 55430 -1530
rect 55230 -1570 55430 -1540
rect 59260 -1540 59320 -1530
rect 59400 -1520 59960 -1470
rect 60080 -1520 61320 -1430
rect 61440 -1520 62680 -1430
rect 62800 -1470 64040 -1430
rect 62800 -1520 63420 -1470
rect 59400 -1530 63420 -1520
rect 59400 -1540 59460 -1530
rect 59260 -1570 59460 -1540
rect 63360 -1540 63420 -1530
rect 63500 -1520 64040 -1470
rect 64160 -1520 65400 -1430
rect 65520 -1520 66760 -1430
rect 66880 -1470 68120 -1430
rect 66880 -1520 67530 -1470
rect 63500 -1530 67530 -1520
rect 63500 -1540 63560 -1530
rect 63360 -1570 63560 -1540
rect 67470 -1540 67530 -1530
rect 67610 -1520 68120 -1470
rect 68240 -1520 69480 -1430
rect 69600 -1520 70840 -1430
rect 70960 -1470 72200 -1430
rect 70960 -1520 71560 -1470
rect 67610 -1530 71560 -1520
rect 67610 -1540 67670 -1530
rect 67470 -1570 67670 -1540
rect 71500 -1540 71560 -1530
rect 71640 -1520 72200 -1470
rect 72320 -1520 73560 -1430
rect 73680 -1520 74920 -1430
rect 75040 -1470 76280 -1430
rect 75040 -1520 75810 -1470
rect 71640 -1530 75810 -1520
rect 71640 -1540 71700 -1530
rect 71500 -1570 71700 -1540
rect 75750 -1540 75810 -1530
rect 75890 -1520 76280 -1470
rect 76400 -1520 77640 -1430
rect 77760 -1520 79000 -1430
rect 79120 -1470 80360 -1430
rect 79120 -1520 79770 -1470
rect 75890 -1530 79770 -1520
rect 75890 -1540 75950 -1530
rect 75750 -1570 75950 -1540
rect 79710 -1540 79770 -1530
rect 79850 -1520 80360 -1470
rect 80480 -1520 81720 -1430
rect 81840 -1520 83080 -1430
rect 83200 -1470 84440 -1430
rect 83200 -1520 83950 -1470
rect 79850 -1530 83950 -1520
rect 79850 -1540 79910 -1530
rect 79710 -1570 79910 -1540
rect 83890 -1540 83950 -1530
rect 84030 -1520 84440 -1470
rect 84560 -1520 85800 -1430
rect 85920 -1474 87320 -1430
rect 85920 -1520 86508 -1474
rect 84030 -1530 86508 -1520
rect 84030 -1540 84090 -1530
rect 83890 -1570 84090 -1540
rect 86450 -1544 86508 -1530
rect 86588 -1530 87320 -1474
rect 86588 -1534 86650 -1530
rect 86588 -1544 86648 -1534
rect 86450 -1572 86648 -1544
rect -490 -1630 -210 -1610
<< via4 >>
rect -460 400 -200 670
rect -470 -1610 -210 -1340
<< metal5 >>
rect -560 670 -140 800
rect -560 400 -460 670
rect -200 400 -140 670
rect -560 -1340 -140 400
rect -560 -1610 -470 -1340
rect -210 -1610 -140 -1340
rect -560 -1820 -140 -1610
<< labels >>
rlabel metal2 370 -100 370 -100 1 in1
rlabel metal2 1460 -90 1460 -90 1 in2
rlabel metal2 4540 -100 4540 -100 1 in2
rlabel metal2 4540 -100 4540 -100 1 in3
rlabel metal2 15720 -90 15720 -90 1 in4
rlabel metal3 59100 -190 59100 -190 1 in5
rlabel metal2 -760 60 -760 60 1 in
rlabel metal4 -740 -910 -740 -910 1 out
rlabel metal4 -102 556 -102 556 1 vdd!
rlabel metal4 -114 -332 -114 -332 1 gnd!
<< end >>
