magic
tech sky130A
timestamp 1640608635
<< nmos >>
rect -5 0 30 720
<< ndiff >>
rect -95 700 -5 720
rect -95 650 -75 700
rect -25 650 -5 700
rect -95 595 -5 650
rect -95 545 -75 595
rect -25 545 -5 595
rect -95 490 -5 545
rect -95 440 -75 490
rect -25 440 -5 490
rect -95 385 -5 440
rect -95 335 -75 385
rect -25 335 -5 385
rect -95 280 -5 335
rect -95 230 -75 280
rect -25 230 -5 280
rect -95 175 -5 230
rect -95 125 -75 175
rect -25 125 -5 175
rect -95 70 -5 125
rect -95 20 -75 70
rect -25 20 -5 70
rect -95 0 -5 20
rect 30 700 120 720
rect 30 650 50 700
rect 100 650 120 700
rect 30 595 120 650
rect 30 545 50 595
rect 100 545 120 595
rect 30 490 120 545
rect 30 440 50 490
rect 100 440 120 490
rect 30 385 120 440
rect 30 335 50 385
rect 100 335 120 385
rect 30 280 120 335
rect 30 230 50 280
rect 100 230 120 280
rect 30 175 120 230
rect 30 125 50 175
rect 100 125 120 175
rect 30 70 120 125
rect 30 20 50 70
rect 100 20 120 70
rect 30 0 120 20
<< ndiffc >>
rect -75 650 -25 700
rect -75 545 -25 595
rect -75 440 -25 490
rect -75 335 -25 385
rect -75 230 -25 280
rect -75 125 -25 175
rect -75 20 -25 70
rect 50 650 100 700
rect 50 545 100 595
rect 50 440 100 490
rect 50 335 100 385
rect 50 230 100 280
rect 50 125 100 175
rect 50 20 100 70
<< poly >>
rect -20 790 50 800
rect -20 740 -10 790
rect 40 740 50 790
rect -20 730 50 740
rect -5 720 30 730
rect -5 -20 30 0
<< polycont >>
rect -10 740 40 790
<< locali >>
rect -20 790 50 800
rect -20 740 -10 790
rect 40 740 50 790
rect -20 730 50 740
rect -85 700 -15 710
rect -85 650 -75 700
rect -25 650 -15 700
rect -85 595 -15 650
rect -85 545 -75 595
rect -25 545 -15 595
rect -85 490 -15 545
rect -85 440 -75 490
rect -25 440 -15 490
rect -85 385 -15 440
rect -85 335 -75 385
rect -25 335 -15 385
rect -85 280 -15 335
rect -85 230 -75 280
rect -25 230 -15 280
rect -85 175 -15 230
rect -85 125 -75 175
rect -25 125 -15 175
rect -85 70 -15 125
rect -85 20 -75 70
rect -25 20 -15 70
rect -85 10 -15 20
rect 40 700 110 710
rect 40 650 50 700
rect 100 650 110 700
rect 40 595 110 650
rect 40 545 50 595
rect 100 545 110 595
rect 40 490 110 545
rect 40 440 50 490
rect 100 440 110 490
rect 40 385 110 440
rect 40 335 50 385
rect 100 335 110 385
rect 40 280 110 335
rect 40 230 50 280
rect 100 230 110 280
rect 40 175 110 230
rect 40 125 50 175
rect 100 125 110 175
rect 40 70 110 125
rect 40 20 50 70
rect 100 20 110 70
rect 40 10 110 20
<< labels >>
rlabel locali 10 795 10 795 1 vcont
rlabel locali -75 705 -75 705 1 vin
rlabel locali 105 705 105 705 1 vout
<< end >>
