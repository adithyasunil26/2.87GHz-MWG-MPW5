magic
tech sky130A
magscale 1 2
timestamp 1641278308
<< nmos >>
rect 350 0 380 500
rect 580 0 610 500
rect 810 0 840 500
rect 1040 0 1070 500
rect 1270 0 1300 500
rect 1500 0 1530 500
rect 1730 0 1760 500
rect 1960 0 1990 500
rect 2190 0 2220 500
rect 2420 0 2450 500
rect 2650 0 2680 500
rect 2880 0 2910 500
rect 3110 0 3140 500
rect 3340 0 3370 500
rect 3570 0 3600 500
rect 3800 0 3830 500
rect 4030 0 4060 500
rect 4260 0 4290 500
rect 4490 0 4520 500
rect 4720 0 4750 500
rect 4950 0 4980 500
rect 5180 0 5210 500
rect 5410 0 5440 500
rect 5640 0 5670 500
rect 5870 0 5900 500
rect 6100 0 6130 500
rect 6330 0 6360 500
rect 6560 0 6590 500
rect 6790 0 6820 500
rect 7020 0 7050 500
rect 350 -710 380 -210
rect 580 -710 610 -210
rect 810 -710 840 -210
rect 1040 -710 1070 -210
rect 1270 -710 1300 -210
rect 1500 -710 1530 -210
rect 1730 -710 1760 -210
rect 1960 -710 1990 -210
rect 2190 -710 2220 -210
rect 2420 -710 2450 -210
rect 2650 -710 2680 -210
rect 2880 -710 2910 -210
rect 3110 -710 3140 -210
rect 3340 -710 3370 -210
rect 3570 -710 3600 -210
rect 3800 -710 3830 -210
rect 4030 -710 4060 -210
rect 4260 -710 4290 -210
rect 4490 -710 4520 -210
rect 4720 -710 4750 -210
rect 4950 -710 4980 -210
rect 5180 -710 5210 -210
rect 5410 -710 5440 -210
rect 5640 -710 5670 -210
rect 5870 -710 5900 -210
rect 6100 -710 6130 -210
rect 6330 -710 6360 -210
rect 6560 -710 6590 -210
rect 6790 -710 6820 -210
rect 7020 -710 7050 -210
<< ndiff >>
rect 150 450 350 500
rect 150 350 200 450
rect 300 350 350 450
rect 150 150 350 350
rect 150 50 200 150
rect 300 50 350 150
rect 150 0 350 50
rect 380 450 580 500
rect 380 350 430 450
rect 530 350 580 450
rect 380 150 580 350
rect 380 50 430 150
rect 530 50 580 150
rect 380 0 580 50
rect 610 450 810 500
rect 610 350 660 450
rect 760 350 810 450
rect 610 150 810 350
rect 610 50 660 150
rect 760 50 810 150
rect 610 0 810 50
rect 840 450 1040 500
rect 840 350 890 450
rect 990 350 1040 450
rect 840 150 1040 350
rect 840 50 890 150
rect 990 50 1040 150
rect 840 0 1040 50
rect 1070 450 1270 500
rect 1070 350 1120 450
rect 1220 350 1270 450
rect 1070 150 1270 350
rect 1070 50 1120 150
rect 1220 50 1270 150
rect 1070 0 1270 50
rect 1300 450 1500 500
rect 1300 350 1350 450
rect 1450 350 1500 450
rect 1300 150 1500 350
rect 1300 50 1350 150
rect 1450 50 1500 150
rect 1300 0 1500 50
rect 1530 450 1730 500
rect 1530 350 1580 450
rect 1680 350 1730 450
rect 1530 150 1730 350
rect 1530 50 1580 150
rect 1680 50 1730 150
rect 1530 0 1730 50
rect 1760 450 1960 500
rect 1760 350 1810 450
rect 1910 350 1960 450
rect 1760 150 1960 350
rect 1760 50 1810 150
rect 1910 50 1960 150
rect 1760 0 1960 50
rect 1990 450 2190 500
rect 1990 350 2040 450
rect 2140 350 2190 450
rect 1990 150 2190 350
rect 1990 50 2040 150
rect 2140 50 2190 150
rect 1990 0 2190 50
rect 2220 450 2420 500
rect 2220 350 2270 450
rect 2370 350 2420 450
rect 2220 150 2420 350
rect 2220 50 2270 150
rect 2370 50 2420 150
rect 2220 0 2420 50
rect 2450 450 2650 500
rect 2450 350 2500 450
rect 2600 350 2650 450
rect 2450 150 2650 350
rect 2450 50 2500 150
rect 2600 50 2650 150
rect 2450 0 2650 50
rect 2680 450 2880 500
rect 2680 350 2730 450
rect 2830 350 2880 450
rect 2680 150 2880 350
rect 2680 50 2730 150
rect 2830 50 2880 150
rect 2680 0 2880 50
rect 2910 450 3110 500
rect 2910 350 2960 450
rect 3060 350 3110 450
rect 2910 150 3110 350
rect 2910 50 2960 150
rect 3060 50 3110 150
rect 2910 0 3110 50
rect 3140 450 3340 500
rect 3140 350 3190 450
rect 3290 350 3340 450
rect 3140 150 3340 350
rect 3140 50 3190 150
rect 3290 50 3340 150
rect 3140 0 3340 50
rect 3370 450 3570 500
rect 3370 350 3420 450
rect 3520 350 3570 450
rect 3370 150 3570 350
rect 3370 50 3420 150
rect 3520 50 3570 150
rect 3370 0 3570 50
rect 3600 450 3800 500
rect 3600 350 3650 450
rect 3750 350 3800 450
rect 3600 150 3800 350
rect 3600 50 3650 150
rect 3750 50 3800 150
rect 3600 0 3800 50
rect 3830 450 4030 500
rect 3830 350 3880 450
rect 3980 350 4030 450
rect 3830 150 4030 350
rect 3830 50 3880 150
rect 3980 50 4030 150
rect 3830 0 4030 50
rect 4060 450 4260 500
rect 4060 350 4110 450
rect 4210 350 4260 450
rect 4060 150 4260 350
rect 4060 50 4110 150
rect 4210 50 4260 150
rect 4060 0 4260 50
rect 4290 450 4490 500
rect 4290 350 4340 450
rect 4440 350 4490 450
rect 4290 150 4490 350
rect 4290 50 4340 150
rect 4440 50 4490 150
rect 4290 0 4490 50
rect 4520 450 4720 500
rect 4520 350 4570 450
rect 4670 350 4720 450
rect 4520 150 4720 350
rect 4520 50 4570 150
rect 4670 50 4720 150
rect 4520 0 4720 50
rect 4750 450 4950 500
rect 4750 350 4800 450
rect 4900 350 4950 450
rect 4750 150 4950 350
rect 4750 50 4800 150
rect 4900 50 4950 150
rect 4750 0 4950 50
rect 4980 450 5180 500
rect 4980 350 5030 450
rect 5130 350 5180 450
rect 4980 150 5180 350
rect 4980 50 5030 150
rect 5130 50 5180 150
rect 4980 0 5180 50
rect 5210 450 5410 500
rect 5210 350 5260 450
rect 5360 350 5410 450
rect 5210 150 5410 350
rect 5210 50 5260 150
rect 5360 50 5410 150
rect 5210 0 5410 50
rect 5440 450 5640 500
rect 5440 350 5490 450
rect 5590 350 5640 450
rect 5440 150 5640 350
rect 5440 50 5490 150
rect 5590 50 5640 150
rect 5440 0 5640 50
rect 5670 450 5870 500
rect 5670 350 5720 450
rect 5820 350 5870 450
rect 5670 150 5870 350
rect 5670 50 5720 150
rect 5820 50 5870 150
rect 5670 0 5870 50
rect 5900 450 6100 500
rect 5900 350 5950 450
rect 6050 350 6100 450
rect 5900 150 6100 350
rect 5900 50 5950 150
rect 6050 50 6100 150
rect 5900 0 6100 50
rect 6130 450 6330 500
rect 6130 350 6180 450
rect 6280 350 6330 450
rect 6130 150 6330 350
rect 6130 50 6180 150
rect 6280 50 6330 150
rect 6130 0 6330 50
rect 6360 450 6560 500
rect 6360 350 6410 450
rect 6510 350 6560 450
rect 6360 150 6560 350
rect 6360 50 6410 150
rect 6510 50 6560 150
rect 6360 0 6560 50
rect 6590 450 6790 500
rect 6590 350 6640 450
rect 6740 350 6790 450
rect 6590 150 6790 350
rect 6590 50 6640 150
rect 6740 50 6790 150
rect 6590 0 6790 50
rect 6820 450 7020 500
rect 6820 350 6870 450
rect 6970 350 7020 450
rect 6820 150 7020 350
rect 6820 50 6870 150
rect 6970 50 7020 150
rect 6820 0 7020 50
rect 7050 450 7250 500
rect 7050 350 7100 450
rect 7200 350 7250 450
rect 7050 150 7250 350
rect 7050 50 7100 150
rect 7200 50 7250 150
rect 7050 0 7250 50
rect 150 -260 350 -210
rect 150 -360 200 -260
rect 300 -360 350 -260
rect 150 -560 350 -360
rect 150 -660 200 -560
rect 300 -660 350 -560
rect 150 -710 350 -660
rect 380 -260 580 -210
rect 380 -360 430 -260
rect 530 -360 580 -260
rect 380 -560 580 -360
rect 380 -660 430 -560
rect 530 -660 580 -560
rect 380 -710 580 -660
rect 610 -260 810 -210
rect 610 -360 660 -260
rect 760 -360 810 -260
rect 610 -560 810 -360
rect 610 -660 660 -560
rect 760 -660 810 -560
rect 610 -710 810 -660
rect 840 -260 1040 -210
rect 840 -360 890 -260
rect 990 -360 1040 -260
rect 840 -560 1040 -360
rect 840 -660 890 -560
rect 990 -660 1040 -560
rect 840 -710 1040 -660
rect 1070 -260 1270 -210
rect 1070 -360 1120 -260
rect 1220 -360 1270 -260
rect 1070 -560 1270 -360
rect 1070 -660 1120 -560
rect 1220 -660 1270 -560
rect 1070 -710 1270 -660
rect 1300 -260 1500 -210
rect 1300 -360 1350 -260
rect 1450 -360 1500 -260
rect 1300 -560 1500 -360
rect 1300 -660 1350 -560
rect 1450 -660 1500 -560
rect 1300 -710 1500 -660
rect 1530 -260 1730 -210
rect 1530 -360 1580 -260
rect 1680 -360 1730 -260
rect 1530 -560 1730 -360
rect 1530 -660 1580 -560
rect 1680 -660 1730 -560
rect 1530 -710 1730 -660
rect 1760 -260 1960 -210
rect 1760 -360 1810 -260
rect 1910 -360 1960 -260
rect 1760 -560 1960 -360
rect 1760 -660 1810 -560
rect 1910 -660 1960 -560
rect 1760 -710 1960 -660
rect 1990 -260 2190 -210
rect 1990 -360 2040 -260
rect 2140 -360 2190 -260
rect 1990 -560 2190 -360
rect 1990 -660 2040 -560
rect 2140 -660 2190 -560
rect 1990 -710 2190 -660
rect 2220 -260 2420 -210
rect 2220 -360 2270 -260
rect 2370 -360 2420 -260
rect 2220 -560 2420 -360
rect 2220 -660 2270 -560
rect 2370 -660 2420 -560
rect 2220 -710 2420 -660
rect 2450 -260 2650 -210
rect 2450 -360 2500 -260
rect 2600 -360 2650 -260
rect 2450 -560 2650 -360
rect 2450 -660 2500 -560
rect 2600 -660 2650 -560
rect 2450 -710 2650 -660
rect 2680 -260 2880 -210
rect 2680 -360 2730 -260
rect 2830 -360 2880 -260
rect 2680 -560 2880 -360
rect 2680 -660 2730 -560
rect 2830 -660 2880 -560
rect 2680 -710 2880 -660
rect 2910 -260 3110 -210
rect 2910 -360 2960 -260
rect 3060 -360 3110 -260
rect 2910 -560 3110 -360
rect 2910 -660 2960 -560
rect 3060 -660 3110 -560
rect 2910 -710 3110 -660
rect 3140 -260 3340 -210
rect 3140 -360 3190 -260
rect 3290 -360 3340 -260
rect 3140 -560 3340 -360
rect 3140 -660 3190 -560
rect 3290 -660 3340 -560
rect 3140 -710 3340 -660
rect 3370 -260 3570 -210
rect 3370 -360 3420 -260
rect 3520 -360 3570 -260
rect 3370 -560 3570 -360
rect 3370 -660 3420 -560
rect 3520 -660 3570 -560
rect 3370 -710 3570 -660
rect 3600 -260 3800 -210
rect 3600 -360 3650 -260
rect 3750 -360 3800 -260
rect 3600 -560 3800 -360
rect 3600 -660 3650 -560
rect 3750 -660 3800 -560
rect 3600 -710 3800 -660
rect 3830 -260 4030 -210
rect 3830 -360 3880 -260
rect 3980 -360 4030 -260
rect 3830 -560 4030 -360
rect 3830 -660 3880 -560
rect 3980 -660 4030 -560
rect 3830 -710 4030 -660
rect 4060 -260 4260 -210
rect 4060 -360 4110 -260
rect 4210 -360 4260 -260
rect 4060 -560 4260 -360
rect 4060 -660 4110 -560
rect 4210 -660 4260 -560
rect 4060 -710 4260 -660
rect 4290 -260 4490 -210
rect 4290 -360 4340 -260
rect 4440 -360 4490 -260
rect 4290 -560 4490 -360
rect 4290 -660 4340 -560
rect 4440 -660 4490 -560
rect 4290 -710 4490 -660
rect 4520 -260 4720 -210
rect 4520 -360 4570 -260
rect 4670 -360 4720 -260
rect 4520 -560 4720 -360
rect 4520 -660 4570 -560
rect 4670 -660 4720 -560
rect 4520 -710 4720 -660
rect 4750 -260 4950 -210
rect 4750 -360 4800 -260
rect 4900 -360 4950 -260
rect 4750 -560 4950 -360
rect 4750 -660 4800 -560
rect 4900 -660 4950 -560
rect 4750 -710 4950 -660
rect 4980 -260 5180 -210
rect 4980 -360 5030 -260
rect 5130 -360 5180 -260
rect 4980 -560 5180 -360
rect 4980 -660 5030 -560
rect 5130 -660 5180 -560
rect 4980 -710 5180 -660
rect 5210 -260 5410 -210
rect 5210 -360 5260 -260
rect 5360 -360 5410 -260
rect 5210 -560 5410 -360
rect 5210 -660 5260 -560
rect 5360 -660 5410 -560
rect 5210 -710 5410 -660
rect 5440 -260 5640 -210
rect 5440 -360 5490 -260
rect 5590 -360 5640 -260
rect 5440 -560 5640 -360
rect 5440 -660 5490 -560
rect 5590 -660 5640 -560
rect 5440 -710 5640 -660
rect 5670 -260 5870 -210
rect 5670 -360 5720 -260
rect 5820 -360 5870 -260
rect 5670 -560 5870 -360
rect 5670 -660 5720 -560
rect 5820 -660 5870 -560
rect 5670 -710 5870 -660
rect 5900 -260 6100 -210
rect 5900 -360 5950 -260
rect 6050 -360 6100 -260
rect 5900 -560 6100 -360
rect 5900 -660 5950 -560
rect 6050 -660 6100 -560
rect 5900 -710 6100 -660
rect 6130 -260 6330 -210
rect 6130 -360 6180 -260
rect 6280 -360 6330 -260
rect 6130 -560 6330 -360
rect 6130 -660 6180 -560
rect 6280 -660 6330 -560
rect 6130 -710 6330 -660
rect 6360 -260 6560 -210
rect 6360 -360 6410 -260
rect 6510 -360 6560 -260
rect 6360 -560 6560 -360
rect 6360 -660 6410 -560
rect 6510 -660 6560 -560
rect 6360 -710 6560 -660
rect 6590 -260 6790 -210
rect 6590 -360 6640 -260
rect 6740 -360 6790 -260
rect 6590 -560 6790 -360
rect 6590 -660 6640 -560
rect 6740 -660 6790 -560
rect 6590 -710 6790 -660
rect 6820 -260 7020 -210
rect 6820 -360 6870 -260
rect 6970 -360 7020 -260
rect 6820 -560 7020 -360
rect 6820 -660 6870 -560
rect 6970 -660 7020 -560
rect 6820 -710 7020 -660
rect 7050 -260 7250 -210
rect 7050 -360 7100 -260
rect 7200 -360 7250 -260
rect 7050 -560 7250 -360
rect 7050 -660 7100 -560
rect 7200 -660 7250 -560
rect 7050 -710 7250 -660
<< ndiffc >>
rect 200 350 300 450
rect 200 50 300 150
rect 430 350 530 450
rect 430 50 530 150
rect 660 350 760 450
rect 660 50 760 150
rect 890 350 990 450
rect 890 50 990 150
rect 1120 350 1220 450
rect 1120 50 1220 150
rect 1350 350 1450 450
rect 1350 50 1450 150
rect 1580 350 1680 450
rect 1580 50 1680 150
rect 1810 350 1910 450
rect 1810 50 1910 150
rect 2040 350 2140 450
rect 2040 50 2140 150
rect 2270 350 2370 450
rect 2270 50 2370 150
rect 2500 350 2600 450
rect 2500 50 2600 150
rect 2730 350 2830 450
rect 2730 50 2830 150
rect 2960 350 3060 450
rect 2960 50 3060 150
rect 3190 350 3290 450
rect 3190 50 3290 150
rect 3420 350 3520 450
rect 3420 50 3520 150
rect 3650 350 3750 450
rect 3650 50 3750 150
rect 3880 350 3980 450
rect 3880 50 3980 150
rect 4110 350 4210 450
rect 4110 50 4210 150
rect 4340 350 4440 450
rect 4340 50 4440 150
rect 4570 350 4670 450
rect 4570 50 4670 150
rect 4800 350 4900 450
rect 4800 50 4900 150
rect 5030 350 5130 450
rect 5030 50 5130 150
rect 5260 350 5360 450
rect 5260 50 5360 150
rect 5490 350 5590 450
rect 5490 50 5590 150
rect 5720 350 5820 450
rect 5720 50 5820 150
rect 5950 350 6050 450
rect 5950 50 6050 150
rect 6180 350 6280 450
rect 6180 50 6280 150
rect 6410 350 6510 450
rect 6410 50 6510 150
rect 6640 350 6740 450
rect 6640 50 6740 150
rect 6870 350 6970 450
rect 6870 50 6970 150
rect 7100 350 7200 450
rect 7100 50 7200 150
rect 200 -360 300 -260
rect 200 -660 300 -560
rect 430 -360 530 -260
rect 430 -660 530 -560
rect 660 -360 760 -260
rect 660 -660 760 -560
rect 890 -360 990 -260
rect 890 -660 990 -560
rect 1120 -360 1220 -260
rect 1120 -660 1220 -560
rect 1350 -360 1450 -260
rect 1350 -660 1450 -560
rect 1580 -360 1680 -260
rect 1580 -660 1680 -560
rect 1810 -360 1910 -260
rect 1810 -660 1910 -560
rect 2040 -360 2140 -260
rect 2040 -660 2140 -560
rect 2270 -360 2370 -260
rect 2270 -660 2370 -560
rect 2500 -360 2600 -260
rect 2500 -660 2600 -560
rect 2730 -360 2830 -260
rect 2730 -660 2830 -560
rect 2960 -360 3060 -260
rect 2960 -660 3060 -560
rect 3190 -360 3290 -260
rect 3190 -660 3290 -560
rect 3420 -360 3520 -260
rect 3420 -660 3520 -560
rect 3650 -360 3750 -260
rect 3650 -660 3750 -560
rect 3880 -360 3980 -260
rect 3880 -660 3980 -560
rect 4110 -360 4210 -260
rect 4110 -660 4210 -560
rect 4340 -360 4440 -260
rect 4340 -660 4440 -560
rect 4570 -360 4670 -260
rect 4570 -660 4670 -560
rect 4800 -360 4900 -260
rect 4800 -660 4900 -560
rect 5030 -360 5130 -260
rect 5030 -660 5130 -560
rect 5260 -360 5360 -260
rect 5260 -660 5360 -560
rect 5490 -360 5590 -260
rect 5490 -660 5590 -560
rect 5720 -360 5820 -260
rect 5720 -660 5820 -560
rect 5950 -360 6050 -260
rect 5950 -660 6050 -560
rect 6180 -360 6280 -260
rect 6180 -660 6280 -560
rect 6410 -360 6510 -260
rect 6410 -660 6510 -560
rect 6640 -360 6740 -260
rect 6640 -660 6740 -560
rect 6870 -360 6970 -260
rect 6870 -660 6970 -560
rect 7100 -360 7200 -260
rect 7100 -660 7200 -560
<< psubdiff >>
rect -1780 1470 -1520 1500
rect -1780 1270 -1750 1470
rect -1550 1270 -1520 1470
rect -1780 1240 -1520 1270
rect -690 1470 -430 1500
rect -690 1270 -660 1470
rect -460 1270 -430 1470
rect -690 1240 -430 1270
rect 310 1470 570 1500
rect 310 1270 340 1470
rect 540 1270 570 1470
rect 310 1240 570 1270
rect 1310 1470 1570 1500
rect 1310 1270 1340 1470
rect 1540 1270 1570 1470
rect 1310 1240 1570 1270
rect 2330 1470 2590 1500
rect 2330 1270 2360 1470
rect 2560 1270 2590 1470
rect 2330 1240 2590 1270
rect 3330 1470 3590 1500
rect 3330 1270 3360 1470
rect 3560 1270 3590 1470
rect 3330 1240 3590 1270
rect 4330 1470 4590 1500
rect 4330 1270 4360 1470
rect 4560 1270 4590 1470
rect 4330 1240 4590 1270
rect 5350 1470 5610 1500
rect 5350 1270 5380 1470
rect 5580 1270 5610 1470
rect 5350 1240 5610 1270
rect 6350 1470 6610 1500
rect 6350 1270 6380 1470
rect 6580 1270 6610 1470
rect 6350 1240 6610 1270
rect 7350 1470 7610 1500
rect 7350 1270 7380 1470
rect 7580 1270 7610 1470
rect 7350 1240 7610 1270
rect -2230 820 -1970 850
rect -2230 620 -2200 820
rect -2000 620 -1970 820
rect 7740 830 8000 860
rect 7740 630 7770 830
rect 7970 630 8000 830
rect -2230 590 -1970 620
rect 7740 600 8000 630
rect -2230 -200 -1970 -170
rect -2230 -400 -2200 -200
rect -2000 -400 -1970 -200
rect 7740 -190 8000 -160
rect -2230 -430 -1970 -400
rect 7740 -390 7770 -190
rect 7970 -390 8000 -190
rect 7740 -420 8000 -390
rect -2230 -1200 -1970 -1170
rect -2230 -1400 -2200 -1200
rect -2000 -1400 -1970 -1200
rect -2230 -1430 -1970 -1400
rect 7740 -1190 8000 -1160
rect 7740 -1390 7770 -1190
rect 7970 -1390 8000 -1190
rect 7740 -1420 8000 -1390
rect -1810 -1470 -1550 -1440
rect -1810 -1670 -1780 -1470
rect -1580 -1670 -1550 -1470
rect -1810 -1700 -1550 -1670
rect -720 -1470 -460 -1440
rect -720 -1670 -690 -1470
rect -490 -1670 -460 -1470
rect -720 -1700 -460 -1670
rect 280 -1470 540 -1440
rect 280 -1670 310 -1470
rect 510 -1670 540 -1470
rect 280 -1700 540 -1670
rect 1280 -1470 1540 -1440
rect 1280 -1670 1310 -1470
rect 1510 -1670 1540 -1470
rect 1280 -1700 1540 -1670
rect 2300 -1470 2560 -1440
rect 2300 -1670 2330 -1470
rect 2530 -1670 2560 -1470
rect 2300 -1700 2560 -1670
rect 3300 -1470 3560 -1440
rect 3300 -1670 3330 -1470
rect 3530 -1670 3560 -1470
rect 3300 -1700 3560 -1670
rect 4300 -1470 4560 -1440
rect 4300 -1670 4330 -1470
rect 4530 -1670 4560 -1470
rect 4300 -1700 4560 -1670
rect 5320 -1470 5580 -1440
rect 5320 -1670 5350 -1470
rect 5550 -1670 5580 -1470
rect 5320 -1700 5580 -1670
rect 6320 -1470 6580 -1440
rect 6320 -1670 6350 -1470
rect 6550 -1670 6580 -1470
rect 6320 -1700 6580 -1670
rect 7320 -1470 7580 -1440
rect 7320 -1670 7350 -1470
rect 7550 -1670 7580 -1470
rect 7320 -1700 7580 -1670
<< psubdiffcont >>
rect -1750 1270 -1550 1470
rect -660 1270 -460 1470
rect 340 1270 540 1470
rect 1340 1270 1540 1470
rect 2360 1270 2560 1470
rect 3360 1270 3560 1470
rect 4360 1270 4560 1470
rect 5380 1270 5580 1470
rect 6380 1270 6580 1470
rect 7380 1270 7580 1470
rect -2200 620 -2000 820
rect 7770 630 7970 830
rect -2200 -400 -2000 -200
rect 7770 -390 7970 -190
rect -2200 -1400 -2000 -1200
rect 7770 -1390 7970 -1190
rect -1780 -1670 -1580 -1470
rect -690 -1670 -490 -1470
rect 310 -1670 510 -1470
rect 1310 -1670 1510 -1470
rect 2330 -1670 2530 -1470
rect 3330 -1670 3530 -1470
rect 4330 -1670 4530 -1470
rect 5350 -1670 5550 -1470
rect 6350 -1670 6550 -1470
rect 7350 -1670 7550 -1470
<< poly >>
rect 310 610 420 630
rect 310 540 330 610
rect 400 540 420 610
rect 310 520 420 540
rect 540 610 650 630
rect 540 540 560 610
rect 630 540 650 610
rect 540 520 650 540
rect 770 610 880 630
rect 770 540 790 610
rect 860 540 880 610
rect 770 520 880 540
rect 1000 610 1110 630
rect 1000 540 1020 610
rect 1090 540 1110 610
rect 1000 520 1110 540
rect 1230 610 1340 630
rect 1230 540 1250 610
rect 1320 540 1340 610
rect 1230 520 1340 540
rect 1460 610 1570 630
rect 1460 540 1480 610
rect 1550 540 1570 610
rect 1460 520 1570 540
rect 1690 610 1800 630
rect 1690 540 1710 610
rect 1780 540 1800 610
rect 1690 520 1800 540
rect 1920 610 2030 630
rect 1920 540 1940 610
rect 2010 540 2030 610
rect 1920 520 2030 540
rect 2150 610 2260 630
rect 2150 540 2170 610
rect 2240 540 2260 610
rect 2150 520 2260 540
rect 2380 610 2490 630
rect 2380 540 2400 610
rect 2470 540 2490 610
rect 2380 520 2490 540
rect 2610 610 2720 630
rect 2610 540 2630 610
rect 2700 540 2720 610
rect 2610 520 2720 540
rect 2840 610 2950 630
rect 2840 540 2860 610
rect 2930 540 2950 610
rect 2840 520 2950 540
rect 3070 610 3180 630
rect 3070 540 3090 610
rect 3160 540 3180 610
rect 3070 520 3180 540
rect 3300 610 3410 630
rect 3300 540 3320 610
rect 3390 540 3410 610
rect 3300 520 3410 540
rect 3530 610 3640 630
rect 3530 540 3550 610
rect 3620 540 3640 610
rect 3530 520 3640 540
rect 3760 610 3870 630
rect 3760 540 3780 610
rect 3850 540 3870 610
rect 3760 520 3870 540
rect 3990 610 4100 630
rect 3990 540 4010 610
rect 4080 540 4100 610
rect 3990 520 4100 540
rect 4220 610 4330 630
rect 4220 540 4240 610
rect 4310 540 4330 610
rect 4220 520 4330 540
rect 4450 610 4560 630
rect 4450 540 4470 610
rect 4540 540 4560 610
rect 4450 520 4560 540
rect 4680 610 4790 630
rect 4680 540 4700 610
rect 4770 540 4790 610
rect 4680 520 4790 540
rect 4910 610 5020 630
rect 4910 540 4930 610
rect 5000 540 5020 610
rect 4910 520 5020 540
rect 5140 610 5250 630
rect 5140 540 5160 610
rect 5230 540 5250 610
rect 5140 520 5250 540
rect 5370 610 5480 630
rect 5370 540 5390 610
rect 5460 540 5480 610
rect 5370 520 5480 540
rect 5600 610 5710 630
rect 5600 540 5620 610
rect 5690 540 5710 610
rect 5600 520 5710 540
rect 5830 610 5940 630
rect 5830 540 5850 610
rect 5920 540 5940 610
rect 5830 520 5940 540
rect 6060 610 6170 630
rect 6060 540 6080 610
rect 6150 540 6170 610
rect 6060 520 6170 540
rect 6290 610 6400 630
rect 6290 540 6310 610
rect 6380 540 6400 610
rect 6290 520 6400 540
rect 6520 610 6630 630
rect 6520 540 6540 610
rect 6610 540 6630 610
rect 6520 520 6630 540
rect 6750 610 6860 630
rect 6750 540 6770 610
rect 6840 540 6860 610
rect 6750 520 6860 540
rect 6980 610 7090 630
rect 6980 540 7000 610
rect 7070 540 7090 610
rect 6980 520 7090 540
rect 350 500 380 520
rect 580 500 610 520
rect 810 500 840 520
rect 1040 500 1070 520
rect 1270 500 1300 520
rect 1500 500 1530 520
rect 1730 500 1760 520
rect 1960 500 1990 520
rect 2190 500 2220 520
rect 2420 500 2450 520
rect 2650 500 2680 520
rect 2880 500 2910 520
rect 3110 500 3140 520
rect 3340 500 3370 520
rect 3570 500 3600 520
rect 3800 500 3830 520
rect 4030 500 4060 520
rect 4260 500 4290 520
rect 4490 500 4520 520
rect 4720 500 4750 520
rect 4950 500 4980 520
rect 5180 500 5210 520
rect 5410 500 5440 520
rect 5640 500 5670 520
rect 5870 500 5900 520
rect 6100 500 6130 520
rect 6330 500 6360 520
rect 6560 500 6590 520
rect 6790 500 6820 520
rect 7020 500 7050 520
rect 350 -30 380 0
rect 580 -30 610 0
rect 810 -30 840 0
rect 1040 -30 1070 0
rect 1270 -30 1300 0
rect 1500 -30 1530 0
rect 1730 -30 1760 0
rect 1960 -30 1990 0
rect 2190 -30 2220 0
rect 2420 -30 2450 0
rect 2650 -30 2680 0
rect 2880 -30 2910 0
rect 3110 -30 3140 0
rect 3340 -30 3370 0
rect 3570 -30 3600 0
rect 3800 -30 3830 0
rect 4030 -30 4060 0
rect 4260 -30 4290 0
rect 4490 -30 4520 0
rect 4720 -30 4750 0
rect 4950 -30 4980 0
rect 5180 -30 5210 0
rect 5410 -30 5440 0
rect 5640 -30 5670 0
rect 5870 -30 5900 0
rect 6100 -30 6130 0
rect 6330 -30 6360 0
rect 6560 -30 6590 0
rect 6790 -30 6820 0
rect 7020 -30 7050 0
rect 350 -210 380 -180
rect 580 -210 610 -180
rect 810 -210 840 -180
rect 1040 -210 1070 -180
rect 1270 -210 1300 -180
rect 1500 -210 1530 -180
rect 1730 -210 1760 -180
rect 1960 -210 1990 -180
rect 2190 -210 2220 -180
rect 2420 -210 2450 -180
rect 2650 -210 2680 -180
rect 2880 -210 2910 -180
rect 3110 -210 3140 -180
rect 3340 -210 3370 -180
rect 3570 -210 3600 -180
rect 3800 -210 3830 -180
rect 4030 -210 4060 -180
rect 4260 -210 4290 -180
rect 4490 -210 4520 -180
rect 4720 -210 4750 -180
rect 4950 -210 4980 -180
rect 5180 -210 5210 -180
rect 5410 -210 5440 -180
rect 5640 -210 5670 -180
rect 5870 -210 5900 -180
rect 6100 -210 6130 -180
rect 6330 -210 6360 -180
rect 6560 -210 6590 -180
rect 6790 -210 6820 -180
rect 7020 -210 7050 -180
rect 350 -730 380 -710
rect 580 -730 610 -710
rect 810 -730 840 -710
rect 1040 -730 1070 -710
rect 1270 -730 1300 -710
rect 1500 -730 1530 -710
rect 1730 -730 1760 -710
rect 1960 -730 1990 -710
rect 2190 -730 2220 -710
rect 2420 -730 2450 -710
rect 2650 -730 2680 -710
rect 2880 -730 2910 -710
rect 3110 -730 3140 -710
rect 3340 -730 3370 -710
rect 3570 -730 3600 -710
rect 3800 -730 3830 -710
rect 4030 -730 4060 -710
rect 4260 -730 4290 -710
rect 4490 -730 4520 -710
rect 4720 -730 4750 -710
rect 4950 -730 4980 -710
rect 5180 -730 5210 -710
rect 5410 -730 5440 -710
rect 5640 -730 5670 -710
rect 5870 -730 5900 -710
rect 6100 -730 6130 -710
rect 6330 -730 6360 -710
rect 6560 -730 6590 -710
rect 6790 -730 6820 -710
rect 7020 -730 7050 -710
rect 310 -750 420 -730
rect 310 -820 330 -750
rect 400 -820 420 -750
rect 310 -840 420 -820
rect 540 -750 650 -730
rect 540 -820 560 -750
rect 630 -820 650 -750
rect 540 -840 650 -820
rect 770 -750 880 -730
rect 770 -820 790 -750
rect 860 -820 880 -750
rect 770 -840 880 -820
rect 1000 -750 1110 -730
rect 1000 -820 1020 -750
rect 1090 -820 1110 -750
rect 1000 -840 1110 -820
rect 1230 -750 1340 -730
rect 1230 -820 1250 -750
rect 1320 -820 1340 -750
rect 1230 -840 1340 -820
rect 1460 -750 1570 -730
rect 1460 -820 1480 -750
rect 1550 -820 1570 -750
rect 1460 -840 1570 -820
rect 1690 -750 1800 -730
rect 1690 -820 1710 -750
rect 1780 -820 1800 -750
rect 1690 -840 1800 -820
rect 1920 -750 2030 -730
rect 1920 -820 1940 -750
rect 2010 -820 2030 -750
rect 1920 -840 2030 -820
rect 2150 -750 2260 -730
rect 2150 -820 2170 -750
rect 2240 -820 2260 -750
rect 2150 -840 2260 -820
rect 2380 -750 2490 -730
rect 2380 -820 2400 -750
rect 2470 -820 2490 -750
rect 2380 -840 2490 -820
rect 2610 -750 2720 -730
rect 2610 -820 2630 -750
rect 2700 -820 2720 -750
rect 2610 -840 2720 -820
rect 2840 -750 2950 -730
rect 2840 -820 2860 -750
rect 2930 -820 2950 -750
rect 2840 -840 2950 -820
rect 3070 -750 3180 -730
rect 3070 -820 3090 -750
rect 3160 -820 3180 -750
rect 3070 -840 3180 -820
rect 3300 -750 3410 -730
rect 3300 -820 3320 -750
rect 3390 -820 3410 -750
rect 3300 -840 3410 -820
rect 3530 -750 3640 -730
rect 3530 -820 3550 -750
rect 3620 -820 3640 -750
rect 3530 -840 3640 -820
rect 3760 -750 3870 -730
rect 3760 -820 3780 -750
rect 3850 -820 3870 -750
rect 3760 -840 3870 -820
rect 3990 -750 4100 -730
rect 3990 -820 4010 -750
rect 4080 -820 4100 -750
rect 3990 -840 4100 -820
rect 4220 -750 4330 -730
rect 4220 -820 4240 -750
rect 4310 -820 4330 -750
rect 4220 -840 4330 -820
rect 4450 -750 4560 -730
rect 4450 -820 4470 -750
rect 4540 -820 4560 -750
rect 4450 -840 4560 -820
rect 4680 -750 4790 -730
rect 4680 -820 4700 -750
rect 4770 -820 4790 -750
rect 4680 -840 4790 -820
rect 4910 -750 5020 -730
rect 4910 -820 4930 -750
rect 5000 -820 5020 -750
rect 4910 -840 5020 -820
rect 5140 -750 5250 -730
rect 5140 -820 5160 -750
rect 5230 -820 5250 -750
rect 5140 -840 5250 -820
rect 5370 -750 5480 -730
rect 5370 -820 5390 -750
rect 5460 -820 5480 -750
rect 5370 -840 5480 -820
rect 5600 -750 5710 -730
rect 5600 -820 5620 -750
rect 5690 -820 5710 -750
rect 5600 -840 5710 -820
rect 5830 -750 5940 -730
rect 5830 -820 5850 -750
rect 5920 -820 5940 -750
rect 5830 -840 5940 -820
rect 6060 -750 6170 -730
rect 6060 -820 6080 -750
rect 6150 -820 6170 -750
rect 6060 -840 6170 -820
rect 6290 -750 6400 -730
rect 6290 -820 6310 -750
rect 6380 -820 6400 -750
rect 6290 -840 6400 -820
rect 6520 -750 6630 -730
rect 6520 -820 6540 -750
rect 6610 -820 6630 -750
rect 6520 -840 6630 -820
rect 6750 -750 6860 -730
rect 6750 -820 6770 -750
rect 6840 -820 6860 -750
rect 6750 -840 6860 -820
rect 6980 -750 7090 -730
rect 6980 -820 7000 -750
rect 7070 -820 7090 -750
rect 6980 -840 7090 -820
<< polycont >>
rect 330 540 400 610
rect 560 540 630 610
rect 790 540 860 610
rect 1020 540 1090 610
rect 1250 540 1320 610
rect 1480 540 1550 610
rect 1710 540 1780 610
rect 1940 540 2010 610
rect 2170 540 2240 610
rect 2400 540 2470 610
rect 2630 540 2700 610
rect 2860 540 2930 610
rect 3090 540 3160 610
rect 3320 540 3390 610
rect 3550 540 3620 610
rect 3780 540 3850 610
rect 4010 540 4080 610
rect 4240 540 4310 610
rect 4470 540 4540 610
rect 4700 540 4770 610
rect 4930 540 5000 610
rect 5160 540 5230 610
rect 5390 540 5460 610
rect 5620 540 5690 610
rect 5850 540 5920 610
rect 6080 540 6150 610
rect 6310 540 6380 610
rect 6540 540 6610 610
rect 6770 540 6840 610
rect 7000 540 7070 610
rect 330 -820 400 -750
rect 560 -820 630 -750
rect 790 -820 860 -750
rect 1020 -820 1090 -750
rect 1250 -820 1320 -750
rect 1480 -820 1550 -750
rect 1710 -820 1780 -750
rect 1940 -820 2010 -750
rect 2170 -820 2240 -750
rect 2400 -820 2470 -750
rect 2630 -820 2700 -750
rect 2860 -820 2930 -750
rect 3090 -820 3160 -750
rect 3320 -820 3390 -750
rect 3550 -820 3620 -750
rect 3780 -820 3850 -750
rect 4010 -820 4080 -750
rect 4240 -820 4310 -750
rect 4470 -820 4540 -750
rect 4700 -820 4770 -750
rect 4930 -820 5000 -750
rect 5160 -820 5230 -750
rect 5390 -820 5460 -750
rect 5620 -820 5690 -750
rect 5850 -820 5920 -750
rect 6080 -820 6150 -750
rect 6310 -820 6380 -750
rect 6540 -820 6610 -750
rect 6770 -820 6840 -750
rect 7000 -820 7070 -750
<< locali >>
rect -2340 1470 8080 1580
rect -2340 1270 -1750 1470
rect -1550 1270 -660 1470
rect -460 1270 340 1470
rect 540 1270 1340 1470
rect 1540 1270 2360 1470
rect 2560 1270 3360 1470
rect 3560 1270 4360 1470
rect 4560 1270 5380 1470
rect 5580 1270 6380 1470
rect 6580 1270 7380 1470
rect 7580 1270 8080 1470
rect -2340 1130 8080 1270
rect -2340 820 -1890 1130
rect -2340 620 -2200 820
rect -2000 620 -1890 820
rect 7630 830 8080 1130
rect 7630 630 7770 830
rect 7970 630 8080 830
rect -2340 -200 -1890 620
rect 310 610 420 630
rect 310 540 330 610
rect 400 540 420 610
rect 310 520 420 540
rect 540 610 650 630
rect 540 540 560 610
rect 630 540 650 610
rect 540 520 650 540
rect 770 610 880 630
rect 770 540 790 610
rect 860 540 880 610
rect 770 520 880 540
rect 1000 610 1110 630
rect 1000 540 1020 610
rect 1090 540 1110 610
rect 1000 520 1110 540
rect 1230 610 1340 630
rect 1230 540 1250 610
rect 1320 540 1340 610
rect 1230 520 1340 540
rect 1460 610 1570 630
rect 1460 540 1480 610
rect 1550 540 1570 610
rect 1460 520 1570 540
rect 1690 610 1800 630
rect 1690 540 1710 610
rect 1780 540 1800 610
rect 1690 520 1800 540
rect 1920 610 2030 630
rect 1920 540 1940 610
rect 2010 540 2030 610
rect 1920 520 2030 540
rect 2150 610 2260 630
rect 2150 540 2170 610
rect 2240 540 2260 610
rect 2150 520 2260 540
rect 2380 610 2490 630
rect 2380 540 2400 610
rect 2470 540 2490 610
rect 2380 520 2490 540
rect 2610 610 2720 630
rect 2610 540 2630 610
rect 2700 540 2720 610
rect 2610 520 2720 540
rect 2840 610 2950 630
rect 2840 540 2860 610
rect 2930 540 2950 610
rect 2840 520 2950 540
rect 3070 610 3180 630
rect 3070 540 3090 610
rect 3160 540 3180 610
rect 3070 520 3180 540
rect 3300 610 3410 630
rect 3300 540 3320 610
rect 3390 540 3410 610
rect 3300 520 3410 540
rect 3530 610 3640 630
rect 3530 540 3550 610
rect 3620 540 3640 610
rect 3530 520 3640 540
rect 3760 610 3870 630
rect 3760 540 3780 610
rect 3850 540 3870 610
rect 3760 520 3870 540
rect 3990 610 4100 630
rect 3990 540 4010 610
rect 4080 540 4100 610
rect 3990 520 4100 540
rect 4220 610 4330 630
rect 4220 540 4240 610
rect 4310 540 4330 610
rect 4220 520 4330 540
rect 4450 610 4560 630
rect 4450 540 4470 610
rect 4540 540 4560 610
rect 4450 520 4560 540
rect 4680 610 4790 630
rect 4680 540 4700 610
rect 4770 540 4790 610
rect 4680 520 4790 540
rect 4910 610 5020 630
rect 4910 540 4930 610
rect 5000 540 5020 610
rect 4910 520 5020 540
rect 5140 610 5250 630
rect 5140 540 5160 610
rect 5230 540 5250 610
rect 5140 520 5250 540
rect 5370 610 5480 630
rect 5370 540 5390 610
rect 5460 540 5480 610
rect 5370 520 5480 540
rect 5600 610 5710 630
rect 5600 540 5620 610
rect 5690 540 5710 610
rect 5600 520 5710 540
rect 5830 610 5940 630
rect 5830 540 5850 610
rect 5920 540 5940 610
rect 5830 520 5940 540
rect 6060 610 6170 630
rect 6060 540 6080 610
rect 6150 540 6170 610
rect 6060 520 6170 540
rect 6290 610 6400 630
rect 6290 540 6310 610
rect 6380 540 6400 610
rect 6290 520 6400 540
rect 6520 610 6630 630
rect 6520 540 6540 610
rect 6610 540 6630 610
rect 6520 520 6630 540
rect 6750 610 6860 630
rect 6750 540 6770 610
rect 6840 540 6860 610
rect 6750 520 6860 540
rect 6980 610 7090 630
rect 6980 540 7000 610
rect 7070 540 7090 610
rect 6980 520 7090 540
rect 180 450 320 470
rect 180 350 200 450
rect 300 350 320 450
rect 180 330 320 350
rect 410 450 550 470
rect 410 350 430 450
rect 530 350 550 450
rect 410 330 550 350
rect 640 450 780 470
rect 640 350 660 450
rect 760 350 780 450
rect 640 330 780 350
rect 870 450 1010 470
rect 870 350 890 450
rect 990 350 1010 450
rect 870 330 1010 350
rect 1100 450 1240 470
rect 1100 350 1120 450
rect 1220 350 1240 450
rect 1100 330 1240 350
rect 1330 450 1470 470
rect 1330 350 1350 450
rect 1450 350 1470 450
rect 1330 330 1470 350
rect 1560 450 1700 470
rect 1560 350 1580 450
rect 1680 350 1700 450
rect 1560 330 1700 350
rect 1790 450 1930 470
rect 1790 350 1810 450
rect 1910 350 1930 450
rect 1790 330 1930 350
rect 2020 450 2160 470
rect 2020 350 2040 450
rect 2140 350 2160 450
rect 2020 330 2160 350
rect 2250 450 2390 470
rect 2250 350 2270 450
rect 2370 350 2390 450
rect 2250 330 2390 350
rect 2480 450 2620 470
rect 2480 350 2500 450
rect 2600 350 2620 450
rect 2480 330 2620 350
rect 2710 450 2850 470
rect 2710 350 2730 450
rect 2830 350 2850 450
rect 2710 330 2850 350
rect 2940 450 3080 470
rect 2940 350 2960 450
rect 3060 350 3080 450
rect 2940 330 3080 350
rect 3170 450 3310 470
rect 3170 350 3190 450
rect 3290 350 3310 450
rect 3170 330 3310 350
rect 3400 450 3540 470
rect 3400 350 3420 450
rect 3520 350 3540 450
rect 3400 330 3540 350
rect 3630 450 3770 470
rect 3630 350 3650 450
rect 3750 350 3770 450
rect 3630 330 3770 350
rect 3860 450 4000 470
rect 3860 350 3880 450
rect 3980 350 4000 450
rect 3860 330 4000 350
rect 4090 450 4230 470
rect 4090 350 4110 450
rect 4210 350 4230 450
rect 4090 330 4230 350
rect 4320 450 4460 470
rect 4320 350 4340 450
rect 4440 350 4460 450
rect 4320 330 4460 350
rect 4550 450 4690 470
rect 4550 350 4570 450
rect 4670 350 4690 450
rect 4550 330 4690 350
rect 4780 450 4920 470
rect 4780 350 4800 450
rect 4900 350 4920 450
rect 4780 330 4920 350
rect 5010 450 5150 470
rect 5010 350 5030 450
rect 5130 350 5150 450
rect 5010 330 5150 350
rect 5240 450 5380 470
rect 5240 350 5260 450
rect 5360 350 5380 450
rect 5240 330 5380 350
rect 5470 450 5610 470
rect 5470 350 5490 450
rect 5590 350 5610 450
rect 5470 330 5610 350
rect 5700 450 5840 470
rect 5700 350 5720 450
rect 5820 350 5840 450
rect 5700 330 5840 350
rect 5930 450 6070 470
rect 5930 350 5950 450
rect 6050 350 6070 450
rect 5930 330 6070 350
rect 6160 450 6300 470
rect 6160 350 6180 450
rect 6280 350 6300 450
rect 6160 330 6300 350
rect 6390 450 6530 470
rect 6390 350 6410 450
rect 6510 350 6530 450
rect 6390 330 6530 350
rect 6620 450 6760 470
rect 6620 350 6640 450
rect 6740 350 6760 450
rect 6620 330 6760 350
rect 6850 450 6990 470
rect 6850 350 6870 450
rect 6970 350 6990 450
rect 6850 330 6990 350
rect 7080 450 7220 470
rect 7080 350 7100 450
rect 7200 350 7220 450
rect 7080 330 7220 350
rect 180 150 320 170
rect 180 50 200 150
rect 300 50 320 150
rect 180 30 320 50
rect 410 150 550 170
rect 410 50 430 150
rect 530 50 550 150
rect 410 30 550 50
rect 640 150 780 170
rect 640 50 660 150
rect 760 50 780 150
rect 640 30 780 50
rect 870 150 1010 170
rect 870 50 890 150
rect 990 50 1010 150
rect 870 30 1010 50
rect 1100 150 1240 170
rect 1100 50 1120 150
rect 1220 50 1240 150
rect 1100 30 1240 50
rect 1330 150 1470 170
rect 1330 50 1350 150
rect 1450 50 1470 150
rect 1330 30 1470 50
rect 1560 150 1700 170
rect 1560 50 1580 150
rect 1680 50 1700 150
rect 1560 30 1700 50
rect 1790 150 1930 170
rect 1790 50 1810 150
rect 1910 50 1930 150
rect 1790 30 1930 50
rect 2020 150 2160 170
rect 2020 50 2040 150
rect 2140 50 2160 150
rect 2020 30 2160 50
rect 2250 150 2390 170
rect 2250 50 2270 150
rect 2370 50 2390 150
rect 2250 30 2390 50
rect 2480 150 2620 170
rect 2480 50 2500 150
rect 2600 50 2620 150
rect 2480 30 2620 50
rect 2710 150 2850 170
rect 2710 50 2730 150
rect 2830 50 2850 150
rect 2710 30 2850 50
rect 2940 150 3080 170
rect 2940 50 2960 150
rect 3060 50 3080 150
rect 2940 30 3080 50
rect 3170 150 3310 170
rect 3170 50 3190 150
rect 3290 50 3310 150
rect 3170 30 3310 50
rect 3400 150 3540 170
rect 3400 50 3420 150
rect 3520 50 3540 150
rect 3400 30 3540 50
rect 3630 150 3770 170
rect 3630 50 3650 150
rect 3750 50 3770 150
rect 3630 30 3770 50
rect 3860 150 4000 170
rect 3860 50 3880 150
rect 3980 50 4000 150
rect 3860 30 4000 50
rect 4090 150 4230 170
rect 4090 50 4110 150
rect 4210 50 4230 150
rect 4090 30 4230 50
rect 4320 150 4460 170
rect 4320 50 4340 150
rect 4440 50 4460 150
rect 4320 30 4460 50
rect 4550 150 4690 170
rect 4550 50 4570 150
rect 4670 50 4690 150
rect 4550 30 4690 50
rect 4780 150 4920 170
rect 4780 50 4800 150
rect 4900 50 4920 150
rect 4780 30 4920 50
rect 5010 150 5150 170
rect 5010 50 5030 150
rect 5130 50 5150 150
rect 5010 30 5150 50
rect 5240 150 5380 170
rect 5240 50 5260 150
rect 5360 50 5380 150
rect 5240 30 5380 50
rect 5470 150 5610 170
rect 5470 50 5490 150
rect 5590 50 5610 150
rect 5470 30 5610 50
rect 5700 150 5840 170
rect 5700 50 5720 150
rect 5820 50 5840 150
rect 5700 30 5840 50
rect 5930 150 6070 170
rect 5930 50 5950 150
rect 6050 50 6070 150
rect 5930 30 6070 50
rect 6160 150 6300 170
rect 6160 50 6180 150
rect 6280 50 6300 150
rect 6160 30 6300 50
rect 6390 150 6530 170
rect 6390 50 6410 150
rect 6510 50 6530 150
rect 6390 30 6530 50
rect 6620 150 6760 170
rect 6620 50 6640 150
rect 6740 50 6760 150
rect 6620 30 6760 50
rect 6850 150 6990 170
rect 6850 50 6870 150
rect 6970 50 6990 150
rect 6850 30 6990 50
rect 7080 150 7220 170
rect 7080 50 7100 150
rect 7200 50 7220 150
rect 7080 30 7220 50
rect -2340 -400 -2200 -200
rect -2000 -400 -1890 -200
rect 7630 -190 8080 630
rect 180 -260 320 -240
rect 180 -360 200 -260
rect 300 -360 320 -260
rect 180 -380 320 -360
rect 410 -260 550 -240
rect 410 -360 430 -260
rect 530 -360 550 -260
rect 410 -380 550 -360
rect 640 -260 780 -240
rect 640 -360 660 -260
rect 760 -360 780 -260
rect 640 -380 780 -360
rect 870 -260 1010 -240
rect 870 -360 890 -260
rect 990 -360 1010 -260
rect 870 -380 1010 -360
rect 1100 -260 1240 -240
rect 1100 -360 1120 -260
rect 1220 -360 1240 -260
rect 1100 -380 1240 -360
rect 1330 -260 1470 -240
rect 1330 -360 1350 -260
rect 1450 -360 1470 -260
rect 1330 -380 1470 -360
rect 1560 -260 1700 -240
rect 1560 -360 1580 -260
rect 1680 -360 1700 -260
rect 1560 -380 1700 -360
rect 1790 -260 1930 -240
rect 1790 -360 1810 -260
rect 1910 -360 1930 -260
rect 1790 -380 1930 -360
rect 2020 -260 2160 -240
rect 2020 -360 2040 -260
rect 2140 -360 2160 -260
rect 2020 -380 2160 -360
rect 2250 -260 2390 -240
rect 2250 -360 2270 -260
rect 2370 -360 2390 -260
rect 2250 -380 2390 -360
rect 2480 -260 2620 -240
rect 2480 -360 2500 -260
rect 2600 -360 2620 -260
rect 2480 -380 2620 -360
rect 2710 -260 2850 -240
rect 2710 -360 2730 -260
rect 2830 -360 2850 -260
rect 2710 -380 2850 -360
rect 2940 -260 3080 -240
rect 2940 -360 2960 -260
rect 3060 -360 3080 -260
rect 2940 -380 3080 -360
rect 3170 -260 3310 -240
rect 3170 -360 3190 -260
rect 3290 -360 3310 -260
rect 3170 -380 3310 -360
rect 3400 -260 3540 -240
rect 3400 -360 3420 -260
rect 3520 -360 3540 -260
rect 3400 -380 3540 -360
rect 3630 -260 3770 -240
rect 3630 -360 3650 -260
rect 3750 -360 3770 -260
rect 3630 -380 3770 -360
rect 3860 -260 4000 -240
rect 3860 -360 3880 -260
rect 3980 -360 4000 -260
rect 3860 -380 4000 -360
rect 4090 -260 4230 -240
rect 4090 -360 4110 -260
rect 4210 -360 4230 -260
rect 4090 -380 4230 -360
rect 4320 -260 4460 -240
rect 4320 -360 4340 -260
rect 4440 -360 4460 -260
rect 4320 -380 4460 -360
rect 4550 -260 4690 -240
rect 4550 -360 4570 -260
rect 4670 -360 4690 -260
rect 4550 -380 4690 -360
rect 4780 -260 4920 -240
rect 4780 -360 4800 -260
rect 4900 -360 4920 -260
rect 4780 -380 4920 -360
rect 5010 -260 5150 -240
rect 5010 -360 5030 -260
rect 5130 -360 5150 -260
rect 5010 -380 5150 -360
rect 5240 -260 5380 -240
rect 5240 -360 5260 -260
rect 5360 -360 5380 -260
rect 5240 -380 5380 -360
rect 5470 -260 5610 -240
rect 5470 -360 5490 -260
rect 5590 -360 5610 -260
rect 5470 -380 5610 -360
rect 5700 -260 5840 -240
rect 5700 -360 5720 -260
rect 5820 -360 5840 -260
rect 5700 -380 5840 -360
rect 5930 -260 6070 -240
rect 5930 -360 5950 -260
rect 6050 -360 6070 -260
rect 5930 -380 6070 -360
rect 6160 -260 6300 -240
rect 6160 -360 6180 -260
rect 6280 -360 6300 -260
rect 6160 -380 6300 -360
rect 6390 -260 6530 -240
rect 6390 -360 6410 -260
rect 6510 -360 6530 -260
rect 6390 -380 6530 -360
rect 6620 -260 6760 -240
rect 6620 -360 6640 -260
rect 6740 -360 6760 -260
rect 6620 -380 6760 -360
rect 6850 -260 6990 -240
rect 6850 -360 6870 -260
rect 6970 -360 6990 -260
rect 6850 -380 6990 -360
rect 7080 -260 7220 -240
rect 7080 -360 7100 -260
rect 7200 -360 7220 -260
rect 7080 -380 7220 -360
rect -2340 -1200 -1890 -400
rect 7630 -390 7770 -190
rect 7970 -390 8080 -190
rect 180 -560 320 -540
rect 180 -660 200 -560
rect 300 -660 320 -560
rect 180 -680 320 -660
rect 410 -560 550 -540
rect 410 -660 430 -560
rect 530 -660 550 -560
rect 410 -680 550 -660
rect 640 -560 780 -540
rect 640 -660 660 -560
rect 760 -660 780 -560
rect 640 -680 780 -660
rect 870 -560 1010 -540
rect 870 -660 890 -560
rect 990 -660 1010 -560
rect 870 -680 1010 -660
rect 1100 -560 1240 -540
rect 1100 -660 1120 -560
rect 1220 -660 1240 -560
rect 1100 -680 1240 -660
rect 1330 -560 1470 -540
rect 1330 -660 1350 -560
rect 1450 -660 1470 -560
rect 1330 -680 1470 -660
rect 1560 -560 1700 -540
rect 1560 -660 1580 -560
rect 1680 -660 1700 -560
rect 1560 -680 1700 -660
rect 1790 -560 1930 -540
rect 1790 -660 1810 -560
rect 1910 -660 1930 -560
rect 1790 -680 1930 -660
rect 2020 -560 2160 -540
rect 2020 -660 2040 -560
rect 2140 -660 2160 -560
rect 2020 -680 2160 -660
rect 2250 -560 2390 -540
rect 2250 -660 2270 -560
rect 2370 -660 2390 -560
rect 2250 -680 2390 -660
rect 2480 -560 2620 -540
rect 2480 -660 2500 -560
rect 2600 -660 2620 -560
rect 2480 -680 2620 -660
rect 2710 -560 2850 -540
rect 2710 -660 2730 -560
rect 2830 -660 2850 -560
rect 2710 -680 2850 -660
rect 2940 -560 3080 -540
rect 2940 -660 2960 -560
rect 3060 -660 3080 -560
rect 2940 -680 3080 -660
rect 3170 -560 3310 -540
rect 3170 -660 3190 -560
rect 3290 -660 3310 -560
rect 3170 -680 3310 -660
rect 3400 -560 3540 -540
rect 3400 -660 3420 -560
rect 3520 -660 3540 -560
rect 3400 -680 3540 -660
rect 3630 -560 3770 -540
rect 3630 -660 3650 -560
rect 3750 -660 3770 -560
rect 3630 -680 3770 -660
rect 3860 -560 4000 -540
rect 3860 -660 3880 -560
rect 3980 -660 4000 -560
rect 3860 -680 4000 -660
rect 4090 -560 4230 -540
rect 4090 -660 4110 -560
rect 4210 -660 4230 -560
rect 4090 -680 4230 -660
rect 4320 -560 4460 -540
rect 4320 -660 4340 -560
rect 4440 -660 4460 -560
rect 4320 -680 4460 -660
rect 4550 -560 4690 -540
rect 4550 -660 4570 -560
rect 4670 -660 4690 -560
rect 4550 -680 4690 -660
rect 4780 -560 4920 -540
rect 4780 -660 4800 -560
rect 4900 -660 4920 -560
rect 4780 -680 4920 -660
rect 5010 -560 5150 -540
rect 5010 -660 5030 -560
rect 5130 -660 5150 -560
rect 5010 -680 5150 -660
rect 5240 -560 5380 -540
rect 5240 -660 5260 -560
rect 5360 -660 5380 -560
rect 5240 -680 5380 -660
rect 5470 -560 5610 -540
rect 5470 -660 5490 -560
rect 5590 -660 5610 -560
rect 5470 -680 5610 -660
rect 5700 -560 5840 -540
rect 5700 -660 5720 -560
rect 5820 -660 5840 -560
rect 5700 -680 5840 -660
rect 5930 -560 6070 -540
rect 5930 -660 5950 -560
rect 6050 -660 6070 -560
rect 5930 -680 6070 -660
rect 6160 -560 6300 -540
rect 6160 -660 6180 -560
rect 6280 -660 6300 -560
rect 6160 -680 6300 -660
rect 6390 -560 6530 -540
rect 6390 -660 6410 -560
rect 6510 -660 6530 -560
rect 6390 -680 6530 -660
rect 6620 -560 6760 -540
rect 6620 -660 6640 -560
rect 6740 -660 6760 -560
rect 6620 -680 6760 -660
rect 6850 -560 6990 -540
rect 6850 -660 6870 -560
rect 6970 -660 6990 -560
rect 6850 -680 6990 -660
rect 7080 -560 7220 -540
rect 7080 -660 7100 -560
rect 7200 -660 7220 -560
rect 7080 -680 7220 -660
rect 310 -750 420 -730
rect 310 -820 330 -750
rect 400 -820 420 -750
rect 310 -840 420 -820
rect 540 -750 650 -730
rect 540 -820 560 -750
rect 630 -820 650 -750
rect 540 -840 650 -820
rect 770 -750 880 -730
rect 770 -820 790 -750
rect 860 -820 880 -750
rect 770 -840 880 -820
rect 1000 -750 1110 -730
rect 1000 -820 1020 -750
rect 1090 -820 1110 -750
rect 1000 -840 1110 -820
rect 1230 -750 1340 -730
rect 1230 -820 1250 -750
rect 1320 -820 1340 -750
rect 1230 -840 1340 -820
rect 1460 -750 1570 -730
rect 1460 -820 1480 -750
rect 1550 -820 1570 -750
rect 1460 -840 1570 -820
rect 1690 -750 1800 -730
rect 1690 -820 1710 -750
rect 1780 -820 1800 -750
rect 1690 -840 1800 -820
rect 1920 -750 2030 -730
rect 1920 -820 1940 -750
rect 2010 -820 2030 -750
rect 1920 -840 2030 -820
rect 2150 -750 2260 -730
rect 2150 -820 2170 -750
rect 2240 -820 2260 -750
rect 2150 -840 2260 -820
rect 2380 -750 2490 -730
rect 2380 -820 2400 -750
rect 2470 -820 2490 -750
rect 2380 -840 2490 -820
rect 2610 -750 2720 -730
rect 2610 -820 2630 -750
rect 2700 -820 2720 -750
rect 2610 -840 2720 -820
rect 2840 -750 2950 -730
rect 2840 -820 2860 -750
rect 2930 -820 2950 -750
rect 2840 -840 2950 -820
rect 3070 -750 3180 -730
rect 3070 -820 3090 -750
rect 3160 -820 3180 -750
rect 3070 -840 3180 -820
rect 3300 -750 3410 -730
rect 3300 -820 3320 -750
rect 3390 -820 3410 -750
rect 3300 -840 3410 -820
rect 3530 -750 3640 -730
rect 3530 -820 3550 -750
rect 3620 -820 3640 -750
rect 3530 -840 3640 -820
rect 3760 -750 3870 -730
rect 3760 -820 3780 -750
rect 3850 -820 3870 -750
rect 3760 -840 3870 -820
rect 3990 -750 4100 -730
rect 3990 -820 4010 -750
rect 4080 -820 4100 -750
rect 3990 -840 4100 -820
rect 4220 -750 4330 -730
rect 4220 -820 4240 -750
rect 4310 -820 4330 -750
rect 4220 -840 4330 -820
rect 4450 -750 4560 -730
rect 4450 -820 4470 -750
rect 4540 -820 4560 -750
rect 4450 -840 4560 -820
rect 4680 -750 4790 -730
rect 4680 -820 4700 -750
rect 4770 -820 4790 -750
rect 4680 -840 4790 -820
rect 4910 -750 5020 -730
rect 4910 -820 4930 -750
rect 5000 -820 5020 -750
rect 4910 -840 5020 -820
rect 5140 -750 5250 -730
rect 5140 -820 5160 -750
rect 5230 -820 5250 -750
rect 5140 -840 5250 -820
rect 5370 -750 5480 -730
rect 5370 -820 5390 -750
rect 5460 -820 5480 -750
rect 5370 -840 5480 -820
rect 5600 -750 5710 -730
rect 5600 -820 5620 -750
rect 5690 -820 5710 -750
rect 5600 -840 5710 -820
rect 5830 -750 5940 -730
rect 5830 -820 5850 -750
rect 5920 -820 5940 -750
rect 5830 -840 5940 -820
rect 6060 -750 6170 -730
rect 6060 -820 6080 -750
rect 6150 -820 6170 -750
rect 6060 -840 6170 -820
rect 6290 -750 6400 -730
rect 6290 -820 6310 -750
rect 6380 -820 6400 -750
rect 6290 -840 6400 -820
rect 6520 -750 6630 -730
rect 6520 -820 6540 -750
rect 6610 -820 6630 -750
rect 6520 -840 6630 -820
rect 6750 -750 6860 -730
rect 6750 -820 6770 -750
rect 6840 -820 6860 -750
rect 6750 -840 6860 -820
rect 6980 -750 7090 -730
rect 6980 -820 7000 -750
rect 7070 -820 7090 -750
rect 6980 -840 7090 -820
rect -2340 -1400 -2200 -1200
rect -2000 -1360 -1890 -1200
rect 7630 -1190 8080 -390
rect 7630 -1360 7770 -1190
rect -2000 -1390 7770 -1360
rect 7970 -1390 8080 -1190
rect -2000 -1400 8080 -1390
rect -2340 -1470 8080 -1400
rect -2340 -1670 -1780 -1470
rect -1580 -1670 -690 -1470
rect -490 -1670 310 -1470
rect 510 -1670 1310 -1470
rect 1510 -1670 2330 -1470
rect 2530 -1670 3330 -1470
rect 3530 -1670 4330 -1470
rect 4530 -1670 5350 -1470
rect 5550 -1670 6350 -1470
rect 6550 -1670 7350 -1470
rect 7550 -1670 8080 -1470
rect -2340 -1810 8080 -1670
<< viali >>
rect 330 540 400 610
rect 560 540 630 610
rect 790 540 860 610
rect 1020 540 1090 610
rect 1250 540 1320 610
rect 1480 540 1550 610
rect 1710 540 1780 610
rect 1940 540 2010 610
rect 2170 540 2240 610
rect 2400 540 2470 610
rect 2630 540 2700 610
rect 2860 540 2930 610
rect 3090 540 3160 610
rect 3320 540 3390 610
rect 3550 540 3620 610
rect 3780 540 3850 610
rect 4010 540 4080 610
rect 4240 540 4310 610
rect 4470 540 4540 610
rect 4700 540 4770 610
rect 4930 540 5000 610
rect 5160 540 5230 610
rect 5390 540 5460 610
rect 5620 540 5690 610
rect 5850 540 5920 610
rect 6080 540 6150 610
rect 6310 540 6380 610
rect 6540 540 6610 610
rect 6770 540 6840 610
rect 7000 540 7070 610
rect 200 350 300 450
rect 660 350 760 450
rect 1120 350 1220 450
rect 1580 350 1680 450
rect 2040 350 2140 450
rect 2500 350 2600 450
rect 2960 350 3060 450
rect 3420 350 3520 450
rect 3880 350 3980 450
rect 4340 350 4440 450
rect 4800 350 4900 450
rect 5260 350 5360 450
rect 5720 350 5820 450
rect 6180 350 6280 450
rect 6640 350 6740 450
rect 7100 350 7200 450
rect 430 50 530 150
rect 890 50 990 150
rect 1350 50 1450 150
rect 1810 50 1910 150
rect 2270 50 2370 150
rect 2730 50 2830 150
rect 3190 50 3290 150
rect 3650 50 3750 150
rect 4110 50 4210 150
rect 4570 50 4670 150
rect 5030 50 5130 150
rect 5490 50 5590 150
rect 5950 50 6050 150
rect 6410 50 6510 150
rect 6870 50 6970 150
rect 430 -360 530 -260
rect 890 -360 990 -260
rect 1350 -360 1450 -260
rect 1810 -360 1910 -260
rect 2270 -360 2370 -260
rect 2730 -360 2830 -260
rect 3190 -360 3290 -260
rect 3650 -360 3750 -260
rect 4110 -360 4210 -260
rect 4570 -360 4670 -260
rect 5030 -360 5130 -260
rect 5490 -360 5590 -260
rect 5950 -360 6050 -260
rect 6410 -360 6510 -260
rect 6870 -360 6970 -260
rect 200 -660 300 -560
rect 660 -660 760 -560
rect 1120 -660 1220 -560
rect 1580 -660 1680 -560
rect 2040 -660 2140 -560
rect 2500 -660 2600 -560
rect 2960 -660 3060 -560
rect 3420 -660 3520 -560
rect 3880 -660 3980 -560
rect 4340 -660 4440 -560
rect 4800 -660 4900 -560
rect 5260 -660 5360 -560
rect 5720 -660 5820 -560
rect 6180 -660 6280 -560
rect 6640 -660 6740 -560
rect 7100 -660 7200 -560
rect 330 -820 400 -750
rect 560 -820 630 -750
rect 790 -820 860 -750
rect 1020 -820 1090 -750
rect 1250 -820 1320 -750
rect 1480 -820 1550 -750
rect 1710 -820 1780 -750
rect 1940 -820 2010 -750
rect 2170 -820 2240 -750
rect 2400 -820 2470 -750
rect 2630 -820 2700 -750
rect 2860 -820 2930 -750
rect 3090 -820 3160 -750
rect 3320 -820 3390 -750
rect 3550 -820 3620 -750
rect 3780 -820 3850 -750
rect 4010 -820 4080 -750
rect 4240 -820 4310 -750
rect 4470 -820 4540 -750
rect 4700 -820 4770 -750
rect 4930 -820 5000 -750
rect 5160 -820 5230 -750
rect 5390 -820 5460 -750
rect 5620 -820 5690 -750
rect 5850 -820 5920 -750
rect 6080 -820 6150 -750
rect 6310 -820 6380 -750
rect 6540 -820 6610 -750
rect 6770 -820 6840 -750
rect 7000 -820 7070 -750
<< metal1 >>
rect 310 610 420 630
rect 310 540 330 610
rect 400 540 420 610
rect 310 520 420 540
rect 540 610 650 630
rect 540 540 560 610
rect 630 540 650 610
rect 540 520 650 540
rect 770 610 880 630
rect 770 540 790 610
rect 860 540 880 610
rect 770 520 880 540
rect 1000 610 1110 630
rect 1000 540 1020 610
rect 1090 540 1110 610
rect 1000 520 1110 540
rect 1230 610 1340 630
rect 1230 540 1250 610
rect 1320 540 1340 610
rect 1230 520 1340 540
rect 1460 610 1570 630
rect 1460 540 1480 610
rect 1550 540 1570 610
rect 1460 520 1570 540
rect 1690 610 1800 630
rect 1690 540 1710 610
rect 1780 540 1800 610
rect 1690 520 1800 540
rect 1920 610 2030 630
rect 1920 540 1940 610
rect 2010 540 2030 610
rect 1920 520 2030 540
rect 2150 610 2260 630
rect 2150 540 2170 610
rect 2240 540 2260 610
rect 2150 520 2260 540
rect 2380 610 2490 630
rect 2380 540 2400 610
rect 2470 540 2490 610
rect 2380 520 2490 540
rect 2610 610 2720 630
rect 2610 540 2630 610
rect 2700 540 2720 610
rect 2610 520 2720 540
rect 2840 610 2950 630
rect 2840 540 2860 610
rect 2930 540 2950 610
rect 2840 520 2950 540
rect 3070 610 3180 630
rect 3070 540 3090 610
rect 3160 540 3180 610
rect 3070 520 3180 540
rect 3300 610 3410 630
rect 3300 540 3320 610
rect 3390 540 3410 610
rect 3300 520 3410 540
rect 3530 610 3640 630
rect 3530 540 3550 610
rect 3620 540 3640 610
rect 3530 520 3640 540
rect 3760 610 3870 630
rect 3760 540 3780 610
rect 3850 540 3870 610
rect 3760 520 3870 540
rect 3990 610 4100 630
rect 3990 540 4010 610
rect 4080 540 4100 610
rect 3990 520 4100 540
rect 4220 610 4330 630
rect 4220 540 4240 610
rect 4310 540 4330 610
rect 4220 520 4330 540
rect 4450 610 4560 630
rect 4450 540 4470 610
rect 4540 540 4560 610
rect 4450 520 4560 540
rect 4680 610 4790 630
rect 4680 540 4700 610
rect 4770 540 4790 610
rect 4680 520 4790 540
rect 4910 610 5020 630
rect 4910 540 4930 610
rect 5000 540 5020 610
rect 4910 520 5020 540
rect 5140 610 5250 630
rect 5140 540 5160 610
rect 5230 540 5250 610
rect 5140 520 5250 540
rect 5370 610 5480 630
rect 5370 540 5390 610
rect 5460 540 5480 610
rect 5370 520 5480 540
rect 5600 610 5710 630
rect 5600 540 5620 610
rect 5690 540 5710 610
rect 5600 520 5710 540
rect 5830 610 5940 630
rect 5830 540 5850 610
rect 5920 540 5940 610
rect 5830 520 5940 540
rect 6060 610 6170 630
rect 6060 540 6080 610
rect 6150 540 6170 610
rect 6060 520 6170 540
rect 6290 610 6400 630
rect 6290 540 6310 610
rect 6380 540 6400 610
rect 6290 520 6400 540
rect 6520 610 6630 630
rect 6520 540 6540 610
rect 6610 540 6630 610
rect 6520 520 6630 540
rect 6750 610 6860 630
rect 6750 540 6770 610
rect 6840 540 6860 610
rect 6750 520 6860 540
rect 6980 610 7090 630
rect 6980 540 7000 610
rect 7070 540 7090 610
rect 6980 520 7090 540
rect 180 450 320 470
rect 180 350 200 450
rect 300 350 320 450
rect 180 330 320 350
rect 640 450 780 470
rect 640 350 660 450
rect 760 350 780 450
rect 640 330 780 350
rect 1100 450 1240 470
rect 1100 350 1120 450
rect 1220 350 1240 450
rect 1100 330 1240 350
rect 1560 450 1700 470
rect 1560 350 1580 450
rect 1680 350 1700 450
rect 1560 330 1700 350
rect 2020 450 2160 470
rect 2020 350 2040 450
rect 2140 350 2160 450
rect 2020 330 2160 350
rect 2480 450 2620 470
rect 2480 350 2500 450
rect 2600 350 2620 450
rect 2480 330 2620 350
rect 2940 450 3080 470
rect 2940 350 2960 450
rect 3060 350 3080 450
rect 2940 330 3080 350
rect 3400 450 3540 470
rect 3400 350 3420 450
rect 3520 350 3540 450
rect 3400 330 3540 350
rect 3860 450 4000 470
rect 3860 350 3880 450
rect 3980 350 4000 450
rect 3860 330 4000 350
rect 4320 450 4460 470
rect 4320 350 4340 450
rect 4440 350 4460 450
rect 4320 330 4460 350
rect 4780 450 4920 470
rect 4780 350 4800 450
rect 4900 350 4920 450
rect 4780 330 4920 350
rect 5240 450 5380 470
rect 5240 350 5260 450
rect 5360 350 5380 450
rect 5240 330 5380 350
rect 5700 450 5840 470
rect 5700 350 5720 450
rect 5820 350 5840 450
rect 5700 330 5840 350
rect 6160 450 6300 470
rect 6160 350 6180 450
rect 6280 350 6300 450
rect 6160 330 6300 350
rect 6620 450 6760 470
rect 6620 350 6640 450
rect 6740 350 6760 450
rect 6620 330 6760 350
rect 7080 450 7220 470
rect 7080 350 7100 450
rect 7200 350 7220 450
rect 7080 330 7220 350
rect 410 150 550 170
rect 410 50 430 150
rect 530 50 550 150
rect 410 30 550 50
rect 870 150 1010 170
rect 870 50 890 150
rect 990 50 1010 150
rect 870 30 1010 50
rect 1330 150 1470 170
rect 1330 50 1350 150
rect 1450 50 1470 150
rect 1330 30 1470 50
rect 1790 150 1930 170
rect 1790 50 1810 150
rect 1910 50 1930 150
rect 1790 30 1930 50
rect 2250 150 2390 170
rect 2250 50 2270 150
rect 2370 50 2390 150
rect 2250 30 2390 50
rect 2710 150 2850 170
rect 2710 50 2730 150
rect 2830 50 2850 150
rect 2710 30 2850 50
rect 3170 150 3310 170
rect 3170 50 3190 150
rect 3290 50 3310 150
rect 3170 30 3310 50
rect 3630 150 3770 170
rect 3630 50 3650 150
rect 3750 50 3770 150
rect 3630 30 3770 50
rect 4090 150 4230 170
rect 4090 50 4110 150
rect 4210 50 4230 150
rect 4090 30 4230 50
rect 4550 150 4690 170
rect 4550 50 4570 150
rect 4670 50 4690 150
rect 4550 30 4690 50
rect 5010 150 5150 170
rect 5010 50 5030 150
rect 5130 50 5150 150
rect 5010 30 5150 50
rect 5470 150 5610 170
rect 5470 50 5490 150
rect 5590 50 5610 150
rect 5470 30 5610 50
rect 5930 150 6070 170
rect 5930 50 5950 150
rect 6050 50 6070 150
rect 5930 30 6070 50
rect 6390 150 6530 170
rect 6390 50 6410 150
rect 6510 50 6530 150
rect 6390 30 6530 50
rect 6850 150 6990 170
rect 6850 50 6870 150
rect 6970 50 6990 150
rect 6850 30 6990 50
rect 410 -260 550 -240
rect 410 -360 430 -260
rect 530 -360 550 -260
rect 410 -380 550 -360
rect 870 -260 1010 -240
rect 870 -360 890 -260
rect 990 -360 1010 -260
rect 870 -380 1010 -360
rect 1330 -260 1470 -240
rect 1330 -360 1350 -260
rect 1450 -360 1470 -260
rect 1330 -380 1470 -360
rect 1790 -260 1930 -240
rect 1790 -360 1810 -260
rect 1910 -360 1930 -260
rect 1790 -380 1930 -360
rect 2250 -260 2390 -240
rect 2250 -360 2270 -260
rect 2370 -360 2390 -260
rect 2250 -380 2390 -360
rect 2710 -260 2850 -240
rect 2710 -360 2730 -260
rect 2830 -360 2850 -260
rect 2710 -380 2850 -360
rect 3170 -260 3310 -240
rect 3170 -360 3190 -260
rect 3290 -360 3310 -260
rect 3170 -380 3310 -360
rect 3630 -260 3770 -240
rect 3630 -360 3650 -260
rect 3750 -360 3770 -260
rect 3630 -380 3770 -360
rect 4090 -260 4230 -240
rect 4090 -360 4110 -260
rect 4210 -360 4230 -260
rect 4090 -380 4230 -360
rect 4550 -260 4690 -240
rect 4550 -360 4570 -260
rect 4670 -360 4690 -260
rect 4550 -380 4690 -360
rect 5010 -260 5150 -240
rect 5010 -360 5030 -260
rect 5130 -360 5150 -260
rect 5010 -380 5150 -360
rect 5470 -260 5610 -240
rect 5470 -360 5490 -260
rect 5590 -360 5610 -260
rect 5470 -380 5610 -360
rect 5930 -260 6070 -240
rect 5930 -360 5950 -260
rect 6050 -360 6070 -260
rect 5930 -380 6070 -360
rect 6390 -260 6530 -240
rect 6390 -360 6410 -260
rect 6510 -360 6530 -260
rect 6390 -380 6530 -360
rect 6850 -260 6990 -240
rect 6850 -360 6870 -260
rect 6970 -360 6990 -260
rect 6850 -380 6990 -360
rect 180 -560 320 -540
rect 180 -660 200 -560
rect 300 -660 320 -560
rect 180 -680 320 -660
rect 640 -560 780 -540
rect 640 -660 660 -560
rect 760 -660 780 -560
rect 640 -680 780 -660
rect 1100 -560 1240 -540
rect 1100 -660 1120 -560
rect 1220 -660 1240 -560
rect 1100 -680 1240 -660
rect 1560 -560 1700 -540
rect 1560 -660 1580 -560
rect 1680 -660 1700 -560
rect 1560 -680 1700 -660
rect 2020 -560 2160 -540
rect 2020 -660 2040 -560
rect 2140 -660 2160 -560
rect 2020 -680 2160 -660
rect 2480 -560 2620 -540
rect 2480 -660 2500 -560
rect 2600 -660 2620 -560
rect 2480 -680 2620 -660
rect 2940 -560 3080 -540
rect 2940 -660 2960 -560
rect 3060 -660 3080 -560
rect 2940 -680 3080 -660
rect 3400 -560 3540 -540
rect 3400 -660 3420 -560
rect 3520 -660 3540 -560
rect 3400 -680 3540 -660
rect 3860 -560 4000 -540
rect 3860 -660 3880 -560
rect 3980 -660 4000 -560
rect 3860 -680 4000 -660
rect 4320 -560 4460 -540
rect 4320 -660 4340 -560
rect 4440 -660 4460 -560
rect 4320 -680 4460 -660
rect 4780 -560 4920 -540
rect 4780 -660 4800 -560
rect 4900 -660 4920 -560
rect 4780 -680 4920 -660
rect 5240 -560 5380 -540
rect 5240 -660 5260 -560
rect 5360 -660 5380 -560
rect 5240 -680 5380 -660
rect 5700 -560 5840 -540
rect 5700 -660 5720 -560
rect 5820 -660 5840 -560
rect 5700 -680 5840 -660
rect 6160 -560 6300 -540
rect 6160 -660 6180 -560
rect 6280 -660 6300 -560
rect 6160 -680 6300 -660
rect 6620 -560 6760 -540
rect 6620 -660 6640 -560
rect 6740 -660 6760 -560
rect 6620 -680 6760 -660
rect 7080 -560 7220 -540
rect 7080 -660 7100 -560
rect 7200 -660 7220 -560
rect 7080 -680 7220 -660
rect 310 -750 420 -730
rect 310 -820 330 -750
rect 400 -820 420 -750
rect 310 -840 420 -820
rect 540 -750 650 -730
rect 540 -820 560 -750
rect 630 -820 650 -750
rect 540 -840 650 -820
rect 770 -750 880 -730
rect 770 -820 790 -750
rect 860 -820 880 -750
rect 770 -840 880 -820
rect 1000 -750 1110 -730
rect 1000 -820 1020 -750
rect 1090 -820 1110 -750
rect 1000 -840 1110 -820
rect 1230 -750 1340 -730
rect 1230 -820 1250 -750
rect 1320 -820 1340 -750
rect 1230 -840 1340 -820
rect 1460 -750 1570 -730
rect 1460 -820 1480 -750
rect 1550 -820 1570 -750
rect 1460 -840 1570 -820
rect 1690 -750 1800 -730
rect 1690 -820 1710 -750
rect 1780 -820 1800 -750
rect 1690 -840 1800 -820
rect 1920 -750 2030 -730
rect 1920 -820 1940 -750
rect 2010 -820 2030 -750
rect 1920 -840 2030 -820
rect 2150 -750 2260 -730
rect 2150 -820 2170 -750
rect 2240 -820 2260 -750
rect 2150 -840 2260 -820
rect 2380 -750 2490 -730
rect 2380 -820 2400 -750
rect 2470 -820 2490 -750
rect 2380 -840 2490 -820
rect 2610 -750 2720 -730
rect 2610 -820 2630 -750
rect 2700 -820 2720 -750
rect 2610 -840 2720 -820
rect 2840 -750 2950 -730
rect 2840 -820 2860 -750
rect 2930 -820 2950 -750
rect 2840 -840 2950 -820
rect 3070 -750 3180 -730
rect 3070 -820 3090 -750
rect 3160 -820 3180 -750
rect 3070 -840 3180 -820
rect 3300 -750 3410 -730
rect 3300 -820 3320 -750
rect 3390 -820 3410 -750
rect 3300 -840 3410 -820
rect 3530 -750 3640 -730
rect 3530 -820 3550 -750
rect 3620 -820 3640 -750
rect 3530 -840 3640 -820
rect 3760 -750 3870 -730
rect 3760 -820 3780 -750
rect 3850 -820 3870 -750
rect 3760 -840 3870 -820
rect 3990 -750 4100 -730
rect 3990 -820 4010 -750
rect 4080 -820 4100 -750
rect 3990 -840 4100 -820
rect 4220 -750 4330 -730
rect 4220 -820 4240 -750
rect 4310 -820 4330 -750
rect 4220 -840 4330 -820
rect 4450 -750 4560 -730
rect 4450 -820 4470 -750
rect 4540 -820 4560 -750
rect 4450 -840 4560 -820
rect 4680 -750 4790 -730
rect 4680 -820 4700 -750
rect 4770 -820 4790 -750
rect 4680 -840 4790 -820
rect 4910 -750 5020 -730
rect 4910 -820 4930 -750
rect 5000 -820 5020 -750
rect 4910 -840 5020 -820
rect 5140 -750 5250 -730
rect 5140 -820 5160 -750
rect 5230 -820 5250 -750
rect 5140 -840 5250 -820
rect 5370 -750 5480 -730
rect 5370 -820 5390 -750
rect 5460 -820 5480 -750
rect 5370 -840 5480 -820
rect 5600 -750 5710 -730
rect 5600 -820 5620 -750
rect 5690 -820 5710 -750
rect 5600 -840 5710 -820
rect 5830 -750 5940 -730
rect 5830 -820 5850 -750
rect 5920 -820 5940 -750
rect 5830 -840 5940 -820
rect 6060 -750 6170 -730
rect 6060 -820 6080 -750
rect 6150 -820 6170 -750
rect 6060 -840 6170 -820
rect 6290 -750 6400 -730
rect 6290 -820 6310 -750
rect 6380 -820 6400 -750
rect 6290 -840 6400 -820
rect 6520 -750 6630 -730
rect 6520 -820 6540 -750
rect 6610 -820 6630 -750
rect 6520 -840 6630 -820
rect 6750 -750 6860 -730
rect 6750 -820 6770 -750
rect 6840 -820 6860 -750
rect 6750 -840 6860 -820
rect 6980 -750 7090 -730
rect 6980 -820 7000 -750
rect 7070 -820 7090 -750
rect 6980 -840 7090 -820
<< via1 >>
rect 330 540 400 610
rect 560 540 630 610
rect 790 540 860 610
rect 1020 540 1090 610
rect 1250 540 1320 610
rect 1480 540 1550 610
rect 1710 540 1780 610
rect 1940 540 2010 610
rect 2170 540 2240 610
rect 2400 540 2470 610
rect 2630 540 2700 610
rect 2860 540 2930 610
rect 3090 540 3160 610
rect 3320 540 3390 610
rect 3550 540 3620 610
rect 3780 540 3850 610
rect 4010 540 4080 610
rect 4240 540 4310 610
rect 4470 540 4540 610
rect 4700 540 4770 610
rect 4930 540 5000 610
rect 5160 540 5230 610
rect 5390 540 5460 610
rect 5620 540 5690 610
rect 5850 540 5920 610
rect 6080 540 6150 610
rect 6310 540 6380 610
rect 6540 540 6610 610
rect 6770 540 6840 610
rect 7000 540 7070 610
rect 200 350 300 450
rect 660 350 760 450
rect 1120 350 1220 450
rect 1580 350 1680 450
rect 2040 350 2140 450
rect 2500 350 2600 450
rect 2960 350 3060 450
rect 3420 350 3520 450
rect 3880 350 3980 450
rect 4340 350 4440 450
rect 4800 350 4900 450
rect 5260 350 5360 450
rect 5720 350 5820 450
rect 6180 350 6280 450
rect 6640 350 6740 450
rect 7100 350 7200 450
rect 430 50 530 150
rect 890 50 990 150
rect 1350 50 1450 150
rect 1810 50 1910 150
rect 2270 50 2370 150
rect 2730 50 2830 150
rect 3190 50 3290 150
rect 3650 50 3750 150
rect 4110 50 4210 150
rect 4570 50 4670 150
rect 5030 50 5130 150
rect 5490 50 5590 150
rect 5950 50 6050 150
rect 6410 50 6510 150
rect 6870 50 6970 150
rect 430 -360 530 -260
rect 890 -360 990 -260
rect 1350 -360 1450 -260
rect 1810 -360 1910 -260
rect 2270 -360 2370 -260
rect 2730 -360 2830 -260
rect 3190 -360 3290 -260
rect 3650 -360 3750 -260
rect 4110 -360 4210 -260
rect 4570 -360 4670 -260
rect 5030 -360 5130 -260
rect 5490 -360 5590 -260
rect 5950 -360 6050 -260
rect 6410 -360 6510 -260
rect 6870 -360 6970 -260
rect 200 -660 300 -560
rect 660 -660 760 -560
rect 1120 -660 1220 -560
rect 1580 -660 1680 -560
rect 2040 -660 2140 -560
rect 2500 -660 2600 -560
rect 2960 -660 3060 -560
rect 3420 -660 3520 -560
rect 3880 -660 3980 -560
rect 4340 -660 4440 -560
rect 4800 -660 4900 -560
rect 5260 -660 5360 -560
rect 5720 -660 5820 -560
rect 6180 -660 6280 -560
rect 6640 -660 6740 -560
rect 7100 -660 7200 -560
rect 330 -820 400 -750
rect 560 -820 630 -750
rect 790 -820 860 -750
rect 1020 -820 1090 -750
rect 1250 -820 1320 -750
rect 1480 -820 1550 -750
rect 1710 -820 1780 -750
rect 1940 -820 2010 -750
rect 2170 -820 2240 -750
rect 2400 -820 2470 -750
rect 2630 -820 2700 -750
rect 2860 -820 2930 -750
rect 3090 -820 3160 -750
rect 3320 -820 3390 -750
rect 3550 -820 3620 -750
rect 3780 -820 3850 -750
rect 4010 -820 4080 -750
rect 4240 -820 4310 -750
rect 4470 -820 4540 -750
rect 4700 -820 4770 -750
rect 4930 -820 5000 -750
rect 5160 -820 5230 -750
rect 5390 -820 5460 -750
rect 5620 -820 5690 -750
rect 5850 -820 5920 -750
rect 6080 -820 6150 -750
rect 6310 -820 6380 -750
rect 6540 -820 6610 -750
rect 6770 -820 6840 -750
rect 7000 -820 7070 -750
<< metal2 >>
rect 310 610 420 630
rect 540 610 650 630
rect 770 610 880 630
rect 1000 610 1110 630
rect 1230 610 1340 630
rect 1460 610 1570 630
rect 310 540 330 610
rect 400 540 560 610
rect 630 540 790 610
rect 860 540 910 610
rect 970 540 1020 610
rect 1090 540 1250 610
rect 1320 540 1480 610
rect 1550 540 1570 610
rect 310 520 420 540
rect 540 520 650 540
rect 770 520 880 540
rect 1000 520 1110 540
rect 1230 520 1340 540
rect 1460 520 1570 540
rect 1690 610 1800 630
rect 1920 610 2030 630
rect 2150 610 2260 630
rect 2380 610 2490 630
rect 2610 610 2720 630
rect 2840 610 2950 630
rect 3070 620 3410 630
rect 3070 610 3200 620
rect 1690 540 1710 610
rect 1780 540 1940 610
rect 2010 540 2170 610
rect 2240 540 2400 610
rect 2470 540 2630 610
rect 2700 540 2860 610
rect 2930 540 3090 610
rect 3160 540 3200 610
rect 1690 520 1800 540
rect 1920 520 2030 540
rect 2150 520 2260 540
rect 2380 520 2490 540
rect 2610 520 2720 540
rect 2840 520 2950 540
rect 3070 530 3200 540
rect 3280 610 3410 620
rect 3530 610 3640 630
rect 3760 610 3870 630
rect 3990 610 4100 630
rect 4220 610 4330 630
rect 4450 620 4790 630
rect 4450 610 4580 620
rect 3280 540 3320 610
rect 3390 540 3550 610
rect 3620 540 3780 610
rect 3850 540 4010 610
rect 4080 540 4240 610
rect 4310 540 4470 610
rect 4540 540 4580 610
rect 3280 530 3410 540
rect 3070 520 3410 530
rect 3530 520 3640 540
rect 3760 520 3870 540
rect 3990 520 4100 540
rect 4220 520 4330 540
rect 4450 530 4580 540
rect 4660 610 4790 620
rect 4910 610 5020 630
rect 5140 610 5250 630
rect 5370 610 5480 630
rect 5600 610 5710 630
rect 5830 610 5940 630
rect 6060 610 6170 630
rect 6290 610 6400 630
rect 6520 610 6630 630
rect 6750 610 6860 630
rect 6980 610 7090 630
rect 4660 540 4700 610
rect 4770 540 4930 610
rect 5000 540 5160 610
rect 5230 540 5390 610
rect 5460 540 5620 610
rect 5690 540 5850 610
rect 5920 540 6080 610
rect 6150 540 6310 610
rect 6380 540 6540 610
rect 6610 540 6770 610
rect 6840 540 7000 610
rect 7070 540 7090 610
rect 4660 530 4790 540
rect 4450 520 4790 530
rect 4910 520 5020 540
rect 5140 520 5250 540
rect 5370 520 5480 540
rect 5600 520 5710 540
rect 5830 520 5940 540
rect 6060 520 6170 540
rect 6290 520 6400 540
rect 6520 520 6630 540
rect 6750 520 6860 540
rect 6980 520 7090 540
rect 180 450 320 470
rect 180 350 200 450
rect 300 430 320 450
rect 640 450 780 470
rect 640 430 660 450
rect 300 370 660 430
rect 300 350 320 370
rect 180 330 320 350
rect 640 350 660 370
rect 760 430 780 450
rect 1100 450 1240 470
rect 1100 430 1120 450
rect 760 370 1120 430
rect 760 350 780 370
rect 640 330 780 350
rect 1100 350 1120 370
rect 1220 430 1240 450
rect 1560 450 1700 470
rect 1560 430 1580 450
rect 1220 370 1580 430
rect 1220 350 1240 370
rect 1100 330 1240 350
rect 1560 350 1580 370
rect 1680 430 1700 450
rect 2020 450 2160 470
rect 2020 430 2040 450
rect 1680 370 2040 430
rect 1680 350 1700 370
rect 1560 330 1700 350
rect 2020 350 2040 370
rect 2140 430 2160 450
rect 2480 450 2620 470
rect 2480 430 2500 450
rect 2140 370 2500 430
rect 2140 350 2160 370
rect 2020 330 2160 350
rect 2480 350 2500 370
rect 2600 430 2620 450
rect 2940 450 3080 470
rect 2940 430 2960 450
rect 2600 370 2960 430
rect 2600 350 2620 370
rect 2480 330 2620 350
rect 2940 350 2960 370
rect 3060 430 3080 450
rect 3400 450 3540 470
rect 3400 430 3420 450
rect 3060 370 3420 430
rect 3060 350 3080 370
rect 2940 330 3080 350
rect 3400 350 3420 370
rect 3520 430 3540 450
rect 3860 450 4000 470
rect 3860 430 3880 450
rect 3520 370 3880 430
rect 3520 350 3540 370
rect 3400 330 3540 350
rect 3860 350 3880 370
rect 3980 430 4000 450
rect 4320 450 4460 470
rect 4320 430 4340 450
rect 3980 370 4340 430
rect 3980 350 4000 370
rect 3860 330 4000 350
rect 4320 350 4340 370
rect 4440 430 4460 450
rect 4780 450 4920 470
rect 4780 430 4800 450
rect 4440 370 4800 430
rect 4440 350 4460 370
rect 4320 330 4460 350
rect 4780 350 4800 370
rect 4900 430 4920 450
rect 5240 450 5380 470
rect 5240 430 5260 450
rect 4900 370 5260 430
rect 4900 350 4920 370
rect 4780 330 4920 350
rect 5240 350 5260 370
rect 5360 430 5380 450
rect 5700 450 5840 470
rect 5700 430 5720 450
rect 5360 370 5720 430
rect 5360 350 5380 370
rect 5240 330 5380 350
rect 5700 350 5720 370
rect 5820 430 5840 450
rect 6160 450 6300 470
rect 6160 430 6180 450
rect 5820 370 6180 430
rect 5820 350 5840 370
rect 5700 330 5840 350
rect 6160 350 6180 370
rect 6280 430 6300 450
rect 6620 450 6760 470
rect 6620 430 6640 450
rect 6280 370 6640 430
rect 6280 350 6300 370
rect 6160 330 6300 350
rect 6620 350 6640 370
rect 6740 430 6760 450
rect 7080 450 7220 470
rect 7080 430 7100 450
rect 6740 370 7100 430
rect 6740 350 6760 370
rect 6620 330 6760 350
rect 7080 350 7100 370
rect 7200 350 7220 450
rect 7080 330 7220 350
rect 410 150 550 170
rect 410 50 430 150
rect 530 130 550 150
rect 870 150 1010 170
rect 870 130 890 150
rect 530 70 890 130
rect 530 50 550 70
rect 410 30 550 50
rect 870 50 890 70
rect 990 130 1010 150
rect 1330 150 1470 170
rect 1330 130 1350 150
rect 990 70 1350 130
rect 990 50 1010 70
rect 870 30 1010 50
rect 1330 50 1350 70
rect 1450 50 1470 150
rect 1790 150 1930 170
rect 1790 130 1810 150
rect 1730 70 1810 130
rect 1330 30 1470 50
rect 1790 50 1810 70
rect 1910 130 1930 150
rect 2250 150 2390 170
rect 2250 130 2270 150
rect 1910 70 2270 130
rect 1910 50 1930 70
rect 1790 30 1930 50
rect 2250 50 2270 70
rect 2370 130 2390 150
rect 2710 150 2850 170
rect 2710 130 2730 150
rect 2370 70 2730 130
rect 2370 50 2390 70
rect 2250 30 2390 50
rect 2710 50 2730 70
rect 2830 130 2850 150
rect 3170 150 3310 170
rect 3170 130 3190 150
rect 2830 70 3190 130
rect 2830 50 2850 70
rect 2710 30 2850 50
rect 3170 50 3190 70
rect 3290 130 3310 150
rect 3630 150 3770 170
rect 3630 130 3650 150
rect 3290 70 3650 130
rect 3290 50 3310 70
rect 3170 30 3310 50
rect 3630 50 3650 70
rect 3750 130 3770 150
rect 4090 150 4230 170
rect 4090 130 4110 150
rect 3750 70 4110 130
rect 3750 50 3770 70
rect 3630 30 3770 50
rect 4090 50 4110 70
rect 4210 130 4230 150
rect 4550 150 4690 170
rect 4550 130 4570 150
rect 4210 70 4570 130
rect 4210 50 4230 70
rect 4090 30 4230 50
rect 4550 50 4570 70
rect 4670 130 4690 150
rect 5010 150 5150 170
rect 5010 130 5030 150
rect 4670 70 5030 130
rect 4670 50 4690 70
rect 4550 30 4690 50
rect 5010 50 5030 70
rect 5130 130 5150 150
rect 5470 150 5610 170
rect 5470 130 5490 150
rect 5130 70 5490 130
rect 5130 50 5150 70
rect 5010 30 5150 50
rect 5470 50 5490 70
rect 5590 130 5610 150
rect 5930 150 6070 170
rect 5930 130 5950 150
rect 5590 70 5950 130
rect 5590 50 5610 70
rect 5470 30 5610 50
rect 5930 50 5950 70
rect 6050 130 6070 150
rect 6390 150 6530 170
rect 6390 130 6410 150
rect 6050 70 6410 130
rect 6050 50 6070 70
rect 5930 30 6070 50
rect 6390 50 6410 70
rect 6510 130 6530 150
rect 6850 150 6990 170
rect 6850 130 6870 150
rect 6510 70 6870 130
rect 6510 50 6530 70
rect 6390 30 6530 50
rect 6850 50 6870 70
rect 6970 130 6990 150
rect 6970 70 7050 130
rect 6970 50 6990 70
rect 6850 30 6990 50
rect 410 -260 550 -240
rect 410 -360 430 -260
rect 530 -280 550 -260
rect 870 -260 1010 -240
rect 870 -280 890 -260
rect 530 -340 890 -280
rect 530 -360 550 -340
rect 410 -380 550 -360
rect 870 -360 890 -340
rect 990 -280 1010 -260
rect 1330 -260 1470 -240
rect 1330 -280 1350 -260
rect 990 -340 1350 -280
rect 990 -360 1010 -340
rect 870 -380 1010 -360
rect 1330 -360 1350 -340
rect 1450 -360 1470 -260
rect 1790 -260 1930 -240
rect 1790 -280 1810 -260
rect 1730 -340 1810 -280
rect 1330 -380 1470 -360
rect 1790 -360 1810 -340
rect 1910 -280 1930 -260
rect 2250 -260 2390 -240
rect 2250 -280 2270 -260
rect 1910 -340 2270 -280
rect 1910 -360 1930 -340
rect 1790 -380 1930 -360
rect 2250 -360 2270 -340
rect 2370 -280 2390 -260
rect 2710 -260 2850 -240
rect 2710 -280 2730 -260
rect 2370 -340 2730 -280
rect 2370 -360 2390 -340
rect 2250 -380 2390 -360
rect 2710 -360 2730 -340
rect 2830 -280 2850 -260
rect 3170 -260 3310 -240
rect 3170 -280 3190 -260
rect 2830 -340 3190 -280
rect 2830 -360 2850 -340
rect 2710 -380 2850 -360
rect 3170 -360 3190 -340
rect 3290 -280 3310 -260
rect 3630 -260 3770 -240
rect 3630 -280 3650 -260
rect 3290 -340 3650 -280
rect 3290 -360 3310 -340
rect 3170 -380 3310 -360
rect 3630 -360 3650 -340
rect 3750 -280 3770 -260
rect 4090 -260 4230 -240
rect 4090 -280 4110 -260
rect 3750 -340 4110 -280
rect 3750 -360 3770 -340
rect 3630 -380 3770 -360
rect 4090 -360 4110 -340
rect 4210 -280 4230 -260
rect 4550 -260 4690 -240
rect 4550 -280 4570 -260
rect 4210 -340 4570 -280
rect 4210 -360 4230 -340
rect 4090 -380 4230 -360
rect 4550 -360 4570 -340
rect 4670 -280 4690 -260
rect 5010 -260 5150 -240
rect 5010 -280 5030 -260
rect 4670 -340 5030 -280
rect 4670 -360 4690 -340
rect 4550 -380 4690 -360
rect 5010 -360 5030 -340
rect 5130 -280 5150 -260
rect 5470 -260 5610 -240
rect 5470 -280 5490 -260
rect 5130 -340 5490 -280
rect 5130 -360 5150 -340
rect 5010 -380 5150 -360
rect 5470 -360 5490 -340
rect 5590 -280 5610 -260
rect 5930 -260 6070 -240
rect 5930 -280 5950 -260
rect 5590 -340 5950 -280
rect 5590 -360 5610 -340
rect 5470 -380 5610 -360
rect 5930 -360 5950 -340
rect 6050 -280 6070 -260
rect 6390 -260 6530 -240
rect 6390 -280 6410 -260
rect 6050 -340 6410 -280
rect 6050 -360 6070 -340
rect 5930 -380 6070 -360
rect 6390 -360 6410 -340
rect 6510 -280 6530 -260
rect 6850 -260 6990 -240
rect 6850 -280 6870 -260
rect 6510 -340 6870 -280
rect 6510 -360 6530 -340
rect 6390 -380 6530 -360
rect 6850 -360 6870 -340
rect 6970 -280 6990 -260
rect 6970 -340 7050 -280
rect 6970 -360 6990 -340
rect 6850 -380 6990 -360
rect 180 -560 320 -540
rect 180 -660 200 -560
rect 300 -580 320 -560
rect 640 -560 780 -540
rect 640 -580 660 -560
rect 300 -640 660 -580
rect 300 -660 320 -640
rect 180 -680 320 -660
rect 640 -660 660 -640
rect 760 -580 780 -560
rect 1100 -560 1240 -540
rect 1100 -580 1120 -560
rect 760 -640 1120 -580
rect 760 -660 780 -640
rect 640 -680 780 -660
rect 1100 -660 1120 -640
rect 1220 -580 1240 -560
rect 1560 -560 1700 -540
rect 1560 -580 1580 -560
rect 1220 -640 1580 -580
rect 1220 -660 1240 -640
rect 1100 -680 1240 -660
rect 1560 -660 1580 -640
rect 1680 -580 1700 -560
rect 2020 -560 2160 -540
rect 2020 -580 2040 -560
rect 1680 -640 2040 -580
rect 1680 -660 1700 -640
rect 1560 -680 1700 -660
rect 2020 -660 2040 -640
rect 2140 -580 2160 -560
rect 2480 -560 2620 -540
rect 2480 -580 2500 -560
rect 2140 -640 2500 -580
rect 2140 -660 2160 -640
rect 2020 -680 2160 -660
rect 2480 -660 2500 -640
rect 2600 -580 2620 -560
rect 2940 -560 3080 -540
rect 2940 -580 2960 -560
rect 2600 -640 2960 -580
rect 2600 -660 2620 -640
rect 2480 -680 2620 -660
rect 2940 -660 2960 -640
rect 3060 -580 3080 -560
rect 3400 -560 3540 -540
rect 3400 -580 3420 -560
rect 3060 -640 3420 -580
rect 3060 -660 3080 -640
rect 2940 -680 3080 -660
rect 3400 -660 3420 -640
rect 3520 -580 3540 -560
rect 3860 -560 4000 -540
rect 3860 -580 3880 -560
rect 3520 -640 3880 -580
rect 3520 -660 3540 -640
rect 3400 -680 3540 -660
rect 3860 -660 3880 -640
rect 3980 -580 4000 -560
rect 4320 -560 4460 -540
rect 4320 -580 4340 -560
rect 3980 -640 4340 -580
rect 3980 -660 4000 -640
rect 3860 -680 4000 -660
rect 4320 -660 4340 -640
rect 4440 -580 4460 -560
rect 4780 -560 4920 -540
rect 4780 -580 4800 -560
rect 4440 -640 4800 -580
rect 4440 -660 4460 -640
rect 4320 -680 4460 -660
rect 4780 -660 4800 -640
rect 4900 -580 4920 -560
rect 5240 -560 5380 -540
rect 5240 -580 5260 -560
rect 4900 -640 5260 -580
rect 4900 -660 4920 -640
rect 4780 -680 4920 -660
rect 5240 -660 5260 -640
rect 5360 -580 5380 -560
rect 5700 -560 5840 -540
rect 5700 -580 5720 -560
rect 5360 -640 5720 -580
rect 5360 -660 5380 -640
rect 5240 -680 5380 -660
rect 5700 -660 5720 -640
rect 5820 -580 5840 -560
rect 6160 -560 6300 -540
rect 6160 -580 6180 -560
rect 5820 -640 6180 -580
rect 5820 -660 5840 -640
rect 5700 -680 5840 -660
rect 6160 -660 6180 -640
rect 6280 -580 6300 -560
rect 6620 -560 6760 -540
rect 6620 -580 6640 -560
rect 6280 -640 6640 -580
rect 6280 -660 6300 -640
rect 6160 -680 6300 -660
rect 6620 -660 6640 -640
rect 6740 -580 6760 -560
rect 7080 -560 7220 -540
rect 7080 -580 7100 -560
rect 6740 -640 7100 -580
rect 6740 -660 6760 -640
rect 6620 -680 6760 -660
rect 7080 -660 7100 -640
rect 7200 -660 7220 -560
rect 7080 -680 7220 -660
rect 310 -750 420 -730
rect 540 -750 650 -730
rect 770 -750 880 -730
rect 1000 -750 1110 -730
rect 1230 -750 1340 -730
rect 1460 -750 1570 -730
rect 310 -820 330 -750
rect 400 -820 560 -750
rect 630 -820 790 -750
rect 860 -820 910 -750
rect 970 -820 1020 -750
rect 1090 -820 1250 -750
rect 1320 -820 1480 -750
rect 1550 -820 1570 -750
rect 310 -840 420 -820
rect 540 -840 650 -820
rect 770 -840 880 -820
rect 1000 -840 1110 -820
rect 1230 -840 1340 -820
rect 1460 -840 1570 -820
rect 1690 -750 1800 -730
rect 1920 -750 2030 -730
rect 2150 -750 2260 -730
rect 2380 -750 2490 -730
rect 2610 -750 2720 -730
rect 2840 -750 2950 -730
rect 3070 -750 3180 -730
rect 3300 -750 3410 -730
rect 3530 -740 3870 -730
rect 3530 -750 3660 -740
rect 1690 -820 1710 -750
rect 1780 -820 1940 -750
rect 2010 -820 2170 -750
rect 2240 -820 2400 -750
rect 2470 -820 2630 -750
rect 2700 -820 2860 -750
rect 2930 -820 3090 -750
rect 3160 -820 3320 -750
rect 3390 -820 3550 -750
rect 3620 -820 3660 -750
rect 1690 -840 1800 -820
rect 1920 -840 2030 -820
rect 2150 -840 2260 -820
rect 2380 -840 2490 -820
rect 2610 -840 2720 -820
rect 2840 -840 2950 -820
rect 3070 -840 3180 -820
rect 3300 -840 3410 -820
rect 3530 -830 3660 -820
rect 3740 -750 3870 -740
rect 3990 -750 4100 -730
rect 4220 -750 4330 -730
rect 4450 -750 4560 -730
rect 4680 -750 4790 -730
rect 4910 -740 5250 -730
rect 4910 -750 5040 -740
rect 3740 -820 3780 -750
rect 3850 -820 4010 -750
rect 4080 -820 4240 -750
rect 4310 -820 4470 -750
rect 4540 -820 4700 -750
rect 4770 -820 4930 -750
rect 5000 -820 5040 -750
rect 3740 -830 3870 -820
rect 3530 -840 3870 -830
rect 3990 -840 4100 -820
rect 4220 -840 4330 -820
rect 4450 -840 4560 -820
rect 4680 -840 4790 -820
rect 4910 -830 5040 -820
rect 5120 -750 5250 -740
rect 5370 -750 5480 -730
rect 5600 -750 5710 -730
rect 5830 -750 5940 -730
rect 6060 -750 6170 -730
rect 6290 -750 6400 -730
rect 6520 -750 6630 -730
rect 6750 -750 6860 -730
rect 6980 -750 7090 -730
rect 5120 -820 5160 -750
rect 5230 -820 5390 -750
rect 5460 -820 5620 -750
rect 5690 -820 5850 -750
rect 5920 -820 6080 -750
rect 6150 -820 6310 -750
rect 6380 -820 6540 -750
rect 6610 -820 6770 -750
rect 6840 -820 7000 -750
rect 7070 -820 7090 -750
rect 5120 -830 5250 -820
rect 4910 -840 5250 -830
rect 5370 -840 5480 -820
rect 5600 -840 5710 -820
rect 5830 -840 5940 -820
rect 6060 -840 6170 -820
rect 6290 -840 6400 -820
rect 6520 -840 6630 -820
rect 6750 -840 6860 -820
rect 6980 -840 7090 -820
<< via2 >>
rect 910 540 970 610
rect 3200 530 3280 620
rect 4580 530 4660 620
rect 200 350 300 450
rect 430 50 530 150
rect 890 50 990 150
rect 1350 50 1450 150
rect 1810 50 1910 150
rect 3650 50 3750 150
rect 4110 50 4210 150
rect 5030 50 5130 150
rect 6870 50 6970 150
rect 430 -360 530 -260
rect 890 -360 990 -260
rect 1350 -360 1450 -260
rect 1810 -360 1910 -260
rect 3190 -360 3290 -260
rect 4110 -360 4210 -260
rect 4570 -360 4670 -260
rect 6870 -360 6970 -260
rect 200 -660 300 -560
rect 910 -820 970 -750
rect 3660 -830 3740 -740
rect 5040 -830 5120 -740
<< metal3 >>
rect -1590 -560 -370 1010
rect 820 790 1060 820
rect 820 710 850 790
rect 930 710 950 790
rect 1030 710 1060 790
rect 820 680 1060 710
rect 1730 800 1970 830
rect 1730 720 1760 800
rect 1840 720 1860 800
rect 1940 720 1970 800
rect 1730 690 1970 720
rect 4030 800 4270 830
rect 4030 720 4060 800
rect 4140 720 4160 800
rect 4240 720 4270 800
rect 4030 690 4270 720
rect 6790 800 7030 830
rect 6790 720 6820 800
rect 6900 720 6920 800
rect 7000 720 7030 800
rect 6790 690 7030 720
rect 910 620 970 680
rect 900 610 980 620
rect 900 540 910 610
rect 970 540 980 610
rect 900 530 980 540
rect 180 450 320 470
rect 180 350 200 450
rect 300 350 320 450
rect 180 330 320 350
rect 1820 170 1900 690
rect 3190 620 3290 630
rect 3190 530 3200 620
rect 3280 530 3290 620
rect 410 150 550 170
rect 410 50 430 150
rect 530 50 550 150
rect 410 30 550 50
rect 870 150 1010 170
rect 870 50 890 150
rect 990 50 1010 150
rect 870 30 1010 50
rect 1330 150 1470 170
rect 1330 50 1350 150
rect 1450 50 1470 150
rect 1330 30 1470 50
rect 1790 150 1930 170
rect 1790 50 1810 150
rect 1910 50 1930 150
rect 1790 30 1930 50
rect 450 -50 510 30
rect 910 -50 970 30
rect 1370 -50 1430 30
rect 430 -60 530 -50
rect 430 -150 440 -60
rect 520 -150 530 -60
rect 430 -160 530 -150
rect 890 -60 990 -50
rect 890 -150 900 -60
rect 980 -150 990 -60
rect 890 -160 990 -150
rect 1350 -60 1450 -50
rect 1350 -150 1360 -60
rect 1440 -150 1450 -60
rect 1350 -160 1450 -150
rect 450 -240 510 -160
rect 910 -240 970 -160
rect 1370 -240 1430 -160
rect 3190 -240 3290 530
rect 4120 170 4200 690
rect 4570 620 4670 630
rect 4570 530 4580 620
rect 4660 530 4670 620
rect 3630 150 3770 170
rect 3630 50 3650 150
rect 3750 50 3770 150
rect 3630 30 3770 50
rect 4090 150 4230 170
rect 4090 50 4110 150
rect 4210 50 4230 150
rect 4090 30 4230 50
rect 410 -260 550 -240
rect 410 -360 430 -260
rect 530 -360 550 -260
rect 410 -380 550 -360
rect 870 -260 1010 -240
rect 870 -360 890 -260
rect 990 -360 1010 -260
rect 870 -380 1010 -360
rect 1330 -260 1470 -240
rect 1330 -360 1350 -260
rect 1450 -360 1470 -260
rect 1330 -380 1470 -360
rect 1790 -260 1930 -240
rect 1790 -360 1810 -260
rect 1910 -360 1930 -260
rect 1790 -380 1930 -360
rect 3170 -260 3310 -240
rect 3170 -360 3190 -260
rect 3290 -360 3310 -260
rect 3170 -380 3310 -360
rect 180 -560 320 -540
rect -1590 -660 200 -560
rect 300 -660 320 -560
rect -1590 -1190 -370 -660
rect 180 -680 320 -660
rect 900 -750 980 -740
rect 900 -820 910 -750
rect 970 -820 980 -750
rect 900 -830 980 -820
rect 910 -890 970 -830
rect 820 -920 1060 -890
rect 1820 -900 1900 -380
rect 3650 -740 3750 30
rect 4570 -240 4670 530
rect 6880 170 6960 690
rect 5010 150 5150 170
rect 5010 50 5030 150
rect 5130 50 5150 150
rect 5010 30 5150 50
rect 6850 150 6990 170
rect 6850 50 6870 150
rect 6970 50 6990 150
rect 6850 30 6990 50
rect 4090 -260 4230 -240
rect 4090 -360 4110 -260
rect 4210 -360 4230 -260
rect 4090 -380 4230 -360
rect 4550 -260 4690 -240
rect 4550 -360 4570 -260
rect 4670 -360 4690 -260
rect 4550 -380 4690 -360
rect 3650 -830 3660 -740
rect 3740 -830 3750 -740
rect 3650 -840 3750 -830
rect 4120 -900 4200 -380
rect 5030 -740 5130 30
rect 6850 -260 6990 -240
rect 6850 -360 6870 -260
rect 6970 -360 6990 -260
rect 6850 -380 6990 -360
rect 5030 -830 5040 -740
rect 5120 -830 5130 -740
rect 5030 -840 5130 -830
rect 6880 -900 6960 -380
rect 820 -1000 850 -920
rect 930 -1000 950 -920
rect 1030 -1000 1060 -920
rect 820 -1030 1060 -1000
rect 1740 -930 1980 -900
rect 1740 -1010 1770 -930
rect 1850 -1010 1870 -930
rect 1950 -1010 1980 -930
rect 1740 -1040 1980 -1010
rect 4040 -930 4280 -900
rect 6800 -930 7040 -900
rect 4040 -1010 4070 -930
rect 4150 -1010 4170 -930
rect 4250 -1000 6830 -930
rect 4250 -1010 4280 -1000
rect 4040 -1040 4280 -1010
rect 6800 -1010 6830 -1000
rect 6910 -1010 6930 -930
rect 7010 -1010 7040 -930
rect 6800 -1040 7040 -1010
<< via3 >>
rect 850 710 930 790
rect 950 710 1030 790
rect 1760 720 1840 800
rect 1860 720 1940 800
rect 4060 720 4140 800
rect 4160 720 4240 800
rect 6820 720 6900 800
rect 6920 720 7000 800
rect 200 350 300 450
rect 440 -150 520 -60
rect 900 -150 980 -60
rect 1360 -150 1440 -60
rect 6870 50 6970 150
rect 6870 -360 6970 -260
rect 850 -1000 930 -920
rect 950 -1000 1030 -920
rect 1770 -1010 1850 -930
rect 1870 -1010 1950 -930
rect 4070 -1010 4150 -930
rect 4170 -1010 4250 -930
rect 6830 -1010 6910 -930
rect 6930 -1010 7010 -930
<< mimcap >>
rect -1490 870 -448 910
rect -1490 -1050 -1450 870
rect -488 -1050 -448 870
rect -1490 -1090 -448 -1050
<< mimcapcontact >>
rect -1450 -1050 -488 870
<< metal4 >>
rect -1451 870 -487 871
rect -1451 -1050 -1450 870
rect -488 450 -487 870
rect 820 790 1060 820
rect 1730 800 1970 830
rect 1730 790 1760 800
rect 820 710 850 790
rect 930 710 950 790
rect 1030 720 1760 790
rect 1840 720 1860 800
rect 1940 790 1970 800
rect 4030 800 4270 830
rect 4030 790 4060 800
rect 1940 720 4060 790
rect 4140 720 4160 800
rect 4240 790 4270 800
rect 6790 800 7030 830
rect 6790 790 6820 800
rect 4240 720 6820 790
rect 6900 720 6920 800
rect 7000 720 7030 800
rect 1030 710 1060 720
rect 820 680 1060 710
rect 1730 690 1970 720
rect 4030 690 4270 720
rect 6790 690 7030 720
rect 180 450 320 470
rect -488 350 200 450
rect 300 350 320 450
rect -488 -1050 -487 350
rect 180 330 320 350
rect 6850 150 6990 170
rect 6850 50 6870 150
rect 6970 130 6990 150
rect 6970 70 7500 130
rect 6970 50 6990 70
rect 6850 30 6990 50
rect 430 -60 530 -50
rect 890 -60 990 -50
rect 1350 -60 1450 -50
rect 130 -150 440 -60
rect 520 -150 900 -60
rect 980 -150 1360 -60
rect 1440 -150 1580 -60
rect 430 -160 530 -150
rect 890 -160 990 -150
rect 1350 -160 1450 -150
rect 6850 -260 6990 -240
rect 6850 -360 6870 -260
rect 6970 -280 6990 -260
rect 6970 -340 7500 -280
rect 6970 -360 6990 -340
rect 6850 -380 6990 -360
rect 820 -920 1060 -890
rect 820 -1000 850 -920
rect 930 -1000 950 -920
rect 1030 -930 1060 -920
rect 1740 -930 1980 -900
rect 4040 -930 4280 -900
rect 6800 -930 7040 -900
rect 1030 -1000 1770 -930
rect 820 -1030 1060 -1000
rect 1740 -1010 1770 -1000
rect 1850 -1010 1870 -930
rect 1950 -1000 4070 -930
rect 1950 -1010 1980 -1000
rect 1740 -1040 1980 -1010
rect 4040 -1010 4070 -1000
rect 4150 -1010 4170 -930
rect 4250 -1000 6830 -930
rect 4250 -1010 4280 -1000
rect 4040 -1040 4280 -1010
rect 6800 -1010 6830 -1000
rect 6910 -1010 6930 -930
rect 7010 -1010 7040 -930
rect 6800 -1040 7040 -1010
rect -1451 -1051 -487 -1050
<< labels >>
rlabel metal4 7430 100 7430 100 1 von
rlabel metal4 7440 -310 7440 -310 1 vop
rlabel via3 470 -110 470 -110 1 Gnd
<< end >>
