magic
tech sky130A
timestamp 1641018497
<< viali >>
rect 4865 645 4885 665
<< metal1 >>
rect 7050 1205 7085 1215
rect 7005 1190 7085 1205
rect 7050 1180 7085 1190
rect 7055 1070 7090 1080
rect 7005 1055 7090 1070
rect 7055 1045 7090 1055
rect 4855 670 4895 675
rect 4855 640 4860 670
rect 4890 640 4895 670
rect 4855 635 4895 640
<< via1 >>
rect 4860 665 4890 670
rect 4860 645 4865 665
rect 4865 645 4885 665
rect 4885 645 4890 665
rect 4860 640 4890 645
<< metal2 >>
rect 5410 1240 5445 1275
rect 245 685 285 695
rect 245 665 315 685
rect 4850 670 4900 680
rect 245 655 285 665
rect 4850 640 4860 670
rect 4890 640 4900 670
rect 4850 630 4900 640
rect 4875 415 4890 630
rect 4875 400 5430 415
use pd  pd_0
timestamp 1640980777
transform 1 0 5535 0 1 855
box -215 -855 1685 810
use divider  divider_0
timestamp 1641018497
transform 1 0 490 0 1 235
box -490 -235 4690 2150
<< end >>
