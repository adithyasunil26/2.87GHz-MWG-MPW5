magic
tech sky130A
timestamp 1647806434
<< locali >>
rect -151 4655 4 4664
rect -151 4633 -137 4655
rect -152 4524 -137 4633
rect -5 4524 4 4655
rect -152 4507 4 4524
rect -152 4037 3 4507
rect -152 3891 3965 4037
rect -42 3886 3965 3891
rect 3805 3537 3955 3886
rect 27 1458 160 2216
rect 27 1334 581 1458
rect 4708 1370 5156 1530
rect 49 1331 581 1334
rect 448 1255 578 1331
rect 3820 250 3950 255
rect -914 -109 -16 -107
rect 3810 -109 3950 250
rect -914 -243 3950 -109
rect -914 -245 3940 -243
rect -914 -254 -16 -245
rect 3810 -248 3940 -245
rect -904 -3082 -762 -254
rect -468 -436 85 -417
rect 5022 -431 5156 1370
rect 2573 -436 5156 -431
rect -468 -437 5156 -436
rect -478 -466 5156 -437
rect -478 -581 5151 -466
rect -478 -586 2593 -581
rect -478 -589 85 -586
rect -478 -1522 -341 -589
rect -198 -1522 5 -1500
rect -488 -1528 5 -1522
rect -488 -1653 -168 -1528
rect -33 -1653 5 -1528
rect -488 -1664 5 -1653
rect -198 -1676 5 -1664
rect -208 -3082 -18 -3069
rect -909 -3085 -18 -3082
rect -909 -3102 -13 -3085
rect -909 -3211 -160 -3102
rect -48 -3211 -13 -3102
rect -909 -3224 -13 -3211
rect -208 -3232 -13 -3224
<< viali >>
rect -137 4524 -5 4655
rect -168 -1653 -33 -1528
rect -160 -3211 -48 -3102
<< metal1 >>
rect -151 4655 4 4664
rect -151 4524 -137 4655
rect -5 4524 4 4655
rect -151 4507 4 4524
rect -198 -1528 5 -1500
rect -198 -1653 -168 -1528
rect -33 -1653 5 -1528
rect -198 -1676 5 -1653
rect -208 -3085 -18 -3069
rect -208 -3102 -13 -3085
rect -208 -3211 -160 -3102
rect -48 -3211 -13 -3102
rect -208 -3232 -13 -3211
<< via1 >>
rect -137 4524 -5 4655
rect -168 -1653 -33 -1528
rect -160 -3211 -48 -3102
<< metal2 >>
rect -151 4655 4 4664
rect -151 4524 -137 4655
rect -5 4524 4 4655
rect -151 4507 4 4524
rect -198 -1528 5 -1500
rect -198 -1653 -168 -1528
rect -33 -1653 5 -1528
rect -198 -1676 5 -1653
rect -208 -3085 -18 -3069
rect -208 -3102 -13 -3085
rect -208 -3211 -160 -3102
rect -48 -3211 -13 -3102
rect -208 -3232 -13 -3211
<< via2 >>
rect -137 4524 -5 4655
rect -168 -1653 -33 -1528
rect -160 -3211 -48 -3102
<< metal3 >>
rect -151 4655 4 4664
rect -151 4524 -137 4655
rect -5 4524 4 4655
rect -151 4507 4 4524
rect -198 -1528 5 -1500
rect -198 -1653 -168 -1528
rect -33 -1653 5 -1528
rect -198 -1676 5 -1653
rect -208 -3085 -18 -3069
rect -208 -3102 -13 -3085
rect -208 -3211 -160 -3102
rect -48 -3211 -13 -3102
rect -208 -3232 -13 -3211
<< via3 >>
rect -137 4524 -5 4655
rect -168 -1653 -33 -1528
rect -160 -3211 -48 -3102
<< metal4 >>
rect -1048 4969 321 4970
rect -1392 4834 321 4969
rect -1381 294 -1184 4834
rect -152 4655 21 4672
rect -152 4524 -137 4655
rect -5 4524 21 4655
rect -152 4518 21 4524
rect -151 4507 4 4518
rect -1381 -1 249 294
rect -1381 -1237 -1184 -1
rect -1381 -1373 344 -1237
rect -1381 -2787 -1184 -1373
rect -198 -1528 5 -1500
rect -198 -1653 -168 -1528
rect -33 -1653 5 -1528
rect -198 -1676 5 -1653
rect -1398 -2923 315 -2787
rect -26 -3069 112 -3064
rect -208 -3102 112 -3069
rect -208 -3211 -160 -3102
rect -48 -3138 112 -3102
rect -48 -3211 96 -3138
rect -208 -3219 96 -3211
rect -208 -3232 -13 -3219
<< via4 >>
rect 265 3605 393 3724
<< metal5 >>
rect 191 3893 410 4220
rect -345 3724 410 3893
rect -345 3705 265 3724
rect -339 -576 -151 3705
rect 191 3605 265 3705
rect 393 3605 410 3724
rect 191 3579 410 3605
rect -339 -753 392 -576
rect -339 -776 386 -753
rect 169 -2019 397 -2008
rect 157 -2373 397 -2019
rect 157 -2384 385 -2373
use cp  cp_0
timestamp 1640911461
transform 1 0 415 0 1 1715
box -415 -1715 4690 2035
use tapered_buf  tapered_buf_0
timestamp 1647784636
transform 1 0 469 0 1 5051
box -470 -910 43675 400
use tapered_buf  tapered_buf_1
timestamp 1647784636
transform 1 0 447 0 1 -1140
box -470 -910 43675 400
use tapered_buf  tapered_buf_2
timestamp 1647784636
transform 1 0 447 0 1 -2688
box -470 -910 43675 400
<< labels >>
rlabel space 5 5096 5 5096 1 up
rlabel space 7 -1106 7 -1106 1 out
rlabel space -11 -2638 -11 -2638 1 down
rlabel metal4 -1257 -2167 -1257 -2167 1 gnd!
rlabel metal5 311 -2207 311 -2207 1 vdd!
<< end >>
