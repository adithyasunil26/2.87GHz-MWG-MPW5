magic
tech sky130A
timestamp 1640997741
<< locali >>
rect 4960 3650 4980 3670
rect 4935 3130 4975 3170
<< viali >>
rect 4940 3650 4960 3670
rect 9555 645 9580 670
<< metal1 >>
rect 4930 3675 4970 3680
rect 4930 3645 4935 3675
rect 4965 3645 4970 3675
rect 4930 3640 4970 3645
rect 9545 675 9590 680
rect 9545 640 9550 675
rect 9585 640 9590 675
rect 9545 635 9590 640
<< via1 >>
rect 4935 3670 4965 3675
rect 4935 3650 4940 3670
rect 4940 3650 4960 3670
rect 4960 3650 4965 3670
rect 4935 3645 4965 3650
rect 9550 670 9585 675
rect 9550 645 9555 670
rect 9555 645 9580 670
rect 9580 645 9585 670
rect 9550 640 9585 645
<< metal2 >>
rect 4055 5985 4675 6105
rect 4650 685 4675 5985
rect 4925 3675 4975 3685
rect 4925 3645 4935 3675
rect 4965 3645 4975 3675
rect 4925 3635 4975 3645
rect 5430 2050 5475 2055
rect 5430 2015 5435 2050
rect 5470 2015 5475 2050
rect 5430 2010 5475 2015
rect 4650 665 5015 685
rect 9540 680 9595 685
rect 9540 635 9545 680
rect 9590 635 9595 680
rect 9540 630 9595 635
<< via2 >>
rect 4935 3645 4965 3675
rect 5435 2015 5470 2050
rect 9545 675 9590 680
rect 9545 640 9550 675
rect 9550 640 9585 675
rect 9585 640 9590 675
rect 9545 635 9590 640
<< metal3 >>
rect 4925 3680 4975 3685
rect 4925 3640 4930 3680
rect 4970 3640 4975 3680
rect 4925 3635 4975 3640
rect 4865 2750 4915 2755
rect 4865 2710 4870 2750
rect 4910 2730 4915 2750
rect 4910 2710 9595 2730
rect 4865 2690 9595 2710
rect 5425 2055 5480 2060
rect 5425 2010 5430 2055
rect 5475 2010 5480 2055
rect 5425 2005 5480 2010
rect 9540 690 9590 2690
rect 9535 680 9600 690
rect 9535 635 9545 680
rect 9590 635 9600 680
rect 9535 625 9600 635
<< via3 >>
rect 4930 3675 4970 3680
rect 4930 3645 4935 3675
rect 4935 3645 4965 3675
rect 4965 3645 4970 3675
rect 4930 3640 4970 3645
rect 4870 2710 4910 2750
rect 5430 2050 5475 2055
rect 5430 2015 5435 2050
rect 5435 2015 5470 2050
rect 5470 2015 5475 2050
rect 5430 2010 5475 2015
<< metal4 >>
rect 4870 3680 4980 3690
rect 4870 3640 4930 3680
rect 4970 3640 4980 3680
rect 4870 3630 4980 3640
rect 4870 2760 4900 3630
rect 4860 2750 4920 2760
rect 4860 2710 4870 2750
rect 4910 2710 4920 2750
rect 4860 2700 4920 2710
rect 5430 2110 5490 2150
rect 5430 2060 5465 2110
rect 5425 2055 5480 2060
rect 5425 2010 5430 2055
rect 5475 2010 5480 2055
rect 5425 2005 5480 2010
use divbuf  divbuf_0
timestamp 1640990631
transform 1 0 5155 0 1 3655
box -460 -1085 31200 495
use divider  divider_0
timestamp 1640980777
transform 1 0 5185 0 1 235
box -490 -235 4690 2150
use ro_complete  ro_complete_0
timestamp 1640997741
transform 1 0 57 0 1 5330
box -57 -5330 4455 1440
<< end >>
