magic
tech sky130A
timestamp 1640957225
<< nwell >>
rect -85 -15 335 475
<< nmos >>
rect -10 -335 5 -135
rect 115 -335 130 -135
rect 240 -335 255 -185
<< pmos >>
rect -10 10 5 270
rect 115 10 130 270
rect 240 10 255 390
<< ndiff >>
rect -50 -165 -10 -135
rect -50 -190 -45 -165
rect -20 -190 -10 -165
rect -50 -210 -10 -190
rect -50 -235 -45 -210
rect -20 -235 -10 -210
rect -50 -255 -10 -235
rect -50 -280 -45 -255
rect -20 -280 -10 -255
rect -50 -300 -10 -280
rect -50 -325 -45 -300
rect -20 -325 -10 -300
rect -50 -335 -10 -325
rect 5 -165 45 -135
rect 5 -190 15 -165
rect 40 -190 45 -165
rect 5 -210 45 -190
rect 5 -235 15 -210
rect 40 -235 45 -210
rect 5 -255 45 -235
rect 5 -280 15 -255
rect 40 -280 45 -255
rect 5 -300 45 -280
rect 5 -325 15 -300
rect 40 -325 45 -300
rect 5 -335 45 -325
rect 75 -165 115 -135
rect 75 -190 80 -165
rect 105 -190 115 -165
rect 75 -210 115 -190
rect 75 -235 80 -210
rect 105 -235 115 -210
rect 75 -255 115 -235
rect 75 -280 80 -255
rect 105 -280 115 -255
rect 75 -300 115 -280
rect 75 -325 80 -300
rect 105 -325 115 -300
rect 75 -335 115 -325
rect 130 -165 170 -135
rect 130 -190 140 -165
rect 165 -190 170 -165
rect 130 -210 170 -190
rect 130 -235 140 -210
rect 165 -235 170 -210
rect 130 -255 170 -235
rect 130 -280 140 -255
rect 165 -280 170 -255
rect 130 -300 170 -280
rect 130 -325 140 -300
rect 165 -325 170 -300
rect 130 -335 170 -325
rect 200 -210 240 -185
rect 200 -235 205 -210
rect 230 -235 240 -210
rect 200 -255 240 -235
rect 200 -280 205 -255
rect 230 -280 240 -255
rect 200 -300 240 -280
rect 200 -325 205 -300
rect 230 -325 240 -300
rect 200 -335 240 -325
rect 255 -210 295 -185
rect 255 -235 265 -210
rect 290 -235 295 -210
rect 255 -255 295 -235
rect 255 -280 265 -255
rect 290 -280 295 -255
rect 255 -300 295 -280
rect 255 -325 265 -300
rect 290 -325 295 -300
rect 255 -335 295 -325
<< pdiff >>
rect 200 360 240 390
rect 200 335 205 360
rect 230 335 240 360
rect 200 315 240 335
rect 200 290 205 315
rect 230 290 240 315
rect 200 270 240 290
rect -50 225 -10 270
rect -50 200 -45 225
rect -20 200 -10 225
rect -50 180 -10 200
rect -50 155 -45 180
rect -20 155 -10 180
rect -50 135 -10 155
rect -50 110 -45 135
rect -20 110 -10 135
rect -50 90 -10 110
rect -50 65 -45 90
rect -20 65 -10 90
rect -50 45 -10 65
rect -50 20 -45 45
rect -20 20 -10 45
rect -50 10 -10 20
rect 5 225 45 270
rect 5 200 15 225
rect 40 200 45 225
rect 5 180 45 200
rect 5 155 15 180
rect 40 155 45 180
rect 5 135 45 155
rect 5 110 15 135
rect 40 110 45 135
rect 5 90 45 110
rect 5 65 15 90
rect 40 65 45 90
rect 5 45 45 65
rect 5 20 15 45
rect 40 20 45 45
rect 5 10 45 20
rect 75 225 115 270
rect 75 200 80 225
rect 105 200 115 225
rect 75 180 115 200
rect 75 155 80 180
rect 105 155 115 180
rect 75 135 115 155
rect 75 110 80 135
rect 105 110 115 135
rect 75 90 115 110
rect 75 65 80 90
rect 105 65 115 90
rect 75 45 115 65
rect 75 20 80 45
rect 105 20 115 45
rect 75 10 115 20
rect 130 225 170 270
rect 130 200 140 225
rect 165 200 170 225
rect 130 180 170 200
rect 130 155 140 180
rect 165 155 170 180
rect 130 135 170 155
rect 130 110 140 135
rect 165 110 170 135
rect 130 90 170 110
rect 130 65 140 90
rect 165 65 170 90
rect 130 45 170 65
rect 130 20 140 45
rect 165 20 170 45
rect 130 10 170 20
rect 200 245 205 270
rect 230 245 240 270
rect 200 225 240 245
rect 200 200 205 225
rect 230 200 240 225
rect 200 180 240 200
rect 200 155 205 180
rect 230 155 240 180
rect 200 135 240 155
rect 200 110 205 135
rect 230 110 240 135
rect 200 90 240 110
rect 200 65 205 90
rect 230 65 240 90
rect 200 45 240 65
rect 200 20 205 45
rect 230 20 240 45
rect 200 10 240 20
rect 255 360 295 390
rect 255 335 265 360
rect 290 335 295 360
rect 255 315 295 335
rect 255 290 265 315
rect 290 290 295 315
rect 255 270 295 290
rect 255 245 265 270
rect 290 245 295 270
rect 255 225 295 245
rect 255 200 265 225
rect 290 200 295 225
rect 255 180 295 200
rect 255 155 265 180
rect 290 155 295 180
rect 255 135 295 155
rect 255 110 265 135
rect 290 110 295 135
rect 255 90 295 110
rect 255 65 265 90
rect 290 65 295 90
rect 255 45 295 65
rect 255 20 265 45
rect 290 20 295 45
rect 255 10 295 20
<< ndiffc >>
rect -45 -190 -20 -165
rect -45 -235 -20 -210
rect -45 -280 -20 -255
rect -45 -325 -20 -300
rect 15 -190 40 -165
rect 15 -235 40 -210
rect 15 -280 40 -255
rect 15 -325 40 -300
rect 80 -190 105 -165
rect 80 -235 105 -210
rect 80 -280 105 -255
rect 80 -325 105 -300
rect 140 -190 165 -165
rect 140 -235 165 -210
rect 140 -280 165 -255
rect 140 -325 165 -300
rect 205 -235 230 -210
rect 205 -280 230 -255
rect 205 -325 230 -300
rect 265 -235 290 -210
rect 265 -280 290 -255
rect 265 -325 290 -300
<< pdiffc >>
rect 205 335 230 360
rect 205 290 230 315
rect -45 200 -20 225
rect -45 155 -20 180
rect -45 110 -20 135
rect -45 65 -20 90
rect -45 20 -20 45
rect 15 200 40 225
rect 15 155 40 180
rect 15 110 40 135
rect 15 65 40 90
rect 15 20 40 45
rect 80 200 105 225
rect 80 155 105 180
rect 80 110 105 135
rect 80 65 105 90
rect 80 20 105 45
rect 140 200 165 225
rect 140 155 165 180
rect 140 110 165 135
rect 140 65 165 90
rect 140 20 165 45
rect 205 245 230 270
rect 205 200 230 225
rect 205 155 230 180
rect 205 110 230 135
rect 205 65 230 90
rect 205 20 230 45
rect 265 335 290 360
rect 265 290 290 315
rect 265 245 290 270
rect 265 200 290 225
rect 265 155 290 180
rect 265 110 290 135
rect 265 65 290 90
rect 265 20 290 45
<< poly >>
rect 240 390 255 410
rect -10 270 5 295
rect 115 270 130 295
rect -10 -75 5 10
rect 115 -75 130 10
rect -50 -85 5 -75
rect -50 -105 -40 -85
rect -20 -105 5 -85
rect -50 -115 5 -105
rect 75 -85 130 -75
rect 240 -80 255 10
rect 75 -105 85 -85
rect 105 -105 130 -85
rect 75 -115 130 -105
rect -10 -135 5 -115
rect 115 -135 130 -115
rect 200 -90 255 -80
rect 200 -110 210 -90
rect 230 -110 255 -90
rect 200 -120 255 -110
rect 240 -185 255 -120
rect -10 -370 5 -335
rect 115 -370 130 -335
rect 240 -370 255 -335
<< polycont >>
rect -40 -105 -20 -85
rect 85 -105 105 -85
rect 210 -110 230 -90
<< locali >>
rect 200 440 205 460
rect 225 440 230 460
rect 200 425 230 440
rect 205 390 230 425
rect 200 360 235 390
rect -45 325 -40 345
rect -45 270 -20 325
rect 75 325 80 345
rect 100 325 105 345
rect 75 310 105 325
rect 80 270 105 310
rect 200 335 205 360
rect 230 335 235 360
rect 200 315 235 335
rect 200 290 205 315
rect 230 290 235 315
rect 200 270 235 290
rect -50 225 -15 270
rect -50 200 -45 225
rect -20 200 -15 225
rect -50 180 -15 200
rect -50 155 -45 180
rect -20 155 -15 180
rect -50 135 -15 155
rect -50 110 -45 135
rect -20 110 -15 135
rect -50 90 -15 110
rect -50 65 -45 90
rect -20 65 -15 90
rect -50 45 -15 65
rect -50 20 -45 45
rect -20 20 -15 45
rect -50 10 -15 20
rect 10 225 45 270
rect 10 200 15 225
rect 40 200 45 225
rect 10 180 45 200
rect 10 155 15 180
rect 40 155 45 180
rect 10 135 45 155
rect 10 110 15 135
rect 40 110 45 135
rect 10 90 45 110
rect 10 65 15 90
rect 40 65 45 90
rect 10 45 45 65
rect 10 20 15 45
rect 40 20 45 45
rect 10 10 45 20
rect 75 225 110 270
rect 75 200 80 225
rect 105 200 110 225
rect 75 180 110 200
rect 75 155 80 180
rect 105 155 110 180
rect 75 135 110 155
rect 75 110 80 135
rect 105 110 110 135
rect 75 90 110 110
rect 75 65 80 90
rect 105 65 110 90
rect 75 45 110 65
rect 75 20 80 45
rect 105 20 110 45
rect 75 10 110 20
rect 135 225 170 270
rect 135 200 140 225
rect 165 200 170 225
rect 135 180 170 200
rect 135 155 140 180
rect 165 155 170 180
rect 135 135 170 155
rect 135 110 140 135
rect 165 110 170 135
rect 135 90 170 110
rect 135 65 140 90
rect 165 65 170 90
rect 135 45 170 65
rect 135 20 140 45
rect 165 20 170 45
rect 135 10 170 20
rect 200 245 205 270
rect 230 245 235 270
rect 200 225 235 245
rect 200 200 205 225
rect 230 200 235 225
rect 200 180 235 200
rect 200 155 205 180
rect 230 155 235 180
rect 200 135 235 155
rect 200 110 205 135
rect 230 110 235 135
rect 200 90 235 110
rect 200 65 205 90
rect 230 65 235 90
rect 200 45 235 65
rect 200 20 205 45
rect 230 20 235 45
rect 200 10 235 20
rect 260 360 295 390
rect 260 335 265 360
rect 290 335 295 360
rect 260 315 295 335
rect 260 290 265 315
rect 290 290 295 315
rect 260 270 295 290
rect 260 245 265 270
rect 290 245 295 270
rect 260 225 295 245
rect 260 200 265 225
rect 290 200 295 225
rect 260 180 295 200
rect 260 155 265 180
rect 290 155 295 180
rect 260 135 295 155
rect 260 110 265 135
rect 290 110 295 135
rect 260 90 295 110
rect 260 65 265 90
rect 290 65 295 90
rect 260 45 295 65
rect 260 20 265 45
rect 290 20 295 45
rect 260 10 295 20
rect 15 -10 40 10
rect 140 -10 165 10
rect 15 -30 165 -10
rect -50 -85 -10 -75
rect 75 -85 115 -75
rect -85 -105 -40 -85
rect -20 -105 -10 -85
rect 65 -105 85 -85
rect 105 -105 115 -85
rect -50 -115 -10 -105
rect 75 -115 115 -105
rect 140 -90 165 -30
rect 200 -90 240 -80
rect 140 -110 210 -90
rect 230 -110 240 -90
rect 140 -135 165 -110
rect 200 -120 240 -110
rect 265 -95 290 10
rect 265 -120 335 -95
rect -50 -165 -15 -135
rect -50 -190 -45 -165
rect -20 -190 -15 -165
rect -50 -210 -15 -190
rect -50 -235 -45 -210
rect -20 -235 -15 -210
rect -50 -255 -15 -235
rect -50 -280 -45 -255
rect -20 -280 -15 -255
rect -50 -300 -15 -280
rect -50 -325 -45 -300
rect -20 -325 -15 -300
rect -50 -335 -15 -325
rect 10 -165 45 -135
rect 10 -190 15 -165
rect 40 -190 45 -165
rect 10 -210 45 -190
rect 75 -165 110 -135
rect 75 -190 80 -165
rect 105 -190 110 -165
rect 75 -210 110 -190
rect 10 -235 15 -210
rect 40 -235 80 -210
rect 105 -235 110 -210
rect 10 -255 45 -235
rect 10 -280 15 -255
rect 40 -280 45 -255
rect 10 -300 45 -280
rect 10 -325 15 -300
rect 40 -325 45 -300
rect 10 -335 45 -325
rect 75 -255 110 -235
rect 75 -280 80 -255
rect 105 -280 110 -255
rect 75 -300 110 -280
rect 75 -325 80 -300
rect 105 -325 110 -300
rect 75 -335 110 -325
rect 135 -165 170 -135
rect 135 -190 140 -165
rect 165 -190 170 -165
rect 265 -185 290 -120
rect 135 -210 170 -190
rect 135 -235 140 -210
rect 165 -235 170 -210
rect 135 -255 170 -235
rect 135 -280 140 -255
rect 165 -280 170 -255
rect 135 -300 170 -280
rect 135 -325 140 -300
rect 165 -325 170 -300
rect 135 -335 170 -325
rect 200 -210 235 -185
rect 200 -235 205 -210
rect 230 -235 235 -210
rect 200 -255 235 -235
rect 200 -280 205 -255
rect 230 -280 235 -255
rect 200 -300 235 -280
rect 200 -325 205 -300
rect 230 -325 235 -300
rect 200 -335 235 -325
rect 260 -210 295 -185
rect 260 -235 265 -210
rect 290 -235 295 -210
rect 260 -255 295 -235
rect 260 -280 265 -255
rect 290 -280 295 -255
rect 260 -300 295 -280
rect 260 -325 265 -300
rect 290 -325 295 -300
rect 260 -335 295 -325
rect -45 -395 -20 -335
rect 205 -375 230 -335
rect -25 -415 -20 -395
rect 200 -395 225 -375
rect 200 -415 205 -395
<< viali >>
rect 205 440 225 460
rect -40 325 -20 345
rect 80 325 100 345
rect 45 -105 65 -85
rect -45 -415 -25 -395
rect 205 -415 225 -395
<< metal1 >>
rect 195 465 235 470
rect 195 435 200 465
rect 230 435 235 465
rect 195 430 235 435
rect -50 350 -10 355
rect -50 320 -45 350
rect -15 320 -10 350
rect -50 315 -10 320
rect 70 350 110 355
rect 70 320 75 350
rect 105 320 110 350
rect 70 315 110 320
rect -85 -60 60 -45
rect 45 -75 60 -60
rect 35 -85 75 -75
rect 35 -105 45 -85
rect 65 -105 75 -85
rect 35 -115 75 -105
rect -55 -390 -15 -385
rect -55 -420 -50 -390
rect -20 -420 -15 -390
rect -55 -425 -15 -420
rect 195 -390 235 -385
rect 195 -420 200 -390
rect 230 -420 235 -390
rect 195 -425 235 -420
<< via1 >>
rect 200 460 230 465
rect 200 440 205 460
rect 205 440 225 460
rect 225 440 230 460
rect 200 435 230 440
rect -45 345 -15 350
rect -45 325 -40 345
rect -40 325 -20 345
rect -20 325 -15 345
rect -45 320 -15 325
rect 75 345 105 350
rect 75 325 80 345
rect 80 325 100 345
rect 100 325 105 345
rect 75 320 105 325
rect -50 -395 -20 -390
rect -50 -415 -45 -395
rect -45 -415 -25 -395
rect -25 -415 -20 -395
rect -50 -420 -20 -415
rect 200 -395 230 -390
rect 200 -415 205 -395
rect 205 -415 225 -395
rect 225 -415 230 -395
rect 200 -420 230 -415
<< metal2 >>
rect 190 470 240 475
rect 190 430 195 470
rect 235 430 240 470
rect 190 425 240 430
rect -55 355 -5 360
rect -55 315 -50 355
rect -10 315 -5 355
rect -55 310 -5 315
rect 65 355 115 360
rect 65 315 70 355
rect 110 315 115 355
rect 65 310 115 315
rect -60 -385 -10 -380
rect -60 -425 -55 -385
rect -15 -425 -10 -385
rect -60 -430 -10 -425
rect 190 -385 240 -380
rect 190 -425 195 -385
rect 235 -425 240 -385
rect 190 -430 240 -425
<< via2 >>
rect 195 465 235 470
rect 195 435 200 465
rect 200 435 230 465
rect 230 435 235 465
rect 195 430 235 435
rect -50 350 -10 355
rect -50 320 -45 350
rect -45 320 -15 350
rect -15 320 -10 350
rect -50 315 -10 320
rect 70 350 110 355
rect 70 320 75 350
rect 75 320 105 350
rect 105 320 110 350
rect 70 315 110 320
rect -55 -390 -15 -385
rect -55 -420 -50 -390
rect -50 -420 -20 -390
rect -20 -420 -15 -390
rect -55 -425 -15 -420
rect 195 -390 235 -385
rect 195 -420 200 -390
rect 200 -420 230 -390
rect 230 -420 235 -390
rect 195 -425 235 -420
<< metal3 >>
rect 190 470 240 475
rect 190 430 195 470
rect 235 430 240 470
rect 190 425 240 430
rect -55 355 -5 360
rect -55 315 -50 355
rect -10 315 -5 355
rect -55 310 -5 315
rect 65 355 115 360
rect 65 315 70 355
rect 110 315 115 355
rect 65 310 115 315
rect -65 -380 -5 -375
rect -65 -430 -60 -380
rect -10 -430 -5 -380
rect -65 -435 -5 -430
rect 185 -380 245 -375
rect 185 -430 190 -380
rect 240 -430 245 -380
rect 185 -435 245 -430
<< via3 >>
rect 195 430 235 470
rect -50 315 -10 355
rect 70 315 110 355
rect -60 -385 -10 -380
rect -60 -425 -55 -385
rect -55 -425 -15 -385
rect -15 -425 -10 -385
rect -60 -430 -10 -425
rect 190 -385 240 -380
rect 190 -425 195 -385
rect 195 -425 235 -385
rect 235 -425 240 -385
rect 190 -430 240 -425
<< metal4 >>
rect 190 470 240 475
rect -85 440 195 470
rect -45 360 -15 440
rect 75 360 105 440
rect 190 430 195 440
rect 235 440 335 470
rect 235 430 240 440
rect 190 425 240 430
rect -55 355 -5 360
rect -55 315 -50 355
rect -10 315 -5 355
rect -55 310 -5 315
rect 65 355 115 360
rect 65 315 70 355
rect 110 315 115 355
rect 65 310 115 315
rect -65 -380 -5 -375
rect -65 -430 -60 -380
rect -10 -385 -5 -380
rect 185 -380 245 -375
rect 185 -385 190 -380
rect -10 -420 190 -385
rect -10 -430 -5 -420
rect -65 -435 -5 -430
rect 185 -430 190 -420
rect 240 -385 245 -380
rect 240 -420 295 -385
rect 240 -430 245 -420
rect 185 -435 245 -430
<< labels >>
rlabel metal4 -55 -420 295 -385 1 GND
rlabel nwell -85 440 335 470 1 VDD
rlabel locali 265 -120 335 -95 1 OUT
rlabel locali -85 -105 -20 -85 1 A
rlabel metal1 -85 -60 60 -45 1 B
rlabel metal1 45 -105 60 -60 1 B
rlabel locali 45 -105 105 -85 1 B
rlabel locali 15 -235 105 -210 1 Z1
rlabel locali 140 -110 230 -90 1 out1
rlabel locali 219 -363 219 -363 1 gnd!
rlabel locali 214 405 214 405 1 vdd!
<< end >>
