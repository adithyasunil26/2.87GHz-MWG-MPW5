magic
tech sky130A
magscale 1 2
timestamp 1647892250
<< locali >>
rect -1330 15702 -928 15778
rect -1330 15440 -1270 15702
rect -1008 15440 -928 15702
rect -1330 15380 -928 15440
rect -332 13768 -18 13796
rect -332 13528 -300 13768
rect -48 13528 -18 13768
rect -332 13502 -18 13528
rect 2892 -60 2996 2750
rect 3862 0 3966 2718
rect 4852 186 4956 2802
rect 2880 -222 3000 -60
rect 2772 -238 3000 -222
rect -4346 -490 3000 -238
rect -4346 -498 2990 -490
rect -4346 -18236 -4128 -498
rect 2772 -500 2990 -498
rect 3854 -670 3966 0
rect 4842 -116 4956 186
rect -3738 -672 3974 -670
rect -3852 -862 3974 -672
rect -3852 -3954 -3678 -862
rect -3404 -1024 -3152 -1004
rect 4842 -1024 4948 -116
rect 5802 -124 5906 2730
rect 6792 -68 6896 2740
rect 7998 380 8102 2874
rect -3404 -1192 4958 -1024
rect -3868 -16426 -3660 -3954
rect -3404 -13796 -3152 -1192
rect -2900 -1330 -2478 -1322
rect 5790 -1330 5906 -124
rect -2900 -1350 5926 -1330
rect -2904 -1540 5926 -1350
rect -2904 -1544 2400 -1540
rect -2904 -1562 -2478 -1544
rect -2904 -10638 -2672 -1562
rect -2412 -1760 -2244 -1754
rect -2412 -1770 5984 -1760
rect 6790 -1770 6910 -68
rect -2412 -1926 6910 -1770
rect -2412 -1936 6906 -1926
rect -2412 -2910 -2244 -1936
rect 7996 -2078 8110 380
rect -2426 -2990 -2244 -2910
rect -2024 -2088 -1874 -2080
rect -288 -2088 8120 -2078
rect -2024 -2274 8120 -2088
rect -2024 -2294 -226 -2274
rect -2426 -6404 -2248 -2990
rect -2024 -4064 -1874 -2294
rect -2024 -4116 -1464 -4064
rect -2024 -4324 -1744 -4116
rect -1500 -4324 -1464 -4116
rect -2024 -4360 -1464 -4324
rect -2426 -7296 -2250 -6404
rect -2426 -7326 -1436 -7296
rect -2426 -7556 -1760 -7326
rect -1532 -7556 -1436 -7326
rect -2426 -7592 -1436 -7556
rect -1796 -7604 -1498 -7592
rect -2916 -10686 -1724 -10638
rect -2916 -10924 -2412 -10686
rect -2162 -10924 -1724 -10686
rect -2916 -10966 -1724 -10924
rect -3404 -13870 -1514 -13796
rect -3404 -14130 -2272 -13870
rect -1988 -14130 -1514 -13870
rect -3404 -14186 -1514 -14130
rect -3868 -17416 -3648 -16426
rect -3868 -17470 -1754 -17416
rect -3868 -17684 -2602 -17470
rect -2366 -17684 -1754 -17470
rect -3868 -17740 -1754 -17684
rect -4356 -18450 -4128 -18236
rect -4356 -20614 -4136 -18450
rect -2910 -20614 -2472 -20592
rect -4366 -20646 -2166 -20614
rect -4366 -20986 -2866 -20646
rect -2526 -20986 -2166 -20646
rect -4366 -21018 -2166 -20986
rect -2910 -21030 -2472 -21018
<< viali >>
rect -1270 15440 -1008 15702
rect -300 13528 -48 13768
rect 1450 13590 1580 13712
rect 66 6308 274 6500
rect -1744 -4324 -1500 -4116
rect -1760 -7556 -1532 -7326
rect -2412 -10924 -2162 -10686
rect -2272 -14130 -1988 -13870
rect -2602 -17684 -2366 -17470
rect -2866 -20986 -2526 -20646
<< metal1 >>
rect -1330 15702 -928 15778
rect -1330 15440 -1270 15702
rect -1008 15440 -928 15702
rect -1330 15380 -928 15440
rect -1256 12298 -1056 15380
rect -332 13782 -18 13796
rect 1274 13782 1626 13796
rect -332 13768 1626 13782
rect -332 13528 -300 13768
rect -48 13712 1626 13768
rect -48 13590 1450 13712
rect 1580 13590 1626 13712
rect -48 13528 1626 13590
rect -332 13516 1626 13528
rect -332 13502 -18 13516
rect 1274 13512 1626 13516
rect -1256 12228 -1008 12298
rect 366 12228 1912 12232
rect -1256 12044 1912 12228
rect -1256 12032 478 12044
rect -1256 12030 256 12032
rect 28 6500 312 6560
rect 28 6308 66 6500
rect 274 6308 312 6500
rect 28 6244 312 6308
rect -1780 -4116 -1438 -4060
rect -1780 -4324 -1744 -4116
rect -1500 -4324 -1438 -4116
rect -1780 -4372 -1438 -4324
rect -1796 -7326 -1498 -7296
rect -1796 -7556 -1760 -7326
rect -1532 -7556 -1498 -7326
rect -1796 -7604 -1498 -7556
rect -2468 -10686 -2100 -10644
rect -2468 -10924 -2412 -10686
rect -2162 -10924 -2100 -10686
rect -2468 -10960 -2100 -10924
rect -2314 -13870 -1946 -13820
rect -2314 -14130 -2272 -13870
rect -1988 -14130 -1946 -13870
rect -2314 -14172 -1946 -14130
rect -2640 -17470 -2322 -17424
rect -2640 -17684 -2602 -17470
rect -2366 -17684 -2322 -17470
rect -2640 -17732 -2322 -17684
rect -2910 -20646 -2472 -20592
rect -2910 -20986 -2866 -20646
rect -2526 -20986 -2472 -20646
rect -2910 -21030 -2472 -20986
<< via1 >>
rect -1270 15440 -1008 15702
rect -300 13528 -48 13768
rect 66 6308 274 6500
rect -1744 -4324 -1500 -4116
rect -1760 -7556 -1532 -7326
rect -2412 -10924 -2162 -10686
rect -2272 -14130 -1988 -13870
rect -2602 -17684 -2366 -17470
rect -2866 -20986 -2526 -20646
<< metal2 >>
rect -2714 19876 -2426 19878
rect -2714 19744 -702 19876
rect -2714 14738 -2426 19744
rect -1330 15702 -928 15778
rect -1330 15440 -1270 15702
rect -1008 15440 -928 15702
rect -1330 15380 -928 15440
rect -1708 14738 8948 14744
rect -2714 14456 8948 14738
rect -2714 14446 3650 14456
rect -2714 14440 -1530 14446
rect -332 13768 -18 13796
rect -332 13528 -300 13768
rect -48 13528 -18 13768
rect -332 13502 -18 13528
rect 8698 12686 8938 14456
rect 28 6500 312 6560
rect 28 6308 66 6500
rect 274 6308 312 6500
rect 28 6244 312 6308
rect -1780 -4116 -1438 -4060
rect -1780 -4324 -1744 -4116
rect -1500 -4324 -1438 -4116
rect -1780 -4372 -1438 -4324
rect -1796 -7326 -1498 -7296
rect -1796 -7556 -1760 -7326
rect -1532 -7556 -1498 -7326
rect -1796 -7604 -1498 -7556
rect -2468 -10686 -2100 -10644
rect -2468 -10924 -2412 -10686
rect -2162 -10924 -2100 -10686
rect -2468 -10960 -2100 -10924
rect -2314 -13870 -1946 -13820
rect -2314 -14130 -2272 -13870
rect -1988 -14130 -1946 -13870
rect -2314 -14172 -1946 -14130
rect -2640 -17470 -2322 -17424
rect -2640 -17684 -2602 -17470
rect -2366 -17684 -2322 -17470
rect -2640 -17732 -2322 -17684
rect -2910 -20646 -2472 -20592
rect -2910 -20986 -2866 -20646
rect -2526 -20986 -2472 -20646
rect -2910 -21030 -2472 -20986
<< via2 >>
rect -1270 15440 -1008 15702
rect -300 13528 -48 13768
rect 66 6308 274 6500
rect -1744 -4324 -1500 -4116
rect -1760 -7556 -1532 -7326
rect -2412 -10924 -2162 -10686
rect -2272 -14130 -1988 -13870
rect -2602 -17684 -2366 -17470
rect -2866 -20986 -2526 -20646
<< metal3 >>
rect -1330 15702 -928 15778
rect -1330 15440 -1270 15702
rect -1008 15440 -928 15702
rect -1330 15380 -928 15440
rect -332 13768 -18 13796
rect -332 13528 -300 13768
rect -48 13528 -18 13768
rect -332 13502 -18 13528
rect 28 6500 312 6560
rect 28 6308 66 6500
rect 274 6308 312 6500
rect 28 6244 312 6308
rect -1780 -4116 -1438 -4060
rect -1780 -4324 -1744 -4116
rect -1500 -4324 -1438 -4116
rect -1780 -4372 -1438 -4324
rect -1796 -7326 -1498 -7296
rect -1796 -7556 -1760 -7326
rect -1532 -7556 -1498 -7326
rect -1796 -7604 -1498 -7556
rect -2468 -10686 -2100 -10644
rect -2468 -10924 -2412 -10686
rect -2162 -10924 -2100 -10686
rect -2468 -10960 -2100 -10924
rect -2314 -13870 -1946 -13820
rect -2314 -14130 -2272 -13870
rect -1988 -14130 -1946 -13870
rect -2314 -14172 -1946 -14130
rect -2640 -17470 -2322 -17424
rect -2640 -17684 -2602 -17470
rect -2366 -17684 -2322 -17470
rect -2640 -17732 -2322 -17684
rect -2910 -20646 -2472 -20592
rect -2910 -20986 -2866 -20646
rect -2526 -20986 -2472 -20646
rect -2910 -21030 -2472 -20986
<< via3 >>
rect -1270 15440 -1008 15702
rect -300 13528 -48 13768
rect 66 6308 274 6500
rect -1744 -4324 -1500 -4116
rect -1760 -7556 -1532 -7326
rect -2412 -10924 -2162 -10686
rect -2272 -14130 -1988 -13870
rect -2602 -17684 -2366 -17470
rect -2866 -20986 -2526 -20646
<< metal4 >>
rect -5924 19302 -138 19582
rect -5924 16298 -5304 19302
rect -1404 16298 -834 16304
rect -5924 16018 -128 16298
rect -5924 6740 -5304 16018
rect -1404 16006 -834 16018
rect -1330 15718 -928 15778
rect -1330 15702 -648 15718
rect -1330 15440 -1270 15702
rect -1008 15456 -648 15702
rect -1008 15440 -928 15456
rect -1330 15380 -928 15440
rect -332 13768 -18 13796
rect -332 13528 -300 13768
rect -48 13528 -18 13768
rect -332 13502 -18 13528
rect -5924 6500 334 6740
rect -5924 6308 66 6500
rect 274 6308 334 6500
rect -5924 6074 334 6308
rect -5924 -3498 -5304 6074
rect -5924 -3760 -728 -3498
rect -5924 -6734 -5304 -3760
rect -1874 -4116 -1308 -4028
rect -1874 -4324 -1744 -4116
rect -1500 -4324 -1308 -4116
rect -1874 -4376 -1308 -4324
rect -2610 -6734 -2426 -6722
rect -5924 -6996 -2426 -6734
rect -5924 -10040 -5304 -6996
rect -2610 -7004 -2426 -6996
rect -2250 -6734 -2004 -6722
rect -2250 -6996 -680 -6734
rect -2250 -7004 -2004 -6996
rect -1900 -7326 -1286 -7290
rect -1900 -7556 -1760 -7326
rect -1532 -7556 -1286 -7326
rect -1900 -7598 -1286 -7556
rect -1796 -7604 -1498 -7598
rect -5924 -10302 -900 -10040
rect -5924 -13292 -5304 -10302
rect -2676 -10686 -1426 -10638
rect -2676 -10924 -2412 -10686
rect -2162 -10924 -1426 -10686
rect -2676 -10966 -1426 -10924
rect -5924 -13554 -824 -13292
rect -5924 -16852 -5304 -13554
rect -2766 -13870 -1344 -13776
rect -2766 -14130 -2272 -13870
rect -1988 -14130 -1344 -13870
rect -2766 -14206 -1344 -14130
rect -5924 -17114 -970 -16852
rect -5924 -20088 -5304 -17114
rect -3326 -17470 -1688 -17384
rect -3326 -17684 -2602 -17470
rect -2366 -17684 -1688 -17470
rect -3326 -17760 -1688 -17684
rect -5924 -20348 -942 -20088
rect -5054 -20350 -942 -20348
rect -3152 -20646 -1542 -20592
rect -3152 -20986 -2866 -20646
rect -2526 -20986 -1542 -20646
rect -3152 -21008 -1542 -20986
rect -2910 -21030 -2472 -21008
<< via4 >>
rect -300 13528 -48 13768
<< metal5 >>
rect -444 17258 46 17998
rect -372 14164 60 14948
rect -418 13768 66 14164
rect -418 13528 -300 13768
rect -48 13528 66 13768
rect -418 13096 66 13528
rect -1220 12634 66 13096
rect -1212 438 -726 12634
rect -1210 122 -734 438
rect -1210 -58 -738 122
rect -1212 -2524 -738 -58
rect -1212 -3030 -1110 -2524
rect -1212 -5040 -726 -5012
rect -1212 -5754 -636 -5040
rect -1212 -6232 -992 -5754
rect -1222 -8206 -1038 -8046
rect -1284 -9104 -676 -8206
rect -1310 -11986 -720 -11610
rect -1370 -12322 -720 -11986
rect -1370 -12790 -1150 -12322
rect -1406 -15360 -762 -14838
rect -1474 -15882 -762 -15360
rect -1474 -16164 -1254 -15882
rect -1432 -18392 -1192 -18378
rect -1432 -18848 -898 -18392
rect -1422 -19118 -898 -18848
rect -1422 -19400 -1202 -19118
use tapered_buf  tapered_buf_3
timestamp 1647889165
transform 1 0 -512 0 1 -6542
box -940 -1820 87350 802
use tapered_buf  tapered_buf_4
timestamp 1647889165
transform 1 0 -750 0 1 -9858
box -940 -1820 87350 802
use tapered_buf  tapered_buf_5
timestamp 1647889165
transform 1 0 -670 0 1 -13096
box -940 -1820 87350 802
use tapered_buf  tapered_buf_6
timestamp 1647889165
transform 1 0 -828 0 1 -16658
box -940 -1820 87350 802
use tapered_buf  tapered_buf_7
timestamp 1647889165
transform 1 0 -748 0 1 -19896
box -940 -1820 87350 802
use ro_complete  ro_complete_0
timestamp 1647892250
transform 1 0 696 0 1 11380
box -696 -11380 9322 2880
use tapered_buf  tapered_buf_2
timestamp 1647889165
transform 1 0 -592 0 1 -3304
box -940 -1820 87350 802
use DIGITAL_BUFFER_v1  DIGITAL_BUFFER_v1_0
timestamp 1647892099
transform 1 0 120 0 1 19734
box -940 -1820 87350 1165
use tapered_buf  tapered_buf_0
timestamp 1647889165
transform 1 0 200 0 1 16504
box -940 -1820 87350 802
<< labels >>
rlabel space -224 20520 -224 20520 1 vdd!
rlabel space -648 16568 -648 16568 1 vcont
rlabel space -676 18818 -676 18818 1 out
rlabel metal4 -5688 6380 -5688 6380 1 gnd!
rlabel space -1638 -19806 -1638 -19806 1 a0
rlabel space -1708 -16560 -1708 -16560 1 a1
rlabel space -1558 -13010 -1558 -13010 1 a2
rlabel space -1596 -9786 -1596 -9786 1 a3
rlabel space -1402 -6462 -1402 -6462 1 a4
rlabel space -1456 -3212 -1456 -3212 1 a5
rlabel space -756 18842 -756 18842 1 out
<< end >>
