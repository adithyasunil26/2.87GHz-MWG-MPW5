magic
tech sky130A
timestamp 1647804540
<< locali >>
rect -458 708 70 709
rect -470 698 70 708
rect -470 594 -458 698
rect -351 594 70 698
rect -470 585 70 594
rect -470 584 -339 585
<< viali >>
rect -458 594 -351 698
<< metal1 >>
rect 2067 1141 2142 1146
rect 1676 1116 2142 1141
rect 1719 998 1745 999
rect 1666 979 1745 998
rect -470 698 -339 708
rect -470 594 -458 698
rect -351 594 -339 698
rect 1719 655 1745 979
rect -470 584 -339 594
rect 1688 61 1760 655
rect 1685 -94 1765 61
rect 2067 7 2142 1116
rect -520 -100 1765 -94
rect -525 -169 1765 -100
rect 2065 -161 2145 7
rect -525 -172 1757 -169
rect -525 -188 32 -172
rect -525 -2102 -380 -188
rect -60 -316 29 -314
rect 2062 -316 2151 -161
rect -60 -397 2151 -316
rect -60 -402 2140 -397
rect -60 -707 29 -402
rect -143 -742 50 -707
rect -143 -873 -108 -742
rect 13 -873 50 -742
rect -143 -897 50 -873
rect -542 -2128 -354 -2102
rect -542 -2252 -518 -2128
rect -384 -2252 -354 -2128
rect -542 -2273 -354 -2252
<< via1 >>
rect -458 594 -351 698
rect -108 -873 13 -742
rect -518 -2252 -384 -2128
<< metal2 >>
rect -271 3561 -120 3578
rect -271 3441 -260 3561
rect -137 3441 -120 3561
rect -271 3427 -120 3441
rect -470 698 -339 708
rect -470 594 -458 698
rect -351 594 -339 698
rect -470 584 -339 594
rect -231 344 -170 3427
rect -91 2196 22 2210
rect -91 2099 -81 2196
rect 13 2099 22 2196
rect -91 2085 22 2099
rect -65 1192 -18 2085
rect -68 1176 127 1192
rect -68 1175 48 1176
rect -65 1173 -18 1175
rect -231 322 130 344
rect -143 -742 50 -707
rect -143 -873 -108 -742
rect 13 -873 50 -742
rect -143 -897 50 -873
rect -542 -2128 -354 -2102
rect -542 -2252 -518 -2128
rect -384 -2150 -354 -2128
rect -384 -2244 56 -2150
rect -384 -2252 -354 -2244
rect -542 -2273 -354 -2252
<< via2 >>
rect -260 3441 -137 3561
rect -458 594 -351 698
rect -81 2099 13 2196
<< metal3 >>
rect -271 3561 -120 3578
rect -271 3441 -260 3561
rect -137 3441 -120 3561
rect -271 3427 -120 3441
rect -88 2196 22 2205
rect -88 2099 -81 2196
rect 13 2099 22 2196
rect -88 2093 22 2099
rect -470 698 -339 708
rect -470 594 -458 698
rect -351 594 -339 698
rect -470 584 -339 594
<< via3 >>
rect -260 3441 -137 3561
rect -81 2099 13 2196
rect -458 594 -351 698
<< metal4 >>
rect -926 3724 308 3859
rect -924 2510 -768 3724
rect -283 3561 70 3587
rect -283 3441 -260 3561
rect -137 3441 70 3561
rect -283 3425 70 3441
rect -924 2366 354 2510
rect -924 713 -768 2366
rect -91 2196 22 2210
rect -91 2099 -81 2196
rect 13 2099 22 2196
rect -91 2085 22 2099
rect -924 698 -329 713
rect -924 594 -458 698
rect -351 594 -329 698
rect -924 577 -329 594
rect -924 -959 -768 577
rect -924 -1134 329 -959
rect -924 -2333 -768 -1134
rect -947 -2508 293 -2333
<< metal5 >>
rect 186 2938 404 3142
rect 145 -1871 363 -1667
use pd  pd_0
timestamp 1647804088
transform 1 0 215 0 1 781
box -215 -855 1685 810
use tapered_buf  tapered_buf_2
timestamp 1647784636
transform 1 0 434 0 1 -881
box -470 -910 43675 400
use tapered_buf  tapered_buf_3
timestamp 1647784636
transform 1 0 429 0 1 -2234
box -470 -910 43675 400
use tapered_buf  tapered_buf_1
timestamp 1647784636
transform 1 0 473 0 1 3958
box -470 -910 43675 400
use tapered_buf  tapered_buf_0
timestamp 1647784636
transform 1 0 468 0 1 2605
box -470 -910 43675 400
<< labels >>
rlabel space 48 2642 48 2642 1 ref
rlabel space 64 3988 64 3988 1 div
rlabel space 40 -1345 40 -1345 1 up
rlabel space -14 -2692 -14 -2692 1 down
<< end >>
