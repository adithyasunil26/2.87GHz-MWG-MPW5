* SPICE3 file created from pd_buffered.ext - technology: sky130A

X0 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X10 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X12 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X14 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X17 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X18 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X19 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X24 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X25 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X26 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X27 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X28 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X30 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X33 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X34 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X35 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X38 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X40 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X43 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X44 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X46 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X47 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X49 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X50 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X51 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X52 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X53 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X54 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X55 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X56 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X57 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X59 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X60 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X61 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X62 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X63 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X64 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X65 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 vdd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X67 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X68 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X69 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X70 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X71 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X72 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X73 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X74 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X75 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X76 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X77 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X78 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X79 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X80 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X81 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X82 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X83 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X84 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X85 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X86 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X87 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X88 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X89 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X90 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X91 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X92 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X93 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X94 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X95 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X96 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X97 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X98 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X99 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X100 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X101 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X102 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X103 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X104 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X105 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X106 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X107 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X108 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X109 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X110 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X111 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X112 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X113 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X114 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X115 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X116 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X117 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X118 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X119 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X120 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X121 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X122 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X123 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X124 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X125 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X126 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X127 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X128 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X129 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X130 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X131 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X132 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X133 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X134 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X135 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X136 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X137 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X138 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X139 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X140 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X141 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X142 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X143 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X144 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X145 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X146 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X147 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X148 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X149 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X150 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X151 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X152 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X153 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X154 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X155 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X156 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X157 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X158 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X159 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X160 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X161 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X162 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X163 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X164 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X165 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X166 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X167 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X168 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X169 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X170 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X171 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X172 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X173 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X174 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X175 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X176 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X177 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X178 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X179 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X180 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X181 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X182 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X183 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X184 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X185 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X186 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X187 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X188 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X189 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X190 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X191 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X192 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X193 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X194 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X195 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X196 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X197 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X198 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X199 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X200 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X201 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X202 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X203 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X204 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X205 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X206 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X207 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X208 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X209 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X210 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X211 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X212 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X213 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X214 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X215 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X216 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X217 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X218 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X219 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X220 tapered_buf_2/a_160_230# pd_0/UP tapered_buf_2/a_n10_230# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X221 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X222 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X223 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X224 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X225 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X226 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X227 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X228 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X229 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X230 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X231 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X232 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X233 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X234 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X235 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X236 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X237 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X238 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X239 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X240 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X241 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X242 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X243 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X244 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X245 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X246 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X247 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X248 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X249 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X250 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X251 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X252 tapered_buf_2/a_580_0# tapered_buf_2/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X253 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X254 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X255 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X256 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X257 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X258 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X259 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X260 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X261 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X262 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X263 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X264 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X265 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X266 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X267 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X268 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X269 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X270 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X271 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X272 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X273 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X274 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X275 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X276 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X277 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X278 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X279 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X280 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X281 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X282 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X283 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X284 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X285 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X286 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X287 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X288 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X289 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X290 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X291 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X292 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X293 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X294 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X295 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X296 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X297 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X298 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X299 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X300 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X301 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X302 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X303 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X304 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X305 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X306 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X307 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X308 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X309 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X310 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X311 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X312 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X313 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X314 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X315 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X316 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X317 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X318 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X319 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X320 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X321 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X322 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X323 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X324 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X325 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X326 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X327 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X328 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X329 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X330 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X331 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X332 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X333 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X334 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X335 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X336 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X337 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X338 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X339 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X340 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X341 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X342 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X343 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X344 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X345 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X346 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X347 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X348 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X349 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X350 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X351 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X352 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X353 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X354 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X355 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X356 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X357 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X358 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X359 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X360 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X361 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X362 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X363 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X364 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X365 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X366 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X367 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X368 gnd tapered_buf_2/a_160_n140# tapered_buf_2/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X369 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X370 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X371 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X372 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X373 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X374 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X375 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X376 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X377 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X378 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X379 vdd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X380 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X381 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X382 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X383 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X384 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X385 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X386 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X387 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X388 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X389 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X390 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X391 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X392 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X393 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X394 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X395 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X396 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X397 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X398 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X399 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X400 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X401 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X402 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X403 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X404 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X405 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X406 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X407 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X408 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X409 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X410 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X411 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X412 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X413 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X414 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X415 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X416 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X417 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X418 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X419 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X420 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X421 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X422 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X423 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X424 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X425 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X426 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X427 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X428 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X429 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X430 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X431 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X432 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X433 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X434 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X435 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X436 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X437 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X438 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X439 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X440 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X441 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X442 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X443 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X444 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X445 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X446 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X447 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X448 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X449 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X450 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X451 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X452 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X453 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X454 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X455 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X456 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X457 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X458 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X459 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X460 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X461 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X462 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X463 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X464 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X465 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X466 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X467 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X468 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X469 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X470 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X471 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X472 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X473 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X474 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X475 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X476 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X477 gnd tapered_buf_2/a_160_n140# tapered_buf_2/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X478 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X479 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X480 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X481 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X482 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X483 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X484 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X485 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X486 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X487 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X488 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X489 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X490 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X491 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X492 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X493 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X494 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X495 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X496 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X497 vdd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X498 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X499 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X500 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X501 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X502 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X503 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X504 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X505 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X506 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X507 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X508 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X509 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X510 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X511 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X512 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X513 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X514 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X515 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X516 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X517 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X518 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X519 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X520 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X521 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X522 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X523 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X524 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X525 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X526 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X527 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X528 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X529 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X530 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X531 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X532 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X533 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X534 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X535 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X536 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X537 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X538 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X539 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X540 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X541 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X542 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X543 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X544 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X545 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X546 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X547 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X548 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X549 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X550 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X551 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X552 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X553 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X554 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X555 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X556 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X557 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X558 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X559 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X560 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X561 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X562 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X563 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X564 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X565 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X566 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X567 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X568 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X569 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X570 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X571 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X572 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X573 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X574 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X575 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X576 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X577 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X578 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X579 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X580 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X581 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X582 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X583 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X584 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X585 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X586 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X587 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X588 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X589 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X590 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X591 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X592 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X593 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X594 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X595 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X596 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X597 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X598 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X599 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X600 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X601 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X602 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X603 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X604 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X605 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X606 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X607 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X608 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X609 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X610 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X611 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X612 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X613 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X614 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X615 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X616 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X617 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X618 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X619 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X620 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X621 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X622 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X623 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X624 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X625 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X626 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X627 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X628 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X629 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X630 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X631 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X632 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X633 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X634 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X635 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X636 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X637 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X638 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X639 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X640 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X641 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X642 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X643 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X644 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X645 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X646 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X647 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X648 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X649 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X650 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X651 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X652 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X653 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X654 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X655 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X656 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X657 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X658 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X659 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X660 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X661 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X662 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X663 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X664 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X665 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X666 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X667 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X668 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X669 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X670 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X671 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X672 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X673 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X674 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X675 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X676 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X677 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X678 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X679 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X680 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X681 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X682 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X683 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X684 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X685 vdd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X686 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X687 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X688 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X689 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X690 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X691 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X692 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X693 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X694 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X695 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X696 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X697 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X698 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X699 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X700 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X701 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X702 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X703 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X704 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X705 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X706 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X707 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X708 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X709 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X710 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X711 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X712 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X713 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X714 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X715 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X716 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X717 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X718 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X719 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X720 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X721 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X722 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X723 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X724 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X725 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X726 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X727 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X728 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X729 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X730 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X731 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X732 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X733 tapered_buf_2/a_580_0# tapered_buf_2/a_160_n140# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X734 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X735 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X736 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X737 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X738 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X739 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X740 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X741 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X742 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X743 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X744 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X745 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X746 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X747 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X748 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X749 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X750 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X751 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X752 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X753 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X754 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X755 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X756 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X757 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X758 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X759 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X760 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X761 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X762 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X763 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X764 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X765 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X766 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X767 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X768 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X769 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X770 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X771 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X772 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X773 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X774 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X775 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X776 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X777 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X778 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X779 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X780 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X781 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X782 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X783 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X784 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X785 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X786 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X787 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X788 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X789 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X790 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X791 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X792 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X793 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X794 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X795 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X796 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X797 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X798 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X799 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X800 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X801 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X802 tapered_buf_2/a_160_n140# pd_0/UP tapered_buf_2/a_n10_n140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X803 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X804 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X805 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X806 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X807 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X808 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X809 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X810 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X811 vdd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X812 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X813 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X814 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X815 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X816 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X817 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X818 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X819 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X820 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X821 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X822 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X823 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X824 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X825 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X826 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X827 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X828 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X829 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X830 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X831 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X832 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X833 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X834 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X835 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X836 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X837 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X838 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X839 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X840 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X841 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X842 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X843 tapered_buf_2/a_580_0# tapered_buf_2/a_160_n140# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X844 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X845 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X846 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X847 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X848 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X849 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X850 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X851 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X852 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X853 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X854 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X855 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X856 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X857 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X858 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X859 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X860 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X861 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X862 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X863 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X864 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X865 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X866 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X867 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X868 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X869 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X870 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X871 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X872 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X873 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X874 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X875 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X876 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X877 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X878 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X879 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X880 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X881 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X882 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X883 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X884 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X885 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X886 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X887 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X888 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X889 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X890 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X891 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X892 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X893 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X894 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X895 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X896 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X897 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X898 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X899 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X900 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X901 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X902 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X903 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X904 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X905 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X906 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X907 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X908 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X909 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X910 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X911 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X912 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X913 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X914 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X915 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X916 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X917 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X918 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X919 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X920 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X921 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X922 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X923 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X924 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X925 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X926 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X927 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X928 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X929 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X930 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X931 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X932 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X933 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X934 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X935 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X936 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X937 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X938 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X939 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X940 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X941 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X942 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X943 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X944 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X945 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X946 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X947 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X948 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X949 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X950 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X951 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X952 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X953 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X954 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X955 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X956 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X957 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X958 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X959 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X960 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X961 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X962 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X963 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X964 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X965 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X966 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X967 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X968 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X969 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X970 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X971 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X972 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X973 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X974 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X975 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X976 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X977 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X978 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X979 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X980 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X981 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X982 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X983 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X984 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X985 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X986 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X987 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X988 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X989 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X990 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X991 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X992 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X993 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X994 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X995 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X996 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X997 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X998 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X999 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1000 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1001 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1002 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1003 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1004 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1005 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1006 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1007 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1008 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1009 vdd tapered_buf_2/a_160_n140# tapered_buf_2/a_580_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1010 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1011 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1012 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1013 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1014 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1015 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1016 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1017 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1018 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1019 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1020 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1021 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1022 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1023 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1024 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1025 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1026 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1027 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1028 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1029 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1030 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1031 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1032 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1033 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1034 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1035 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1036 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1037 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1038 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1039 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1040 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1041 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1042 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1043 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1044 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1045 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1046 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1047 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1048 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1049 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1050 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1051 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1052 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1053 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1054 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1055 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1056 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1057 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1058 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1059 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1060 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1061 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1062 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1063 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1064 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1065 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1066 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1067 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1068 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1069 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1070 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1071 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1072 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1073 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1074 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1075 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1076 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1077 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1078 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1079 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1080 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1081 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1082 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1083 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1084 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1085 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1086 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1087 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1088 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1089 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1090 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1091 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1092 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1093 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1094 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1095 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1096 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1097 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1098 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1099 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1100 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1101 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1102 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1103 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1104 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1105 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1106 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1107 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1108 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1109 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1110 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1111 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1112 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1113 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1114 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1115 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1116 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1117 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1118 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1119 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1120 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1121 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1122 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1123 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1124 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1125 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1126 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1127 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1128 vdd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1129 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1130 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1131 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1132 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1133 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1134 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1135 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1136 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1137 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1138 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1139 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1140 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1141 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1142 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1143 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1144 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1145 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1146 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1147 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1148 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1149 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1150 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1151 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1152 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1153 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1154 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1155 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1156 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1157 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1158 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1159 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1160 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1161 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1162 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1163 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1164 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1165 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1166 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1167 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1168 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1169 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1170 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1171 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1172 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1173 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1174 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1175 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1176 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1177 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1178 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1179 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1180 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1181 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1182 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1183 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1184 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1185 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1186 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1187 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1188 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1189 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1190 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1191 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1192 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1193 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1194 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1195 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1196 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1197 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1198 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1199 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1200 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1201 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1202 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1203 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1204 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1205 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1206 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1207 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1208 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1209 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1210 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1211 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1212 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1213 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1214 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1215 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1216 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1217 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1218 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1219 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1220 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1221 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1222 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1223 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1224 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1225 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1226 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1227 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1228 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1229 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1230 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1231 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1232 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1233 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1234 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1235 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1236 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1237 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1238 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1239 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1240 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1241 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1242 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1243 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1244 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1245 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1246 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1247 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1248 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1249 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1250 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1251 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1252 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1253 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1254 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1255 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1256 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1257 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1258 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1259 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1260 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1261 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1262 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1263 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1264 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1265 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1266 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1267 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1268 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1269 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1270 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1271 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1272 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1273 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1274 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1275 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1276 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1277 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1278 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1279 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1280 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1281 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1282 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1283 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1284 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1285 vdd tapered_buf_2/a_160_n140# tapered_buf_2/a_580_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1286 tapered_buf_2/a_580_0# tapered_buf_2/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1287 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1288 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1289 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1290 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1291 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1292 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1293 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1294 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1295 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1296 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1297 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1298 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1299 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1300 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1301 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1302 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1303 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1304 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1305 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1306 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1307 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1308 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1309 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1310 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1311 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1312 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1313 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1314 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1315 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1316 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1317 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1318 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1319 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1320 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1321 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1322 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1323 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1324 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1325 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1326 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1327 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1328 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1329 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1330 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1331 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1332 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1333 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1334 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1335 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1336 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1337 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1338 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1339 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1340 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1341 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1342 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1343 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1344 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1345 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1346 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1347 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1348 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1349 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1350 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1351 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1352 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1353 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1354 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1355 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1356 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1357 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1358 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1359 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1360 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1361 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1362 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1363 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1364 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1365 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1366 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1367 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1368 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1369 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1370 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1371 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1372 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1373 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1374 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1375 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1376 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1377 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1378 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1379 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1380 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1381 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1382 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1383 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1384 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1385 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1386 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1387 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1388 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1389 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1390 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1391 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1392 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1393 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1394 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1395 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1396 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1397 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1398 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1399 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1400 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1401 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1402 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1403 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1404 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1405 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1406 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1407 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1408 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1409 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1410 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1411 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1412 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1413 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1414 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1415 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1416 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1417 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1418 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1419 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1420 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1421 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1422 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1423 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1424 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1425 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1426 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1427 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1428 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1429 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1430 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1431 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1432 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1433 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1434 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1435 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1436 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1437 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1438 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1439 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1440 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1441 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1442 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1443 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1444 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1445 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1446 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1447 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1448 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1449 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1450 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1451 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1452 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1453 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1454 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1455 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1456 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1457 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1458 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1459 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1460 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1461 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1462 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1463 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1464 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1465 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1466 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1467 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1468 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1469 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1470 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1471 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1472 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1473 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1474 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1475 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1476 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1477 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1478 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1479 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1480 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1481 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1482 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1483 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1484 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1485 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1486 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1487 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1488 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1489 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1490 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1491 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1492 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1493 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1494 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1495 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1496 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1497 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1498 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1499 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1500 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1501 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1502 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1503 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1504 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1505 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1506 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1507 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1508 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1509 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1510 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1511 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1512 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1513 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1514 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1515 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1516 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1517 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1518 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1519 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1520 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1521 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1522 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1523 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1524 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1525 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1526 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1527 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1528 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1529 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1530 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1531 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1532 vdd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1533 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1534 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1535 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1536 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1537 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1538 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1539 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1540 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1541 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1542 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1543 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1544 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1545 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1546 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1547 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1548 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1549 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1550 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1551 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1552 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1553 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1554 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1555 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1556 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1557 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1558 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1559 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1560 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1561 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1562 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1563 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1564 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1565 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1566 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1567 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1568 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1569 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1570 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1571 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1572 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1573 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1574 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1575 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1576 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1577 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1578 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1579 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1580 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1581 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1582 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1583 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1584 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1585 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1586 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1587 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1588 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1589 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1590 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1591 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1592 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1593 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1594 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1595 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1596 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1597 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1598 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1599 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1600 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1601 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1602 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1603 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1604 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1605 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1606 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1607 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1608 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1609 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1610 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1611 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1612 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1613 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1614 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1615 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1616 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1617 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1618 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1619 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1620 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1621 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1622 gnd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1623 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1624 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1625 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1626 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1627 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1628 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1629 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1630 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1631 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1632 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1633 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1634 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1635 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1636 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1637 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1638 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1639 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1640 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1641 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1642 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1643 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1644 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1645 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1646 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1647 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1648 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1649 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1650 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1651 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1652 vdd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1653 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1654 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1655 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1656 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1657 tapered_buf_2/a_1650_0# tapered_buf_2/a_580_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1658 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1659 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1660 vdd tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1661 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1662 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1663 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1664 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1665 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1666 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1667 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1668 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1669 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1670 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1671 gnd tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1672 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1673 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1674 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1675 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1676 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1677 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1678 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1679 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1680 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1681 vdd tapered_buf_2/a_210_n610# tapered_buf_2/out tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1682 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1683 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1684 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1685 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1686 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1687 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1688 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1689 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1690 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1691 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1692 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1693 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1694 gnd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1695 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1696 gnd tapered_buf_2/a_210_n610# tapered_buf_2/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1697 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1698 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# vdd tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1699 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1700 vdd tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# tapered_buf_2/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1701 tapered_buf_2/out tapered_buf_2/a_210_n610# vdd tapered_buf_2/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1702 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1703 tapered_buf_2/a_210_n610# tapered_buf_2/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1704 tapered_buf_2/out tapered_buf_2/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1705 tapered_buf_2/a_4670_0# tapered_buf_2/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1706 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1707 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1708 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1709 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1710 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1711 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1712 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1713 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1714 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1715 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1716 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1717 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1718 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1719 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1720 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1721 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1722 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1723 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1724 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1725 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1726 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1727 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1728 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1729 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1730 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1731 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1732 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1733 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1734 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1735 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1736 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1737 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1738 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1739 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1740 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1741 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1742 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1743 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1744 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1745 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1746 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1747 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1748 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1749 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1750 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1751 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1752 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1753 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1754 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1755 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1756 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1757 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1758 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1759 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1760 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1761 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1762 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1763 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1764 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1765 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1766 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1767 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1768 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1769 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1770 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1771 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1772 vdd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1773 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1774 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1775 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1776 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1777 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1778 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1779 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1780 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1781 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1782 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1783 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1784 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1785 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1786 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1787 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1788 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1789 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1790 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1791 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1792 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1793 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1794 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1795 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1796 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1797 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1798 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1799 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1800 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1801 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1802 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1803 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1804 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1805 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1806 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1807 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1808 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1809 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1810 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1811 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1812 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1813 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1814 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1815 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1816 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1817 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1818 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1819 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1820 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1821 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1822 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1823 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1824 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1825 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1826 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1827 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1828 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1829 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1830 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1831 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1832 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1833 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1834 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1835 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1836 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1837 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1838 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1839 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1840 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1841 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1842 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1843 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1844 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1845 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1846 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1847 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1848 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1849 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1850 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1851 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1852 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1853 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1854 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1855 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1856 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1857 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1858 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1859 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1860 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1861 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1862 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1863 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1864 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1865 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1866 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1867 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1868 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1869 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1870 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1871 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1872 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1873 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1874 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1875 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1876 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1877 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1878 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1879 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1880 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1881 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1882 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1883 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1884 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1885 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1886 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1887 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1888 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1889 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1890 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1891 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1892 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1893 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1894 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1895 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1896 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1897 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1898 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1899 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1900 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1901 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1902 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1903 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1904 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1905 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1906 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1907 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1908 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1909 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1910 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1911 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1912 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1913 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1914 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1915 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1916 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1917 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1918 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1919 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1920 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1921 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1922 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1923 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1924 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1925 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1926 tapered_buf_3/a_160_230# pd_0/DOWN tapered_buf_3/a_n10_230# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1927 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1928 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1929 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1930 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1931 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1932 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1933 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1934 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1935 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1936 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1937 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1938 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1939 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1940 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1941 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1942 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1943 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1944 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1945 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1946 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1947 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1948 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1949 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1950 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1951 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1952 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1953 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1954 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1955 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1956 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1957 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1958 tapered_buf_3/a_580_0# tapered_buf_3/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1959 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1960 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1961 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1962 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1963 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1964 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1965 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1966 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1967 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1968 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1969 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1970 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1971 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1972 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1973 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1974 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1975 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1976 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1977 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1978 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1979 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1980 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1981 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1982 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1983 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1984 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1985 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1986 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1987 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1988 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1989 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1990 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1991 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1992 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1993 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1994 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1995 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1996 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1997 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1998 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1999 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2000 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2001 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2002 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2003 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2004 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2005 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2006 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2007 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2008 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2009 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2010 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2011 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2012 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2013 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2014 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2015 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2016 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2017 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2018 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2019 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2020 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2021 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2022 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2023 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2024 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2025 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2026 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2027 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2028 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2029 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2030 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2031 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2032 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2033 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2034 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2035 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2036 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2037 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2038 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2039 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2040 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2041 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2042 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2043 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2044 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2045 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2046 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2047 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2048 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2049 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2050 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2051 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2052 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2053 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2054 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2055 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2056 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2057 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2058 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2059 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2060 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2061 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2062 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2063 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2064 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2065 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2066 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2067 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2068 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2069 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2070 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2071 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2072 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2073 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2074 gnd tapered_buf_3/a_160_n140# tapered_buf_3/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2075 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2076 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2077 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2078 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2079 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2080 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2081 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2082 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2083 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2084 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2085 vdd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2086 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2087 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2088 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2089 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2090 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2091 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2092 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2093 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2094 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2095 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2096 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2097 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2098 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2099 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2100 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2101 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2102 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2103 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2104 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2105 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2106 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2107 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2108 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2109 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2110 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2111 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2112 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2113 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2114 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2115 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2116 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2117 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2118 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2119 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2120 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2121 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2122 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2123 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2124 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2125 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2126 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2127 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2128 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2129 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2130 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2131 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2132 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2133 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2134 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2135 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2136 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2137 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2138 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2139 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2140 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2141 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2142 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2143 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2144 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2145 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2146 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2147 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2148 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2149 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2150 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2151 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2152 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2153 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2154 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2155 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2156 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2157 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2158 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2159 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2160 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2161 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2162 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2163 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2164 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2165 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2166 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2167 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2168 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2169 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2170 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2171 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2172 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2173 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2174 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2175 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2176 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2177 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2178 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2179 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2180 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2181 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2182 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2183 gnd tapered_buf_3/a_160_n140# tapered_buf_3/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2184 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2185 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2186 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2187 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2188 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2189 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2190 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2191 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2192 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2193 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2194 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2195 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2196 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2197 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2198 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2199 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2200 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2201 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2202 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2203 vdd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2204 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2205 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2206 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2207 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2208 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2209 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2210 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2211 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2212 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2213 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2214 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2215 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2216 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2217 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2218 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2219 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2220 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2221 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2222 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2223 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2224 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2225 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2226 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2227 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2228 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2229 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2230 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2231 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2232 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2233 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2234 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2235 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2236 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2237 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2238 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2239 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2240 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2241 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2242 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2243 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2244 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2245 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2246 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2247 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2248 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2249 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2250 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2251 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2252 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2253 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2254 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2255 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2256 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2257 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2258 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2259 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2260 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2261 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2262 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2263 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2264 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2265 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2266 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2267 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2268 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2269 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2270 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2271 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2272 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2273 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2274 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2275 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2276 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2277 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2278 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2279 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2280 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2281 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2282 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2283 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2284 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2285 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2286 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2287 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2288 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2289 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2290 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2291 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2292 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2293 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2294 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2295 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2296 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2297 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2298 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2299 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2300 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2301 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2302 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2303 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2304 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2305 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2306 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2307 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2308 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2309 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2310 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2311 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2312 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2313 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2314 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2315 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2316 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2317 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2318 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2319 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2320 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2321 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2322 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2323 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2324 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2325 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2326 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2327 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2328 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2329 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2330 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2331 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2332 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2333 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2334 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2335 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2336 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2337 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2338 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2339 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2340 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2341 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2342 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2343 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2344 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2345 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2346 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2347 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2348 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2349 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2350 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2351 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2352 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2353 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2354 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2355 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2356 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2357 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2358 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2359 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2360 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2361 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2362 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2363 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2364 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2365 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2366 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2367 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2368 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2369 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2370 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2371 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2372 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2373 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2374 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2375 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2376 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2377 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2378 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2379 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2380 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2381 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2382 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2383 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2384 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2385 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2386 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2387 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2388 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2389 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2390 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2391 vdd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2392 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2393 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2394 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2395 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2396 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2397 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2398 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2399 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2400 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2401 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2402 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2403 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2404 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2405 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2406 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2407 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2408 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2409 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2410 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2411 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2412 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2413 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2414 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2415 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2416 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2417 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2418 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2419 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2420 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2421 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2422 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2423 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2424 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2425 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2426 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2427 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2428 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2429 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2430 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2431 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2432 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2433 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2434 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2435 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2436 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2437 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2438 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2439 tapered_buf_3/a_580_0# tapered_buf_3/a_160_n140# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2440 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2441 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2442 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2443 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2444 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2445 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2446 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2447 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2448 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2449 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2450 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2451 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2452 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2453 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2454 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2455 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2456 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2457 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2458 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2459 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2460 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2461 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2462 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2463 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2464 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2465 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2466 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2467 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2468 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2469 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2470 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2471 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2472 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2473 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2474 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2475 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2476 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2477 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2478 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2479 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2480 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2481 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2482 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2483 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2484 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2485 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2486 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2487 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2488 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2489 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2490 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2491 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2492 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2493 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2494 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2495 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2496 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2497 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2498 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2499 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2500 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2501 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2502 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2503 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2504 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2505 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2506 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2507 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2508 tapered_buf_3/a_160_n140# pd_0/DOWN tapered_buf_3/a_n10_n140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2509 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2510 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2511 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2512 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2513 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2514 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2515 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2516 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2517 vdd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2518 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2519 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2520 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2521 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2522 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2523 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2524 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2525 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2526 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2527 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2528 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2529 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2530 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2531 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2532 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2533 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2534 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2535 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2536 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2537 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2538 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2539 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2540 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2541 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2542 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2543 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2544 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2545 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2546 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2547 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2548 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2549 tapered_buf_3/a_580_0# tapered_buf_3/a_160_n140# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2550 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2551 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2552 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2553 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2554 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2555 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2556 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2557 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2558 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2559 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2560 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2561 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2562 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2563 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2564 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2565 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2566 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2567 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2568 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2569 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2570 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2571 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2572 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2573 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2574 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2575 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2576 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2577 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2578 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2579 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2580 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2581 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2582 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2583 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2584 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2585 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2586 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2587 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2588 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2589 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2590 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2591 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2592 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2593 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2594 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2595 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2596 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2597 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2598 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2599 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2600 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2601 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2602 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2603 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2604 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2605 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2606 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2607 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2608 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2609 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2610 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2611 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2612 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2613 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2614 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2615 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2616 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2617 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2618 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2619 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2620 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2621 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2622 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2623 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2624 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2625 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2626 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2627 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2628 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2629 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2630 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2631 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2632 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2633 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2634 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2635 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2636 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2637 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2638 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2639 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2640 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2641 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2642 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2643 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2644 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2645 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2646 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2647 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2648 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2649 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2650 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2651 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2652 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2653 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2654 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2655 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2656 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2657 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2658 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2659 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2660 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2661 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2662 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2663 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2664 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2665 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2666 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2667 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2668 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2669 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2670 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2671 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2672 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2673 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2674 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2675 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2676 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2677 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2678 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2679 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2680 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2681 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2682 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2683 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2684 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2685 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2686 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2687 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2688 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2689 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2690 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2691 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2692 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2693 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2694 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2695 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2696 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2697 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2698 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2699 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2700 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2701 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2702 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2703 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2704 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2705 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2706 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2707 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2708 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2709 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2710 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2711 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2712 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2713 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2714 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2715 vdd tapered_buf_3/a_160_n140# tapered_buf_3/a_580_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2716 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2717 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2718 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2719 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2720 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2721 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2722 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2723 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2724 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2725 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2726 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2727 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2728 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2729 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2730 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2731 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2732 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2733 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2734 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2735 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2736 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2737 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2738 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2739 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2740 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2741 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2742 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2743 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2744 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2745 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2746 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2747 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2748 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2749 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2750 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2751 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2752 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2753 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2754 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2755 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2756 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2757 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2758 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2759 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2760 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2761 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2762 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2763 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2764 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2765 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2766 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2767 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2768 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2769 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2770 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2771 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2772 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2773 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2774 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2775 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2776 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2777 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2778 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2779 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2780 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2781 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2782 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2783 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2784 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2785 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2786 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2787 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2788 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2789 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2790 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2791 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2792 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2793 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2794 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2795 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2796 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2797 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2798 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2799 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2800 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2801 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2802 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2803 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2804 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2805 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2806 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2807 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2808 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2809 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2810 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2811 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2812 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2813 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2814 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2815 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2816 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2817 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2818 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2819 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2820 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2821 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2822 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2823 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2824 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2825 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2826 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2827 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2828 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2829 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2830 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2831 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2832 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2833 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2834 vdd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2835 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2836 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2837 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2838 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2839 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2840 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2841 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2842 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2843 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2844 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2845 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2846 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2847 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2848 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2849 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2850 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2851 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2852 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2853 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2854 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2855 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2856 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2857 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2858 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2859 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2860 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2861 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2862 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2863 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2864 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2865 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2866 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2867 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2868 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2869 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2870 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2871 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2872 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2873 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2874 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2875 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2876 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2877 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2878 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2879 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2880 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2881 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2882 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2883 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2884 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2885 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2886 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2887 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2888 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2889 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2890 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2891 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2892 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2893 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2894 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2895 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2896 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2897 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2898 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2899 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2900 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2901 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2902 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2903 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2904 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2905 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2906 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2907 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2908 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2909 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2910 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2911 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2912 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2913 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2914 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2915 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2916 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2917 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2918 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2919 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2920 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2921 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2922 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2923 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2924 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2925 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2926 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2927 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2928 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2929 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2930 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2931 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2932 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2933 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2934 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2935 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2936 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2937 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2938 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2939 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2940 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2941 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2942 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2943 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2944 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2945 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2946 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2947 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2948 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2949 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2950 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2951 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2952 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2953 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2954 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2955 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2956 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2957 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2958 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2959 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2960 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2961 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2962 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2963 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2964 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2965 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2966 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2967 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2968 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2969 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2970 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2971 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2972 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2973 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2974 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2975 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2976 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2977 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2978 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2979 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2980 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2981 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2982 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2983 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2984 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2985 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2986 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2987 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2988 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2989 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2990 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2991 vdd tapered_buf_3/a_160_n140# tapered_buf_3/a_580_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2992 tapered_buf_3/a_580_0# tapered_buf_3/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2993 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2994 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2995 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2996 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2997 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2998 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2999 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3000 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3001 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3002 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3003 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3004 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3005 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3006 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3007 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3008 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3009 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3010 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3011 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3012 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3013 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3014 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3015 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3016 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3017 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3018 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3019 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3020 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3021 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3022 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3023 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3024 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3025 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3026 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3027 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3028 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3029 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3030 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3031 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3032 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3033 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3034 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3035 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3036 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3037 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3038 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3039 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3040 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3041 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3042 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3043 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3044 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3045 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3046 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3047 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3048 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3049 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3050 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3051 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3052 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3053 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3054 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3055 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3056 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3057 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3058 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3059 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3060 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3061 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3062 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3063 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3064 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3065 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3066 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3067 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3068 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3069 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3070 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3071 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3072 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3073 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3074 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3075 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3076 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3077 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3078 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3079 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3080 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3081 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3082 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3083 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3084 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3085 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3086 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3087 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3088 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3089 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3090 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3091 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3092 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3093 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3094 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3095 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3096 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3097 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3098 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3099 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3100 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3101 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3102 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3103 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3104 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3105 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3106 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3107 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3108 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3109 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3110 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3111 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3112 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3113 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3114 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3115 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3116 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3117 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3118 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3119 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3120 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3121 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3122 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3123 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3124 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3125 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3126 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3127 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3128 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3129 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3130 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3131 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3132 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3133 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3134 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3135 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3136 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3137 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3138 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3139 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3140 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3141 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3142 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3143 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3144 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3145 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3146 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3147 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3148 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3149 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3150 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3151 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3152 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3153 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3154 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3155 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3156 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3157 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3158 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3159 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3160 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3161 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3162 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3163 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3164 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3165 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3166 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3167 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3168 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3169 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3170 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3171 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3172 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3173 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3174 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3175 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3176 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3177 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3178 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3179 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3180 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3181 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3182 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3183 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3184 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3185 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3186 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3187 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3188 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3189 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3190 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3191 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3192 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3193 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3194 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3195 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3196 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3197 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3198 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3199 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3200 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3201 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3202 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3203 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3204 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3205 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3206 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3207 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3208 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3209 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3210 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3211 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3212 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3213 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3214 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3215 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3216 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3217 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3218 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3219 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3220 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3221 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3222 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3223 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3224 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3225 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3226 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3227 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3228 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3229 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3230 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3231 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3232 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3233 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3234 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3235 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3236 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3237 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3238 vdd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3239 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3240 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3241 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3242 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3243 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3244 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3245 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3246 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3247 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3248 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3249 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3250 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3251 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3252 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3253 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3254 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3255 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3256 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3257 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3258 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3259 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3260 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3261 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3262 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3263 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3264 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3265 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3266 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3267 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3268 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3269 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3270 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3271 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3272 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3273 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3274 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3275 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3276 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3277 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3278 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3279 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3280 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3281 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3282 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3283 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3284 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3285 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3286 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3287 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3288 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3289 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3290 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3291 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3292 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3293 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3294 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3295 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3296 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3297 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3298 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3299 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3300 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3301 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3302 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3303 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3304 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3305 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3306 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3307 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3308 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3309 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3310 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3311 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3312 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3313 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3314 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3315 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3316 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3317 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3318 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3319 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3320 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3321 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3322 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3323 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3324 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3325 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3326 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3327 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3328 gnd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3329 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3330 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3331 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3332 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3333 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3334 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3335 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3336 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3337 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3338 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3339 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3340 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3341 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3342 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3343 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3344 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3345 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3346 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3347 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3348 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3349 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3350 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3351 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3352 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3353 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3354 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3355 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3356 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3357 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3358 vdd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3359 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3360 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3361 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3362 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3363 tapered_buf_3/a_1650_0# tapered_buf_3/a_580_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3364 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3365 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3366 vdd tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3367 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3368 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3369 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3370 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3371 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3372 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3373 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3374 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3375 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3376 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3377 gnd tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3378 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3379 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3380 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3381 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3382 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3383 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3384 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3385 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3386 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3387 vdd tapered_buf_3/a_210_n610# tapered_buf_3/out tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3388 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3389 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3390 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3391 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3392 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3393 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3394 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3395 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3396 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3397 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3398 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3399 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3400 gnd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3401 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3402 gnd tapered_buf_3/a_210_n610# tapered_buf_3/out gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3403 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3404 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# vdd tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3405 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3406 vdd tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# tapered_buf_3/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3407 tapered_buf_3/out tapered_buf_3/a_210_n610# vdd tapered_buf_3/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3408 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3409 tapered_buf_3/a_210_n610# tapered_buf_3/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3410 tapered_buf_3/out tapered_buf_3/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3411 tapered_buf_3/a_4670_0# tapered_buf_3/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3412 pd_0/UP pd_0/tspc_r_0/Qbar1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3413 pd_0/tspc_r_0/Qbar pd_0/UP gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3414 pd_0/tspc_r_0/Z1 vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3415 pd_0/UP pd_0/tspc_r_0/Qbar1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3416 pd_0/tspc_r_0/Qbar1 pd_0/REF pd_0/tspc_r_0/z5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3417 pd_0/tspc_r_0/z5 pd_0/tspc_r_0/Z3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3418 pd_0/tspc_r_0/Z3 pd_0/REF vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3419 pd_0/tspc_r_0/Z2 pd_0/REF pd_0/tspc_r_0/Z1 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3420 pd_0/tspc_r_0/Z3 pd_0/tspc_r_0/Z2 pd_0/tspc_r_0/Z4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3421 pd_0/tspc_r_0/Z4 pd_0/REF gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3422 pd_0/tspc_r_0/Z3 pd_0/R gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3423 pd_0/tspc_r_0/Qbar pd_0/UP vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3424 pd_0/tspc_r_0/Qbar1 pd_0/tspc_r_0/Z3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3425 pd_0/tspc_r_0/Z2 vdd gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3426 pd_0/DOWN pd_0/tspc_r_1/Qbar1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3427 pd_0/tspc_r_1/Qbar pd_0/DOWN gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3428 pd_0/tspc_r_1/Z1 vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3429 pd_0/DOWN pd_0/tspc_r_1/Qbar1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3430 pd_0/tspc_r_1/Qbar1 pd_0/DIV pd_0/tspc_r_1/z5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3431 pd_0/tspc_r_1/z5 pd_0/tspc_r_1/Z3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3432 pd_0/tspc_r_1/Z3 pd_0/DIV vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3433 pd_0/tspc_r_1/Z2 pd_0/DIV pd_0/tspc_r_1/Z1 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3434 pd_0/tspc_r_1/Z3 pd_0/tspc_r_1/Z2 pd_0/tspc_r_1/Z4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3435 pd_0/tspc_r_1/Z4 pd_0/DIV gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3436 pd_0/tspc_r_1/Z3 pd_0/R gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3437 pd_0/tspc_r_1/Qbar pd_0/DOWN vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3438 pd_0/tspc_r_1/Qbar1 pd_0/tspc_r_1/Z3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3439 pd_0/tspc_r_1/Z2 vdd gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3440 pd_0/R pd_0/and_pd_0/Out1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3441 pd_0/and_pd_0/Out1 pd_0/UP pd_0/and_pd_0/Z1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3442 pd_0/and_pd_0/Out1 pd_0/UP vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3443 pd_0/and_pd_0/Z1 pd_0/DOWN gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3444 pd_0/and_pd_0/Out1 pd_0/DOWN vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X3445 pd_0/R pd_0/and_pd_0/Out1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=150000u
X3446 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3447 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3448 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3449 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3450 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3451 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3452 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3453 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3454 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3455 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3456 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3457 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3458 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3459 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3460 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3461 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3462 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3463 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3464 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3465 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3466 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3467 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3468 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3469 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3470 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3471 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3472 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3473 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3474 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3475 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3476 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3477 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3478 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3479 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3480 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3481 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3482 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3483 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3484 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3485 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3486 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3487 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3488 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3489 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3490 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3491 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3492 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3493 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3494 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3495 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3496 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3497 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3498 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3499 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3500 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3501 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3502 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3503 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3504 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3505 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3506 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3507 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3508 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3509 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3510 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3511 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3512 vdd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3513 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3514 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3515 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3516 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3517 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3518 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3519 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3520 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3521 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3522 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3523 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3524 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3525 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3526 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3527 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3528 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3529 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3530 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3531 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3532 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3533 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3534 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3535 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3536 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3537 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3538 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3539 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3540 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3541 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3542 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3543 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3544 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3545 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3546 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3547 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3548 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3549 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3550 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3551 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3552 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3553 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3554 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3555 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3556 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3557 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3558 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3559 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3560 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3561 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3562 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3563 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3564 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3565 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3566 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3567 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3568 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3569 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3570 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3571 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3572 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3573 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3574 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3575 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3576 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3577 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3578 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3579 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3580 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3581 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3582 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3583 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3584 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3585 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3586 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3587 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3588 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3589 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3590 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3591 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3592 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3593 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3594 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3595 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3596 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3597 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3598 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3599 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3600 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3601 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3602 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3603 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3604 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3605 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3606 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3607 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3608 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3609 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3610 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3611 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3612 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3613 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3614 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3615 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3616 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3617 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3618 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3619 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3620 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3621 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3622 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3623 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3624 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3625 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3626 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3627 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3628 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3629 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3630 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3631 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3632 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3633 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3634 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3635 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3636 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3637 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3638 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3639 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3640 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3641 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3642 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3643 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3644 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3645 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3646 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3647 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3648 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3649 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3650 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3651 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3652 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3653 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3654 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3655 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3656 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3657 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3658 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3659 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3660 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3661 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3662 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3663 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3664 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3665 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3666 tapered_buf_0/a_160_230# tapered_buf_0/in tapered_buf_0/a_n10_230# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3667 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3668 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3669 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3670 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3671 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3672 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3673 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3674 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3675 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3676 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3677 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3678 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3679 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3680 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3681 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3682 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3683 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3684 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3685 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3686 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3687 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3688 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3689 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3690 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3691 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3692 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3693 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3694 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3695 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3696 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3697 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3698 tapered_buf_0/a_580_0# tapered_buf_0/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3699 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3700 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3701 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3702 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3703 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3704 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3705 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3706 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3707 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3708 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3709 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3710 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3711 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3712 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3713 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3714 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3715 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3716 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3717 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3718 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3719 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3720 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3721 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3722 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3723 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3724 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3725 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3726 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3727 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3728 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3729 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3730 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3731 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3732 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3733 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3734 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3735 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3736 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3737 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3738 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3739 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3740 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3741 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3742 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3743 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3744 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3745 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3746 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3747 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3748 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3749 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3750 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3751 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3752 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3753 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3754 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3755 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3756 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3757 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3758 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3759 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3760 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3761 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3762 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3763 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3764 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3765 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3766 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3767 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3768 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3769 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3770 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3771 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3772 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3773 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3774 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3775 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3776 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3777 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3778 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3779 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3780 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3781 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3782 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3783 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3784 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3785 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3786 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3787 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3788 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3789 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3790 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3791 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3792 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3793 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3794 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3795 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3796 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3797 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3798 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3799 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3800 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3801 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3802 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3803 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3804 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3805 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3806 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3807 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3808 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3809 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3810 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3811 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3812 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3813 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3814 gnd tapered_buf_0/a_160_n140# tapered_buf_0/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3815 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3816 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3817 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3818 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3819 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3820 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3821 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3822 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3823 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3824 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3825 vdd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3826 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3827 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3828 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3829 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3830 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3831 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3832 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3833 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3834 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3835 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3836 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3837 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3838 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3839 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3840 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3841 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3842 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3843 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3844 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3845 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3846 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3847 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3848 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3849 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3850 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3851 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3852 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3853 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3854 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3855 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3856 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3857 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3858 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3859 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3860 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3861 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3862 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3863 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3864 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3865 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3866 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3867 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3868 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3869 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3870 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3871 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3872 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3873 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3874 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3875 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3876 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3877 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3878 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3879 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3880 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3881 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3882 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3883 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3884 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3885 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3886 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3887 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3888 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3889 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3890 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3891 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3892 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3893 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3894 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3895 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3896 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3897 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3898 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3899 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3900 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3901 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3902 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3903 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3904 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3905 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3906 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3907 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3908 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3909 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3910 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3911 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3912 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3913 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3914 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3915 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3916 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3917 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3918 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3919 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3920 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3921 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3922 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3923 gnd tapered_buf_0/a_160_n140# tapered_buf_0/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3924 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3925 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3926 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3927 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3928 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3929 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3930 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3931 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3932 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3933 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3934 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3935 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3936 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3937 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3938 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3939 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3940 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3941 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3942 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3943 vdd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3944 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3945 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3946 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3947 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3948 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3949 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3950 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3951 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3952 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3953 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3954 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3955 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3956 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3957 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3958 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3959 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3960 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3961 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3962 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3963 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3964 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3965 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3966 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3967 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3968 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3969 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3970 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3971 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3972 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3973 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3974 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3975 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3976 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3977 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3978 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3979 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3980 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3981 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3982 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3983 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3984 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3985 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3986 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3987 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3988 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3989 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3990 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3991 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3992 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3993 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3994 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3995 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3996 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3997 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3998 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3999 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4000 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4001 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4002 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4003 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4004 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4005 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4006 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4007 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4008 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4009 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4010 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4011 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4012 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4013 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4014 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4015 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4016 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4017 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4018 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4019 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4020 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4021 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4022 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4023 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4024 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4025 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4026 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4027 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4028 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4029 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4030 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4031 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4032 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4033 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4034 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4035 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4036 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4037 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4038 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4039 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4040 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4041 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4042 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4043 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4044 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4045 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4046 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4047 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4048 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4049 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4050 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4051 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4052 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4053 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4054 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4055 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4056 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4057 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4058 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4059 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4060 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4061 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4062 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4063 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4064 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4065 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4066 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4067 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4068 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4069 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4070 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4071 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4072 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4073 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4074 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4075 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4076 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4077 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4078 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4079 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4080 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4081 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4082 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4083 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4084 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4085 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4086 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4087 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4088 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4089 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4090 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4091 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4092 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4093 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4094 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4095 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4096 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4097 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4098 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4099 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4100 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4101 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4102 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4103 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4104 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4105 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4106 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4107 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4108 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4109 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4110 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4111 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4112 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4113 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4114 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4115 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4116 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4117 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4118 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4119 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4120 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4121 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4122 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4123 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4124 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4125 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4126 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4127 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4128 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4129 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4130 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4131 vdd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4132 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4133 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4134 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4135 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4136 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4137 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4138 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4139 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4140 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4141 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4142 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4143 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4144 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4145 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4146 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4147 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4148 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4149 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4150 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4151 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4152 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4153 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4154 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4155 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4156 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4157 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4158 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4159 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4160 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4161 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4162 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4163 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4164 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4165 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4166 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4167 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4168 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4169 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4170 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4171 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4172 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4173 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4174 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4175 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4176 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4177 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4178 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4179 tapered_buf_0/a_580_0# tapered_buf_0/a_160_n140# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4180 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4181 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4182 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4183 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4184 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4185 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4186 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4187 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4188 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4189 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4190 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4191 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4192 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4193 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4194 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4195 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4196 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4197 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4198 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4199 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4200 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4201 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4202 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4203 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4204 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4205 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4206 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4207 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4208 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4209 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4210 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4211 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4212 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4213 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4214 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4215 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4216 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4217 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4218 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4219 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4220 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4221 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4222 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4223 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4224 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4225 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4226 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4227 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4228 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4229 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4230 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4231 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4232 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4233 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4234 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4235 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4236 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4237 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4238 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4239 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4240 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4241 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4242 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4243 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4244 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4245 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4246 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4247 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4248 tapered_buf_0/a_160_n140# tapered_buf_0/in tapered_buf_0/a_n10_n140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4249 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4250 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4251 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4252 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4253 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4254 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4255 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4256 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4257 vdd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4258 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4259 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4260 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4261 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4262 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4263 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4264 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4265 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4266 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4267 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4268 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4269 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4270 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4271 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4272 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4273 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4274 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4275 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4276 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4277 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4278 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4279 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4280 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4281 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4282 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4283 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4284 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4285 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4286 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4287 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4288 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4289 tapered_buf_0/a_580_0# tapered_buf_0/a_160_n140# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4290 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4291 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4292 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4293 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4294 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4295 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4296 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4297 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4298 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4299 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4300 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4301 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4302 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4303 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4304 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4305 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4306 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4307 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4308 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4309 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4310 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4311 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4312 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4313 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4314 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4315 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4316 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4317 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4318 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4319 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4320 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4321 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4322 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4323 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4324 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4325 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4326 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4327 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4328 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4329 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4330 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4331 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4332 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4333 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4334 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4335 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4336 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4337 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4338 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4339 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4340 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4341 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4342 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4343 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4344 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4345 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4346 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4347 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4348 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4349 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4350 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4351 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4352 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4353 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4354 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4355 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4356 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4357 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4358 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4359 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4360 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4361 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4362 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4363 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4364 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4365 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4366 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4367 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4368 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4369 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4370 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4371 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4372 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4373 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4374 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4375 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4376 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4377 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4378 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4379 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4380 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4381 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4382 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4383 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4384 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4385 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4386 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4387 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4388 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4389 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4390 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4391 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4392 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4393 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4394 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4395 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4396 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4397 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4398 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4399 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4400 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4401 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4402 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4403 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4404 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4405 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4406 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4407 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4408 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4409 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4410 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4411 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4412 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4413 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4414 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4415 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4416 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4417 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4418 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4419 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4420 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4421 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4422 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4423 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4424 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4425 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4426 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4427 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4428 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4429 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4430 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4431 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4432 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4433 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4434 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4435 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4436 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4437 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4438 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4439 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4440 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4441 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4442 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4443 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4444 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4445 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4446 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4447 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4448 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4449 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4450 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4451 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4452 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4453 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4454 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4455 vdd tapered_buf_0/a_160_n140# tapered_buf_0/a_580_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4456 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4457 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4458 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4459 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4460 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4461 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4462 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4463 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4464 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4465 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4466 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4467 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4468 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4469 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4470 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4471 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4472 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4473 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4474 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4475 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4476 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4477 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4478 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4479 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4480 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4481 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4482 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4483 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4484 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4485 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4486 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4487 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4488 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4489 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4490 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4491 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4492 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4493 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4494 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4495 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4496 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4497 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4498 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4499 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4500 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4501 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4502 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4503 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4504 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4505 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4506 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4507 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4508 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4509 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4510 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4511 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4512 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4513 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4514 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4515 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4516 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4517 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4518 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4519 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4520 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4521 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4522 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4523 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4524 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4525 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4526 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4527 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4528 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4529 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4530 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4531 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4532 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4533 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4534 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4535 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4536 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4537 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4538 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4539 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4540 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4541 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4542 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4543 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4544 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4545 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4546 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4547 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4548 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4549 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4550 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4551 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4552 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4553 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4554 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4555 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4556 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4557 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4558 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4559 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4560 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4561 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4562 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4563 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4564 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4565 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4566 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4567 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4568 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4569 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4570 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4571 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4572 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4573 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4574 vdd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4575 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4576 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4577 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4578 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4579 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4580 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4581 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4582 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4583 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4584 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4585 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4586 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4587 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4588 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4589 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4590 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4591 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4592 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4593 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4594 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4595 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4596 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4597 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4598 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4599 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4600 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4601 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4602 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4603 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4604 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4605 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4606 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4607 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4608 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4609 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4610 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4611 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4612 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4613 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4614 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4615 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4616 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4617 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4618 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4619 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4620 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4621 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4622 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4623 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4624 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4625 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4626 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4627 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4628 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4629 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4630 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4631 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4632 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4633 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4634 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4635 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4636 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4637 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4638 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4639 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4640 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4641 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4642 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4643 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4644 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4645 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4646 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4647 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4648 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4649 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4650 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4651 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4652 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4653 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4654 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4655 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4656 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4657 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4658 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4659 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4660 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4661 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4662 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4663 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4664 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4665 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4666 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4667 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4668 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4669 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4670 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4671 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4672 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4673 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4674 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4675 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4676 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4677 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4678 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4679 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4680 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4681 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4682 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4683 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4684 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4685 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4686 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4687 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4688 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4689 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4690 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4691 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4692 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4693 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4694 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4695 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4696 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4697 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4698 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4699 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4700 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4701 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4702 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4703 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4704 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4705 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4706 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4707 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4708 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4709 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4710 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4711 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4712 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4713 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4714 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4715 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4716 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4717 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4718 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4719 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4720 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4721 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4722 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4723 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4724 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4725 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4726 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4727 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4728 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4729 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4730 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4731 vdd tapered_buf_0/a_160_n140# tapered_buf_0/a_580_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4732 tapered_buf_0/a_580_0# tapered_buf_0/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4733 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4734 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4735 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4736 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4737 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4738 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4739 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4740 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4741 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4742 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4743 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4744 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4745 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4746 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4747 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4748 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4749 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4750 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4751 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4752 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4753 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4754 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4755 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4756 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4757 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4758 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4759 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4760 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4761 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4762 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4763 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4764 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4765 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4766 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4767 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4768 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4769 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4770 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4771 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4772 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4773 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4774 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4775 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4776 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4777 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4778 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4779 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4780 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4781 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4782 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4783 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4784 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4785 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4786 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4787 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4788 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4789 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4790 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4791 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4792 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4793 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4794 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4795 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4796 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4797 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4798 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4799 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4800 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4801 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4802 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4803 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4804 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4805 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4806 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4807 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4808 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4809 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4810 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4811 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4812 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4813 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4814 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4815 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4816 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4817 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4818 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4819 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4820 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4821 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4822 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4823 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4824 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4825 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4826 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4827 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4828 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4829 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4830 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4831 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4832 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4833 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4834 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4835 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4836 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4837 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4838 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4839 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4840 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4841 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4842 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4843 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4844 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4845 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4846 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4847 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4848 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4849 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4850 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4851 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4852 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4853 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4854 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4855 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4856 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4857 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4858 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4859 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4860 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4861 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4862 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4863 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4864 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4865 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4866 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4867 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4868 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4869 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4870 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4871 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4872 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4873 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4874 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4875 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4876 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4877 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4878 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4879 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4880 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4881 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4882 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4883 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4884 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4885 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4886 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4887 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4888 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4889 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4890 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4891 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4892 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4893 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4894 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4895 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4896 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4897 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4898 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4899 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4900 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4901 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4902 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4903 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4904 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4905 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4906 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4907 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4908 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4909 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4910 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4911 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4912 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4913 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4914 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4915 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4916 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4917 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4918 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4919 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4920 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4921 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4922 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4923 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4924 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4925 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4926 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4927 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4928 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4929 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4930 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4931 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4932 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4933 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4934 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4935 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4936 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4937 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4938 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4939 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4940 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4941 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4942 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4943 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4944 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4945 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4946 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4947 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4948 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4949 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4950 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4951 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4952 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4953 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4954 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4955 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4956 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4957 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4958 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4959 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4960 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4961 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4962 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4963 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4964 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4965 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4966 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4967 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4968 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4969 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4970 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4971 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4972 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4973 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4974 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4975 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4976 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4977 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4978 vdd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4979 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4980 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4981 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4982 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4983 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4984 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4985 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4986 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4987 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4988 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4989 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4990 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4991 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4992 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4993 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4994 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4995 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X4996 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4997 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4998 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4999 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5000 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5001 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5002 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5003 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5004 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5005 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5006 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5007 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5008 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5009 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5010 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5011 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5012 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5013 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5014 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5015 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5016 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5017 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5018 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5019 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5020 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5021 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5022 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5023 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5024 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5025 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5026 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5027 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5028 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5029 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5030 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5031 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5032 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5033 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5034 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5035 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5036 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5037 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5038 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5039 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5040 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5041 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5042 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5043 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5044 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5045 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5046 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5047 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5048 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5049 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5050 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5051 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5052 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5053 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5054 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5055 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5056 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5057 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5058 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5059 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5060 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5061 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5062 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5063 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5064 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5065 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5066 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5067 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5068 gnd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5069 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5070 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5071 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5072 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5073 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5074 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5075 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5076 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5077 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5078 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5079 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5080 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5081 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5082 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5083 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5084 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5085 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5086 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5087 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5088 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5089 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5090 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5091 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5092 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5093 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5094 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5095 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5096 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5097 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5098 vdd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5099 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5100 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5101 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5102 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5103 tapered_buf_0/a_1650_0# tapered_buf_0/a_580_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5104 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5105 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5106 vdd tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5107 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5108 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5109 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5110 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5111 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5112 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5113 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5114 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5115 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5116 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5117 gnd tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5118 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5119 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5120 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5121 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5122 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5123 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5124 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5125 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5126 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5127 vdd tapered_buf_0/a_210_n610# pd_0/REF tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5128 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5129 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5130 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5131 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5132 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5133 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5134 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5135 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5136 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5137 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5138 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5139 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5140 gnd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5141 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5142 gnd tapered_buf_0/a_210_n610# pd_0/REF gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5143 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5144 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# vdd tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5145 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5146 vdd tapered_buf_0/a_4670_0# tapered_buf_0/a_210_n610# tapered_buf_0/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5147 pd_0/REF tapered_buf_0/a_210_n610# vdd tapered_buf_0/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5148 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5149 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5150 pd_0/REF tapered_buf_0/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5151 tapered_buf_0/a_4670_0# tapered_buf_0/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5152 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5153 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5154 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5155 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5156 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5157 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5158 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5159 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5160 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5161 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5162 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5163 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5164 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5165 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5166 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5167 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5168 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5169 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5170 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5171 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5172 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5173 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5174 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5175 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5176 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5177 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5178 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5179 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5180 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5181 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5182 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5183 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5184 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5185 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5186 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5187 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5188 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5189 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5190 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5191 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5192 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5193 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5194 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5195 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5196 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5197 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5198 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5199 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5200 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5201 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5202 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5203 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5204 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5205 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5206 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5207 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5208 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5209 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5210 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5211 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5212 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5213 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5214 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5215 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5216 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5217 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5218 vdd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5219 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5220 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5221 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5222 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5223 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5224 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5225 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5226 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5227 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5228 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5229 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5230 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5231 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5232 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5233 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5234 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5235 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5236 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5237 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5238 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5239 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5240 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5241 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5242 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5243 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5244 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5245 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5246 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5247 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5248 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5249 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5250 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5251 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5252 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5253 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5254 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5255 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5256 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5257 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5258 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5259 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5260 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5261 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5262 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5263 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5264 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5265 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5266 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5267 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5268 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5269 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5270 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5271 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5272 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5273 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5274 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5275 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5276 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5277 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5278 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5279 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5280 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5281 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5282 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5283 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5284 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5285 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5286 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5287 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5288 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5289 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5290 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5291 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5292 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5293 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5294 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5295 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5296 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5297 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5298 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5299 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5300 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5301 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5302 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5303 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5304 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5305 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5306 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5307 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5308 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5309 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5310 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5311 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5312 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5313 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5314 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5315 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5316 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5317 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5318 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5319 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5320 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5321 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5322 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5323 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5324 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5325 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5326 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5327 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5328 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5329 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5330 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5331 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5332 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5333 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5334 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5335 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5336 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5337 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5338 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5339 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5340 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5341 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5342 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5343 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5344 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5345 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5346 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5347 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5348 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5349 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5350 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5351 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5352 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5353 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5354 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5355 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5356 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5357 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5358 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5359 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5360 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5361 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5362 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5363 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5364 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5365 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5366 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5367 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5368 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5369 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5370 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5371 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5372 tapered_buf_1/a_160_230# tapered_buf_1/in tapered_buf_1/a_n10_230# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5373 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5374 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5375 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5376 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5377 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5378 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5379 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5380 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5381 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5382 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5383 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5384 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5385 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5386 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5387 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5388 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5389 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5390 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5391 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5392 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5393 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5394 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5395 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5396 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5397 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5398 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5399 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5400 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5401 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5402 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5403 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5404 tapered_buf_1/a_580_0# tapered_buf_1/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5405 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5406 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5407 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5408 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5409 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5410 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5411 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5412 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5413 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5414 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5415 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5416 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5417 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5418 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5419 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5420 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5421 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5422 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5423 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5424 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5425 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5426 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5427 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5428 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5429 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5430 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5431 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5432 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5433 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5434 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5435 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5436 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5437 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5438 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5439 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5440 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5441 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5442 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5443 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5444 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5445 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5446 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5447 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5448 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5449 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5450 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5451 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5452 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5453 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5454 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5455 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5456 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5457 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5458 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5459 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5460 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5461 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5462 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5463 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5464 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5465 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5466 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5467 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5468 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5469 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5470 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5471 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5472 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5473 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5474 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5475 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5476 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5477 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5478 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5479 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5480 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5481 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5482 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5483 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5484 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5485 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5486 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5487 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5488 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5489 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5490 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5491 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5492 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5493 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5494 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5495 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5496 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5497 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5498 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5499 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5500 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5501 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5502 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5503 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5504 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5505 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5506 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5507 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5508 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5509 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5510 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5511 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5512 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5513 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5514 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5515 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5516 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5517 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5518 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5519 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5520 gnd tapered_buf_1/a_160_n140# tapered_buf_1/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5521 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5522 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5523 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5524 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5525 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5526 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5527 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5528 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5529 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5530 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5531 vdd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5532 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5533 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5534 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5535 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5536 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5537 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5538 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5539 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5540 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5541 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5542 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5543 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5544 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5545 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5546 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5547 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5548 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5549 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5550 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5551 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5552 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5553 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5554 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5555 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5556 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5557 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5558 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5559 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5560 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5561 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5562 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5563 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5564 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5565 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5566 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5567 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5568 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5569 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5570 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5571 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5572 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5573 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5574 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5575 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5576 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5577 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5578 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5579 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5580 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5581 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5582 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5583 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5584 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5585 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5586 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5587 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5588 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5589 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5590 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5591 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5592 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5593 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5594 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5595 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5596 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5597 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5598 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5599 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5600 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5601 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5602 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5603 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5604 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5605 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5606 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5607 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5608 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5609 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5610 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5611 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5612 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5613 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5614 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5615 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5616 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5617 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5618 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5619 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5620 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5621 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5622 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5623 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5624 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5625 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5626 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5627 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5628 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5629 gnd tapered_buf_1/a_160_n140# tapered_buf_1/a_580_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5630 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5631 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5632 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5633 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5634 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5635 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5636 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5637 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5638 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5639 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5640 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5641 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5642 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5643 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5644 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5645 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5646 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5647 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5648 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5649 vdd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5650 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5651 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5652 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5653 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5654 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5655 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5656 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5657 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5658 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5659 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5660 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5661 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5662 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5663 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5664 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5665 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5666 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5667 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5668 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5669 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5670 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5671 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5672 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5673 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5674 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5675 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5676 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5677 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5678 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5679 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5680 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5681 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5682 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5683 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5684 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5685 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5686 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5687 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5688 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5689 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5690 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5691 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5692 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5693 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5694 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5695 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5696 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5697 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5698 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5699 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5700 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5701 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5702 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5703 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5704 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5705 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5706 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5707 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5708 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5709 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5710 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5711 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5712 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5713 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5714 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5715 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5716 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5717 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5718 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5719 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5720 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5721 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5722 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5723 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5724 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5725 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5726 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5727 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5728 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5729 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5730 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5731 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5732 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5733 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5734 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5735 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5736 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5737 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5738 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5739 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5740 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5741 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5742 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5743 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5744 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5745 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5746 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5747 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5748 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5749 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5750 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5751 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5752 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5753 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5754 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5755 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5756 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5757 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5758 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5759 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5760 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5761 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5762 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5763 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5764 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5765 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5766 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5767 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5768 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5769 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5770 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5771 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5772 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5773 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5774 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5775 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5776 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5777 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5778 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5779 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5780 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5781 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5782 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5783 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5784 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5785 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5786 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5787 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5788 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5789 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5790 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5791 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5792 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5793 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5794 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5795 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5796 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5797 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5798 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5799 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5800 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5801 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5802 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5803 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5804 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5805 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5806 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5807 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5808 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5809 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5810 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5811 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5812 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5813 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5814 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5815 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5816 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5817 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5818 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5819 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5820 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5821 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5822 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5823 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5824 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5825 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5826 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5827 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5828 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5829 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5830 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5831 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5832 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5833 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5834 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5835 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5836 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5837 vdd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5838 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5839 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5840 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5841 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5842 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5843 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5844 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5845 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5846 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5847 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5848 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5849 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5850 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5851 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5852 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5853 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5854 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5855 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5856 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5857 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5858 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5859 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5860 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5861 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5862 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5863 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5864 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5865 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5866 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5867 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5868 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5869 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5870 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5871 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5872 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5873 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5874 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5875 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5876 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5877 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5878 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5879 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5880 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5881 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5882 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5883 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5884 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5885 tapered_buf_1/a_580_0# tapered_buf_1/a_160_n140# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5886 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5887 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5888 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5889 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5890 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5891 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5892 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5893 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5894 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5895 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5896 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5897 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5898 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5899 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5900 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5901 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5902 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5903 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5904 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5905 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5906 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5907 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5908 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5909 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5910 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5911 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5912 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5913 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5914 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5915 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5916 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5917 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5918 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5919 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5920 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5921 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5922 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5923 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5924 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5925 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5926 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5927 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5928 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5929 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5930 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5931 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5932 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5933 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5934 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5935 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5936 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5937 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5938 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5939 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5940 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5941 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5942 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5943 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5944 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5945 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5946 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5947 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5948 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5949 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5950 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5951 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5952 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5953 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5954 tapered_buf_1/a_160_n140# tapered_buf_1/in tapered_buf_1/a_n10_n140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5955 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5956 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5957 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5958 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5959 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5960 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5961 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5962 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5963 vdd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5964 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5965 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5966 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5967 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5968 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5969 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5970 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5971 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5972 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5973 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5974 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5975 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5976 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5977 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5978 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5979 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5980 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5981 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5982 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5983 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5984 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5985 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5986 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5987 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5988 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5989 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5990 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5991 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X5992 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5993 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5994 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5995 tapered_buf_1/a_580_0# tapered_buf_1/a_160_n140# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5996 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5997 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5998 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5999 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6000 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6001 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6002 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6003 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6004 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6005 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6006 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6007 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6008 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6009 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6010 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6011 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6012 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6013 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6014 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6015 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6016 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6017 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6018 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6019 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6020 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6021 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6022 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6023 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6024 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6025 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6026 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6027 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6028 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6029 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6030 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6031 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6032 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6033 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6034 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6035 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6036 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6037 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6038 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6039 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6040 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6041 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6042 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6043 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6044 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6045 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6046 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6047 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6048 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6049 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6050 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6051 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6052 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6053 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6054 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6055 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6056 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6057 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6058 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6059 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6060 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6061 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6062 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6063 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6064 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6065 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6066 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6067 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6068 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6069 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6070 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6071 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6072 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6073 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6074 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6075 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6076 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6077 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6078 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6079 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6080 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6081 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6082 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6083 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6084 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6085 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6086 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6087 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6088 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6089 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6090 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6091 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6092 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6093 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6094 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6095 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6096 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6097 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6098 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6099 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6100 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6101 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6102 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6103 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6104 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6105 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6106 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6107 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6108 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6109 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6110 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6111 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6112 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6113 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6114 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6115 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6116 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6117 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6118 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6119 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6120 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6121 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6122 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6123 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6124 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6125 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6126 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6127 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6128 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6129 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6130 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6131 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6132 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6133 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6134 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6135 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6136 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6137 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6138 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6139 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6140 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6141 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6142 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6143 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6144 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6145 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6146 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6147 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6148 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6149 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6150 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6151 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6152 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6153 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6154 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6155 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6156 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6157 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6158 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6159 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6160 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6161 vdd tapered_buf_1/a_160_n140# tapered_buf_1/a_580_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6162 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6163 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6164 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6165 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6166 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6167 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6168 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6169 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6170 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6171 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6172 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6173 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6174 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6175 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6176 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6177 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6178 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6179 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6180 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6181 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6182 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6183 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6184 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6185 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6186 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6187 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6188 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6189 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6190 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6191 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6192 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6193 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6194 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6195 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6196 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6197 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6198 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6199 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6200 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6201 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6202 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6203 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6204 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6205 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6206 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6207 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6208 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6209 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6210 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6211 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6212 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6213 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6214 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6215 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6216 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6217 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6218 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6219 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6220 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6221 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6222 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6223 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6224 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6225 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6226 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6227 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6228 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6229 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6230 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6231 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6232 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6233 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6234 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6235 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6236 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6237 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6238 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6239 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6240 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6241 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6242 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6243 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6244 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6245 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6246 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6247 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6248 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6249 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6250 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6251 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6252 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6253 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6254 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6255 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6256 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6257 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6258 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6259 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6260 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6261 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6262 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6263 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6264 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6265 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6266 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6267 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6268 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6269 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6270 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6271 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6272 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6273 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6274 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6275 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6276 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6277 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6278 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6279 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6280 vdd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6281 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6282 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6283 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6284 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6285 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6286 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6287 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6288 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6289 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6290 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6291 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6292 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6293 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6294 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6295 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6296 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6297 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6298 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6299 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6300 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6301 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6302 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6303 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6304 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6305 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6306 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6307 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6308 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6309 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6310 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6311 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6312 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6313 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6314 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6315 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6316 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6317 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6318 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6319 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6320 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6321 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6322 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6323 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6324 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6325 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6326 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6327 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6328 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6329 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6330 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6331 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6332 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6333 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6334 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6335 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6336 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6337 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6338 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6339 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6340 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6341 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6342 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6343 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6344 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6345 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6346 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6347 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6348 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6349 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6350 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6351 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6352 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6353 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6354 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6355 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6356 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6357 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6358 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6359 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6360 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6361 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6362 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6363 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6364 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6365 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6366 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6367 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6368 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6369 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6370 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6371 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6372 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6373 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6374 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6375 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6376 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6377 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6378 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6379 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6380 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6381 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6382 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6383 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6384 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6385 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6386 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6387 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6388 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6389 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6390 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6391 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6392 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6393 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6394 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6395 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6396 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6397 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6398 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6399 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6400 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6401 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6402 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6403 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6404 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6405 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6406 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6407 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6408 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6409 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6410 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6411 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6412 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6413 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6414 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6415 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6416 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6417 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6418 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6419 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6420 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6421 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6422 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6423 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6424 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6425 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6426 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6427 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6428 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6429 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6430 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6431 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6432 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6433 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6434 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6435 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6436 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6437 vdd tapered_buf_1/a_160_n140# tapered_buf_1/a_580_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6438 tapered_buf_1/a_580_0# tapered_buf_1/a_160_n140# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6439 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6440 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6441 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6442 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6443 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6444 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6445 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6446 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6447 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6448 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6449 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6450 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6451 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6452 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6453 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6454 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6455 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6456 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6457 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6458 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6459 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6460 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6461 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6462 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6463 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6464 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6465 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6466 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6467 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6468 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6469 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6470 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6471 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6472 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6473 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6474 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6475 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6476 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6477 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6478 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6479 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6480 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6481 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6482 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6483 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6484 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6485 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6486 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6487 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6488 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6489 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6490 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6491 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6492 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6493 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6494 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6495 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6496 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6497 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6498 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6499 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6500 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6501 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6502 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6503 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6504 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6505 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6506 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6507 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6508 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6509 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6510 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6511 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6512 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6513 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6514 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6515 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6516 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6517 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6518 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6519 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6520 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6521 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6522 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6523 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6524 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6525 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6526 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6527 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6528 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6529 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6530 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6531 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6532 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6533 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6534 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6535 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6536 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6537 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6538 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6539 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6540 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6541 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6542 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6543 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6544 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6545 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6546 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6547 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6548 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6549 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6550 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6551 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6552 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6553 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6554 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6555 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6556 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6557 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6558 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6559 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6560 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6561 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6562 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6563 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6564 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6565 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6566 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6567 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6568 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6569 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6570 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6571 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6572 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6573 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6574 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6575 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6576 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6577 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6578 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6579 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6580 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6581 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6582 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6583 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6584 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6585 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6586 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6587 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6588 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6589 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6590 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6591 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6592 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6593 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6594 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6595 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6596 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6597 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6598 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6599 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6600 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6601 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6602 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6603 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6604 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6605 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6606 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6607 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6608 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6609 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6610 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6611 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6612 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6613 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6614 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6615 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6616 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6617 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6618 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6619 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6620 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6621 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6622 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6623 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6624 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6625 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6626 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6627 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6628 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6629 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6630 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6631 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6632 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6633 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6634 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6635 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6636 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6637 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6638 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6639 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6640 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6641 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6642 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6643 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6644 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6645 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6646 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6647 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6648 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6649 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6650 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6651 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6652 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6653 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6654 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6655 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6656 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6657 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6658 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6659 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6660 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6661 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6662 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6663 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6664 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6665 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6666 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6667 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6668 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6669 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6670 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6671 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6672 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6673 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6674 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6675 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6676 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6677 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6678 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6679 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6680 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6681 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6682 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6683 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6684 vdd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6685 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6686 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6687 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6688 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6689 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6690 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6691 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6692 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6693 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6694 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6695 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6696 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6697 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6698 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6699 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6700 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6701 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6702 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6703 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6704 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6705 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6706 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6707 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6708 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6709 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6710 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6711 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6712 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6713 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6714 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6715 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6716 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6717 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6718 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6719 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6720 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6721 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6722 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6723 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6724 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6725 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6726 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6727 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6728 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6729 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6730 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6731 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6732 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6733 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6734 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6735 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6736 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6737 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6738 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6739 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6740 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6741 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6742 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6743 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6744 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6745 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6746 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6747 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6748 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6749 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6750 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6751 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6752 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6753 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6754 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6755 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6756 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6757 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6758 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6759 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6760 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6761 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6762 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6763 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6764 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6765 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6766 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6767 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6768 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6769 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6770 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6771 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6772 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6773 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6774 gnd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6775 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6776 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6777 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6778 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6779 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6780 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6781 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6782 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6783 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6784 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6785 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6786 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6787 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6788 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6789 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6790 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6791 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6792 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6793 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6794 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6795 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6796 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6797 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6798 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6799 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6800 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6801 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6802 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6803 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6804 vdd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6805 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6806 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6807 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6808 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6809 tapered_buf_1/a_1650_0# tapered_buf_1/a_580_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6810 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6811 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6812 vdd tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6813 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6814 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6815 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6816 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6817 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6818 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6819 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6820 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6821 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6822 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6823 gnd tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6824 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6825 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6826 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6827 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6828 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6829 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6830 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6831 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6832 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6833 vdd tapered_buf_1/a_210_n610# pd_0/DIV tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6834 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6835 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6836 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6837 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6838 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6839 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6840 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6841 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6842 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6843 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6844 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6845 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6846 gnd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6847 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6848 gnd tapered_buf_1/a_210_n610# pd_0/DIV gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6849 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6850 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# vdd tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6851 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6852 vdd tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# tapered_buf_1/w_n70_170# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6853 pd_0/DIV tapered_buf_1/a_210_n610# vdd tapered_buf_1/w_70_n1420# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X6854 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6855 tapered_buf_1/a_210_n610# tapered_buf_1/a_4670_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6856 pd_0/DIV tapered_buf_1/a_210_n610# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6857 tapered_buf_1/a_4670_0# tapered_buf_1/a_1650_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
C0 pd_0/REF pd_0/DIV 0.51fF
C1 pd_0/tspc_r_1/Qbar1 pd_0/tspc_r_1/Qbar 0.01fF
C2 pd_0/tspc_r_1/Z3 pd_0/R 0.28fF
C3 tapered_buf_3/a_580_0# tapered_buf_3/a_210_n610# 0.84fF
C4 pd_0/tspc_r_0/Z3 pd_0/UP 0.03fF
C5 tapered_buf_3/a_160_n140# pd_0/DOWN 0.19fF
C6 tapered_buf_1/a_n10_230# tapered_buf_1/a_160_230# 0.09fF
C7 tapered_buf_1/a_1650_0# tapered_buf_1/a_210_n610# 2.89fF
C8 tapered_buf_1/a_160_n140# tapered_buf_1/a_n10_n140# 0.05fF
C9 tapered_buf_2/a_580_0# tapered_buf_2/a_1650_0# 1.27fF
C10 tapered_buf_0/in pd_0/DIV 0.02fF
C11 tapered_buf_0/a_160_n140# tapered_buf_0/a_580_0# 0.35fF
C12 tapered_buf_0/in tapered_buf_0/a_n10_n140# 0.04fF
C13 tapered_buf_0/a_580_0# tapered_buf_0/a_1650_0# 1.27fF
C14 pd_0/DOWN pd_0/R 0.36fF
C15 pd_0/tspc_r_1/Z3 pd_0/tspc_r_1/Z4 0.20fF
C16 pd_0/DIV pd_0/tspc_r_1/z5 0.04fF
C17 pd_0/tspc_r_1/Z1 pd_0/tspc_r_1/Z2 0.71fF
C18 tapered_buf_3/a_4670_0# tapered_buf_3/a_210_n610# 29.21fF
C19 tapered_buf_0/a_1650_0# tapered_buf_0/a_4670_0# 4.78fF
C20 tapered_buf_0/a_160_230# tapered_buf_0/a_580_0# 0.02fF
C21 pd_0/tspc_r_0/Z3 pd_0/tspc_r_0/Z1 0.09fF
C22 pd_0/REF pd_0/tspc_r_0/Z2 0.19fF
C23 tapered_buf_2/a_160_n140# tapered_buf_2/a_160_230# 0.17fF
C24 tapered_buf_2/a_1650_0# tapered_buf_2/a_4670_0# 4.78fF
C25 pd_0/tspc_r_0/Qbar pd_0/R 0.03fF
C26 pd_0/R pd_0/and_pd_0/Out1 0.33fF
C27 pd_0/tspc_r_1/Qbar1 pd_0/tspc_r_1/z5 0.20fF
C28 tapered_buf_0/a_210_n610# tapered_buf_0/a_580_0# 0.84fF
C29 tapered_buf_3/a_n10_230# pd_0/DOWN 0.02fF
C30 tapered_buf_1/a_n10_230# tapered_buf_1/a_n10_n140# 0.01fF
C31 tapered_buf_2/a_160_n140# tapered_buf_2/a_210_n610# 0.22fF
C32 tapered_buf_0/a_210_n610# tapered_buf_0/a_4670_0# 29.21fF
C33 pd_0/DIV pd_0/tspc_r_1/Qbar1 0.12fF
C34 tapered_buf_3/a_160_n140# tapered_buf_3/a_580_0# 0.35fF
C35 tapered_buf_0/a_160_n140# tapered_buf_0/in 0.19fF
C36 pd_0/UP pd_0/DOWN 1.06fF
C37 pd_0/tspc_r_0/Z4 pd_0/tspc_r_0/z5 0.04fF
C38 pd_0/REF pd_0/tspc_r_0/Z4 0.02fF
C39 pd_0/UP pd_0/tspc_r_0/Qbar 0.21fF
C40 tapered_buf_2/a_n10_230# tapered_buf_2/a_160_230# 0.09fF
C41 tapered_buf_2/a_1650_0# tapered_buf_2/a_210_n610# 2.89fF
C42 tapered_buf_2/a_160_n140# tapered_buf_2/a_n10_n140# 0.05fF
C43 pd_0/UP pd_0/and_pd_0/Out1 0.33fF
C44 pd_0/tspc_r_1/Z3 pd_0/DOWN 0.03fF
C45 tapered_buf_3/a_580_0# tapered_buf_3/a_1650_0# 1.27fF
C46 pd_0/R pd_0/and_pd_0/Z1 0.02fF
C47 tapered_buf_0/a_210_n610# pd_0/REF 26.29fF
C48 pd_0/REF pd_0/R 0.61fF
C49 tapered_buf_0/in tapered_buf_0/a_n10_230# 0.02fF
C50 pd_0/tspc_r_0/Z3 pd_0/tspc_r_0/z5 0.11fF
C51 tapered_buf_0/a_160_n140# tapered_buf_0/a_n10_n140# 0.05fF
C52 pd_0/tspc_r_1/Z3 pd_0/tspc_r_1/Z1 0.09fF
C53 pd_0/DIV pd_0/tspc_r_1/Z2 0.19fF
C54 tapered_buf_3/a_160_n140# tapered_buf_3/a_160_230# 0.17fF
C55 tapered_buf_3/a_1650_0# tapered_buf_3/a_4670_0# 4.78fF
C56 pd_0/REF pd_0/tspc_r_0/Z3 0.65fF
C57 tapered_buf_1/a_580_0# tapered_buf_1/a_160_230# 0.02fF
C58 pd_0/tspc_r_0/Qbar pd_0/DOWN 0.02fF
C59 pd_0/tspc_r_0/Qbar1 pd_0/R 0.30fF
C60 pd_0/DOWN pd_0/and_pd_0/Out1 0.12fF
C61 pd_0/UP pd_0/tspc_r_0/z5 0.03fF
C62 tapered_buf_2/a_n10_230# tapered_buf_2/a_n10_n140# 0.01fF
C63 pd_0/tspc_r_0/Qbar pd_0/and_pd_0/Out1 0.05fF
C64 pd_0/UP pd_0/and_pd_0/Z1 0.06fF
C65 pd_0/DIV pd_0/R 0.51fF
C66 tapered_buf_3/a_160_n140# tapered_buf_3/a_210_n610# 0.22fF
C67 tapered_buf_0/a_n10_n140# tapered_buf_0/a_n10_230# 0.01fF
C68 pd_0/tspc_r_0/Z3 pd_0/tspc_r_0/Qbar1 0.38fF
C69 tapered_buf_1/a_580_0# tapered_buf_1/a_210_n610# 0.84fF
C70 tapered_buf_1/in tapered_buf_1/a_n10_n140# 0.04fF
C71 pd_0/tspc_r_1/Z4 pd_0/tspc_r_1/z5 0.04fF
C72 pd_0/tspc_r_0/Z2 pd_0/tspc_r_0/Z4 0.14fF
C73 pd_0/tspc_r_1/Qbar1 pd_0/R 0.01fF
C74 pd_0/DIV pd_0/tspc_r_1/Z4 0.02fF
C75 pd_0/DOWN pd_0/tspc_r_1/Qbar 0.21fF
C76 tapered_buf_3/a_n10_230# tapered_buf_3/a_160_230# 0.09fF
C77 tapered_buf_3/a_1650_0# tapered_buf_3/a_210_n610# 2.89fF
C78 tapered_buf_3/a_160_n140# tapered_buf_3/a_n10_n140# 0.05fF
C79 tapered_buf_0/a_160_230# tapered_buf_0/a_160_n140# 0.17fF
C80 pd_0/REF pd_0/tspc_r_0/Z1 0.17fF
C81 pd_0/tspc_r_0/Qbar1 pd_0/UP 0.11fF
C82 tapered_buf_1/a_4670_0# tapered_buf_1/a_210_n610# 29.21fF
C83 pd_0/tspc_r_0/Z2 pd_0/R 0.21fF
C84 pd_0/DOWN pd_0/and_pd_0/Z1 0.06fF
C85 tapered_buf_1/in tapered_buf_1/a_160_n140# 0.19fF
C86 tapered_buf_2/a_210_n610# tapered_buf_2/out 26.29fF
C87 pd_0/tspc_r_0/Qbar pd_0/and_pd_0/Z1 0.02fF
C88 pd_0/tspc_r_1/Z3 pd_0/tspc_r_1/z5 0.11fF
C89 tapered_buf_2/a_n10_n140# pd_0/UP 0.04fF
C90 pd_0/and_pd_0/Out1 pd_0/and_pd_0/Z1 0.18fF
C91 tapered_buf_0/a_210_n610# tapered_buf_0/a_160_n140# 0.22fF
C92 pd_0/tspc_r_0/Z3 pd_0/tspc_r_0/Z2 0.25fF
C93 tapered_buf_2/a_580_0# tapered_buf_2/a_160_230# 0.02fF
C94 tapered_buf_0/a_160_230# tapered_buf_0/a_n10_230# 0.09fF
C95 tapered_buf_0/a_210_n610# tapered_buf_0/a_1650_0# 2.89fF
C96 pd_0/DIV pd_0/tspc_r_1/Z3 0.65fF
C97 tapered_buf_1/a_160_n140# tapered_buf_1/a_580_0# 0.35fF
C98 pd_0/DOWN pd_0/tspc_r_1/z5 0.03fF
C99 pd_0/tspc_r_1/Z2 pd_0/R 0.21fF
C100 tapered_buf_3/a_n10_230# tapered_buf_3/a_n10_n140# 0.01fF
C101 pd_0/tspc_r_0/Qbar1 pd_0/tspc_r_0/Qbar 0.01fF
C102 tapered_buf_2/a_580_0# tapered_buf_2/a_210_n610# 0.84fF
C103 pd_0/tspc_r_1/Z3 pd_0/tspc_r_1/Qbar1 0.38fF
C104 tapered_buf_2/a_160_n140# pd_0/UP 0.19fF
C105 tapered_buf_1/in tapered_buf_1/a_n10_230# 0.02fF
C106 tapered_buf_1/a_580_0# tapered_buf_1/a_1650_0# 1.27fF
C107 pd_0/tspc_r_1/Z2 pd_0/tspc_r_1/Z4 0.14fF
C108 pd_0/tspc_r_0/Z3 pd_0/tspc_r_0/Z4 0.20fF
C109 pd_0/REF pd_0/tspc_r_0/z5 0.04fF
C110 pd_0/tspc_r_0/Z1 pd_0/tspc_r_0/Z2 0.71fF
C111 tapered_buf_2/a_4670_0# tapered_buf_2/a_210_n610# 29.21fF
C112 pd_0/tspc_r_0/Z4 pd_0/tspc_r_1/Z4 0.02fF
C113 pd_0/DIV pd_0/tspc_r_1/Z1 0.17fF
C114 pd_0/tspc_r_1/Qbar1 pd_0/DOWN 0.11fF
C115 tapered_buf_1/a_160_n140# tapered_buf_1/a_160_230# 0.17fF
C116 tapered_buf_1/a_1650_0# tapered_buf_1/a_4670_0# 4.78fF
C117 pd_0/tspc_r_0/Z3 pd_0/R 0.29fF
C118 tapered_buf_3/a_210_n610# tapered_buf_3/out 26.29fF
C119 pd_0/tspc_r_0/Qbar1 pd_0/tspc_r_0/z5 0.20fF
C120 tapered_buf_3/a_n10_n140# pd_0/DOWN 0.04fF
C121 pd_0/tspc_r_0/z5 pd_0/tspc_r_1/z5 0.02fF
C122 pd_0/tspc_r_1/Z3 pd_0/tspc_r_1/Z2 0.25fF
C123 tapered_buf_3/a_580_0# tapered_buf_3/a_160_230# 0.02fF
C124 tapered_buf_2/a_n10_230# pd_0/UP 0.02fF
C125 pd_0/DIV tapered_buf_1/a_210_n610# 26.29fF
C126 pd_0/REF pd_0/tspc_r_0/Qbar1 0.12fF
C127 tapered_buf_1/a_160_n140# tapered_buf_1/a_210_n610# 0.22fF
C128 tapered_buf_2/a_160_n140# tapered_buf_2/a_580_0# 0.35fF
C129 pd_0/UP pd_0/R 0.45fF
C130 tapered_buf_1/a_n10_n140# tapered_buf_1/w_70_n1420# 0.06fF
C131 tapered_buf_1/a_210_n610# tapered_buf_1/w_70_n1420# 588.54fF
C132 tapered_buf_1/a_160_230# tapered_buf_1/w_70_n1420# 0.15fF
C133 tapered_buf_1/a_n10_230# tapered_buf_1/w_70_n1420# 0.13fF
C134 tapered_buf_1/a_4670_0# tapered_buf_1/w_70_n1420# 250.63fF
C135 tapered_buf_1/a_1650_0# tapered_buf_1/w_70_n1420# 63.04fF
C136 tapered_buf_1/a_580_0# tapered_buf_1/w_70_n1420# 16.64fF
C137 tapered_buf_1/a_160_n140# tapered_buf_1/w_70_n1420# 4.00fF
C138 tapered_buf_1/in tapered_buf_1/w_70_n1420# 1.13fF
C139 tapered_buf_0/a_n10_n140# tapered_buf_1/w_70_n1420# 0.06fF
C140 tapered_buf_0/a_210_n610# tapered_buf_1/w_70_n1420# 588.54fF
C141 tapered_buf_0/a_160_230# tapered_buf_1/w_70_n1420# 0.15fF
C142 tapered_buf_0/a_n10_230# tapered_buf_1/w_70_n1420# 0.13fF
C143 tapered_buf_0/a_4670_0# tapered_buf_1/w_70_n1420# 250.63fF
C144 tapered_buf_0/a_1650_0# tapered_buf_1/w_70_n1420# 63.04fF
C145 tapered_buf_0/a_580_0# tapered_buf_1/w_70_n1420# 16.64fF
C146 tapered_buf_0/a_160_n140# tapered_buf_1/w_70_n1420# 4.00fF
C147 tapered_buf_0/in tapered_buf_1/w_70_n1420# 1.13fF
C148 pd_0/and_pd_0/Z1 tapered_buf_1/w_70_n1420# 0.39fF
C149 pd_0/and_pd_0/Out1 tapered_buf_1/w_70_n1420# 2.22fF
C150 pd_0/tspc_r_1/z5 tapered_buf_1/w_70_n1420# 1.10fF
C151 pd_0/tspc_r_1/Z4 tapered_buf_1/w_70_n1420# 1.07fF
C152 pd_0/R tapered_buf_1/w_70_n1420# 3.06fF
C153 pd_0/tspc_r_1/Qbar tapered_buf_1/w_70_n1420# 0.79fF
C154 pd_0/tspc_r_1/Z2 tapered_buf_1/w_70_n1420# 1.22fF
C155 pd_0/tspc_r_1/Z1 tapered_buf_1/w_70_n1420# 0.67fF
C156 pd_0/DOWN tapered_buf_1/w_70_n1420# 9.89fF
C157 pd_0/tspc_r_1/Qbar1 tapered_buf_1/w_70_n1420# 1.34fF
C158 pd_0/tspc_r_1/Z3 tapered_buf_1/w_70_n1420# 2.12fF
C159 pd_0/DIV tapered_buf_1/w_70_n1420# 390.02fF
C160 pd_0/tspc_r_0/z5 tapered_buf_1/w_70_n1420# 1.10fF
C161 pd_0/tspc_r_0/Z4 tapered_buf_1/w_70_n1420# 1.07fF
C162 pd_0/tspc_r_0/Qbar tapered_buf_1/w_70_n1420# 0.88fF
C163 pd_0/tspc_r_0/Z2 tapered_buf_1/w_70_n1420# 1.22fF
C164 pd_0/tspc_r_0/Z1 tapered_buf_1/w_70_n1420# 0.67fF
C165 pd_0/UP tapered_buf_1/w_70_n1420# 5.50fF
C166 pd_0/tspc_r_0/Qbar1 tapered_buf_1/w_70_n1420# 1.34fF
C167 pd_0/tspc_r_0/Z3 tapered_buf_1/w_70_n1420# 2.12fF
C168 pd_0/REF tapered_buf_1/w_70_n1420# 388.78fF
C169 tapered_buf_3/out tapered_buf_1/w_70_n1420# 385.17fF
C170 tapered_buf_3/a_n10_n140# tapered_buf_1/w_70_n1420# 0.06fF
C171 tapered_buf_3/a_210_n610# tapered_buf_1/w_70_n1420# 588.54fF
C172 tapered_buf_3/a_160_230# tapered_buf_1/w_70_n1420# 0.15fF
C173 tapered_buf_3/a_n10_230# tapered_buf_1/w_70_n1420# 0.13fF
C174 tapered_buf_3/a_4670_0# tapered_buf_1/w_70_n1420# 250.63fF
C175 tapered_buf_3/a_1650_0# tapered_buf_1/w_70_n1420# 63.04fF
C176 tapered_buf_3/a_580_0# tapered_buf_1/w_70_n1420# 16.64fF
C177 tapered_buf_3/a_160_n140# tapered_buf_1/w_70_n1420# 4.00fF
C178 tapered_buf_2/out tapered_buf_1/w_70_n1420# 385.14fF
C179 tapered_buf_2/a_n10_n140# tapered_buf_1/w_70_n1420# 0.06fF
C180 tapered_buf_2/a_210_n610# tapered_buf_1/w_70_n1420# 588.54fF
C181 tapered_buf_2/a_160_230# tapered_buf_1/w_70_n1420# 0.15fF
C182 tapered_buf_2/a_n10_230# tapered_buf_1/w_70_n1420# 0.13fF
C183 tapered_buf_2/a_4670_0# tapered_buf_1/w_70_n1420# 250.63fF
C184 tapered_buf_2/a_1650_0# tapered_buf_1/w_70_n1420# 63.04fF
C185 tapered_buf_2/a_580_0# tapered_buf_1/w_70_n1420# 16.64fF
C186 tapered_buf_2/a_160_n140# tapered_buf_1/w_70_n1420# 4.00fF
