magic
tech sky130A
timestamp 1644270303
<< nwell >>
rect 26424 264625 26589 264812
rect 23497 264291 23832 264611
<< psubdiff >>
rect 69510 340048 70875 340158
rect 69510 338866 69629 340048
rect 70753 338866 70875 340048
rect 69510 338763 70875 338866
rect 76427 340046 77792 340156
rect 76427 338864 76546 340046
rect 77670 338864 77792 340046
rect 76427 338761 77792 338864
rect 83392 340047 84757 340157
rect 83392 338865 83511 340047
rect 84635 338865 84757 340047
rect 83392 338762 84757 338865
rect 90350 340048 91715 340158
rect 90350 338866 90469 340048
rect 91593 338866 91715 340048
rect 90350 338763 91715 338866
rect 97168 340027 98533 340137
rect 97168 338845 97287 340027
rect 98411 338845 98533 340027
rect 97168 338742 98533 338845
rect 104133 340028 105498 340138
rect 104133 338846 104252 340028
rect 105376 338846 105498 340028
rect 104133 338743 105498 338846
rect 111091 340029 112456 340139
rect 111091 338847 111210 340029
rect 112334 338847 112456 340029
rect 111091 338744 112456 338847
rect 118011 340028 119376 340138
rect 118011 338846 118130 340028
rect 119254 338846 119376 340028
rect 118011 338743 119376 338846
rect 124976 340029 126341 340139
rect 124976 338847 125095 340029
rect 126219 338847 126341 340029
rect 124976 338744 126341 338847
rect 131934 340030 133299 340140
rect 131934 338848 132053 340030
rect 133177 338848 133299 340030
rect 131934 338745 133299 338848
rect 138851 340034 140216 340144
rect 138851 338852 138970 340034
rect 140094 338852 140216 340034
rect 138851 338749 140216 338852
rect 145816 340035 147181 340145
rect 145816 338853 145935 340035
rect 147059 338853 147181 340035
rect 145816 338750 147181 338853
rect 152774 340036 154139 340146
rect 152774 338854 152893 340036
rect 154017 338854 154139 340036
rect 152774 338751 154139 338854
rect 159691 340034 161056 340144
rect 159691 338852 159810 340034
rect 160934 338852 161056 340034
rect 159691 338749 161056 338852
rect 166656 340035 168021 340145
rect 166656 338853 166775 340035
rect 167899 338853 168021 340035
rect 166656 338750 168021 338853
rect 173614 340036 174979 340146
rect 173614 338854 173733 340036
rect 174857 338854 174979 340036
rect 173614 338751 174979 338854
rect 180419 340029 181784 340139
rect 180419 338847 180538 340029
rect 181662 338847 181784 340029
rect 180419 338744 181784 338847
rect 187384 340030 188749 340140
rect 187384 338848 187503 340030
rect 188627 338848 188749 340030
rect 187384 338745 188749 338848
rect 194342 340031 195707 340141
rect 194342 338849 194461 340031
rect 195585 338849 195707 340031
rect 194342 338746 195707 338849
rect 201262 340030 202627 340140
rect 201262 338848 201381 340030
rect 202505 338848 202627 340030
rect 201262 338745 202627 338848
rect 208227 340031 209592 340141
rect 208227 338849 208346 340031
rect 209470 338849 209592 340031
rect 208227 338746 209592 338849
rect 215185 340032 216550 340142
rect 215185 338850 215304 340032
rect 216428 338850 216550 340032
rect 215185 338747 216550 338850
rect 69236 332918 70601 333028
rect 69236 331736 69355 332918
rect 70479 331736 70601 332918
rect 69236 331633 70601 331736
rect 76153 332916 77518 333026
rect 76153 331734 76272 332916
rect 77396 331734 77518 332916
rect 76153 331631 77518 331734
rect 83118 332917 84483 333027
rect 83118 331735 83237 332917
rect 84361 331735 84483 332917
rect 83118 331632 84483 331735
rect 90076 332918 91441 333028
rect 90076 331736 90195 332918
rect 91319 331736 91441 332918
rect 90076 331633 91441 331736
rect 96894 332897 98259 333007
rect 96894 331715 97013 332897
rect 98137 331715 98259 332897
rect 96894 331612 98259 331715
rect 103859 332898 105224 333008
rect 103859 331716 103978 332898
rect 105102 331716 105224 332898
rect 103859 331613 105224 331716
rect 110817 332899 112182 333009
rect 110817 331717 110936 332899
rect 112060 331717 112182 332899
rect 110817 331614 112182 331717
rect 117737 332898 119102 333008
rect 117737 331716 117856 332898
rect 118980 331716 119102 332898
rect 117737 331613 119102 331716
rect 124702 332899 126067 333009
rect 124702 331717 124821 332899
rect 125945 331717 126067 332899
rect 124702 331614 126067 331717
rect 131660 332900 133025 333010
rect 131660 331718 131779 332900
rect 132903 331718 133025 332900
rect 131660 331615 133025 331718
rect 138577 332904 139942 333014
rect 138577 331722 138696 332904
rect 139820 331722 139942 332904
rect 138577 331619 139942 331722
rect 145542 332905 146907 333015
rect 145542 331723 145661 332905
rect 146785 331723 146907 332905
rect 145542 331620 146907 331723
rect 152500 332906 153865 333016
rect 152500 331724 152619 332906
rect 153743 331724 153865 332906
rect 152500 331621 153865 331724
rect 159417 332904 160782 333014
rect 159417 331722 159536 332904
rect 160660 331722 160782 332904
rect 159417 331619 160782 331722
rect 166382 332905 167747 333015
rect 166382 331723 166501 332905
rect 167625 331723 167747 332905
rect 166382 331620 167747 331723
rect 173340 332906 174705 333016
rect 173340 331724 173459 332906
rect 174583 331724 174705 332906
rect 173340 331621 174705 331724
rect 180145 332899 181510 333009
rect 180145 331717 180264 332899
rect 181388 331717 181510 332899
rect 180145 331614 181510 331717
rect 187110 332900 188475 333010
rect 187110 331718 187229 332900
rect 188353 331718 188475 332900
rect 187110 331615 188475 331718
rect 194068 332901 195433 333011
rect 194068 331719 194187 332901
rect 195311 331719 195433 332901
rect 194068 331616 195433 331719
rect 200988 332900 202353 333010
rect 200988 331718 201107 332900
rect 202231 331718 202353 332900
rect 200988 331615 202353 331718
rect 207953 332901 209318 333011
rect 207953 331719 208072 332901
rect 209196 331719 209318 332901
rect 207953 331616 209318 331719
rect 214911 332902 216276 333012
rect 214911 331720 215030 332902
rect 216154 331720 216276 332902
rect 214911 331617 216276 331720
rect 69510 326590 70875 326700
rect 69510 325408 69629 326590
rect 70753 325408 70875 326590
rect 69510 325305 70875 325408
rect 76427 326588 77792 326698
rect 76427 325406 76546 326588
rect 77670 325406 77792 326588
rect 76427 325303 77792 325406
rect 83392 326589 84757 326699
rect 83392 325407 83511 326589
rect 84635 325407 84757 326589
rect 83392 325304 84757 325407
rect 90350 326590 91715 326700
rect 90350 325408 90469 326590
rect 91593 325408 91715 326590
rect 90350 325305 91715 325408
rect 97168 326569 98533 326679
rect 97168 325387 97287 326569
rect 98411 325387 98533 326569
rect 97168 325284 98533 325387
rect 104133 326570 105498 326680
rect 104133 325388 104252 326570
rect 105376 325388 105498 326570
rect 104133 325285 105498 325388
rect 111091 326571 112456 326681
rect 111091 325389 111210 326571
rect 112334 325389 112456 326571
rect 111091 325286 112456 325389
rect 118011 326570 119376 326680
rect 118011 325388 118130 326570
rect 119254 325388 119376 326570
rect 118011 325285 119376 325388
rect 124976 326571 126341 326681
rect 124976 325389 125095 326571
rect 126219 325389 126341 326571
rect 124976 325286 126341 325389
rect 131934 326572 133299 326682
rect 131934 325390 132053 326572
rect 133177 325390 133299 326572
rect 131934 325287 133299 325390
rect 138851 326576 140216 326686
rect 138851 325394 138970 326576
rect 140094 325394 140216 326576
rect 138851 325291 140216 325394
rect 145816 326577 147181 326687
rect 145816 325395 145935 326577
rect 147059 325395 147181 326577
rect 145816 325292 147181 325395
rect 152774 326578 154139 326688
rect 152774 325396 152893 326578
rect 154017 325396 154139 326578
rect 152774 325293 154139 325396
rect 159691 326576 161056 326686
rect 159691 325394 159810 326576
rect 160934 325394 161056 326576
rect 159691 325291 161056 325394
rect 166656 326577 168021 326687
rect 166656 325395 166775 326577
rect 167899 325395 168021 326577
rect 166656 325292 168021 325395
rect 173614 326578 174979 326688
rect 173614 325396 173733 326578
rect 174857 325396 174979 326578
rect 173614 325293 174979 325396
rect 180419 326571 181784 326681
rect 180419 325389 180538 326571
rect 181662 325389 181784 326571
rect 180419 325286 181784 325389
rect 187384 326572 188749 326682
rect 187384 325390 187503 326572
rect 188627 325390 188749 326572
rect 187384 325287 188749 325390
rect 194342 326573 195707 326683
rect 194342 325391 194461 326573
rect 195585 325391 195707 326573
rect 194342 325288 195707 325391
rect 201262 326572 202627 326682
rect 201262 325390 201381 326572
rect 202505 325390 202627 326572
rect 201262 325287 202627 325390
rect 208227 326573 209592 326683
rect 208227 325391 208346 326573
rect 209470 325391 209592 326573
rect 208227 325288 209592 325391
rect 215185 326574 216550 326684
rect 215185 325392 215304 326574
rect 216428 325392 216550 326574
rect 215185 325289 216550 325392
rect 69236 319460 70601 319570
rect 69236 318278 69355 319460
rect 70479 318278 70601 319460
rect 69236 318175 70601 318278
rect 76153 319458 77518 319568
rect 76153 318276 76272 319458
rect 77396 318276 77518 319458
rect 76153 318173 77518 318276
rect 83118 319459 84483 319569
rect 83118 318277 83237 319459
rect 84361 318277 84483 319459
rect 83118 318174 84483 318277
rect 90076 319460 91441 319570
rect 90076 318278 90195 319460
rect 91319 318278 91441 319460
rect 90076 318175 91441 318278
rect 96894 319439 98259 319549
rect 96894 318257 97013 319439
rect 98137 318257 98259 319439
rect 96894 318154 98259 318257
rect 103859 319440 105224 319550
rect 103859 318258 103978 319440
rect 105102 318258 105224 319440
rect 103859 318155 105224 318258
rect 110817 319441 112182 319551
rect 110817 318259 110936 319441
rect 112060 318259 112182 319441
rect 110817 318156 112182 318259
rect 117737 319440 119102 319550
rect 117737 318258 117856 319440
rect 118980 318258 119102 319440
rect 117737 318155 119102 318258
rect 124702 319441 126067 319551
rect 124702 318259 124821 319441
rect 125945 318259 126067 319441
rect 124702 318156 126067 318259
rect 131660 319442 133025 319552
rect 131660 318260 131779 319442
rect 132903 318260 133025 319442
rect 131660 318157 133025 318260
rect 138577 319446 139942 319556
rect 138577 318264 138696 319446
rect 139820 318264 139942 319446
rect 138577 318161 139942 318264
rect 145542 319447 146907 319557
rect 145542 318265 145661 319447
rect 146785 318265 146907 319447
rect 145542 318162 146907 318265
rect 152500 319448 153865 319558
rect 152500 318266 152619 319448
rect 153743 318266 153865 319448
rect 152500 318163 153865 318266
rect 159417 319446 160782 319556
rect 159417 318264 159536 319446
rect 160660 318264 160782 319446
rect 159417 318161 160782 318264
rect 166382 319447 167747 319557
rect 166382 318265 166501 319447
rect 167625 318265 167747 319447
rect 166382 318162 167747 318265
rect 173340 319448 174705 319558
rect 173340 318266 173459 319448
rect 174583 318266 174705 319448
rect 173340 318163 174705 318266
rect 180145 319441 181510 319551
rect 180145 318259 180264 319441
rect 181388 318259 181510 319441
rect 180145 318156 181510 318259
rect 187110 319442 188475 319552
rect 187110 318260 187229 319442
rect 188353 318260 188475 319442
rect 187110 318157 188475 318260
rect 194068 319443 195433 319553
rect 194068 318261 194187 319443
rect 195311 318261 195433 319443
rect 194068 318158 195433 318261
rect 200988 319442 202353 319552
rect 200988 318260 201107 319442
rect 202231 318260 202353 319442
rect 200988 318157 202353 318260
rect 207953 319443 209318 319553
rect 207953 318261 208072 319443
rect 209196 318261 209318 319443
rect 207953 318158 209318 318261
rect 214911 319444 216276 319554
rect 214911 318262 215030 319444
rect 216154 318262 216276 319444
rect 214911 318159 216276 318262
rect 20875 312321 22240 312431
rect 20875 311139 20994 312321
rect 22118 311139 22240 312321
rect 20875 311036 22240 311139
rect 27833 312322 29198 312432
rect 27833 311140 27952 312322
rect 29076 311140 29198 312322
rect 27833 311037 29198 311140
rect 34753 312321 36118 312431
rect 34753 311139 34872 312321
rect 35996 311139 36118 312321
rect 34753 311036 36118 311139
rect 41718 312322 43083 312432
rect 41718 311140 41837 312322
rect 42961 311140 43083 312322
rect 41718 311037 43083 311140
rect 48676 312323 50041 312433
rect 48676 311141 48795 312323
rect 49919 311141 50041 312323
rect 48676 311038 50041 311141
rect 55593 312327 56958 312437
rect 55593 311145 55712 312327
rect 56836 311145 56958 312327
rect 55593 311042 56958 311145
rect 62558 312328 63923 312438
rect 62558 311146 62677 312328
rect 63801 311146 63923 312328
rect 62558 311043 63923 311146
rect 69516 312329 70881 312439
rect 69516 311147 69635 312329
rect 70759 311147 70881 312329
rect 69516 311044 70881 311147
rect 76433 312327 77798 312437
rect 76433 311145 76552 312327
rect 77676 311145 77798 312327
rect 76433 311042 77798 311145
rect 83398 312328 84763 312438
rect 83398 311146 83517 312328
rect 84641 311146 84763 312328
rect 83398 311043 84763 311146
rect 90356 312329 91721 312439
rect 90356 311147 90475 312329
rect 91599 311147 91721 312329
rect 90356 311044 91721 311147
rect 97174 312308 98539 312418
rect 97174 311126 97293 312308
rect 98417 311126 98539 312308
rect 97174 311023 98539 311126
rect 104139 312309 105504 312419
rect 104139 311127 104258 312309
rect 105382 311127 105504 312309
rect 104139 311024 105504 311127
rect 111097 312310 112462 312420
rect 111097 311128 111216 312310
rect 112340 311128 112462 312310
rect 111097 311025 112462 311128
rect 118017 312309 119382 312419
rect 118017 311127 118136 312309
rect 119260 311127 119382 312309
rect 118017 311024 119382 311127
rect 124982 312310 126347 312420
rect 124982 311128 125101 312310
rect 126225 311128 126347 312310
rect 124982 311025 126347 311128
rect 131940 312311 133305 312421
rect 131940 311129 132059 312311
rect 133183 311129 133305 312311
rect 131940 311026 133305 311129
rect 138857 312315 140222 312425
rect 138857 311133 138976 312315
rect 140100 311133 140222 312315
rect 138857 311030 140222 311133
rect 145822 312316 147187 312426
rect 145822 311134 145941 312316
rect 147065 311134 147187 312316
rect 145822 311031 147187 311134
rect 152780 312317 154145 312427
rect 152780 311135 152899 312317
rect 154023 311135 154145 312317
rect 152780 311032 154145 311135
rect 159697 312315 161062 312425
rect 159697 311133 159816 312315
rect 160940 311133 161062 312315
rect 159697 311030 161062 311133
rect 166662 312316 168027 312426
rect 166662 311134 166781 312316
rect 167905 311134 168027 312316
rect 166662 311031 168027 311134
rect 173620 312317 174985 312427
rect 173620 311135 173739 312317
rect 174863 311135 174985 312317
rect 173620 311032 174985 311135
rect 180425 312310 181790 312420
rect 180425 311128 180544 312310
rect 181668 311128 181790 312310
rect 180425 311025 181790 311128
rect 187390 312311 188755 312421
rect 187390 311129 187509 312311
rect 188633 311129 188755 312311
rect 187390 311026 188755 311129
rect 194348 312312 195713 312422
rect 194348 311130 194467 312312
rect 195591 311130 195713 312312
rect 194348 311027 195713 311130
rect 201268 312311 202633 312421
rect 201268 311129 201387 312311
rect 202511 311129 202633 312311
rect 201268 311026 202633 311129
rect 208233 312312 209598 312422
rect 208233 311130 208352 312312
rect 209476 311130 209598 312312
rect 208233 311027 209598 311130
rect 215191 312313 216556 312423
rect 215191 311131 215310 312313
rect 216434 311131 216556 312313
rect 215191 311028 216556 311131
rect 20601 305191 21966 305301
rect 20601 304009 20720 305191
rect 21844 304009 21966 305191
rect 20601 303906 21966 304009
rect 27559 305192 28924 305302
rect 27559 304010 27678 305192
rect 28802 304010 28924 305192
rect 27559 303907 28924 304010
rect 34479 305191 35844 305301
rect 34479 304009 34598 305191
rect 35722 304009 35844 305191
rect 34479 303906 35844 304009
rect 41444 305192 42809 305302
rect 41444 304010 41563 305192
rect 42687 304010 42809 305192
rect 41444 303907 42809 304010
rect 48402 305193 49767 305303
rect 48402 304011 48521 305193
rect 49645 304011 49767 305193
rect 48402 303908 49767 304011
rect 55319 305197 56684 305307
rect 55319 304015 55438 305197
rect 56562 304015 56684 305197
rect 55319 303912 56684 304015
rect 62284 305198 63649 305308
rect 62284 304016 62403 305198
rect 63527 304016 63649 305198
rect 62284 303913 63649 304016
rect 69242 305199 70607 305309
rect 69242 304017 69361 305199
rect 70485 304017 70607 305199
rect 69242 303914 70607 304017
rect 76159 305197 77524 305307
rect 76159 304015 76278 305197
rect 77402 304015 77524 305197
rect 76159 303912 77524 304015
rect 83124 305198 84489 305308
rect 83124 304016 83243 305198
rect 84367 304016 84489 305198
rect 83124 303913 84489 304016
rect 90082 305199 91447 305309
rect 90082 304017 90201 305199
rect 91325 304017 91447 305199
rect 90082 303914 91447 304017
rect 96900 305178 98265 305288
rect 96900 303996 97019 305178
rect 98143 303996 98265 305178
rect 96900 303893 98265 303996
rect 103865 305179 105230 305289
rect 103865 303997 103984 305179
rect 105108 303997 105230 305179
rect 103865 303894 105230 303997
rect 110823 305180 112188 305290
rect 110823 303998 110942 305180
rect 112066 303998 112188 305180
rect 110823 303895 112188 303998
rect 117743 305179 119108 305289
rect 117743 303997 117862 305179
rect 118986 303997 119108 305179
rect 117743 303894 119108 303997
rect 124708 305180 126073 305290
rect 124708 303998 124827 305180
rect 125951 303998 126073 305180
rect 124708 303895 126073 303998
rect 131666 305181 133031 305291
rect 131666 303999 131785 305181
rect 132909 303999 133031 305181
rect 131666 303896 133031 303999
rect 138583 305185 139948 305295
rect 138583 304003 138702 305185
rect 139826 304003 139948 305185
rect 138583 303900 139948 304003
rect 145548 305186 146913 305296
rect 145548 304004 145667 305186
rect 146791 304004 146913 305186
rect 145548 303901 146913 304004
rect 152506 305187 153871 305297
rect 152506 304005 152625 305187
rect 153749 304005 153871 305187
rect 152506 303902 153871 304005
rect 159423 305185 160788 305295
rect 159423 304003 159542 305185
rect 160666 304003 160788 305185
rect 159423 303900 160788 304003
rect 166388 305186 167753 305296
rect 166388 304004 166507 305186
rect 167631 304004 167753 305186
rect 166388 303901 167753 304004
rect 173346 305187 174711 305297
rect 173346 304005 173465 305187
rect 174589 304005 174711 305187
rect 173346 303902 174711 304005
rect 180151 305180 181516 305290
rect 180151 303998 180270 305180
rect 181394 303998 181516 305180
rect 180151 303895 181516 303998
rect 187116 305181 188481 305291
rect 187116 303999 187235 305181
rect 188359 303999 188481 305181
rect 187116 303896 188481 303999
rect 194074 305182 195439 305292
rect 194074 304000 194193 305182
rect 195317 304000 195439 305182
rect 194074 303897 195439 304000
rect 200994 305181 202359 305291
rect 200994 303999 201113 305181
rect 202237 303999 202359 305181
rect 200994 303896 202359 303999
rect 207959 305182 209324 305292
rect 207959 304000 208078 305182
rect 209202 304000 209324 305182
rect 207959 303897 209324 304000
rect 214917 305183 216282 305293
rect 214917 304001 215036 305183
rect 216160 304001 216282 305183
rect 214917 303898 216282 304001
rect 20964 295962 22329 296072
rect 20964 294780 21083 295962
rect 22207 294780 22329 295962
rect 20964 294677 22329 294780
rect 27922 295963 29287 296073
rect 27922 294781 28041 295963
rect 29165 294781 29287 295963
rect 27922 294678 29287 294781
rect 34842 295962 36207 296072
rect 34842 294780 34961 295962
rect 36085 294780 36207 295962
rect 34842 294677 36207 294780
rect 41807 295963 43172 296073
rect 41807 294781 41926 295963
rect 43050 294781 43172 295963
rect 41807 294678 43172 294781
rect 48765 295964 50130 296074
rect 48765 294782 48884 295964
rect 50008 294782 50130 295964
rect 48765 294679 50130 294782
rect 55682 295968 57047 296078
rect 55682 294786 55801 295968
rect 56925 294786 57047 295968
rect 55682 294683 57047 294786
rect 62647 295969 64012 296079
rect 62647 294787 62766 295969
rect 63890 294787 64012 295969
rect 62647 294684 64012 294787
rect 69605 295970 70970 296080
rect 69605 294788 69724 295970
rect 70848 294788 70970 295970
rect 69605 294685 70970 294788
rect 76522 295968 77887 296078
rect 76522 294786 76641 295968
rect 77765 294786 77887 295968
rect 76522 294683 77887 294786
rect 83487 295969 84852 296079
rect 83487 294787 83606 295969
rect 84730 294787 84852 295969
rect 83487 294684 84852 294787
rect 90445 295970 91810 296080
rect 90445 294788 90564 295970
rect 91688 294788 91810 295970
rect 90445 294685 91810 294788
rect 97263 295949 98628 296059
rect 97263 294767 97382 295949
rect 98506 294767 98628 295949
rect 97263 294664 98628 294767
rect 104228 295950 105593 296060
rect 104228 294768 104347 295950
rect 105471 294768 105593 295950
rect 104228 294665 105593 294768
rect 111186 295951 112551 296061
rect 111186 294769 111305 295951
rect 112429 294769 112551 295951
rect 111186 294666 112551 294769
rect 118106 295950 119471 296060
rect 118106 294768 118225 295950
rect 119349 294768 119471 295950
rect 118106 294665 119471 294768
rect 125071 295951 126436 296061
rect 125071 294769 125190 295951
rect 126314 294769 126436 295951
rect 125071 294666 126436 294769
rect 132029 295952 133394 296062
rect 132029 294770 132148 295952
rect 133272 294770 133394 295952
rect 132029 294667 133394 294770
rect 138946 295956 140311 296066
rect 138946 294774 139065 295956
rect 140189 294774 140311 295956
rect 138946 294671 140311 294774
rect 145911 295957 147276 296067
rect 145911 294775 146030 295957
rect 147154 294775 147276 295957
rect 145911 294672 147276 294775
rect 152869 295958 154234 296068
rect 152869 294776 152988 295958
rect 154112 294776 154234 295958
rect 152869 294673 154234 294776
rect 159786 295956 161151 296066
rect 159786 294774 159905 295956
rect 161029 294774 161151 295956
rect 159786 294671 161151 294774
rect 166751 295957 168116 296067
rect 166751 294775 166870 295957
rect 167994 294775 168116 295957
rect 166751 294672 168116 294775
rect 173709 295958 175074 296068
rect 173709 294776 173828 295958
rect 174952 294776 175074 295958
rect 173709 294673 175074 294776
rect 180514 295951 181879 296061
rect 180514 294769 180633 295951
rect 181757 294769 181879 295951
rect 180514 294666 181879 294769
rect 187479 295952 188844 296062
rect 187479 294770 187598 295952
rect 188722 294770 188844 295952
rect 187479 294667 188844 294770
rect 194437 295953 195802 296063
rect 194437 294771 194556 295953
rect 195680 294771 195802 295953
rect 194437 294668 195802 294771
rect 201357 295952 202722 296062
rect 201357 294770 201476 295952
rect 202600 294770 202722 295952
rect 201357 294667 202722 294770
rect 208322 295953 209687 296063
rect 208322 294771 208441 295953
rect 209565 294771 209687 295953
rect 208322 294668 209687 294771
rect 215280 295954 216645 296064
rect 215280 294772 215399 295954
rect 216523 294772 216645 295954
rect 215280 294669 216645 294772
rect 222197 295958 223562 296068
rect 222197 294776 222316 295958
rect 223440 294776 223562 295958
rect 222197 294673 223562 294776
rect 229162 295959 230527 296069
rect 229162 294777 229281 295959
rect 230405 294777 230527 295959
rect 229162 294674 230527 294777
rect 236120 295960 237485 296070
rect 236120 294778 236239 295960
rect 237363 294778 237485 295960
rect 236120 294675 237485 294778
rect 243037 295958 244402 296068
rect 243037 294776 243156 295958
rect 244280 294776 244402 295958
rect 243037 294673 244402 294776
rect 250002 295959 251367 296069
rect 250002 294777 250121 295959
rect 251245 294777 251367 295959
rect 250002 294674 251367 294777
rect 256960 295960 258325 296070
rect 256960 294778 257079 295960
rect 258203 294778 258325 295960
rect 256960 294675 258325 294778
rect 264100 295960 265465 296070
rect 264100 294778 264219 295960
rect 265343 294778 265465 295960
rect 264100 294675 265465 294778
rect 271058 295961 272423 296071
rect 271058 294779 271177 295961
rect 272301 294779 272423 295961
rect 271058 294676 272423 294779
rect 278194 295951 279559 296061
rect 278194 294769 278313 295951
rect 279437 294769 279559 295951
rect 278194 294666 279559 294769
rect 20690 288832 22055 288942
rect 20690 287650 20809 288832
rect 21933 287650 22055 288832
rect 20690 287547 22055 287650
rect 27648 288833 29013 288943
rect 27648 287651 27767 288833
rect 28891 287651 29013 288833
rect 27648 287548 29013 287651
rect 34568 288832 35933 288942
rect 34568 287650 34687 288832
rect 35811 287650 35933 288832
rect 34568 287547 35933 287650
rect 41533 288833 42898 288943
rect 41533 287651 41652 288833
rect 42776 287651 42898 288833
rect 41533 287548 42898 287651
rect 48491 288834 49856 288944
rect 48491 287652 48610 288834
rect 49734 287652 49856 288834
rect 48491 287549 49856 287652
rect 55408 288838 56773 288948
rect 55408 287656 55527 288838
rect 56651 287656 56773 288838
rect 55408 287553 56773 287656
rect 62373 288839 63738 288949
rect 62373 287657 62492 288839
rect 63616 287657 63738 288839
rect 62373 287554 63738 287657
rect 69331 288840 70696 288950
rect 69331 287658 69450 288840
rect 70574 287658 70696 288840
rect 69331 287555 70696 287658
rect 76248 288838 77613 288948
rect 76248 287656 76367 288838
rect 77491 287656 77613 288838
rect 76248 287553 77613 287656
rect 83213 288839 84578 288949
rect 83213 287657 83332 288839
rect 84456 287657 84578 288839
rect 83213 287554 84578 287657
rect 90171 288840 91536 288950
rect 90171 287658 90290 288840
rect 91414 287658 91536 288840
rect 90171 287555 91536 287658
rect 96989 288819 98354 288929
rect 96989 287637 97108 288819
rect 98232 287637 98354 288819
rect 96989 287534 98354 287637
rect 103954 288820 105319 288930
rect 103954 287638 104073 288820
rect 105197 287638 105319 288820
rect 103954 287535 105319 287638
rect 110912 288821 112277 288931
rect 110912 287639 111031 288821
rect 112155 287639 112277 288821
rect 110912 287536 112277 287639
rect 117832 288820 119197 288930
rect 117832 287638 117951 288820
rect 119075 287638 119197 288820
rect 117832 287535 119197 287638
rect 124797 288821 126162 288931
rect 124797 287639 124916 288821
rect 126040 287639 126162 288821
rect 124797 287536 126162 287639
rect 131755 288822 133120 288932
rect 131755 287640 131874 288822
rect 132998 287640 133120 288822
rect 131755 287537 133120 287640
rect 138672 288826 140037 288936
rect 138672 287644 138791 288826
rect 139915 287644 140037 288826
rect 138672 287541 140037 287644
rect 145637 288827 147002 288937
rect 145637 287645 145756 288827
rect 146880 287645 147002 288827
rect 145637 287542 147002 287645
rect 152595 288828 153960 288938
rect 152595 287646 152714 288828
rect 153838 287646 153960 288828
rect 152595 287543 153960 287646
rect 159512 288826 160877 288936
rect 159512 287644 159631 288826
rect 160755 287644 160877 288826
rect 159512 287541 160877 287644
rect 166477 288827 167842 288937
rect 166477 287645 166596 288827
rect 167720 287645 167842 288827
rect 166477 287542 167842 287645
rect 173435 288828 174800 288938
rect 173435 287646 173554 288828
rect 174678 287646 174800 288828
rect 173435 287543 174800 287646
rect 180240 288821 181605 288931
rect 180240 287639 180359 288821
rect 181483 287639 181605 288821
rect 180240 287536 181605 287639
rect 187205 288822 188570 288932
rect 187205 287640 187324 288822
rect 188448 287640 188570 288822
rect 187205 287537 188570 287640
rect 194163 288823 195528 288933
rect 194163 287641 194282 288823
rect 195406 287641 195528 288823
rect 194163 287538 195528 287641
rect 201083 288822 202448 288932
rect 201083 287640 201202 288822
rect 202326 287640 202448 288822
rect 201083 287537 202448 287640
rect 208048 288823 209413 288933
rect 208048 287641 208167 288823
rect 209291 287641 209413 288823
rect 208048 287538 209413 287641
rect 215006 288824 216371 288934
rect 215006 287642 215125 288824
rect 216249 287642 216371 288824
rect 215006 287539 216371 287642
rect 221923 288828 223288 288938
rect 221923 287646 222042 288828
rect 223166 287646 223288 288828
rect 221923 287543 223288 287646
rect 228888 288829 230253 288939
rect 228888 287647 229007 288829
rect 230131 287647 230253 288829
rect 228888 287544 230253 287647
rect 235846 288830 237211 288940
rect 235846 287648 235965 288830
rect 237089 287648 237211 288830
rect 235846 287545 237211 287648
rect 242763 288828 244128 288938
rect 242763 287646 242882 288828
rect 244006 287646 244128 288828
rect 242763 287543 244128 287646
rect 249728 288829 251093 288939
rect 249728 287647 249847 288829
rect 250971 287647 251093 288829
rect 249728 287544 251093 287647
rect 256686 288830 258051 288940
rect 256686 287648 256805 288830
rect 257929 287648 258051 288830
rect 256686 287545 258051 287648
rect 263826 288830 265191 288940
rect 263826 287648 263945 288830
rect 265069 287648 265191 288830
rect 263826 287545 265191 287648
rect 270784 288831 272149 288941
rect 270784 287649 270903 288831
rect 272027 287649 272149 288831
rect 270784 287546 272149 287649
rect 277920 288821 279285 288931
rect 277920 287639 278039 288821
rect 279163 287639 279285 288821
rect 277920 287536 279285 287639
rect 20798 282419 22163 282529
rect 20798 281237 20917 282419
rect 22041 281237 22163 282419
rect 20798 281134 22163 281237
rect 27756 282420 29121 282530
rect 27756 281238 27875 282420
rect 28999 281238 29121 282420
rect 27756 281135 29121 281238
rect 34676 282419 36041 282529
rect 34676 281237 34795 282419
rect 35919 281237 36041 282419
rect 34676 281134 36041 281237
rect 41641 282420 43006 282530
rect 41641 281238 41760 282420
rect 42884 281238 43006 282420
rect 41641 281135 43006 281238
rect 48599 282421 49964 282531
rect 48599 281239 48718 282421
rect 49842 281239 49964 282421
rect 48599 281136 49964 281239
rect 55516 282425 56881 282535
rect 55516 281243 55635 282425
rect 56759 281243 56881 282425
rect 55516 281140 56881 281243
rect 62481 282426 63846 282536
rect 62481 281244 62600 282426
rect 63724 281244 63846 282426
rect 62481 281141 63846 281244
rect 69439 282427 70804 282537
rect 69439 281245 69558 282427
rect 70682 281245 70804 282427
rect 69439 281142 70804 281245
rect 76356 282425 77721 282535
rect 76356 281243 76475 282425
rect 77599 281243 77721 282425
rect 76356 281140 77721 281243
rect 83321 282426 84686 282536
rect 83321 281244 83440 282426
rect 84564 281244 84686 282426
rect 83321 281141 84686 281244
rect 90279 282427 91644 282537
rect 90279 281245 90398 282427
rect 91522 281245 91644 282427
rect 90279 281142 91644 281245
rect 97097 282406 98462 282516
rect 97097 281224 97216 282406
rect 98340 281224 98462 282406
rect 97097 281121 98462 281224
rect 104062 282407 105427 282517
rect 104062 281225 104181 282407
rect 105305 281225 105427 282407
rect 104062 281122 105427 281225
rect 111020 282408 112385 282518
rect 111020 281226 111139 282408
rect 112263 281226 112385 282408
rect 111020 281123 112385 281226
rect 117940 282407 119305 282517
rect 117940 281225 118059 282407
rect 119183 281225 119305 282407
rect 117940 281122 119305 281225
rect 124905 282408 126270 282518
rect 124905 281226 125024 282408
rect 126148 281226 126270 282408
rect 124905 281123 126270 281226
rect 131863 282409 133228 282519
rect 131863 281227 131982 282409
rect 133106 281227 133228 282409
rect 131863 281124 133228 281227
rect 138780 282413 140145 282523
rect 138780 281231 138899 282413
rect 140023 281231 140145 282413
rect 138780 281128 140145 281231
rect 145745 282414 147110 282524
rect 145745 281232 145864 282414
rect 146988 281232 147110 282414
rect 145745 281129 147110 281232
rect 152703 282415 154068 282525
rect 152703 281233 152822 282415
rect 153946 281233 154068 282415
rect 152703 281130 154068 281233
rect 159620 282413 160985 282523
rect 159620 281231 159739 282413
rect 160863 281231 160985 282413
rect 159620 281128 160985 281231
rect 166585 282414 167950 282524
rect 166585 281232 166704 282414
rect 167828 281232 167950 282414
rect 166585 281129 167950 281232
rect 173543 282415 174908 282525
rect 173543 281233 173662 282415
rect 174786 281233 174908 282415
rect 173543 281130 174908 281233
rect 180348 282408 181713 282518
rect 180348 281226 180467 282408
rect 181591 281226 181713 282408
rect 180348 281123 181713 281226
rect 187313 282409 188678 282519
rect 187313 281227 187432 282409
rect 188556 281227 188678 282409
rect 187313 281124 188678 281227
rect 194271 282410 195636 282520
rect 194271 281228 194390 282410
rect 195514 281228 195636 282410
rect 194271 281125 195636 281228
rect 201191 282409 202556 282519
rect 201191 281227 201310 282409
rect 202434 281227 202556 282409
rect 201191 281124 202556 281227
rect 208156 282410 209521 282520
rect 208156 281228 208275 282410
rect 209399 281228 209521 282410
rect 208156 281125 209521 281228
rect 215114 282411 216479 282521
rect 215114 281229 215233 282411
rect 216357 281229 216479 282411
rect 215114 281126 216479 281229
rect 222031 282415 223396 282525
rect 222031 281233 222150 282415
rect 223274 281233 223396 282415
rect 222031 281130 223396 281233
rect 228996 282416 230361 282526
rect 228996 281234 229115 282416
rect 230239 281234 230361 282416
rect 228996 281131 230361 281234
rect 235954 282417 237319 282527
rect 235954 281235 236073 282417
rect 237197 281235 237319 282417
rect 235954 281132 237319 281235
rect 242871 282415 244236 282525
rect 242871 281233 242990 282415
rect 244114 281233 244236 282415
rect 242871 281130 244236 281233
rect 249836 282416 251201 282526
rect 249836 281234 249955 282416
rect 251079 281234 251201 282416
rect 249836 281131 251201 281234
rect 256794 282417 258159 282527
rect 256794 281235 256913 282417
rect 258037 281235 258159 282417
rect 256794 281132 258159 281235
rect 263934 282417 265299 282527
rect 263934 281235 264053 282417
rect 265177 281235 265299 282417
rect 263934 281132 265299 281235
rect 270892 282418 272257 282528
rect 270892 281236 271011 282418
rect 272135 281236 272257 282418
rect 270892 281133 272257 281236
rect 278028 282408 279393 282518
rect 278028 281226 278147 282408
rect 279271 281226 279393 282408
rect 278028 281123 279393 281226
rect 69656 273562 71021 273672
rect 69656 272380 69775 273562
rect 70899 272380 71021 273562
rect 69656 272277 71021 272380
rect 76573 273560 77938 273670
rect 76573 272378 76692 273560
rect 77816 272378 77938 273560
rect 76573 272275 77938 272378
rect 83538 273561 84903 273671
rect 83538 272379 83657 273561
rect 84781 272379 84903 273561
rect 83538 272276 84903 272379
rect 90496 273562 91861 273672
rect 90496 272380 90615 273562
rect 91739 272380 91861 273562
rect 90496 272277 91861 272380
rect 97314 273541 98679 273651
rect 97314 272359 97433 273541
rect 98557 272359 98679 273541
rect 97314 272256 98679 272359
rect 104279 273542 105644 273652
rect 104279 272360 104398 273542
rect 105522 272360 105644 273542
rect 104279 272257 105644 272360
rect 111237 273543 112602 273653
rect 111237 272361 111356 273543
rect 112480 272361 112602 273543
rect 111237 272258 112602 272361
rect 118157 273542 119522 273652
rect 118157 272360 118276 273542
rect 119400 272360 119522 273542
rect 118157 272257 119522 272360
rect 125122 273543 126487 273653
rect 125122 272361 125241 273543
rect 126365 272361 126487 273543
rect 125122 272258 126487 272361
rect 132080 273544 133445 273654
rect 132080 272362 132199 273544
rect 133323 272362 133445 273544
rect 132080 272259 133445 272362
rect 138997 273548 140362 273658
rect 138997 272366 139116 273548
rect 140240 272366 140362 273548
rect 138997 272263 140362 272366
rect 145962 273549 147327 273659
rect 145962 272367 146081 273549
rect 147205 272367 147327 273549
rect 145962 272264 147327 272367
rect 152920 273550 154285 273660
rect 152920 272368 153039 273550
rect 154163 272368 154285 273550
rect 152920 272265 154285 272368
rect 159837 273548 161202 273658
rect 159837 272366 159956 273548
rect 161080 272366 161202 273548
rect 159837 272263 161202 272366
rect 166802 273549 168167 273659
rect 166802 272367 166921 273549
rect 168045 272367 168167 273549
rect 166802 272264 168167 272367
rect 173760 273550 175125 273660
rect 173760 272368 173879 273550
rect 175003 272368 175125 273550
rect 173760 272265 175125 272368
rect 180565 273543 181930 273653
rect 180565 272361 180684 273543
rect 181808 272361 181930 273543
rect 180565 272258 181930 272361
rect 187530 273544 188895 273654
rect 187530 272362 187649 273544
rect 188773 272362 188895 273544
rect 187530 272259 188895 272362
rect 194488 273545 195853 273655
rect 194488 272363 194607 273545
rect 195731 272363 195853 273545
rect 194488 272260 195853 272363
rect 201408 273544 202773 273654
rect 201408 272362 201527 273544
rect 202651 272362 202773 273544
rect 201408 272259 202773 272362
rect 208373 273545 209738 273655
rect 208373 272363 208492 273545
rect 209616 272363 209738 273545
rect 208373 272260 209738 272363
rect 215331 273546 216696 273656
rect 215331 272364 215450 273546
rect 216574 272364 216696 273546
rect 215331 272261 216696 272364
rect 222248 273550 223613 273660
rect 222248 272368 222367 273550
rect 223491 272368 223613 273550
rect 222248 272265 223613 272368
rect 69382 266432 70747 266542
rect 69382 265250 69501 266432
rect 70625 265250 70747 266432
rect 69382 265147 70747 265250
rect 76299 266430 77664 266540
rect 76299 265248 76418 266430
rect 77542 265248 77664 266430
rect 76299 265145 77664 265248
rect 83264 266431 84629 266541
rect 83264 265249 83383 266431
rect 84507 265249 84629 266431
rect 83264 265146 84629 265249
rect 90222 266432 91587 266542
rect 90222 265250 90341 266432
rect 91465 265250 91587 266432
rect 90222 265147 91587 265250
rect 97040 266411 98405 266521
rect 97040 265229 97159 266411
rect 98283 265229 98405 266411
rect 97040 265126 98405 265229
rect 104005 266412 105370 266522
rect 104005 265230 104124 266412
rect 105248 265230 105370 266412
rect 104005 265127 105370 265230
rect 110963 266413 112328 266523
rect 110963 265231 111082 266413
rect 112206 265231 112328 266413
rect 110963 265128 112328 265231
rect 117883 266412 119248 266522
rect 117883 265230 118002 266412
rect 119126 265230 119248 266412
rect 117883 265127 119248 265230
rect 124848 266413 126213 266523
rect 124848 265231 124967 266413
rect 126091 265231 126213 266413
rect 124848 265128 126213 265231
rect 131806 266414 133171 266524
rect 131806 265232 131925 266414
rect 133049 265232 133171 266414
rect 131806 265129 133171 265232
rect 138723 266418 140088 266528
rect 138723 265236 138842 266418
rect 139966 265236 140088 266418
rect 138723 265133 140088 265236
rect 145688 266419 147053 266529
rect 145688 265237 145807 266419
rect 146931 265237 147053 266419
rect 145688 265134 147053 265237
rect 152646 266420 154011 266530
rect 152646 265238 152765 266420
rect 153889 265238 154011 266420
rect 152646 265135 154011 265238
rect 159563 266418 160928 266528
rect 159563 265236 159682 266418
rect 160806 265236 160928 266418
rect 159563 265133 160928 265236
rect 166528 266419 167893 266529
rect 166528 265237 166647 266419
rect 167771 265237 167893 266419
rect 166528 265134 167893 265237
rect 173486 266420 174851 266530
rect 173486 265238 173605 266420
rect 174729 265238 174851 266420
rect 173486 265135 174851 265238
rect 180291 266413 181656 266523
rect 180291 265231 180410 266413
rect 181534 265231 181656 266413
rect 180291 265128 181656 265231
rect 187256 266414 188621 266524
rect 187256 265232 187375 266414
rect 188499 265232 188621 266414
rect 187256 265129 188621 265232
rect 194214 266415 195579 266525
rect 194214 265233 194333 266415
rect 195457 265233 195579 266415
rect 194214 265130 195579 265233
rect 201134 266414 202499 266524
rect 201134 265232 201253 266414
rect 202377 265232 202499 266414
rect 201134 265129 202499 265232
rect 208099 266415 209464 266525
rect 208099 265233 208218 266415
rect 209342 265233 209464 266415
rect 208099 265130 209464 265233
rect 215057 266416 216422 266526
rect 215057 265234 215176 266416
rect 216300 265234 216422 266416
rect 215057 265131 216422 265234
rect 221974 266420 223339 266530
rect 221974 265238 222093 266420
rect 223217 265238 223339 266420
rect 221974 265135 223339 265238
rect 69490 260019 70855 260129
rect 69490 258837 69609 260019
rect 70733 258837 70855 260019
rect 69490 258734 70855 258837
rect 76407 260017 77772 260127
rect 76407 258835 76526 260017
rect 77650 258835 77772 260017
rect 76407 258732 77772 258835
rect 83372 260018 84737 260128
rect 83372 258836 83491 260018
rect 84615 258836 84737 260018
rect 83372 258733 84737 258836
rect 90330 260019 91695 260129
rect 90330 258837 90449 260019
rect 91573 258837 91695 260019
rect 90330 258734 91695 258837
rect 97148 259998 98513 260108
rect 97148 258816 97267 259998
rect 98391 258816 98513 259998
rect 97148 258713 98513 258816
rect 104113 259999 105478 260109
rect 104113 258817 104232 259999
rect 105356 258817 105478 259999
rect 104113 258714 105478 258817
rect 111071 260000 112436 260110
rect 111071 258818 111190 260000
rect 112314 258818 112436 260000
rect 111071 258715 112436 258818
rect 117991 259999 119356 260109
rect 117991 258817 118110 259999
rect 119234 258817 119356 259999
rect 117991 258714 119356 258817
rect 124956 260000 126321 260110
rect 124956 258818 125075 260000
rect 126199 258818 126321 260000
rect 124956 258715 126321 258818
rect 131914 260001 133279 260111
rect 131914 258819 132033 260001
rect 133157 258819 133279 260001
rect 131914 258716 133279 258819
rect 138831 260005 140196 260115
rect 138831 258823 138950 260005
rect 140074 258823 140196 260005
rect 138831 258720 140196 258823
rect 145796 260006 147161 260116
rect 145796 258824 145915 260006
rect 147039 258824 147161 260006
rect 145796 258721 147161 258824
rect 152754 260007 154119 260117
rect 152754 258825 152873 260007
rect 153997 258825 154119 260007
rect 152754 258722 154119 258825
rect 159671 260005 161036 260115
rect 159671 258823 159790 260005
rect 160914 258823 161036 260005
rect 159671 258720 161036 258823
rect 166636 260006 168001 260116
rect 166636 258824 166755 260006
rect 167879 258824 168001 260006
rect 166636 258721 168001 258824
rect 173594 260007 174959 260117
rect 173594 258825 173713 260007
rect 174837 258825 174959 260007
rect 173594 258722 174959 258825
rect 180399 260000 181764 260110
rect 180399 258818 180518 260000
rect 181642 258818 181764 260000
rect 180399 258715 181764 258818
rect 187364 260001 188729 260111
rect 187364 258819 187483 260001
rect 188607 258819 188729 260001
rect 187364 258716 188729 258819
rect 194322 260002 195687 260112
rect 194322 258820 194441 260002
rect 195565 258820 195687 260002
rect 194322 258717 195687 258820
rect 201242 260001 202607 260111
rect 201242 258819 201361 260001
rect 202485 258819 202607 260001
rect 201242 258716 202607 258819
rect 208207 260002 209572 260112
rect 208207 258820 208326 260002
rect 209450 258820 209572 260002
rect 208207 258717 209572 258820
rect 215165 260003 216530 260113
rect 215165 258821 215284 260003
rect 216408 258821 216530 260003
rect 215165 258718 216530 258821
rect 222082 260007 223447 260117
rect 222082 258825 222201 260007
rect 223325 258825 223447 260007
rect 222082 258722 223447 258825
rect 83569 249307 84934 249417
rect 83569 248125 83688 249307
rect 84812 248125 84934 249307
rect 83569 248022 84934 248125
rect 90527 249308 91892 249418
rect 90527 248126 90646 249308
rect 91770 248126 91892 249308
rect 90527 248023 91892 248126
rect 97345 249287 98710 249397
rect 97345 248105 97464 249287
rect 98588 248105 98710 249287
rect 97345 248002 98710 248105
rect 104310 249288 105675 249398
rect 104310 248106 104429 249288
rect 105553 248106 105675 249288
rect 104310 248003 105675 248106
rect 111268 249289 112633 249399
rect 111268 248107 111387 249289
rect 112511 248107 112633 249289
rect 111268 248004 112633 248107
rect 118188 249288 119553 249398
rect 118188 248106 118307 249288
rect 119431 248106 119553 249288
rect 118188 248003 119553 248106
rect 125153 249289 126518 249399
rect 125153 248107 125272 249289
rect 126396 248107 126518 249289
rect 125153 248004 126518 248107
rect 132111 249290 133476 249400
rect 132111 248108 132230 249290
rect 133354 248108 133476 249290
rect 132111 248005 133476 248108
rect 139028 249294 140393 249404
rect 139028 248112 139147 249294
rect 140271 248112 140393 249294
rect 139028 248009 140393 248112
rect 145993 249295 147358 249405
rect 145993 248113 146112 249295
rect 147236 248113 147358 249295
rect 145993 248010 147358 248113
rect 152951 249296 154316 249406
rect 152951 248114 153070 249296
rect 154194 248114 154316 249296
rect 152951 248011 154316 248114
rect 159868 249294 161233 249404
rect 159868 248112 159987 249294
rect 161111 248112 161233 249294
rect 159868 248009 161233 248112
rect 166833 249295 168198 249405
rect 166833 248113 166952 249295
rect 168076 248113 168198 249295
rect 166833 248010 168198 248113
rect 173791 249296 175156 249406
rect 173791 248114 173910 249296
rect 175034 248114 175156 249296
rect 173791 248011 175156 248114
rect 180596 249289 181961 249399
rect 180596 248107 180715 249289
rect 181839 248107 181961 249289
rect 180596 248004 181961 248107
rect 187561 249290 188926 249400
rect 187561 248108 187680 249290
rect 188804 248108 188926 249290
rect 187561 248005 188926 248108
rect 194519 249291 195884 249401
rect 194519 248109 194638 249291
rect 195762 248109 195884 249291
rect 194519 248006 195884 248109
rect 201439 249290 202804 249400
rect 201439 248108 201558 249290
rect 202682 248108 202804 249290
rect 201439 248005 202804 248108
rect 208404 249291 209769 249401
rect 208404 248109 208523 249291
rect 209647 248109 209769 249291
rect 208404 248006 209769 248109
rect 215362 249292 216727 249402
rect 215362 248110 215481 249292
rect 216605 248110 216727 249292
rect 215362 248007 216727 248110
rect 222279 249296 223644 249406
rect 222279 248114 222398 249296
rect 223522 248114 223644 249296
rect 222279 248011 223644 248114
rect 83295 242177 84660 242287
rect 83295 240995 83414 242177
rect 84538 240995 84660 242177
rect 83295 240892 84660 240995
rect 90253 242178 91618 242288
rect 90253 240996 90372 242178
rect 91496 240996 91618 242178
rect 90253 240893 91618 240996
rect 97071 242157 98436 242267
rect 97071 240975 97190 242157
rect 98314 240975 98436 242157
rect 97071 240872 98436 240975
rect 104036 242158 105401 242268
rect 104036 240976 104155 242158
rect 105279 240976 105401 242158
rect 104036 240873 105401 240976
rect 110994 242159 112359 242269
rect 110994 240977 111113 242159
rect 112237 240977 112359 242159
rect 110994 240874 112359 240977
rect 117914 242158 119279 242268
rect 117914 240976 118033 242158
rect 119157 240976 119279 242158
rect 117914 240873 119279 240976
rect 124879 242159 126244 242269
rect 124879 240977 124998 242159
rect 126122 240977 126244 242159
rect 124879 240874 126244 240977
rect 131837 242160 133202 242270
rect 131837 240978 131956 242160
rect 133080 240978 133202 242160
rect 131837 240875 133202 240978
rect 138754 242164 140119 242274
rect 138754 240982 138873 242164
rect 139997 240982 140119 242164
rect 138754 240879 140119 240982
rect 145719 242165 147084 242275
rect 145719 240983 145838 242165
rect 146962 240983 147084 242165
rect 145719 240880 147084 240983
rect 152677 242166 154042 242276
rect 152677 240984 152796 242166
rect 153920 240984 154042 242166
rect 152677 240881 154042 240984
rect 159594 242164 160959 242274
rect 159594 240982 159713 242164
rect 160837 240982 160959 242164
rect 159594 240879 160959 240982
rect 166559 242165 167924 242275
rect 166559 240983 166678 242165
rect 167802 240983 167924 242165
rect 166559 240880 167924 240983
rect 173517 242166 174882 242276
rect 173517 240984 173636 242166
rect 174760 240984 174882 242166
rect 173517 240881 174882 240984
rect 180322 242159 181687 242269
rect 180322 240977 180441 242159
rect 181565 240977 181687 242159
rect 180322 240874 181687 240977
rect 187287 242160 188652 242270
rect 187287 240978 187406 242160
rect 188530 240978 188652 242160
rect 187287 240875 188652 240978
rect 194245 242161 195610 242271
rect 194245 240979 194364 242161
rect 195488 240979 195610 242161
rect 194245 240876 195610 240979
rect 201165 242160 202530 242270
rect 201165 240978 201284 242160
rect 202408 240978 202530 242160
rect 201165 240875 202530 240978
rect 208130 242161 209495 242271
rect 208130 240979 208249 242161
rect 209373 240979 209495 242161
rect 208130 240876 209495 240979
rect 215088 242162 216453 242272
rect 215088 240980 215207 242162
rect 216331 240980 216453 242162
rect 215088 240877 216453 240980
rect 222005 242166 223370 242276
rect 222005 240984 222124 242166
rect 223248 240984 223370 242166
rect 222005 240881 223370 240984
rect 83403 235764 84768 235874
rect 83403 234582 83522 235764
rect 84646 234582 84768 235764
rect 83403 234479 84768 234582
rect 90361 235765 91726 235875
rect 90361 234583 90480 235765
rect 91604 234583 91726 235765
rect 90361 234480 91726 234583
rect 97179 235744 98544 235854
rect 97179 234562 97298 235744
rect 98422 234562 98544 235744
rect 97179 234459 98544 234562
rect 104144 235745 105509 235855
rect 104144 234563 104263 235745
rect 105387 234563 105509 235745
rect 104144 234460 105509 234563
rect 111102 235746 112467 235856
rect 111102 234564 111221 235746
rect 112345 234564 112467 235746
rect 111102 234461 112467 234564
rect 118022 235745 119387 235855
rect 118022 234563 118141 235745
rect 119265 234563 119387 235745
rect 118022 234460 119387 234563
rect 124987 235746 126352 235856
rect 124987 234564 125106 235746
rect 126230 234564 126352 235746
rect 124987 234461 126352 234564
rect 131945 235747 133310 235857
rect 131945 234565 132064 235747
rect 133188 234565 133310 235747
rect 131945 234462 133310 234565
rect 138862 235751 140227 235861
rect 138862 234569 138981 235751
rect 140105 234569 140227 235751
rect 138862 234466 140227 234569
rect 145827 235752 147192 235862
rect 145827 234570 145946 235752
rect 147070 234570 147192 235752
rect 145827 234467 147192 234570
rect 152785 235753 154150 235863
rect 152785 234571 152904 235753
rect 154028 234571 154150 235753
rect 152785 234468 154150 234571
rect 159702 235751 161067 235861
rect 159702 234569 159821 235751
rect 160945 234569 161067 235751
rect 159702 234466 161067 234569
rect 166667 235752 168032 235862
rect 166667 234570 166786 235752
rect 167910 234570 168032 235752
rect 166667 234467 168032 234570
rect 173625 235753 174990 235863
rect 173625 234571 173744 235753
rect 174868 234571 174990 235753
rect 173625 234468 174990 234571
rect 180430 235746 181795 235856
rect 180430 234564 180549 235746
rect 181673 234564 181795 235746
rect 180430 234461 181795 234564
rect 187395 235747 188760 235857
rect 187395 234565 187514 235747
rect 188638 234565 188760 235747
rect 187395 234462 188760 234565
rect 194353 235748 195718 235858
rect 194353 234566 194472 235748
rect 195596 234566 195718 235748
rect 194353 234463 195718 234566
rect 201273 235747 202638 235857
rect 201273 234565 201392 235747
rect 202516 234565 202638 235747
rect 201273 234462 202638 234565
rect 208238 235748 209603 235858
rect 208238 234566 208357 235748
rect 209481 234566 209603 235748
rect 208238 234463 209603 234566
rect 215196 235749 216561 235859
rect 215196 234567 215315 235749
rect 216439 234567 216561 235749
rect 215196 234464 216561 234567
rect 222113 235753 223478 235863
rect 222113 234571 222232 235753
rect 223356 234571 223478 235753
rect 222113 234468 223478 234571
rect 48971 229036 50336 229146
rect 48971 227854 49090 229036
rect 50214 227854 50336 229036
rect 48971 227751 50336 227854
rect 55888 229040 57253 229150
rect 55888 227858 56007 229040
rect 57131 227858 57253 229040
rect 55888 227755 57253 227858
rect 62853 229041 64218 229151
rect 62853 227859 62972 229041
rect 64096 227859 64218 229041
rect 62853 227756 64218 227859
rect 69811 229042 71176 229152
rect 69811 227860 69930 229042
rect 71054 227860 71176 229042
rect 69811 227757 71176 227860
rect 76728 229040 78093 229150
rect 76728 227858 76847 229040
rect 77971 227858 78093 229040
rect 76728 227755 78093 227858
rect 83693 229041 85058 229151
rect 83693 227859 83812 229041
rect 84936 227859 85058 229041
rect 83693 227756 85058 227859
rect 90651 229042 92016 229152
rect 90651 227860 90770 229042
rect 91894 227860 92016 229042
rect 90651 227757 92016 227860
rect 97469 229021 98834 229131
rect 97469 227839 97588 229021
rect 98712 227839 98834 229021
rect 97469 227736 98834 227839
rect 104434 229022 105799 229132
rect 104434 227840 104553 229022
rect 105677 227840 105799 229022
rect 104434 227737 105799 227840
rect 111392 229023 112757 229133
rect 111392 227841 111511 229023
rect 112635 227841 112757 229023
rect 111392 227738 112757 227841
rect 118312 229022 119677 229132
rect 118312 227840 118431 229022
rect 119555 227840 119677 229022
rect 118312 227737 119677 227840
rect 125277 229023 126642 229133
rect 125277 227841 125396 229023
rect 126520 227841 126642 229023
rect 125277 227738 126642 227841
rect 132235 229024 133600 229134
rect 132235 227842 132354 229024
rect 133478 227842 133600 229024
rect 132235 227739 133600 227842
rect 139152 229028 140517 229138
rect 139152 227846 139271 229028
rect 140395 227846 140517 229028
rect 139152 227743 140517 227846
rect 146117 229029 147482 229139
rect 146117 227847 146236 229029
rect 147360 227847 147482 229029
rect 146117 227744 147482 227847
rect 153075 229030 154440 229140
rect 153075 227848 153194 229030
rect 154318 227848 154440 229030
rect 153075 227745 154440 227848
rect 159992 229028 161357 229138
rect 159992 227846 160111 229028
rect 161235 227846 161357 229028
rect 159992 227743 161357 227846
rect 166957 229029 168322 229139
rect 166957 227847 167076 229029
rect 168200 227847 168322 229029
rect 166957 227744 168322 227847
rect 173915 229030 175280 229140
rect 173915 227848 174034 229030
rect 175158 227848 175280 229030
rect 173915 227745 175280 227848
rect 180720 229023 182085 229133
rect 180720 227841 180839 229023
rect 181963 227841 182085 229023
rect 180720 227738 182085 227841
rect 187685 229024 189050 229134
rect 187685 227842 187804 229024
rect 188928 227842 189050 229024
rect 187685 227739 189050 227842
rect 194643 229025 196008 229135
rect 194643 227843 194762 229025
rect 195886 227843 196008 229025
rect 194643 227740 196008 227843
rect 201563 229024 202928 229134
rect 201563 227842 201682 229024
rect 202806 227842 202928 229024
rect 201563 227739 202928 227842
rect 208528 229025 209893 229135
rect 208528 227843 208647 229025
rect 209771 227843 209893 229025
rect 208528 227740 209893 227843
rect 215486 229026 216851 229136
rect 215486 227844 215605 229026
rect 216729 227844 216851 229026
rect 215486 227741 216851 227844
rect 222403 229030 223768 229140
rect 222403 227848 222522 229030
rect 223646 227848 223768 229030
rect 222403 227745 223768 227848
rect 229368 229031 230733 229141
rect 229368 227849 229487 229031
rect 230611 227849 230733 229031
rect 229368 227746 230733 227849
rect 236326 229032 237691 229142
rect 236326 227850 236445 229032
rect 237569 227850 237691 229032
rect 236326 227747 237691 227850
rect 243243 229030 244608 229140
rect 243243 227848 243362 229030
rect 244486 227848 244608 229030
rect 243243 227745 244608 227848
rect 250208 229031 251573 229141
rect 250208 227849 250327 229031
rect 251451 227849 251573 229031
rect 250208 227746 251573 227849
rect 257166 229032 258531 229142
rect 257166 227850 257285 229032
rect 258409 227850 258531 229032
rect 257166 227747 258531 227850
rect 264306 229032 265671 229142
rect 264306 227850 264425 229032
rect 265549 227850 265671 229032
rect 264306 227747 265671 227850
rect 271264 229033 272629 229143
rect 271264 227851 271383 229033
rect 272507 227851 272629 229033
rect 271264 227748 272629 227851
rect 278400 229023 279765 229133
rect 278400 227841 278519 229023
rect 279643 227841 279765 229023
rect 278400 227738 279765 227841
rect 48951 223174 50316 223284
rect 48951 221992 49070 223174
rect 50194 221992 50316 223174
rect 48951 221889 50316 221992
rect 55868 223178 57233 223288
rect 55868 221996 55987 223178
rect 57111 221996 57233 223178
rect 55868 221893 57233 221996
rect 62833 223179 64198 223289
rect 62833 221997 62952 223179
rect 64076 221997 64198 223179
rect 62833 221894 64198 221997
rect 69791 223180 71156 223290
rect 69791 221998 69910 223180
rect 71034 221998 71156 223180
rect 69791 221895 71156 221998
rect 76708 223178 78073 223288
rect 76708 221996 76827 223178
rect 77951 221996 78073 223178
rect 76708 221893 78073 221996
rect 83673 223179 85038 223289
rect 83673 221997 83792 223179
rect 84916 221997 85038 223179
rect 83673 221894 85038 221997
rect 90631 223180 91996 223290
rect 90631 221998 90750 223180
rect 91874 221998 91996 223180
rect 90631 221895 91996 221998
rect 97449 223159 98814 223269
rect 97449 221977 97568 223159
rect 98692 221977 98814 223159
rect 97449 221874 98814 221977
rect 104414 223160 105779 223270
rect 104414 221978 104533 223160
rect 105657 221978 105779 223160
rect 104414 221875 105779 221978
rect 111372 223161 112737 223271
rect 111372 221979 111491 223161
rect 112615 221979 112737 223161
rect 111372 221876 112737 221979
rect 118292 223160 119657 223270
rect 118292 221978 118411 223160
rect 119535 221978 119657 223160
rect 118292 221875 119657 221978
rect 125257 223161 126622 223271
rect 125257 221979 125376 223161
rect 126500 221979 126622 223161
rect 125257 221876 126622 221979
rect 132215 223162 133580 223272
rect 132215 221980 132334 223162
rect 133458 221980 133580 223162
rect 132215 221877 133580 221980
rect 139132 223166 140497 223276
rect 139132 221984 139251 223166
rect 140375 221984 140497 223166
rect 139132 221881 140497 221984
rect 146097 223167 147462 223277
rect 146097 221985 146216 223167
rect 147340 221985 147462 223167
rect 146097 221882 147462 221985
rect 153055 223168 154420 223278
rect 153055 221986 153174 223168
rect 154298 221986 154420 223168
rect 153055 221883 154420 221986
rect 159972 223166 161337 223276
rect 159972 221984 160091 223166
rect 161215 221984 161337 223166
rect 159972 221881 161337 221984
rect 166937 223167 168302 223277
rect 166937 221985 167056 223167
rect 168180 221985 168302 223167
rect 166937 221882 168302 221985
rect 173895 223168 175260 223278
rect 173895 221986 174014 223168
rect 175138 221986 175260 223168
rect 173895 221883 175260 221986
rect 180700 223161 182065 223271
rect 180700 221979 180819 223161
rect 181943 221979 182065 223161
rect 180700 221876 182065 221979
rect 187665 223162 189030 223272
rect 187665 221980 187784 223162
rect 188908 221980 189030 223162
rect 187665 221877 189030 221980
rect 194623 223163 195988 223273
rect 194623 221981 194742 223163
rect 195866 221981 195988 223163
rect 194623 221878 195988 221981
rect 201543 223162 202908 223272
rect 201543 221980 201662 223162
rect 202786 221980 202908 223162
rect 201543 221877 202908 221980
rect 208508 223163 209873 223273
rect 208508 221981 208627 223163
rect 209751 221981 209873 223163
rect 208508 221878 209873 221981
rect 215466 223164 216831 223274
rect 215466 221982 215585 223164
rect 216709 221982 216831 223164
rect 215466 221879 216831 221982
rect 222383 223168 223748 223278
rect 222383 221986 222502 223168
rect 223626 221986 223748 223168
rect 222383 221883 223748 221986
rect 229348 223169 230713 223279
rect 229348 221987 229467 223169
rect 230591 221987 230713 223169
rect 229348 221884 230713 221987
rect 236306 223170 237671 223280
rect 236306 221988 236425 223170
rect 237549 221988 237671 223170
rect 236306 221885 237671 221988
rect 243223 223168 244588 223278
rect 243223 221986 243342 223168
rect 244466 221986 244588 223168
rect 243223 221883 244588 221986
rect 250188 223169 251553 223279
rect 250188 221987 250307 223169
rect 251431 221987 251553 223169
rect 250188 221884 251553 221987
rect 257146 223170 258511 223280
rect 257146 221988 257265 223170
rect 258389 221988 258511 223170
rect 257146 221885 258511 221988
rect 264286 223170 265651 223280
rect 264286 221988 264405 223170
rect 265529 221988 265651 223170
rect 264286 221885 265651 221988
rect 271244 223171 272609 223281
rect 271244 221989 271363 223171
rect 272487 221989 272609 223171
rect 271244 221886 272609 221989
rect 278380 223161 279745 223271
rect 278380 221979 278499 223161
rect 279623 221979 279745 223161
rect 278380 221876 279745 221979
rect 21190 211109 22555 211219
rect 21190 209927 21309 211109
rect 22433 209927 22555 211109
rect 21190 209824 22555 209927
rect 28148 211110 29513 211220
rect 28148 209928 28267 211110
rect 29391 209928 29513 211110
rect 28148 209825 29513 209928
rect 35068 211109 36433 211219
rect 35068 209927 35187 211109
rect 36311 209927 36433 211109
rect 35068 209824 36433 209927
rect 42033 211110 43398 211220
rect 42033 209928 42152 211110
rect 43276 209928 43398 211110
rect 42033 209825 43398 209928
rect 48991 211111 50356 211221
rect 48991 209929 49110 211111
rect 50234 209929 50356 211111
rect 48991 209826 50356 209929
rect 55908 211115 57273 211225
rect 55908 209933 56027 211115
rect 57151 209933 57273 211115
rect 55908 209830 57273 209933
rect 62873 211116 64238 211226
rect 62873 209934 62992 211116
rect 64116 209934 64238 211116
rect 62873 209831 64238 209934
rect 69831 211117 71196 211227
rect 69831 209935 69950 211117
rect 71074 209935 71196 211117
rect 69831 209832 71196 209935
rect 76748 211115 78113 211225
rect 76748 209933 76867 211115
rect 77991 209933 78113 211115
rect 76748 209830 78113 209933
rect 83713 211116 85078 211226
rect 83713 209934 83832 211116
rect 84956 209934 85078 211116
rect 83713 209831 85078 209934
rect 90671 211117 92036 211227
rect 90671 209935 90790 211117
rect 91914 209935 92036 211117
rect 90671 209832 92036 209935
rect 97489 211096 98854 211206
rect 97489 209914 97608 211096
rect 98732 209914 98854 211096
rect 97489 209811 98854 209914
rect 104454 211097 105819 211207
rect 104454 209915 104573 211097
rect 105697 209915 105819 211097
rect 104454 209812 105819 209915
rect 111412 211098 112777 211208
rect 111412 209916 111531 211098
rect 112655 209916 112777 211098
rect 111412 209813 112777 209916
rect 118332 211097 119697 211207
rect 118332 209915 118451 211097
rect 119575 209915 119697 211097
rect 118332 209812 119697 209915
rect 125297 211098 126662 211208
rect 125297 209916 125416 211098
rect 126540 209916 126662 211098
rect 125297 209813 126662 209916
rect 132255 211099 133620 211209
rect 132255 209917 132374 211099
rect 133498 209917 133620 211099
rect 132255 209814 133620 209917
rect 139172 211103 140537 211213
rect 139172 209921 139291 211103
rect 140415 209921 140537 211103
rect 139172 209818 140537 209921
rect 146137 211104 147502 211214
rect 146137 209922 146256 211104
rect 147380 209922 147502 211104
rect 146137 209819 147502 209922
rect 153095 211105 154460 211215
rect 153095 209923 153214 211105
rect 154338 209923 154460 211105
rect 153095 209820 154460 209923
rect 160012 211103 161377 211213
rect 160012 209921 160131 211103
rect 161255 209921 161377 211103
rect 160012 209818 161377 209921
rect 166977 211104 168342 211214
rect 166977 209922 167096 211104
rect 168220 209922 168342 211104
rect 166977 209819 168342 209922
rect 173935 211105 175300 211215
rect 173935 209923 174054 211105
rect 175178 209923 175300 211105
rect 173935 209820 175300 209923
rect 180740 211098 182105 211208
rect 180740 209916 180859 211098
rect 181983 209916 182105 211098
rect 180740 209813 182105 209916
rect 187705 211099 189070 211209
rect 187705 209917 187824 211099
rect 188948 209917 189070 211099
rect 187705 209814 189070 209917
rect 194663 211100 196028 211210
rect 194663 209918 194782 211100
rect 195906 209918 196028 211100
rect 194663 209815 196028 209918
rect 201583 211099 202948 211209
rect 201583 209917 201702 211099
rect 202826 209917 202948 211099
rect 201583 209814 202948 209917
rect 208548 211100 209913 211210
rect 208548 209918 208667 211100
rect 209791 209918 209913 211100
rect 208548 209815 209913 209918
rect 215506 211101 216871 211211
rect 215506 209919 215625 211101
rect 216749 209919 216871 211101
rect 215506 209816 216871 209919
rect 222423 211105 223788 211215
rect 222423 209923 222542 211105
rect 223666 209923 223788 211105
rect 222423 209820 223788 209923
rect 229388 211106 230753 211216
rect 229388 209924 229507 211106
rect 230631 209924 230753 211106
rect 229388 209821 230753 209924
rect 236346 211107 237711 211217
rect 236346 209925 236465 211107
rect 237589 209925 237711 211107
rect 236346 209822 237711 209925
rect 243263 211105 244628 211215
rect 243263 209923 243382 211105
rect 244506 209923 244628 211105
rect 243263 209820 244628 209923
rect 250228 211106 251593 211216
rect 250228 209924 250347 211106
rect 251471 209924 251593 211106
rect 250228 209821 251593 209924
rect 257186 211107 258551 211217
rect 257186 209925 257305 211107
rect 258429 209925 258551 211107
rect 257186 209822 258551 209925
rect 264326 211107 265691 211217
rect 264326 209925 264445 211107
rect 265569 209925 265691 211107
rect 264326 209822 265691 209925
rect 271284 211108 272649 211218
rect 271284 209926 271403 211108
rect 272527 209926 272649 211108
rect 271284 209823 272649 209926
rect 278420 211098 279785 211208
rect 278420 209916 278539 211098
rect 279663 209916 279785 211098
rect 278420 209813 279785 209916
rect 20916 203979 22281 204089
rect 20916 202797 21035 203979
rect 22159 202797 22281 203979
rect 20916 202694 22281 202797
rect 27874 203980 29239 204090
rect 27874 202798 27993 203980
rect 29117 202798 29239 203980
rect 27874 202695 29239 202798
rect 34794 203979 36159 204089
rect 34794 202797 34913 203979
rect 36037 202797 36159 203979
rect 34794 202694 36159 202797
rect 41759 203980 43124 204090
rect 41759 202798 41878 203980
rect 43002 202798 43124 203980
rect 41759 202695 43124 202798
rect 48717 203981 50082 204091
rect 48717 202799 48836 203981
rect 49960 202799 50082 203981
rect 48717 202696 50082 202799
rect 55634 203985 56999 204095
rect 55634 202803 55753 203985
rect 56877 202803 56999 203985
rect 55634 202700 56999 202803
rect 62599 203986 63964 204096
rect 62599 202804 62718 203986
rect 63842 202804 63964 203986
rect 62599 202701 63964 202804
rect 69557 203987 70922 204097
rect 69557 202805 69676 203987
rect 70800 202805 70922 203987
rect 69557 202702 70922 202805
rect 76474 203985 77839 204095
rect 76474 202803 76593 203985
rect 77717 202803 77839 203985
rect 76474 202700 77839 202803
rect 83439 203986 84804 204096
rect 83439 202804 83558 203986
rect 84682 202804 84804 203986
rect 83439 202701 84804 202804
rect 90397 203987 91762 204097
rect 90397 202805 90516 203987
rect 91640 202805 91762 203987
rect 90397 202702 91762 202805
rect 97215 203966 98580 204076
rect 97215 202784 97334 203966
rect 98458 202784 98580 203966
rect 97215 202681 98580 202784
rect 104180 203967 105545 204077
rect 104180 202785 104299 203967
rect 105423 202785 105545 203967
rect 104180 202682 105545 202785
rect 111138 203968 112503 204078
rect 111138 202786 111257 203968
rect 112381 202786 112503 203968
rect 111138 202683 112503 202786
rect 118058 203967 119423 204077
rect 118058 202785 118177 203967
rect 119301 202785 119423 203967
rect 118058 202682 119423 202785
rect 125023 203968 126388 204078
rect 125023 202786 125142 203968
rect 126266 202786 126388 203968
rect 125023 202683 126388 202786
rect 131981 203969 133346 204079
rect 131981 202787 132100 203969
rect 133224 202787 133346 203969
rect 131981 202684 133346 202787
rect 138898 203973 140263 204083
rect 138898 202791 139017 203973
rect 140141 202791 140263 203973
rect 138898 202688 140263 202791
rect 145863 203974 147228 204084
rect 145863 202792 145982 203974
rect 147106 202792 147228 203974
rect 145863 202689 147228 202792
rect 152821 203975 154186 204085
rect 152821 202793 152940 203975
rect 154064 202793 154186 203975
rect 152821 202690 154186 202793
rect 159738 203973 161103 204083
rect 159738 202791 159857 203973
rect 160981 202791 161103 203973
rect 159738 202688 161103 202791
rect 166703 203974 168068 204084
rect 166703 202792 166822 203974
rect 167946 202792 168068 203974
rect 166703 202689 168068 202792
rect 173661 203975 175026 204085
rect 173661 202793 173780 203975
rect 174904 202793 175026 203975
rect 173661 202690 175026 202793
rect 180466 203968 181831 204078
rect 180466 202786 180585 203968
rect 181709 202786 181831 203968
rect 180466 202683 181831 202786
rect 187431 203969 188796 204079
rect 187431 202787 187550 203969
rect 188674 202787 188796 203969
rect 187431 202684 188796 202787
rect 194389 203970 195754 204080
rect 194389 202788 194508 203970
rect 195632 202788 195754 203970
rect 194389 202685 195754 202788
rect 201309 203969 202674 204079
rect 201309 202787 201428 203969
rect 202552 202787 202674 203969
rect 201309 202684 202674 202787
rect 208274 203970 209639 204080
rect 208274 202788 208393 203970
rect 209517 202788 209639 203970
rect 208274 202685 209639 202788
rect 215232 203971 216597 204081
rect 215232 202789 215351 203971
rect 216475 202789 216597 203971
rect 215232 202686 216597 202789
rect 222149 203975 223514 204085
rect 222149 202793 222268 203975
rect 223392 202793 223514 203975
rect 222149 202690 223514 202793
rect 229114 203976 230479 204086
rect 229114 202794 229233 203976
rect 230357 202794 230479 203976
rect 229114 202691 230479 202794
rect 236072 203977 237437 204087
rect 236072 202795 236191 203977
rect 237315 202795 237437 203977
rect 236072 202692 237437 202795
rect 242989 203975 244354 204085
rect 242989 202793 243108 203975
rect 244232 202793 244354 203975
rect 242989 202690 244354 202793
rect 249954 203976 251319 204086
rect 249954 202794 250073 203976
rect 251197 202794 251319 203976
rect 249954 202691 251319 202794
rect 256912 203977 258277 204087
rect 256912 202795 257031 203977
rect 258155 202795 258277 203977
rect 256912 202692 258277 202795
rect 264052 203977 265417 204087
rect 264052 202795 264171 203977
rect 265295 202795 265417 203977
rect 264052 202692 265417 202795
rect 271010 203978 272375 204088
rect 271010 202796 271129 203978
rect 272253 202796 272375 203978
rect 271010 202693 272375 202796
rect 278146 203968 279511 204078
rect 278146 202786 278265 203968
rect 279389 202786 279511 203968
rect 278146 202683 279511 202786
rect 21024 197566 22389 197676
rect 21024 196384 21143 197566
rect 22267 196384 22389 197566
rect 21024 196281 22389 196384
rect 27982 197567 29347 197677
rect 27982 196385 28101 197567
rect 29225 196385 29347 197567
rect 27982 196282 29347 196385
rect 34902 197566 36267 197676
rect 34902 196384 35021 197566
rect 36145 196384 36267 197566
rect 34902 196281 36267 196384
rect 41867 197567 43232 197677
rect 41867 196385 41986 197567
rect 43110 196385 43232 197567
rect 41867 196282 43232 196385
rect 48825 197568 50190 197678
rect 48825 196386 48944 197568
rect 50068 196386 50190 197568
rect 48825 196283 50190 196386
rect 55742 197572 57107 197682
rect 55742 196390 55861 197572
rect 56985 196390 57107 197572
rect 55742 196287 57107 196390
rect 62707 197573 64072 197683
rect 62707 196391 62826 197573
rect 63950 196391 64072 197573
rect 62707 196288 64072 196391
rect 69665 197574 71030 197684
rect 69665 196392 69784 197574
rect 70908 196392 71030 197574
rect 69665 196289 71030 196392
rect 76582 197572 77947 197682
rect 76582 196390 76701 197572
rect 77825 196390 77947 197572
rect 76582 196287 77947 196390
rect 83547 197573 84912 197683
rect 83547 196391 83666 197573
rect 84790 196391 84912 197573
rect 83547 196288 84912 196391
rect 90505 197574 91870 197684
rect 90505 196392 90624 197574
rect 91748 196392 91870 197574
rect 90505 196289 91870 196392
rect 97323 197553 98688 197663
rect 97323 196371 97442 197553
rect 98566 196371 98688 197553
rect 97323 196268 98688 196371
rect 104288 197554 105653 197664
rect 104288 196372 104407 197554
rect 105531 196372 105653 197554
rect 104288 196269 105653 196372
rect 111246 197555 112611 197665
rect 111246 196373 111365 197555
rect 112489 196373 112611 197555
rect 111246 196270 112611 196373
rect 118166 197554 119531 197664
rect 118166 196372 118285 197554
rect 119409 196372 119531 197554
rect 118166 196269 119531 196372
rect 125131 197555 126496 197665
rect 125131 196373 125250 197555
rect 126374 196373 126496 197555
rect 125131 196270 126496 196373
rect 132089 197556 133454 197666
rect 132089 196374 132208 197556
rect 133332 196374 133454 197556
rect 132089 196271 133454 196374
rect 139006 197560 140371 197670
rect 139006 196378 139125 197560
rect 140249 196378 140371 197560
rect 139006 196275 140371 196378
rect 145971 197561 147336 197671
rect 145971 196379 146090 197561
rect 147214 196379 147336 197561
rect 145971 196276 147336 196379
rect 152929 197562 154294 197672
rect 152929 196380 153048 197562
rect 154172 196380 154294 197562
rect 152929 196277 154294 196380
rect 159846 197560 161211 197670
rect 159846 196378 159965 197560
rect 161089 196378 161211 197560
rect 159846 196275 161211 196378
rect 166811 197561 168176 197671
rect 166811 196379 166930 197561
rect 168054 196379 168176 197561
rect 166811 196276 168176 196379
rect 173769 197562 175134 197672
rect 173769 196380 173888 197562
rect 175012 196380 175134 197562
rect 173769 196277 175134 196380
rect 180574 197555 181939 197665
rect 180574 196373 180693 197555
rect 181817 196373 181939 197555
rect 180574 196270 181939 196373
rect 187539 197556 188904 197666
rect 187539 196374 187658 197556
rect 188782 196374 188904 197556
rect 187539 196271 188904 196374
rect 194497 197557 195862 197667
rect 194497 196375 194616 197557
rect 195740 196375 195862 197557
rect 194497 196272 195862 196375
rect 201417 197556 202782 197666
rect 201417 196374 201536 197556
rect 202660 196374 202782 197556
rect 201417 196271 202782 196374
rect 208382 197557 209747 197667
rect 208382 196375 208501 197557
rect 209625 196375 209747 197557
rect 208382 196272 209747 196375
rect 215340 197558 216705 197668
rect 215340 196376 215459 197558
rect 216583 196376 216705 197558
rect 215340 196273 216705 196376
rect 222257 197562 223622 197672
rect 222257 196380 222376 197562
rect 223500 196380 223622 197562
rect 222257 196277 223622 196380
rect 229222 197563 230587 197673
rect 229222 196381 229341 197563
rect 230465 196381 230587 197563
rect 229222 196278 230587 196381
rect 236180 197564 237545 197674
rect 236180 196382 236299 197564
rect 237423 196382 237545 197564
rect 236180 196279 237545 196382
rect 243097 197562 244462 197672
rect 243097 196380 243216 197562
rect 244340 196380 244462 197562
rect 243097 196277 244462 196380
rect 250062 197563 251427 197673
rect 250062 196381 250181 197563
rect 251305 196381 251427 197563
rect 250062 196278 251427 196381
rect 257020 197564 258385 197674
rect 257020 196382 257139 197564
rect 258263 196382 258385 197564
rect 257020 196279 258385 196382
rect 264160 197564 265525 197674
rect 264160 196382 264279 197564
rect 265403 196382 265525 197564
rect 264160 196279 265525 196382
rect 271118 197565 272483 197675
rect 271118 196383 271237 197565
rect 272361 196383 272483 197565
rect 271118 196280 272483 196383
rect 278254 197555 279619 197665
rect 278254 196373 278373 197555
rect 279497 196373 279619 197555
rect 278254 196270 279619 196373
rect 76735 193222 78100 193332
rect 76735 192040 76854 193222
rect 77978 192040 78100 193222
rect 76735 191937 78100 192040
rect 83700 193223 85065 193333
rect 83700 192041 83819 193223
rect 84943 192041 85065 193223
rect 83700 191938 85065 192041
rect 90658 193224 92023 193334
rect 90658 192042 90777 193224
rect 91901 192042 92023 193224
rect 90658 191939 92023 192042
rect 97476 193203 98841 193313
rect 97476 192021 97595 193203
rect 98719 192021 98841 193203
rect 97476 191918 98841 192021
rect 104441 193204 105806 193314
rect 104441 192022 104560 193204
rect 105684 192022 105806 193204
rect 104441 191919 105806 192022
rect 111399 193205 112764 193315
rect 111399 192023 111518 193205
rect 112642 192023 112764 193205
rect 111399 191920 112764 192023
rect 118319 193204 119684 193314
rect 118319 192022 118438 193204
rect 119562 192022 119684 193204
rect 118319 191919 119684 192022
rect 125284 193205 126649 193315
rect 125284 192023 125403 193205
rect 126527 192023 126649 193205
rect 125284 191920 126649 192023
rect 132242 193206 133607 193316
rect 132242 192024 132361 193206
rect 133485 192024 133607 193206
rect 132242 191921 133607 192024
rect 139159 193210 140524 193320
rect 139159 192028 139278 193210
rect 140402 192028 140524 193210
rect 139159 191925 140524 192028
rect 146124 193211 147489 193321
rect 146124 192029 146243 193211
rect 147367 192029 147489 193211
rect 146124 191926 147489 192029
rect 153082 193212 154447 193322
rect 153082 192030 153201 193212
rect 154325 192030 154447 193212
rect 153082 191927 154447 192030
rect 159999 193210 161364 193320
rect 159999 192028 160118 193210
rect 161242 192028 161364 193210
rect 159999 191925 161364 192028
rect 166964 193211 168329 193321
rect 166964 192029 167083 193211
rect 168207 192029 168329 193211
rect 166964 191926 168329 192029
rect 173922 193212 175287 193322
rect 173922 192030 174041 193212
rect 175165 192030 175287 193212
rect 173922 191927 175287 192030
rect 180727 193205 182092 193315
rect 180727 192023 180846 193205
rect 181970 192023 182092 193205
rect 180727 191920 182092 192023
rect 187692 193206 189057 193316
rect 187692 192024 187811 193206
rect 188935 192024 189057 193206
rect 187692 191921 189057 192024
rect 194650 193207 196015 193317
rect 194650 192025 194769 193207
rect 195893 192025 196015 193207
rect 194650 191922 196015 192025
rect 201570 193206 202935 193316
rect 201570 192024 201689 193206
rect 202813 192024 202935 193206
rect 201570 191921 202935 192024
rect 208535 193207 209900 193317
rect 208535 192025 208654 193207
rect 209778 192025 209900 193207
rect 208535 191922 209900 192025
rect 215493 193208 216858 193318
rect 215493 192026 215612 193208
rect 216736 192026 216858 193208
rect 215493 191923 216858 192026
rect 222410 193212 223775 193322
rect 222410 192030 222529 193212
rect 223653 192030 223775 193212
rect 222410 191927 223775 192030
rect 229375 193213 230740 193323
rect 229375 192031 229494 193213
rect 230618 192031 230740 193213
rect 229375 191928 230740 192031
rect 236333 193214 237698 193324
rect 236333 192032 236452 193214
rect 237576 192032 237698 193214
rect 236333 191929 237698 192032
rect 243250 193212 244615 193322
rect 243250 192030 243369 193212
rect 244493 192030 244615 193212
rect 243250 191927 244615 192030
rect 250215 193213 251580 193323
rect 250215 192031 250334 193213
rect 251458 192031 251580 193213
rect 250215 191928 251580 192031
rect 257173 193214 258538 193324
rect 257173 192032 257292 193214
rect 258416 192032 258538 193214
rect 257173 191929 258538 192032
rect 264313 193214 265678 193324
rect 264313 192032 264432 193214
rect 265556 192032 265678 193214
rect 264313 191929 265678 192032
rect 271271 193215 272636 193325
rect 271271 192033 271390 193215
rect 272514 192033 272636 193215
rect 271271 191930 272636 192033
rect 278407 193205 279772 193315
rect 278407 192023 278526 193205
rect 279650 192023 279772 193205
rect 278407 191920 279772 192023
rect 76461 186092 77826 186202
rect 76461 184910 76580 186092
rect 77704 184910 77826 186092
rect 76461 184807 77826 184910
rect 83426 186093 84791 186203
rect 83426 184911 83545 186093
rect 84669 184911 84791 186093
rect 83426 184808 84791 184911
rect 90384 186094 91749 186204
rect 90384 184912 90503 186094
rect 91627 184912 91749 186094
rect 90384 184809 91749 184912
rect 97202 186073 98567 186183
rect 97202 184891 97321 186073
rect 98445 184891 98567 186073
rect 97202 184788 98567 184891
rect 104167 186074 105532 186184
rect 104167 184892 104286 186074
rect 105410 184892 105532 186074
rect 104167 184789 105532 184892
rect 111125 186075 112490 186185
rect 111125 184893 111244 186075
rect 112368 184893 112490 186075
rect 111125 184790 112490 184893
rect 118045 186074 119410 186184
rect 118045 184892 118164 186074
rect 119288 184892 119410 186074
rect 118045 184789 119410 184892
rect 125010 186075 126375 186185
rect 125010 184893 125129 186075
rect 126253 184893 126375 186075
rect 125010 184790 126375 184893
rect 131968 186076 133333 186186
rect 131968 184894 132087 186076
rect 133211 184894 133333 186076
rect 131968 184791 133333 184894
rect 138885 186080 140250 186190
rect 138885 184898 139004 186080
rect 140128 184898 140250 186080
rect 138885 184795 140250 184898
rect 145850 186081 147215 186191
rect 145850 184899 145969 186081
rect 147093 184899 147215 186081
rect 145850 184796 147215 184899
rect 152808 186082 154173 186192
rect 152808 184900 152927 186082
rect 154051 184900 154173 186082
rect 152808 184797 154173 184900
rect 159725 186080 161090 186190
rect 159725 184898 159844 186080
rect 160968 184898 161090 186080
rect 159725 184795 161090 184898
rect 166690 186081 168055 186191
rect 166690 184899 166809 186081
rect 167933 184899 168055 186081
rect 166690 184796 168055 184899
rect 173648 186082 175013 186192
rect 173648 184900 173767 186082
rect 174891 184900 175013 186082
rect 173648 184797 175013 184900
rect 180453 186075 181818 186185
rect 180453 184893 180572 186075
rect 181696 184893 181818 186075
rect 180453 184790 181818 184893
rect 187418 186076 188783 186186
rect 187418 184894 187537 186076
rect 188661 184894 188783 186076
rect 187418 184791 188783 184894
rect 194376 186077 195741 186187
rect 194376 184895 194495 186077
rect 195619 184895 195741 186077
rect 194376 184792 195741 184895
rect 201296 186076 202661 186186
rect 201296 184894 201415 186076
rect 202539 184894 202661 186076
rect 201296 184791 202661 184894
rect 208261 186077 209626 186187
rect 208261 184895 208380 186077
rect 209504 184895 209626 186077
rect 208261 184792 209626 184895
rect 215219 186078 216584 186188
rect 215219 184896 215338 186078
rect 216462 184896 216584 186078
rect 215219 184793 216584 184896
rect 222136 186082 223501 186192
rect 222136 184900 222255 186082
rect 223379 184900 223501 186082
rect 222136 184797 223501 184900
rect 229101 186083 230466 186193
rect 229101 184901 229220 186083
rect 230344 184901 230466 186083
rect 229101 184798 230466 184901
rect 236059 186084 237424 186194
rect 236059 184902 236178 186084
rect 237302 184902 237424 186084
rect 236059 184799 237424 184902
rect 242976 186082 244341 186192
rect 242976 184900 243095 186082
rect 244219 184900 244341 186082
rect 242976 184797 244341 184900
rect 249941 186083 251306 186193
rect 249941 184901 250060 186083
rect 251184 184901 251306 186083
rect 249941 184798 251306 184901
rect 256899 186084 258264 186194
rect 256899 184902 257018 186084
rect 258142 184902 258264 186084
rect 256899 184799 258264 184902
rect 264039 186084 265404 186194
rect 264039 184902 264158 186084
rect 265282 184902 265404 186084
rect 264039 184799 265404 184902
rect 270997 186085 272362 186195
rect 270997 184903 271116 186085
rect 272240 184903 272362 186085
rect 270997 184800 272362 184903
rect 278133 186075 279498 186185
rect 278133 184893 278252 186075
rect 279376 184893 279498 186075
rect 278133 184790 279498 184893
rect 76569 179679 77934 179789
rect 76569 178497 76688 179679
rect 77812 178497 77934 179679
rect 76569 178394 77934 178497
rect 83534 179680 84899 179790
rect 83534 178498 83653 179680
rect 84777 178498 84899 179680
rect 83534 178395 84899 178498
rect 90492 179681 91857 179791
rect 90492 178499 90611 179681
rect 91735 178499 91857 179681
rect 90492 178396 91857 178499
rect 97310 179660 98675 179770
rect 97310 178478 97429 179660
rect 98553 178478 98675 179660
rect 97310 178375 98675 178478
rect 104275 179661 105640 179771
rect 104275 178479 104394 179661
rect 105518 178479 105640 179661
rect 104275 178376 105640 178479
rect 111233 179662 112598 179772
rect 111233 178480 111352 179662
rect 112476 178480 112598 179662
rect 111233 178377 112598 178480
rect 118153 179661 119518 179771
rect 118153 178479 118272 179661
rect 119396 178479 119518 179661
rect 118153 178376 119518 178479
rect 125118 179662 126483 179772
rect 125118 178480 125237 179662
rect 126361 178480 126483 179662
rect 125118 178377 126483 178480
rect 132076 179663 133441 179773
rect 132076 178481 132195 179663
rect 133319 178481 133441 179663
rect 132076 178378 133441 178481
rect 138993 179667 140358 179777
rect 138993 178485 139112 179667
rect 140236 178485 140358 179667
rect 138993 178382 140358 178485
rect 145958 179668 147323 179778
rect 145958 178486 146077 179668
rect 147201 178486 147323 179668
rect 145958 178383 147323 178486
rect 152916 179669 154281 179779
rect 152916 178487 153035 179669
rect 154159 178487 154281 179669
rect 152916 178384 154281 178487
rect 159833 179667 161198 179777
rect 159833 178485 159952 179667
rect 161076 178485 161198 179667
rect 159833 178382 161198 178485
rect 166798 179668 168163 179778
rect 166798 178486 166917 179668
rect 168041 178486 168163 179668
rect 166798 178383 168163 178486
rect 173756 179669 175121 179779
rect 173756 178487 173875 179669
rect 174999 178487 175121 179669
rect 173756 178384 175121 178487
rect 180561 179662 181926 179772
rect 180561 178480 180680 179662
rect 181804 178480 181926 179662
rect 180561 178377 181926 178480
rect 187526 179663 188891 179773
rect 187526 178481 187645 179663
rect 188769 178481 188891 179663
rect 187526 178378 188891 178481
rect 194484 179664 195849 179774
rect 194484 178482 194603 179664
rect 195727 178482 195849 179664
rect 194484 178379 195849 178482
rect 201404 179663 202769 179773
rect 201404 178481 201523 179663
rect 202647 178481 202769 179663
rect 201404 178378 202769 178481
rect 208369 179664 209734 179774
rect 208369 178482 208488 179664
rect 209612 178482 209734 179664
rect 208369 178379 209734 178482
rect 215327 179665 216692 179775
rect 215327 178483 215446 179665
rect 216570 178483 216692 179665
rect 215327 178380 216692 178483
rect 222244 179669 223609 179779
rect 222244 178487 222363 179669
rect 223487 178487 223609 179669
rect 222244 178384 223609 178487
rect 229209 179670 230574 179780
rect 229209 178488 229328 179670
rect 230452 178488 230574 179670
rect 229209 178385 230574 178488
rect 236167 179671 237532 179781
rect 236167 178489 236286 179671
rect 237410 178489 237532 179671
rect 236167 178386 237532 178489
rect 243084 179669 244449 179779
rect 243084 178487 243203 179669
rect 244327 178487 244449 179669
rect 243084 178384 244449 178487
rect 250049 179670 251414 179780
rect 250049 178488 250168 179670
rect 251292 178488 251414 179670
rect 250049 178385 251414 178488
rect 257007 179671 258372 179781
rect 257007 178489 257126 179671
rect 258250 178489 258372 179671
rect 257007 178386 258372 178489
rect 264147 179671 265512 179781
rect 264147 178489 264266 179671
rect 265390 178489 265512 179671
rect 264147 178386 265512 178489
rect 271105 179672 272470 179782
rect 271105 178490 271224 179672
rect 272348 178490 272470 179672
rect 271105 178387 272470 178490
rect 278241 179662 279606 179772
rect 278241 178480 278360 179662
rect 279484 178480 279606 179662
rect 278241 178377 279606 178480
rect 48527 173761 49892 173871
rect 48527 172579 48646 173761
rect 49770 172579 49892 173761
rect 48527 172476 49892 172579
rect 55444 173765 56809 173875
rect 55444 172583 55563 173765
rect 56687 172583 56809 173765
rect 55444 172480 56809 172583
rect 62409 173766 63774 173876
rect 62409 172584 62528 173766
rect 63652 172584 63774 173766
rect 62409 172481 63774 172584
rect 69367 173767 70732 173877
rect 69367 172585 69486 173767
rect 70610 172585 70732 173767
rect 69367 172482 70732 172585
rect 76284 173765 77649 173875
rect 76284 172583 76403 173765
rect 77527 172583 77649 173765
rect 76284 172480 77649 172583
rect 83249 173766 84614 173876
rect 83249 172584 83368 173766
rect 84492 172584 84614 173766
rect 83249 172481 84614 172584
rect 90207 173767 91572 173877
rect 90207 172585 90326 173767
rect 91450 172585 91572 173767
rect 90207 172482 91572 172585
rect 97025 173746 98390 173856
rect 97025 172564 97144 173746
rect 98268 172564 98390 173746
rect 97025 172461 98390 172564
rect 103990 173747 105355 173857
rect 103990 172565 104109 173747
rect 105233 172565 105355 173747
rect 103990 172462 105355 172565
rect 110948 173748 112313 173858
rect 110948 172566 111067 173748
rect 112191 172566 112313 173748
rect 110948 172463 112313 172566
rect 117868 173747 119233 173857
rect 117868 172565 117987 173747
rect 119111 172565 119233 173747
rect 117868 172462 119233 172565
rect 124833 173748 126198 173858
rect 124833 172566 124952 173748
rect 126076 172566 126198 173748
rect 124833 172463 126198 172566
rect 131791 173749 133156 173859
rect 131791 172567 131910 173749
rect 133034 172567 133156 173749
rect 131791 172464 133156 172567
rect 138708 173753 140073 173863
rect 138708 172571 138827 173753
rect 139951 172571 140073 173753
rect 138708 172468 140073 172571
rect 145673 173754 147038 173864
rect 145673 172572 145792 173754
rect 146916 172572 147038 173754
rect 145673 172469 147038 172572
rect 152631 173755 153996 173865
rect 152631 172573 152750 173755
rect 153874 172573 153996 173755
rect 152631 172470 153996 172573
rect 159548 173753 160913 173863
rect 159548 172571 159667 173753
rect 160791 172571 160913 173753
rect 159548 172468 160913 172571
rect 166513 173754 167878 173864
rect 166513 172572 166632 173754
rect 167756 172572 167878 173754
rect 166513 172469 167878 172572
rect 173471 173755 174836 173865
rect 173471 172573 173590 173755
rect 174714 172573 174836 173755
rect 173471 172470 174836 172573
rect 180276 173748 181641 173858
rect 180276 172566 180395 173748
rect 181519 172566 181641 173748
rect 180276 172463 181641 172566
rect 187241 173749 188606 173859
rect 187241 172567 187360 173749
rect 188484 172567 188606 173749
rect 187241 172464 188606 172567
rect 194199 173750 195564 173860
rect 194199 172568 194318 173750
rect 195442 172568 195564 173750
rect 194199 172465 195564 172568
rect 201119 173749 202484 173859
rect 201119 172567 201238 173749
rect 202362 172567 202484 173749
rect 201119 172464 202484 172567
rect 208084 173750 209449 173860
rect 208084 172568 208203 173750
rect 209327 172568 209449 173750
rect 208084 172465 209449 172568
rect 215042 173751 216407 173861
rect 215042 172569 215161 173751
rect 216285 172569 216407 173751
rect 215042 172466 216407 172569
rect 221959 173755 223324 173865
rect 221959 172573 222078 173755
rect 223202 172573 223324 173755
rect 221959 172470 223324 172573
rect 228924 173756 230289 173866
rect 228924 172574 229043 173756
rect 230167 172574 230289 173756
rect 228924 172471 230289 172574
rect 235882 173757 237247 173867
rect 235882 172575 236001 173757
rect 237125 172575 237247 173757
rect 235882 172472 237247 172575
rect 242799 173755 244164 173865
rect 242799 172573 242918 173755
rect 244042 172573 244164 173755
rect 242799 172470 244164 172573
rect 249764 173756 251129 173866
rect 249764 172574 249883 173756
rect 251007 172574 251129 173756
rect 249764 172471 251129 172574
rect 256722 173757 258087 173867
rect 256722 172575 256841 173757
rect 257965 172575 258087 173757
rect 256722 172472 258087 172575
rect 263862 173757 265227 173867
rect 263862 172575 263981 173757
rect 265105 172575 265227 173757
rect 263862 172472 265227 172575
rect 270820 173758 272185 173868
rect 270820 172576 270939 173758
rect 272063 172576 272185 173758
rect 270820 172473 272185 172576
rect 277956 173748 279321 173858
rect 277956 172566 278075 173748
rect 279199 172566 279321 173748
rect 277956 172463 279321 172566
rect 48635 167348 50000 167458
rect 48635 166166 48754 167348
rect 49878 166166 50000 167348
rect 48635 166063 50000 166166
rect 55552 167352 56917 167462
rect 55552 166170 55671 167352
rect 56795 166170 56917 167352
rect 55552 166067 56917 166170
rect 62517 167353 63882 167463
rect 62517 166171 62636 167353
rect 63760 166171 63882 167353
rect 62517 166068 63882 166171
rect 69475 167354 70840 167464
rect 69475 166172 69594 167354
rect 70718 166172 70840 167354
rect 69475 166069 70840 166172
rect 76392 167352 77757 167462
rect 76392 166170 76511 167352
rect 77635 166170 77757 167352
rect 76392 166067 77757 166170
rect 83357 167353 84722 167463
rect 83357 166171 83476 167353
rect 84600 166171 84722 167353
rect 83357 166068 84722 166171
rect 90315 167354 91680 167464
rect 90315 166172 90434 167354
rect 91558 166172 91680 167354
rect 90315 166069 91680 166172
rect 97133 167333 98498 167443
rect 97133 166151 97252 167333
rect 98376 166151 98498 167333
rect 97133 166048 98498 166151
rect 104098 167334 105463 167444
rect 104098 166152 104217 167334
rect 105341 166152 105463 167334
rect 104098 166049 105463 166152
rect 111056 167335 112421 167445
rect 111056 166153 111175 167335
rect 112299 166153 112421 167335
rect 111056 166050 112421 166153
rect 117976 167334 119341 167444
rect 117976 166152 118095 167334
rect 119219 166152 119341 167334
rect 117976 166049 119341 166152
rect 124941 167335 126306 167445
rect 124941 166153 125060 167335
rect 126184 166153 126306 167335
rect 124941 166050 126306 166153
rect 131899 167336 133264 167446
rect 131899 166154 132018 167336
rect 133142 166154 133264 167336
rect 131899 166051 133264 166154
rect 138816 167340 140181 167450
rect 138816 166158 138935 167340
rect 140059 166158 140181 167340
rect 138816 166055 140181 166158
rect 145781 167341 147146 167451
rect 145781 166159 145900 167341
rect 147024 166159 147146 167341
rect 145781 166056 147146 166159
rect 152739 167342 154104 167452
rect 152739 166160 152858 167342
rect 153982 166160 154104 167342
rect 152739 166057 154104 166160
rect 159656 167340 161021 167450
rect 159656 166158 159775 167340
rect 160899 166158 161021 167340
rect 159656 166055 161021 166158
rect 166621 167341 167986 167451
rect 166621 166159 166740 167341
rect 167864 166159 167986 167341
rect 166621 166056 167986 166159
rect 173579 167342 174944 167452
rect 173579 166160 173698 167342
rect 174822 166160 174944 167342
rect 173579 166057 174944 166160
rect 180384 167335 181749 167445
rect 180384 166153 180503 167335
rect 181627 166153 181749 167335
rect 180384 166050 181749 166153
rect 187349 167336 188714 167446
rect 187349 166154 187468 167336
rect 188592 166154 188714 167336
rect 187349 166051 188714 166154
rect 194307 167337 195672 167447
rect 194307 166155 194426 167337
rect 195550 166155 195672 167337
rect 194307 166052 195672 166155
rect 201227 167336 202592 167446
rect 201227 166154 201346 167336
rect 202470 166154 202592 167336
rect 201227 166051 202592 166154
rect 208192 167337 209557 167447
rect 208192 166155 208311 167337
rect 209435 166155 209557 167337
rect 208192 166052 209557 166155
rect 215150 167338 216515 167448
rect 215150 166156 215269 167338
rect 216393 166156 216515 167338
rect 215150 166053 216515 166156
rect 222067 167342 223432 167452
rect 222067 166160 222186 167342
rect 223310 166160 223432 167342
rect 222067 166057 223432 166160
rect 229032 167343 230397 167453
rect 229032 166161 229151 167343
rect 230275 166161 230397 167343
rect 229032 166058 230397 166161
rect 235990 167344 237355 167454
rect 235990 166162 236109 167344
rect 237233 166162 237355 167344
rect 235990 166059 237355 166162
rect 242907 167342 244272 167452
rect 242907 166160 243026 167342
rect 244150 166160 244272 167342
rect 242907 166057 244272 166160
rect 249872 167343 251237 167453
rect 249872 166161 249991 167343
rect 251115 166161 251237 167343
rect 249872 166058 251237 166161
rect 256830 167344 258195 167454
rect 256830 166162 256949 167344
rect 258073 166162 258195 167344
rect 256830 166059 258195 166162
rect 263970 167344 265335 167454
rect 263970 166162 264089 167344
rect 265213 166162 265335 167344
rect 263970 166059 265335 166162
rect 270928 167345 272293 167455
rect 270928 166163 271047 167345
rect 272171 166163 272293 167345
rect 270928 166060 272293 166163
rect 278064 167335 279429 167445
rect 278064 166153 278183 167335
rect 279307 166153 279429 167335
rect 278064 166050 279429 166153
rect 21601 160007 22966 160117
rect 21601 158825 21720 160007
rect 22844 158825 22966 160007
rect 21601 158722 22966 158825
rect 28559 160008 29924 160118
rect 28559 158826 28678 160008
rect 29802 158826 29924 160008
rect 28559 158723 29924 158826
rect 35479 160007 36844 160117
rect 35479 158825 35598 160007
rect 36722 158825 36844 160007
rect 35479 158722 36844 158825
rect 42444 160008 43809 160118
rect 42444 158826 42563 160008
rect 43687 158826 43809 160008
rect 42444 158723 43809 158826
rect 49402 160009 50767 160119
rect 49402 158827 49521 160009
rect 50645 158827 50767 160009
rect 49402 158724 50767 158827
rect 56319 160013 57684 160123
rect 56319 158831 56438 160013
rect 57562 158831 57684 160013
rect 56319 158728 57684 158831
rect 63284 160014 64649 160124
rect 63284 158832 63403 160014
rect 64527 158832 64649 160014
rect 63284 158729 64649 158832
rect 70242 160015 71607 160125
rect 70242 158833 70361 160015
rect 71485 158833 71607 160015
rect 70242 158730 71607 158833
rect 77159 160013 78524 160123
rect 77159 158831 77278 160013
rect 78402 158831 78524 160013
rect 77159 158728 78524 158831
rect 84124 160014 85489 160124
rect 84124 158832 84243 160014
rect 85367 158832 85489 160014
rect 84124 158729 85489 158832
rect 91082 160015 92447 160125
rect 91082 158833 91201 160015
rect 92325 158833 92447 160015
rect 91082 158730 92447 158833
rect 97900 159994 99265 160104
rect 97900 158812 98019 159994
rect 99143 158812 99265 159994
rect 97900 158709 99265 158812
rect 104865 159995 106230 160105
rect 104865 158813 104984 159995
rect 106108 158813 106230 159995
rect 104865 158710 106230 158813
rect 111823 159996 113188 160106
rect 111823 158814 111942 159996
rect 113066 158814 113188 159996
rect 111823 158711 113188 158814
rect 118743 159995 120108 160105
rect 118743 158813 118862 159995
rect 119986 158813 120108 159995
rect 118743 158710 120108 158813
rect 125708 159996 127073 160106
rect 125708 158814 125827 159996
rect 126951 158814 127073 159996
rect 125708 158711 127073 158814
rect 132666 159997 134031 160107
rect 132666 158815 132785 159997
rect 133909 158815 134031 159997
rect 132666 158712 134031 158815
rect 139583 160001 140948 160111
rect 139583 158819 139702 160001
rect 140826 158819 140948 160001
rect 139583 158716 140948 158819
rect 146548 160002 147913 160112
rect 146548 158820 146667 160002
rect 147791 158820 147913 160002
rect 146548 158717 147913 158820
rect 153506 160003 154871 160113
rect 153506 158821 153625 160003
rect 154749 158821 154871 160003
rect 153506 158718 154871 158821
rect 160423 160001 161788 160111
rect 160423 158819 160542 160001
rect 161666 158819 161788 160001
rect 160423 158716 161788 158819
rect 167388 160002 168753 160112
rect 167388 158820 167507 160002
rect 168631 158820 168753 160002
rect 167388 158717 168753 158820
rect 174346 160003 175711 160113
rect 174346 158821 174465 160003
rect 175589 158821 175711 160003
rect 174346 158718 175711 158821
rect 181151 159996 182516 160106
rect 181151 158814 181270 159996
rect 182394 158814 182516 159996
rect 181151 158711 182516 158814
rect 188116 159997 189481 160107
rect 188116 158815 188235 159997
rect 189359 158815 189481 159997
rect 188116 158712 189481 158815
rect 195074 159998 196439 160108
rect 195074 158816 195193 159998
rect 196317 158816 196439 159998
rect 195074 158713 196439 158816
rect 201994 159997 203359 160107
rect 201994 158815 202113 159997
rect 203237 158815 203359 159997
rect 201994 158712 203359 158815
rect 208959 159998 210324 160108
rect 208959 158816 209078 159998
rect 210202 158816 210324 159998
rect 208959 158713 210324 158816
rect 215917 159999 217282 160109
rect 215917 158817 216036 159999
rect 217160 158817 217282 159999
rect 215917 158714 217282 158817
rect 222834 160003 224199 160113
rect 222834 158821 222953 160003
rect 224077 158821 224199 160003
rect 222834 158718 224199 158821
rect 229673 159998 231038 160108
rect 229673 158816 229792 159998
rect 230916 158816 231038 159998
rect 229673 158713 231038 158816
rect 236638 159999 238003 160109
rect 236638 158817 236757 159999
rect 237881 158817 238003 159999
rect 236638 158714 238003 158817
rect 243596 160000 244961 160110
rect 243596 158818 243715 160000
rect 244839 158818 244961 160000
rect 243596 158715 244961 158818
rect 250513 160004 251878 160114
rect 250513 158822 250632 160004
rect 251756 158822 251878 160004
rect 250513 158719 251878 158822
rect 257405 159987 258770 160097
rect 257405 158805 257524 159987
rect 258648 158805 258770 159987
rect 257405 158702 258770 158805
rect 264370 159988 265735 160098
rect 264370 158806 264489 159988
rect 265613 158806 265735 159988
rect 264370 158703 265735 158806
rect 271328 159989 272693 160099
rect 271328 158807 271447 159989
rect 272571 158807 272693 159989
rect 271328 158704 272693 158807
rect 278245 159993 279610 160103
rect 278245 158811 278364 159993
rect 279488 158811 279610 159993
rect 278245 158708 279610 158811
rect 21886 155174 23251 155284
rect 21886 153992 22005 155174
rect 23129 153992 23251 155174
rect 21886 153889 23251 153992
rect 28844 155175 30209 155285
rect 28844 153993 28963 155175
rect 30087 153993 30209 155175
rect 28844 153890 30209 153993
rect 35764 155174 37129 155284
rect 35764 153992 35883 155174
rect 37007 153992 37129 155174
rect 35764 153889 37129 153992
rect 42729 155175 44094 155285
rect 42729 153993 42848 155175
rect 43972 153993 44094 155175
rect 42729 153890 44094 153993
rect 49687 155176 51052 155286
rect 49687 153994 49806 155176
rect 50930 153994 51052 155176
rect 49687 153891 51052 153994
rect 56604 155180 57969 155290
rect 56604 153998 56723 155180
rect 57847 153998 57969 155180
rect 56604 153895 57969 153998
rect 63569 155181 64934 155291
rect 63569 153999 63688 155181
rect 64812 153999 64934 155181
rect 63569 153896 64934 153999
rect 70527 155182 71892 155292
rect 70527 154000 70646 155182
rect 71770 154000 71892 155182
rect 70527 153897 71892 154000
rect 77444 155180 78809 155290
rect 77444 153998 77563 155180
rect 78687 153998 78809 155180
rect 77444 153895 78809 153998
rect 84409 155181 85774 155291
rect 84409 153999 84528 155181
rect 85652 153999 85774 155181
rect 84409 153896 85774 153999
rect 91367 155182 92732 155292
rect 91367 154000 91486 155182
rect 92610 154000 92732 155182
rect 91367 153897 92732 154000
rect 98185 155161 99550 155271
rect 98185 153979 98304 155161
rect 99428 153979 99550 155161
rect 98185 153876 99550 153979
rect 105150 155162 106515 155272
rect 105150 153980 105269 155162
rect 106393 153980 106515 155162
rect 105150 153877 106515 153980
rect 112108 155163 113473 155273
rect 112108 153981 112227 155163
rect 113351 153981 113473 155163
rect 112108 153878 113473 153981
rect 119028 155162 120393 155272
rect 119028 153980 119147 155162
rect 120271 153980 120393 155162
rect 119028 153877 120393 153980
rect 125993 155163 127358 155273
rect 125993 153981 126112 155163
rect 127236 153981 127358 155163
rect 125993 153878 127358 153981
rect 132951 155164 134316 155274
rect 132951 153982 133070 155164
rect 134194 153982 134316 155164
rect 132951 153879 134316 153982
rect 139868 155168 141233 155278
rect 139868 153986 139987 155168
rect 141111 153986 141233 155168
rect 139868 153883 141233 153986
rect 146833 155169 148198 155279
rect 146833 153987 146952 155169
rect 148076 153987 148198 155169
rect 146833 153884 148198 153987
rect 153791 155170 155156 155280
rect 153791 153988 153910 155170
rect 155034 153988 155156 155170
rect 153791 153885 155156 153988
rect 160708 155168 162073 155278
rect 160708 153986 160827 155168
rect 161951 153986 162073 155168
rect 160708 153883 162073 153986
rect 167673 155169 169038 155279
rect 167673 153987 167792 155169
rect 168916 153987 169038 155169
rect 167673 153884 169038 153987
rect 174631 155170 175996 155280
rect 174631 153988 174750 155170
rect 175874 153988 175996 155170
rect 174631 153885 175996 153988
rect 181436 155163 182801 155273
rect 181436 153981 181555 155163
rect 182679 153981 182801 155163
rect 181436 153878 182801 153981
rect 188401 155164 189766 155274
rect 188401 153982 188520 155164
rect 189644 153982 189766 155164
rect 188401 153879 189766 153982
rect 195359 155165 196724 155275
rect 195359 153983 195478 155165
rect 196602 153983 196724 155165
rect 195359 153880 196724 153983
rect 202279 155164 203644 155274
rect 202279 153982 202398 155164
rect 203522 153982 203644 155164
rect 202279 153879 203644 153982
rect 209244 155165 210609 155275
rect 209244 153983 209363 155165
rect 210487 153983 210609 155165
rect 209244 153880 210609 153983
rect 216202 155166 217567 155276
rect 216202 153984 216321 155166
rect 217445 153984 217567 155166
rect 216202 153881 217567 153984
rect 223119 155170 224484 155280
rect 223119 153988 223238 155170
rect 224362 153988 224484 155170
rect 223119 153885 224484 153988
rect 229958 155165 231323 155275
rect 229958 153983 230077 155165
rect 231201 153983 231323 155165
rect 229958 153880 231323 153983
rect 236923 155166 238288 155276
rect 236923 153984 237042 155166
rect 238166 153984 238288 155166
rect 236923 153881 238288 153984
rect 243881 155167 245246 155277
rect 243881 153985 244000 155167
rect 245124 153985 245246 155167
rect 243881 153882 245246 153985
rect 250798 155171 252163 155281
rect 250798 153989 250917 155171
rect 252041 153989 252163 155171
rect 250798 153886 252163 153989
rect 257690 155154 259055 155264
rect 257690 153972 257809 155154
rect 258933 153972 259055 155154
rect 257690 153869 259055 153972
rect 264655 155155 266020 155265
rect 264655 153973 264774 155155
rect 265898 153973 266020 155155
rect 264655 153870 266020 153973
rect 271613 155156 272978 155266
rect 271613 153974 271732 155156
rect 272856 153974 272978 155156
rect 271613 153871 272978 153974
rect 278530 155160 279895 155270
rect 278530 153978 278649 155160
rect 279773 153978 279895 155160
rect 278530 153875 279895 153978
rect 21957 149914 23322 150024
rect 21957 148732 22076 149914
rect 23200 148732 23322 149914
rect 21957 148629 23322 148732
rect 28915 149915 30280 150025
rect 28915 148733 29034 149915
rect 30158 148733 30280 149915
rect 28915 148630 30280 148733
rect 35835 149914 37200 150024
rect 35835 148732 35954 149914
rect 37078 148732 37200 149914
rect 35835 148629 37200 148732
rect 42800 149915 44165 150025
rect 42800 148733 42919 149915
rect 44043 148733 44165 149915
rect 42800 148630 44165 148733
rect 49758 149916 51123 150026
rect 49758 148734 49877 149916
rect 51001 148734 51123 149916
rect 49758 148631 51123 148734
rect 56675 149920 58040 150030
rect 56675 148738 56794 149920
rect 57918 148738 58040 149920
rect 56675 148635 58040 148738
rect 63640 149921 65005 150031
rect 63640 148739 63759 149921
rect 64883 148739 65005 149921
rect 63640 148636 65005 148739
rect 70598 149922 71963 150032
rect 70598 148740 70717 149922
rect 71841 148740 71963 149922
rect 70598 148637 71963 148740
rect 77515 149920 78880 150030
rect 77515 148738 77634 149920
rect 78758 148738 78880 149920
rect 77515 148635 78880 148738
rect 84480 149921 85845 150031
rect 84480 148739 84599 149921
rect 85723 148739 85845 149921
rect 84480 148636 85845 148739
rect 91438 149922 92803 150032
rect 91438 148740 91557 149922
rect 92681 148740 92803 149922
rect 91438 148637 92803 148740
rect 98256 149901 99621 150011
rect 98256 148719 98375 149901
rect 99499 148719 99621 149901
rect 98256 148616 99621 148719
rect 105221 149902 106586 150012
rect 105221 148720 105340 149902
rect 106464 148720 106586 149902
rect 105221 148617 106586 148720
rect 112179 149903 113544 150013
rect 112179 148721 112298 149903
rect 113422 148721 113544 149903
rect 112179 148618 113544 148721
rect 119099 149902 120464 150012
rect 119099 148720 119218 149902
rect 120342 148720 120464 149902
rect 119099 148617 120464 148720
rect 126064 149903 127429 150013
rect 126064 148721 126183 149903
rect 127307 148721 127429 149903
rect 126064 148618 127429 148721
rect 133022 149904 134387 150014
rect 133022 148722 133141 149904
rect 134265 148722 134387 149904
rect 133022 148619 134387 148722
rect 139939 149908 141304 150018
rect 139939 148726 140058 149908
rect 141182 148726 141304 149908
rect 139939 148623 141304 148726
rect 146904 149909 148269 150019
rect 146904 148727 147023 149909
rect 148147 148727 148269 149909
rect 146904 148624 148269 148727
rect 153862 149910 155227 150020
rect 153862 148728 153981 149910
rect 155105 148728 155227 149910
rect 153862 148625 155227 148728
rect 160779 149908 162144 150018
rect 160779 148726 160898 149908
rect 162022 148726 162144 149908
rect 160779 148623 162144 148726
rect 167744 149909 169109 150019
rect 167744 148727 167863 149909
rect 168987 148727 169109 149909
rect 167744 148624 169109 148727
rect 174702 149910 176067 150020
rect 174702 148728 174821 149910
rect 175945 148728 176067 149910
rect 174702 148625 176067 148728
rect 181507 149903 182872 150013
rect 181507 148721 181626 149903
rect 182750 148721 182872 149903
rect 181507 148618 182872 148721
rect 188472 149904 189837 150014
rect 188472 148722 188591 149904
rect 189715 148722 189837 149904
rect 188472 148619 189837 148722
rect 195430 149905 196795 150015
rect 195430 148723 195549 149905
rect 196673 148723 196795 149905
rect 195430 148620 196795 148723
rect 202350 149904 203715 150014
rect 202350 148722 202469 149904
rect 203593 148722 203715 149904
rect 202350 148619 203715 148722
rect 209315 149905 210680 150015
rect 209315 148723 209434 149905
rect 210558 148723 210680 149905
rect 209315 148620 210680 148723
rect 216273 149906 217638 150016
rect 216273 148724 216392 149906
rect 217516 148724 217638 149906
rect 216273 148621 217638 148724
rect 223190 149910 224555 150020
rect 223190 148728 223309 149910
rect 224433 148728 224555 149910
rect 223190 148625 224555 148728
rect 230029 149905 231394 150015
rect 230029 148723 230148 149905
rect 231272 148723 231394 149905
rect 230029 148620 231394 148723
rect 236994 149906 238359 150016
rect 236994 148724 237113 149906
rect 238237 148724 238359 149906
rect 236994 148621 238359 148724
rect 243952 149907 245317 150017
rect 243952 148725 244071 149907
rect 245195 148725 245317 149907
rect 243952 148622 245317 148725
rect 250869 149911 252234 150021
rect 250869 148729 250988 149911
rect 252112 148729 252234 149911
rect 250869 148626 252234 148729
rect 257761 149894 259126 150004
rect 257761 148712 257880 149894
rect 259004 148712 259126 149894
rect 257761 148609 259126 148712
rect 264726 149895 266091 150005
rect 264726 148713 264845 149895
rect 265969 148713 266091 149895
rect 264726 148610 266091 148713
rect 271684 149896 273049 150006
rect 271684 148714 271803 149896
rect 272927 148714 273049 149896
rect 271684 148611 273049 148714
rect 278601 149900 279966 150010
rect 278601 148718 278720 149900
rect 279844 148718 279966 149900
rect 278601 148615 279966 148718
rect 21886 144440 23251 144550
rect 21886 143258 22005 144440
rect 23129 143258 23251 144440
rect 21886 143155 23251 143258
rect 28844 144441 30209 144551
rect 28844 143259 28963 144441
rect 30087 143259 30209 144441
rect 28844 143156 30209 143259
rect 35764 144440 37129 144550
rect 35764 143258 35883 144440
rect 37007 143258 37129 144440
rect 35764 143155 37129 143258
rect 42729 144441 44094 144551
rect 42729 143259 42848 144441
rect 43972 143259 44094 144441
rect 42729 143156 44094 143259
rect 49687 144442 51052 144552
rect 49687 143260 49806 144442
rect 50930 143260 51052 144442
rect 49687 143157 51052 143260
rect 56604 144446 57969 144556
rect 56604 143264 56723 144446
rect 57847 143264 57969 144446
rect 56604 143161 57969 143264
rect 63569 144447 64934 144557
rect 63569 143265 63688 144447
rect 64812 143265 64934 144447
rect 63569 143162 64934 143265
rect 70527 144448 71892 144558
rect 70527 143266 70646 144448
rect 71770 143266 71892 144448
rect 70527 143163 71892 143266
rect 77444 144446 78809 144556
rect 77444 143264 77563 144446
rect 78687 143264 78809 144446
rect 77444 143161 78809 143264
rect 84409 144447 85774 144557
rect 84409 143265 84528 144447
rect 85652 143265 85774 144447
rect 84409 143162 85774 143265
rect 91367 144448 92732 144558
rect 91367 143266 91486 144448
rect 92610 143266 92732 144448
rect 91367 143163 92732 143266
rect 98185 144427 99550 144537
rect 98185 143245 98304 144427
rect 99428 143245 99550 144427
rect 98185 143142 99550 143245
rect 105150 144428 106515 144538
rect 105150 143246 105269 144428
rect 106393 143246 106515 144428
rect 105150 143143 106515 143246
rect 112108 144429 113473 144539
rect 112108 143247 112227 144429
rect 113351 143247 113473 144429
rect 112108 143144 113473 143247
rect 119028 144428 120393 144538
rect 119028 143246 119147 144428
rect 120271 143246 120393 144428
rect 119028 143143 120393 143246
rect 125993 144429 127358 144539
rect 125993 143247 126112 144429
rect 127236 143247 127358 144429
rect 125993 143144 127358 143247
rect 132951 144430 134316 144540
rect 132951 143248 133070 144430
rect 134194 143248 134316 144430
rect 132951 143145 134316 143248
rect 139868 144434 141233 144544
rect 139868 143252 139987 144434
rect 141111 143252 141233 144434
rect 139868 143149 141233 143252
rect 146833 144435 148198 144545
rect 146833 143253 146952 144435
rect 148076 143253 148198 144435
rect 146833 143150 148198 143253
rect 153791 144436 155156 144546
rect 153791 143254 153910 144436
rect 155034 143254 155156 144436
rect 153791 143151 155156 143254
rect 160708 144434 162073 144544
rect 160708 143252 160827 144434
rect 161951 143252 162073 144434
rect 160708 143149 162073 143252
rect 167673 144435 169038 144545
rect 167673 143253 167792 144435
rect 168916 143253 169038 144435
rect 167673 143150 169038 143253
rect 174631 144436 175996 144546
rect 174631 143254 174750 144436
rect 175874 143254 175996 144436
rect 174631 143151 175996 143254
rect 181436 144429 182801 144539
rect 181436 143247 181555 144429
rect 182679 143247 182801 144429
rect 181436 143144 182801 143247
rect 188401 144430 189766 144540
rect 188401 143248 188520 144430
rect 189644 143248 189766 144430
rect 188401 143145 189766 143248
rect 195359 144431 196724 144541
rect 195359 143249 195478 144431
rect 196602 143249 196724 144431
rect 195359 143146 196724 143249
rect 202279 144430 203644 144540
rect 202279 143248 202398 144430
rect 203522 143248 203644 144430
rect 202279 143145 203644 143248
rect 209244 144431 210609 144541
rect 209244 143249 209363 144431
rect 210487 143249 210609 144431
rect 209244 143146 210609 143249
rect 216202 144432 217567 144542
rect 216202 143250 216321 144432
rect 217445 143250 217567 144432
rect 216202 143147 217567 143250
rect 223119 144436 224484 144546
rect 223119 143254 223238 144436
rect 224362 143254 224484 144436
rect 223119 143151 224484 143254
rect 22028 138328 23393 138438
rect 22028 137146 22147 138328
rect 23271 137146 23393 138328
rect 22028 137043 23393 137146
rect 28986 138329 30351 138439
rect 28986 137147 29105 138329
rect 30229 137147 30351 138329
rect 28986 137044 30351 137147
rect 35906 138328 37271 138438
rect 35906 137146 36025 138328
rect 37149 137146 37271 138328
rect 35906 137043 37271 137146
rect 42871 138329 44236 138439
rect 42871 137147 42990 138329
rect 44114 137147 44236 138329
rect 42871 137044 44236 137147
rect 49829 138330 51194 138440
rect 49829 137148 49948 138330
rect 51072 137148 51194 138330
rect 49829 137045 51194 137148
rect 56746 138334 58111 138444
rect 56746 137152 56865 138334
rect 57989 137152 58111 138334
rect 56746 137049 58111 137152
rect 63711 138335 65076 138445
rect 63711 137153 63830 138335
rect 64954 137153 65076 138335
rect 63711 137050 65076 137153
rect 70669 138336 72034 138446
rect 70669 137154 70788 138336
rect 71912 137154 72034 138336
rect 70669 137051 72034 137154
rect 77586 138334 78951 138444
rect 77586 137152 77705 138334
rect 78829 137152 78951 138334
rect 77586 137049 78951 137152
rect 84551 138335 85916 138445
rect 84551 137153 84670 138335
rect 85794 137153 85916 138335
rect 84551 137050 85916 137153
rect 91509 138336 92874 138446
rect 91509 137154 91628 138336
rect 92752 137154 92874 138336
rect 91509 137051 92874 137154
rect 98327 138315 99692 138425
rect 98327 137133 98446 138315
rect 99570 137133 99692 138315
rect 98327 137030 99692 137133
rect 105292 138316 106657 138426
rect 105292 137134 105411 138316
rect 106535 137134 106657 138316
rect 105292 137031 106657 137134
rect 112250 138317 113615 138427
rect 112250 137135 112369 138317
rect 113493 137135 113615 138317
rect 112250 137032 113615 137135
rect 119170 138316 120535 138426
rect 119170 137134 119289 138316
rect 120413 137134 120535 138316
rect 119170 137031 120535 137134
rect 126135 138317 127500 138427
rect 126135 137135 126254 138317
rect 127378 137135 127500 138317
rect 126135 137032 127500 137135
rect 133093 138318 134458 138428
rect 133093 137136 133212 138318
rect 134336 137136 134458 138318
rect 133093 137033 134458 137136
rect 140010 138322 141375 138432
rect 140010 137140 140129 138322
rect 141253 137140 141375 138322
rect 140010 137037 141375 137140
rect 146975 138323 148340 138433
rect 146975 137141 147094 138323
rect 148218 137141 148340 138323
rect 146975 137038 148340 137141
rect 153933 138324 155298 138434
rect 153933 137142 154052 138324
rect 155176 137142 155298 138324
rect 153933 137039 155298 137142
rect 160850 138322 162215 138432
rect 160850 137140 160969 138322
rect 162093 137140 162215 138322
rect 160850 137037 162215 137140
rect 167815 138323 169180 138433
rect 167815 137141 167934 138323
rect 169058 137141 169180 138323
rect 167815 137038 169180 137141
rect 174773 138324 176138 138434
rect 174773 137142 174892 138324
rect 176016 137142 176138 138324
rect 174773 137039 176138 137142
rect 181578 138317 182943 138427
rect 181578 137135 181697 138317
rect 182821 137135 182943 138317
rect 181578 137032 182943 137135
rect 188543 138318 189908 138428
rect 188543 137136 188662 138318
rect 189786 137136 189908 138318
rect 188543 137033 189908 137136
rect 195501 138319 196866 138429
rect 195501 137137 195620 138319
rect 196744 137137 196866 138319
rect 195501 137034 196866 137137
rect 202421 138318 203786 138428
rect 202421 137136 202540 138318
rect 203664 137136 203786 138318
rect 202421 137033 203786 137136
rect 209386 138319 210751 138429
rect 209386 137137 209505 138319
rect 210629 137137 210751 138319
rect 209386 137034 210751 137137
rect 216344 138320 217709 138430
rect 216344 137138 216463 138320
rect 217587 137138 217709 138320
rect 216344 137035 217709 137138
rect 223261 138324 224626 138434
rect 223261 137142 223380 138324
rect 224504 137142 224626 138324
rect 223261 137039 224626 137142
rect 21818 130454 23183 130564
rect 21818 129272 21937 130454
rect 23061 129272 23183 130454
rect 21818 129169 23183 129272
rect 28776 130455 30141 130565
rect 28776 129273 28895 130455
rect 30019 129273 30141 130455
rect 28776 129170 30141 129273
rect 35696 130454 37061 130564
rect 35696 129272 35815 130454
rect 36939 129272 37061 130454
rect 35696 129169 37061 129272
rect 42661 130455 44026 130565
rect 42661 129273 42780 130455
rect 43904 129273 44026 130455
rect 42661 129170 44026 129273
rect 49619 130456 50984 130566
rect 49619 129274 49738 130456
rect 50862 129274 50984 130456
rect 49619 129171 50984 129274
rect 56536 130460 57901 130570
rect 56536 129278 56655 130460
rect 57779 129278 57901 130460
rect 56536 129175 57901 129278
rect 63501 130461 64866 130571
rect 63501 129279 63620 130461
rect 64744 129279 64866 130461
rect 63501 129176 64866 129279
rect 70459 130462 71824 130572
rect 70459 129280 70578 130462
rect 71702 129280 71824 130462
rect 70459 129177 71824 129280
rect 77376 130460 78741 130570
rect 77376 129278 77495 130460
rect 78619 129278 78741 130460
rect 77376 129175 78741 129278
rect 84341 130461 85706 130571
rect 84341 129279 84460 130461
rect 85584 129279 85706 130461
rect 84341 129176 85706 129279
rect 91299 130462 92664 130572
rect 91299 129280 91418 130462
rect 92542 129280 92664 130462
rect 91299 129177 92664 129280
rect 98117 130441 99482 130551
rect 98117 129259 98236 130441
rect 99360 129259 99482 130441
rect 98117 129156 99482 129259
rect 105082 130442 106447 130552
rect 105082 129260 105201 130442
rect 106325 129260 106447 130442
rect 105082 129157 106447 129260
rect 112040 130443 113405 130553
rect 112040 129261 112159 130443
rect 113283 129261 113405 130443
rect 112040 129158 113405 129261
rect 118960 130442 120325 130552
rect 118960 129260 119079 130442
rect 120203 129260 120325 130442
rect 118960 129157 120325 129260
rect 125925 130443 127290 130553
rect 125925 129261 126044 130443
rect 127168 129261 127290 130443
rect 125925 129158 127290 129261
rect 132883 130444 134248 130554
rect 132883 129262 133002 130444
rect 134126 129262 134248 130444
rect 132883 129159 134248 129262
rect 139800 130448 141165 130558
rect 139800 129266 139919 130448
rect 141043 129266 141165 130448
rect 139800 129163 141165 129266
rect 146765 130449 148130 130559
rect 146765 129267 146884 130449
rect 148008 129267 148130 130449
rect 146765 129164 148130 129267
rect 153723 130450 155088 130560
rect 153723 129268 153842 130450
rect 154966 129268 155088 130450
rect 153723 129165 155088 129268
rect 160640 130448 162005 130558
rect 160640 129266 160759 130448
rect 161883 129266 162005 130448
rect 160640 129163 162005 129266
rect 167605 130449 168970 130559
rect 167605 129267 167724 130449
rect 168848 129267 168970 130449
rect 167605 129164 168970 129267
rect 174563 130450 175928 130560
rect 174563 129268 174682 130450
rect 175806 129268 175928 130450
rect 174563 129165 175928 129268
rect 181368 130443 182733 130553
rect 181368 129261 181487 130443
rect 182611 129261 182733 130443
rect 181368 129158 182733 129261
rect 188333 130444 189698 130554
rect 188333 129262 188452 130444
rect 189576 129262 189698 130444
rect 188333 129159 189698 129262
rect 195291 130445 196656 130555
rect 195291 129263 195410 130445
rect 196534 129263 196656 130445
rect 195291 129160 196656 129263
rect 202211 130444 203576 130554
rect 202211 129262 202330 130444
rect 203454 129262 203576 130444
rect 202211 129159 203576 129262
rect 209176 130445 210541 130555
rect 209176 129263 209295 130445
rect 210419 129263 210541 130445
rect 209176 129160 210541 129263
rect 216134 130446 217499 130556
rect 216134 129264 216253 130446
rect 217377 129264 217499 130446
rect 216134 129161 217499 129264
rect 223051 130450 224416 130560
rect 223051 129268 223170 130450
rect 224294 129268 224416 130450
rect 223051 129165 224416 129268
rect 21335 119138 22700 119248
rect 21335 117956 21454 119138
rect 22578 117956 22700 119138
rect 21335 117853 22700 117956
rect 28293 119139 29658 119249
rect 28293 117957 28412 119139
rect 29536 117957 29658 119139
rect 28293 117854 29658 117957
rect 35213 119138 36578 119248
rect 35213 117956 35332 119138
rect 36456 117956 36578 119138
rect 35213 117853 36578 117956
rect 42178 119139 43543 119249
rect 42178 117957 42297 119139
rect 43421 117957 43543 119139
rect 42178 117854 43543 117957
rect 49136 119140 50501 119250
rect 49136 117958 49255 119140
rect 50379 117958 50501 119140
rect 49136 117855 50501 117958
rect 56053 119144 57418 119254
rect 56053 117962 56172 119144
rect 57296 117962 57418 119144
rect 56053 117859 57418 117962
rect 63018 119145 64383 119255
rect 63018 117963 63137 119145
rect 64261 117963 64383 119145
rect 63018 117860 64383 117963
rect 69976 119146 71341 119256
rect 69976 117964 70095 119146
rect 71219 117964 71341 119146
rect 69976 117861 71341 117964
rect 76893 119144 78258 119254
rect 76893 117962 77012 119144
rect 78136 117962 78258 119144
rect 76893 117859 78258 117962
rect 83858 119145 85223 119255
rect 83858 117963 83977 119145
rect 85101 117963 85223 119145
rect 83858 117860 85223 117963
rect 90816 119146 92181 119256
rect 90816 117964 90935 119146
rect 92059 117964 92181 119146
rect 90816 117861 92181 117964
rect 97634 119125 98999 119235
rect 97634 117943 97753 119125
rect 98877 117943 98999 119125
rect 97634 117840 98999 117943
rect 104599 119126 105964 119236
rect 104599 117944 104718 119126
rect 105842 117944 105964 119126
rect 104599 117841 105964 117944
rect 111557 119127 112922 119237
rect 111557 117945 111676 119127
rect 112800 117945 112922 119127
rect 111557 117842 112922 117945
rect 118477 119126 119842 119236
rect 118477 117944 118596 119126
rect 119720 117944 119842 119126
rect 118477 117841 119842 117944
rect 125442 119127 126807 119237
rect 125442 117945 125561 119127
rect 126685 117945 126807 119127
rect 125442 117842 126807 117945
rect 132400 119128 133765 119238
rect 132400 117946 132519 119128
rect 133643 117946 133765 119128
rect 132400 117843 133765 117946
rect 139317 119132 140682 119242
rect 139317 117950 139436 119132
rect 140560 117950 140682 119132
rect 139317 117847 140682 117950
rect 146282 119133 147647 119243
rect 146282 117951 146401 119133
rect 147525 117951 147647 119133
rect 146282 117848 147647 117951
rect 153240 119134 154605 119244
rect 153240 117952 153359 119134
rect 154483 117952 154605 119134
rect 153240 117849 154605 117952
rect 160157 119132 161522 119242
rect 160157 117950 160276 119132
rect 161400 117950 161522 119132
rect 160157 117847 161522 117950
rect 167122 119133 168487 119243
rect 167122 117951 167241 119133
rect 168365 117951 168487 119133
rect 167122 117848 168487 117951
rect 174080 119134 175445 119244
rect 174080 117952 174199 119134
rect 175323 117952 175445 119134
rect 174080 117849 175445 117952
rect 180885 119127 182250 119237
rect 180885 117945 181004 119127
rect 182128 117945 182250 119127
rect 180885 117842 182250 117945
rect 187850 119128 189215 119238
rect 187850 117946 187969 119128
rect 189093 117946 189215 119128
rect 187850 117843 189215 117946
rect 194808 119129 196173 119239
rect 194808 117947 194927 119129
rect 196051 117947 196173 119129
rect 194808 117844 196173 117947
rect 201728 119128 203093 119238
rect 201728 117946 201847 119128
rect 202971 117946 203093 119128
rect 201728 117843 203093 117946
rect 208693 119129 210058 119239
rect 208693 117947 208812 119129
rect 209936 117947 210058 119129
rect 208693 117844 210058 117947
rect 215651 119130 217016 119240
rect 215651 117948 215770 119130
rect 216894 117948 217016 119130
rect 215651 117845 217016 117948
rect 222568 119134 223933 119244
rect 222568 117952 222687 119134
rect 223811 117952 223933 119134
rect 222568 117849 223933 117952
rect 229533 119135 230898 119245
rect 229533 117953 229652 119135
rect 230776 117953 230898 119135
rect 229533 117850 230898 117953
rect 236491 119136 237856 119246
rect 236491 117954 236610 119136
rect 237734 117954 237856 119136
rect 236491 117851 237856 117954
rect 243408 119134 244773 119244
rect 243408 117952 243527 119134
rect 244651 117952 244773 119134
rect 243408 117849 244773 117952
rect 250373 119135 251738 119245
rect 250373 117953 250492 119135
rect 251616 117953 251738 119135
rect 250373 117850 251738 117953
rect 257331 119136 258696 119246
rect 257331 117954 257450 119136
rect 258574 117954 258696 119136
rect 257331 117851 258696 117954
rect 264471 119136 265836 119246
rect 264471 117954 264590 119136
rect 265714 117954 265836 119136
rect 264471 117851 265836 117954
rect 271429 119137 272794 119247
rect 271429 117955 271548 119137
rect 272672 117955 272794 119137
rect 271429 117852 272794 117955
rect 278565 119127 279930 119237
rect 278565 117945 278684 119127
rect 279808 117945 279930 119127
rect 278565 117842 279930 117945
rect 21540 111186 22905 111296
rect 21540 110004 21659 111186
rect 22783 110004 22905 111186
rect 21540 109901 22905 110004
rect 28498 111187 29863 111297
rect 28498 110005 28617 111187
rect 29741 110005 29863 111187
rect 28498 109902 29863 110005
rect 35418 111186 36783 111296
rect 35418 110004 35537 111186
rect 36661 110004 36783 111186
rect 35418 109901 36783 110004
rect 42383 111187 43748 111297
rect 42383 110005 42502 111187
rect 43626 110005 43748 111187
rect 42383 109902 43748 110005
rect 49341 111188 50706 111298
rect 49341 110006 49460 111188
rect 50584 110006 50706 111188
rect 49341 109903 50706 110006
rect 56258 111192 57623 111302
rect 56258 110010 56377 111192
rect 57501 110010 57623 111192
rect 56258 109907 57623 110010
rect 63223 111193 64588 111303
rect 63223 110011 63342 111193
rect 64466 110011 64588 111193
rect 63223 109908 64588 110011
rect 70181 111194 71546 111304
rect 70181 110012 70300 111194
rect 71424 110012 71546 111194
rect 70181 109909 71546 110012
rect 77098 111192 78463 111302
rect 77098 110010 77217 111192
rect 78341 110010 78463 111192
rect 77098 109907 78463 110010
rect 84063 111193 85428 111303
rect 84063 110011 84182 111193
rect 85306 110011 85428 111193
rect 84063 109908 85428 110011
rect 91021 111194 92386 111304
rect 91021 110012 91140 111194
rect 92264 110012 92386 111194
rect 91021 109909 92386 110012
rect 97839 111173 99204 111283
rect 97839 109991 97958 111173
rect 99082 109991 99204 111173
rect 97839 109888 99204 109991
rect 104804 111174 106169 111284
rect 104804 109992 104923 111174
rect 106047 109992 106169 111174
rect 104804 109889 106169 109992
rect 111762 111175 113127 111285
rect 111762 109993 111881 111175
rect 113005 109993 113127 111175
rect 111762 109890 113127 109993
rect 118682 111174 120047 111284
rect 118682 109992 118801 111174
rect 119925 109992 120047 111174
rect 118682 109889 120047 109992
rect 125647 111175 127012 111285
rect 125647 109993 125766 111175
rect 126890 109993 127012 111175
rect 125647 109890 127012 109993
rect 132605 111176 133970 111286
rect 132605 109994 132724 111176
rect 133848 109994 133970 111176
rect 132605 109891 133970 109994
rect 139522 111180 140887 111290
rect 139522 109998 139641 111180
rect 140765 109998 140887 111180
rect 139522 109895 140887 109998
rect 146487 111181 147852 111291
rect 146487 109999 146606 111181
rect 147730 109999 147852 111181
rect 146487 109896 147852 109999
rect 153445 111182 154810 111292
rect 153445 110000 153564 111182
rect 154688 110000 154810 111182
rect 153445 109897 154810 110000
rect 160362 111180 161727 111290
rect 160362 109998 160481 111180
rect 161605 109998 161727 111180
rect 160362 109895 161727 109998
rect 167327 111181 168692 111291
rect 167327 109999 167446 111181
rect 168570 109999 168692 111181
rect 167327 109896 168692 109999
rect 174285 111182 175650 111292
rect 174285 110000 174404 111182
rect 175528 110000 175650 111182
rect 174285 109897 175650 110000
rect 181090 111175 182455 111285
rect 181090 109993 181209 111175
rect 182333 109993 182455 111175
rect 181090 109890 182455 109993
rect 188055 111176 189420 111286
rect 188055 109994 188174 111176
rect 189298 109994 189420 111176
rect 188055 109891 189420 109994
rect 195013 111177 196378 111287
rect 195013 109995 195132 111177
rect 196256 109995 196378 111177
rect 195013 109892 196378 109995
rect 201933 111176 203298 111286
rect 201933 109994 202052 111176
rect 203176 109994 203298 111176
rect 201933 109891 203298 109994
rect 208898 111177 210263 111287
rect 208898 109995 209017 111177
rect 210141 109995 210263 111177
rect 208898 109892 210263 109995
rect 215856 111178 217221 111288
rect 215856 109996 215975 111178
rect 217099 109996 217221 111178
rect 215856 109893 217221 109996
rect 222773 111182 224138 111292
rect 222773 110000 222892 111182
rect 224016 110000 224138 111182
rect 222773 109897 224138 110000
rect 229738 111183 231103 111293
rect 229738 110001 229857 111183
rect 230981 110001 231103 111183
rect 229738 109898 231103 110001
rect 236696 111184 238061 111294
rect 236696 110002 236815 111184
rect 237939 110002 238061 111184
rect 236696 109899 238061 110002
rect 243613 111182 244978 111292
rect 243613 110000 243732 111182
rect 244856 110000 244978 111182
rect 243613 109897 244978 110000
rect 250578 111183 251943 111293
rect 250578 110001 250697 111183
rect 251821 110001 251943 111183
rect 250578 109898 251943 110001
rect 257536 111184 258901 111294
rect 257536 110002 257655 111184
rect 258779 110002 258901 111184
rect 257536 109899 258901 110002
rect 264676 111184 266041 111294
rect 264676 110002 264795 111184
rect 265919 110002 266041 111184
rect 264676 109899 266041 110002
rect 271634 111185 272999 111295
rect 271634 110003 271753 111185
rect 272877 110003 272999 111185
rect 271634 109900 272999 110003
rect 278770 111175 280135 111285
rect 278770 109993 278889 111175
rect 280013 109993 280135 111175
rect 278770 109890 280135 109993
rect 21540 102960 22905 103070
rect 21540 101778 21659 102960
rect 22783 101778 22905 102960
rect 21540 101675 22905 101778
rect 28498 102961 29863 103071
rect 28498 101779 28617 102961
rect 29741 101779 29863 102961
rect 28498 101676 29863 101779
rect 35418 102960 36783 103070
rect 35418 101778 35537 102960
rect 36661 101778 36783 102960
rect 35418 101675 36783 101778
rect 42383 102961 43748 103071
rect 42383 101779 42502 102961
rect 43626 101779 43748 102961
rect 42383 101676 43748 101779
rect 49341 102962 50706 103072
rect 49341 101780 49460 102962
rect 50584 101780 50706 102962
rect 49341 101677 50706 101780
rect 56258 102966 57623 103076
rect 56258 101784 56377 102966
rect 57501 101784 57623 102966
rect 56258 101681 57623 101784
rect 63223 102967 64588 103077
rect 63223 101785 63342 102967
rect 64466 101785 64588 102967
rect 63223 101682 64588 101785
rect 70181 102968 71546 103078
rect 70181 101786 70300 102968
rect 71424 101786 71546 102968
rect 70181 101683 71546 101786
rect 77098 102966 78463 103076
rect 77098 101784 77217 102966
rect 78341 101784 78463 102966
rect 77098 101681 78463 101784
rect 84063 102967 85428 103077
rect 84063 101785 84182 102967
rect 85306 101785 85428 102967
rect 84063 101682 85428 101785
rect 91021 102968 92386 103078
rect 91021 101786 91140 102968
rect 92264 101786 92386 102968
rect 91021 101683 92386 101786
rect 97839 102947 99204 103057
rect 97839 101765 97958 102947
rect 99082 101765 99204 102947
rect 97839 101662 99204 101765
rect 104804 102948 106169 103058
rect 104804 101766 104923 102948
rect 106047 101766 106169 102948
rect 104804 101663 106169 101766
rect 111762 102949 113127 103059
rect 111762 101767 111881 102949
rect 113005 101767 113127 102949
rect 111762 101664 113127 101767
rect 118682 102948 120047 103058
rect 118682 101766 118801 102948
rect 119925 101766 120047 102948
rect 118682 101663 120047 101766
rect 125647 102949 127012 103059
rect 125647 101767 125766 102949
rect 126890 101767 127012 102949
rect 125647 101664 127012 101767
rect 132605 102950 133970 103060
rect 132605 101768 132724 102950
rect 133848 101768 133970 102950
rect 132605 101665 133970 101768
rect 139522 102954 140887 103064
rect 139522 101772 139641 102954
rect 140765 101772 140887 102954
rect 139522 101669 140887 101772
rect 146487 102955 147852 103065
rect 146487 101773 146606 102955
rect 147730 101773 147852 102955
rect 146487 101670 147852 101773
rect 153445 102956 154810 103066
rect 153445 101774 153564 102956
rect 154688 101774 154810 102956
rect 153445 101671 154810 101774
rect 160362 102954 161727 103064
rect 160362 101772 160481 102954
rect 161605 101772 161727 102954
rect 160362 101669 161727 101772
rect 167327 102955 168692 103065
rect 167327 101773 167446 102955
rect 168570 101773 168692 102955
rect 167327 101670 168692 101773
rect 174285 102956 175650 103066
rect 174285 101774 174404 102956
rect 175528 101774 175650 102956
rect 174285 101671 175650 101774
rect 181090 102949 182455 103059
rect 181090 101767 181209 102949
rect 182333 101767 182455 102949
rect 181090 101664 182455 101767
rect 188055 102950 189420 103060
rect 188055 101768 188174 102950
rect 189298 101768 189420 102950
rect 188055 101665 189420 101768
rect 195013 102951 196378 103061
rect 195013 101769 195132 102951
rect 196256 101769 196378 102951
rect 195013 101666 196378 101769
rect 201933 102950 203298 103060
rect 201933 101768 202052 102950
rect 203176 101768 203298 102950
rect 201933 101665 203298 101768
rect 208898 102951 210263 103061
rect 208898 101769 209017 102951
rect 210141 101769 210263 102951
rect 208898 101666 210263 101769
rect 215856 102952 217221 103062
rect 215856 101770 215975 102952
rect 217099 101770 217221 102952
rect 215856 101667 217221 101770
rect 222773 102956 224138 103066
rect 222773 101774 222892 102956
rect 224016 101774 224138 102956
rect 222773 101671 224138 101774
rect 229738 102957 231103 103067
rect 229738 101775 229857 102957
rect 230981 101775 231103 102957
rect 229738 101672 231103 101775
rect 236696 102958 238061 103068
rect 236696 101776 236815 102958
rect 237939 101776 238061 102958
rect 236696 101673 238061 101776
rect 243613 102956 244978 103066
rect 243613 101774 243732 102956
rect 244856 101774 244978 102956
rect 243613 101671 244978 101774
rect 250578 102957 251943 103067
rect 250578 101775 250697 102957
rect 251821 101775 251943 102957
rect 250578 101672 251943 101775
rect 257536 102958 258901 103068
rect 257536 101776 257655 102958
rect 258779 101776 258901 102958
rect 257536 101673 258901 101776
rect 264676 102958 266041 103068
rect 264676 101776 264795 102958
rect 265919 101776 266041 102958
rect 264676 101673 266041 101776
rect 271634 102959 272999 103069
rect 271634 101777 271753 102959
rect 272877 101777 272999 102959
rect 271634 101674 272999 101777
rect 278770 102949 280135 103059
rect 278770 101767 278889 102949
rect 280013 101767 280135 102949
rect 278770 101664 280135 101767
rect 21335 95556 22700 95666
rect 21335 94374 21454 95556
rect 22578 94374 22700 95556
rect 21335 94271 22700 94374
rect 28293 95557 29658 95667
rect 28293 94375 28412 95557
rect 29536 94375 29658 95557
rect 28293 94272 29658 94375
rect 35213 95556 36578 95666
rect 35213 94374 35332 95556
rect 36456 94374 36578 95556
rect 35213 94271 36578 94374
rect 42178 95557 43543 95667
rect 42178 94375 42297 95557
rect 43421 94375 43543 95557
rect 42178 94272 43543 94375
rect 49136 95558 50501 95668
rect 49136 94376 49255 95558
rect 50379 94376 50501 95558
rect 49136 94273 50501 94376
rect 56053 95562 57418 95672
rect 56053 94380 56172 95562
rect 57296 94380 57418 95562
rect 56053 94277 57418 94380
rect 63018 95563 64383 95673
rect 63018 94381 63137 95563
rect 64261 94381 64383 95563
rect 63018 94278 64383 94381
rect 69976 95564 71341 95674
rect 69976 94382 70095 95564
rect 71219 94382 71341 95564
rect 69976 94279 71341 94382
rect 76893 95562 78258 95672
rect 76893 94380 77012 95562
rect 78136 94380 78258 95562
rect 76893 94277 78258 94380
rect 83858 95563 85223 95673
rect 83858 94381 83977 95563
rect 85101 94381 85223 95563
rect 83858 94278 85223 94381
rect 90816 95564 92181 95674
rect 90816 94382 90935 95564
rect 92059 94382 92181 95564
rect 90816 94279 92181 94382
rect 97634 95543 98999 95653
rect 97634 94361 97753 95543
rect 98877 94361 98999 95543
rect 97634 94258 98999 94361
rect 104599 95544 105964 95654
rect 104599 94362 104718 95544
rect 105842 94362 105964 95544
rect 104599 94259 105964 94362
rect 111557 95545 112922 95655
rect 111557 94363 111676 95545
rect 112800 94363 112922 95545
rect 111557 94260 112922 94363
rect 118477 95544 119842 95654
rect 118477 94362 118596 95544
rect 119720 94362 119842 95544
rect 118477 94259 119842 94362
rect 125442 95545 126807 95655
rect 125442 94363 125561 95545
rect 126685 94363 126807 95545
rect 125442 94260 126807 94363
rect 132400 95546 133765 95656
rect 132400 94364 132519 95546
rect 133643 94364 133765 95546
rect 132400 94261 133765 94364
rect 139317 95550 140682 95660
rect 139317 94368 139436 95550
rect 140560 94368 140682 95550
rect 139317 94265 140682 94368
rect 146282 95551 147647 95661
rect 146282 94369 146401 95551
rect 147525 94369 147647 95551
rect 146282 94266 147647 94369
rect 153240 95552 154605 95662
rect 153240 94370 153359 95552
rect 154483 94370 154605 95552
rect 153240 94267 154605 94370
rect 160157 95550 161522 95660
rect 160157 94368 160276 95550
rect 161400 94368 161522 95550
rect 160157 94265 161522 94368
rect 167122 95551 168487 95661
rect 167122 94369 167241 95551
rect 168365 94369 168487 95551
rect 167122 94266 168487 94369
rect 174080 95552 175445 95662
rect 174080 94370 174199 95552
rect 175323 94370 175445 95552
rect 174080 94267 175445 94370
rect 180885 95545 182250 95655
rect 180885 94363 181004 95545
rect 182128 94363 182250 95545
rect 180885 94260 182250 94363
rect 187850 95546 189215 95656
rect 187850 94364 187969 95546
rect 189093 94364 189215 95546
rect 187850 94261 189215 94364
rect 194808 95547 196173 95657
rect 194808 94365 194927 95547
rect 196051 94365 196173 95547
rect 194808 94262 196173 94365
rect 201728 95546 203093 95656
rect 201728 94364 201847 95546
rect 202971 94364 203093 95546
rect 201728 94261 203093 94364
rect 208693 95547 210058 95657
rect 208693 94365 208812 95547
rect 209936 94365 210058 95547
rect 208693 94262 210058 94365
rect 215651 95548 217016 95658
rect 215651 94366 215770 95548
rect 216894 94366 217016 95548
rect 215651 94263 217016 94366
rect 222568 95552 223933 95662
rect 222568 94370 222687 95552
rect 223811 94370 223933 95552
rect 222568 94267 223933 94370
rect 229533 95553 230898 95663
rect 229533 94371 229652 95553
rect 230776 94371 230898 95553
rect 229533 94268 230898 94371
rect 236491 95554 237856 95664
rect 236491 94372 236610 95554
rect 237734 94372 237856 95554
rect 236491 94269 237856 94372
rect 243408 95552 244773 95662
rect 243408 94370 243527 95552
rect 244651 94370 244773 95552
rect 243408 94267 244773 94370
rect 250373 95553 251738 95663
rect 250373 94371 250492 95553
rect 251616 94371 251738 95553
rect 250373 94268 251738 94371
rect 257331 95554 258696 95664
rect 257331 94372 257450 95554
rect 258574 94372 258696 95554
rect 257331 94269 258696 94372
rect 264471 95554 265836 95664
rect 264471 94372 264590 95554
rect 265714 94372 265836 95554
rect 264471 94269 265836 94372
rect 271429 95555 272794 95665
rect 271429 94373 271548 95555
rect 272672 94373 272794 95555
rect 271429 94270 272794 94373
rect 278565 95545 279930 95655
rect 278565 94363 278684 95545
rect 279808 94363 279930 95545
rect 278565 94260 279930 94363
rect 21061 88426 22426 88536
rect 21061 87244 21180 88426
rect 22304 87244 22426 88426
rect 21061 87141 22426 87244
rect 28019 88427 29384 88537
rect 28019 87245 28138 88427
rect 29262 87245 29384 88427
rect 28019 87142 29384 87245
rect 34939 88426 36304 88536
rect 34939 87244 35058 88426
rect 36182 87244 36304 88426
rect 34939 87141 36304 87244
rect 41904 88427 43269 88537
rect 41904 87245 42023 88427
rect 43147 87245 43269 88427
rect 41904 87142 43269 87245
rect 48862 88428 50227 88538
rect 48862 87246 48981 88428
rect 50105 87246 50227 88428
rect 48862 87143 50227 87246
rect 55779 88432 57144 88542
rect 55779 87250 55898 88432
rect 57022 87250 57144 88432
rect 55779 87147 57144 87250
rect 62744 88433 64109 88543
rect 62744 87251 62863 88433
rect 63987 87251 64109 88433
rect 62744 87148 64109 87251
rect 69702 88434 71067 88544
rect 69702 87252 69821 88434
rect 70945 87252 71067 88434
rect 69702 87149 71067 87252
rect 76619 88432 77984 88542
rect 76619 87250 76738 88432
rect 77862 87250 77984 88432
rect 76619 87147 77984 87250
rect 83584 88433 84949 88543
rect 83584 87251 83703 88433
rect 84827 87251 84949 88433
rect 83584 87148 84949 87251
rect 90542 88434 91907 88544
rect 90542 87252 90661 88434
rect 91785 87252 91907 88434
rect 90542 87149 91907 87252
rect 97360 88413 98725 88523
rect 97360 87231 97479 88413
rect 98603 87231 98725 88413
rect 97360 87128 98725 87231
rect 104325 88414 105690 88524
rect 104325 87232 104444 88414
rect 105568 87232 105690 88414
rect 104325 87129 105690 87232
rect 111283 88415 112648 88525
rect 111283 87233 111402 88415
rect 112526 87233 112648 88415
rect 111283 87130 112648 87233
rect 118203 88414 119568 88524
rect 118203 87232 118322 88414
rect 119446 87232 119568 88414
rect 118203 87129 119568 87232
rect 125168 88415 126533 88525
rect 125168 87233 125287 88415
rect 126411 87233 126533 88415
rect 125168 87130 126533 87233
rect 132126 88416 133491 88526
rect 132126 87234 132245 88416
rect 133369 87234 133491 88416
rect 132126 87131 133491 87234
rect 139043 88420 140408 88530
rect 139043 87238 139162 88420
rect 140286 87238 140408 88420
rect 139043 87135 140408 87238
rect 146008 88421 147373 88531
rect 146008 87239 146127 88421
rect 147251 87239 147373 88421
rect 146008 87136 147373 87239
rect 152966 88422 154331 88532
rect 152966 87240 153085 88422
rect 154209 87240 154331 88422
rect 152966 87137 154331 87240
rect 159883 88420 161248 88530
rect 159883 87238 160002 88420
rect 161126 87238 161248 88420
rect 159883 87135 161248 87238
rect 166848 88421 168213 88531
rect 166848 87239 166967 88421
rect 168091 87239 168213 88421
rect 166848 87136 168213 87239
rect 173806 88422 175171 88532
rect 173806 87240 173925 88422
rect 175049 87240 175171 88422
rect 173806 87137 175171 87240
rect 180611 88415 181976 88525
rect 180611 87233 180730 88415
rect 181854 87233 181976 88415
rect 180611 87130 181976 87233
rect 187576 88416 188941 88526
rect 187576 87234 187695 88416
rect 188819 87234 188941 88416
rect 187576 87131 188941 87234
rect 194534 88417 195899 88527
rect 194534 87235 194653 88417
rect 195777 87235 195899 88417
rect 194534 87132 195899 87235
rect 201454 88416 202819 88526
rect 201454 87234 201573 88416
rect 202697 87234 202819 88416
rect 201454 87131 202819 87234
rect 208419 88417 209784 88527
rect 208419 87235 208538 88417
rect 209662 87235 209784 88417
rect 208419 87132 209784 87235
rect 215377 88418 216742 88528
rect 215377 87236 215496 88418
rect 216620 87236 216742 88418
rect 215377 87133 216742 87236
rect 222294 88422 223659 88532
rect 222294 87240 222413 88422
rect 223537 87240 223659 88422
rect 222294 87137 223659 87240
rect 229259 88423 230624 88533
rect 229259 87241 229378 88423
rect 230502 87241 230624 88423
rect 229259 87138 230624 87241
rect 236217 88424 237582 88534
rect 236217 87242 236336 88424
rect 237460 87242 237582 88424
rect 236217 87139 237582 87242
rect 243134 88422 244499 88532
rect 243134 87240 243253 88422
rect 244377 87240 244499 88422
rect 243134 87137 244499 87240
rect 250099 88423 251464 88533
rect 250099 87241 250218 88423
rect 251342 87241 251464 88423
rect 250099 87138 251464 87241
rect 257057 88424 258422 88534
rect 257057 87242 257176 88424
rect 258300 87242 258422 88424
rect 257057 87139 258422 87242
rect 264197 88424 265562 88534
rect 264197 87242 264316 88424
rect 265440 87242 265562 88424
rect 264197 87139 265562 87242
rect 271155 88425 272520 88535
rect 271155 87243 271274 88425
rect 272398 87243 272520 88425
rect 271155 87140 272520 87243
rect 278291 88415 279656 88525
rect 278291 87233 278410 88415
rect 279534 87233 279656 88415
rect 278291 87130 279656 87233
rect 21169 82013 22534 82123
rect 21169 80831 21288 82013
rect 22412 80831 22534 82013
rect 21169 80728 22534 80831
rect 28127 82014 29492 82124
rect 28127 80832 28246 82014
rect 29370 80832 29492 82014
rect 28127 80729 29492 80832
rect 35047 82013 36412 82123
rect 35047 80831 35166 82013
rect 36290 80831 36412 82013
rect 35047 80728 36412 80831
rect 42012 82014 43377 82124
rect 42012 80832 42131 82014
rect 43255 80832 43377 82014
rect 42012 80729 43377 80832
rect 48970 82015 50335 82125
rect 48970 80833 49089 82015
rect 50213 80833 50335 82015
rect 48970 80730 50335 80833
rect 55887 82019 57252 82129
rect 55887 80837 56006 82019
rect 57130 80837 57252 82019
rect 55887 80734 57252 80837
rect 62852 82020 64217 82130
rect 62852 80838 62971 82020
rect 64095 80838 64217 82020
rect 62852 80735 64217 80838
rect 69810 82021 71175 82131
rect 69810 80839 69929 82021
rect 71053 80839 71175 82021
rect 69810 80736 71175 80839
rect 76727 82019 78092 82129
rect 76727 80837 76846 82019
rect 77970 80837 78092 82019
rect 76727 80734 78092 80837
rect 83692 82020 85057 82130
rect 83692 80838 83811 82020
rect 84935 80838 85057 82020
rect 83692 80735 85057 80838
rect 90650 82021 92015 82131
rect 90650 80839 90769 82021
rect 91893 80839 92015 82021
rect 90650 80736 92015 80839
rect 97468 82000 98833 82110
rect 97468 80818 97587 82000
rect 98711 80818 98833 82000
rect 97468 80715 98833 80818
rect 104433 82001 105798 82111
rect 104433 80819 104552 82001
rect 105676 80819 105798 82001
rect 104433 80716 105798 80819
rect 111391 82002 112756 82112
rect 111391 80820 111510 82002
rect 112634 80820 112756 82002
rect 111391 80717 112756 80820
rect 118311 82001 119676 82111
rect 118311 80819 118430 82001
rect 119554 80819 119676 82001
rect 118311 80716 119676 80819
rect 125276 82002 126641 82112
rect 125276 80820 125395 82002
rect 126519 80820 126641 82002
rect 125276 80717 126641 80820
rect 132234 82003 133599 82113
rect 132234 80821 132353 82003
rect 133477 80821 133599 82003
rect 132234 80718 133599 80821
rect 139151 82007 140516 82117
rect 139151 80825 139270 82007
rect 140394 80825 140516 82007
rect 139151 80722 140516 80825
rect 146116 82008 147481 82118
rect 146116 80826 146235 82008
rect 147359 80826 147481 82008
rect 146116 80723 147481 80826
rect 153074 82009 154439 82119
rect 153074 80827 153193 82009
rect 154317 80827 154439 82009
rect 153074 80724 154439 80827
rect 159991 82007 161356 82117
rect 159991 80825 160110 82007
rect 161234 80825 161356 82007
rect 159991 80722 161356 80825
rect 166956 82008 168321 82118
rect 166956 80826 167075 82008
rect 168199 80826 168321 82008
rect 166956 80723 168321 80826
rect 173914 82009 175279 82119
rect 173914 80827 174033 82009
rect 175157 80827 175279 82009
rect 173914 80724 175279 80827
rect 180719 82002 182084 82112
rect 180719 80820 180838 82002
rect 181962 80820 182084 82002
rect 180719 80717 182084 80820
rect 187684 82003 189049 82113
rect 187684 80821 187803 82003
rect 188927 80821 189049 82003
rect 187684 80718 189049 80821
rect 194642 82004 196007 82114
rect 194642 80822 194761 82004
rect 195885 80822 196007 82004
rect 194642 80719 196007 80822
rect 201562 82003 202927 82113
rect 201562 80821 201681 82003
rect 202805 80821 202927 82003
rect 201562 80718 202927 80821
rect 208527 82004 209892 82114
rect 208527 80822 208646 82004
rect 209770 80822 209892 82004
rect 208527 80719 209892 80822
rect 215485 82005 216850 82115
rect 215485 80823 215604 82005
rect 216728 80823 216850 82005
rect 215485 80720 216850 80823
rect 222402 82009 223767 82119
rect 222402 80827 222521 82009
rect 223645 80827 223767 82009
rect 222402 80724 223767 80827
rect 229367 82010 230732 82120
rect 229367 80828 229486 82010
rect 230610 80828 230732 82010
rect 229367 80725 230732 80828
rect 236325 82011 237690 82121
rect 236325 80829 236444 82011
rect 237568 80829 237690 82011
rect 236325 80726 237690 80829
rect 243242 82009 244607 82119
rect 243242 80827 243361 82009
rect 244485 80827 244607 82009
rect 243242 80724 244607 80827
rect 250207 82010 251572 82120
rect 250207 80828 250326 82010
rect 251450 80828 251572 82010
rect 250207 80725 251572 80828
rect 257165 82011 258530 82121
rect 257165 80829 257284 82011
rect 258408 80829 258530 82011
rect 257165 80726 258530 80829
rect 264305 82011 265670 82121
rect 264305 80829 264424 82011
rect 265548 80829 265670 82011
rect 264305 80726 265670 80829
rect 271263 82012 272628 82122
rect 271263 80830 271382 82012
rect 272506 80830 272628 82012
rect 271263 80727 272628 80830
rect 278399 82002 279764 82112
rect 278399 80820 278518 82002
rect 279642 80820 279764 82002
rect 278399 80717 279764 80820
rect 21035 70833 22400 70943
rect 21035 69651 21154 70833
rect 22278 69651 22400 70833
rect 21035 69548 22400 69651
rect 27993 70834 29358 70944
rect 27993 69652 28112 70834
rect 29236 69652 29358 70834
rect 27993 69549 29358 69652
rect 34913 70833 36278 70943
rect 34913 69651 35032 70833
rect 36156 69651 36278 70833
rect 34913 69548 36278 69651
rect 41878 70834 43243 70944
rect 41878 69652 41997 70834
rect 43121 69652 43243 70834
rect 41878 69549 43243 69652
rect 48836 70835 50201 70945
rect 48836 69653 48955 70835
rect 50079 69653 50201 70835
rect 48836 69550 50201 69653
rect 55753 70839 57118 70949
rect 55753 69657 55872 70839
rect 56996 69657 57118 70839
rect 55753 69554 57118 69657
rect 62718 70840 64083 70950
rect 62718 69658 62837 70840
rect 63961 69658 64083 70840
rect 62718 69555 64083 69658
rect 69676 70841 71041 70951
rect 69676 69659 69795 70841
rect 70919 69659 71041 70841
rect 69676 69556 71041 69659
rect 76593 70839 77958 70949
rect 76593 69657 76712 70839
rect 77836 69657 77958 70839
rect 76593 69554 77958 69657
rect 83558 70840 84923 70950
rect 83558 69658 83677 70840
rect 84801 69658 84923 70840
rect 83558 69555 84923 69658
rect 90516 70841 91881 70951
rect 90516 69659 90635 70841
rect 91759 69659 91881 70841
rect 90516 69556 91881 69659
rect 97334 70820 98699 70930
rect 97334 69638 97453 70820
rect 98577 69638 98699 70820
rect 97334 69535 98699 69638
rect 104299 70821 105664 70931
rect 104299 69639 104418 70821
rect 105542 69639 105664 70821
rect 104299 69536 105664 69639
rect 111257 70822 112622 70932
rect 111257 69640 111376 70822
rect 112500 69640 112622 70822
rect 111257 69537 112622 69640
rect 118177 70821 119542 70931
rect 118177 69639 118296 70821
rect 119420 69639 119542 70821
rect 118177 69536 119542 69639
rect 125142 70822 126507 70932
rect 125142 69640 125261 70822
rect 126385 69640 126507 70822
rect 125142 69537 126507 69640
rect 132100 70823 133465 70933
rect 132100 69641 132219 70823
rect 133343 69641 133465 70823
rect 132100 69538 133465 69641
rect 139017 70827 140382 70937
rect 139017 69645 139136 70827
rect 140260 69645 140382 70827
rect 139017 69542 140382 69645
rect 145982 70828 147347 70938
rect 145982 69646 146101 70828
rect 147225 69646 147347 70828
rect 145982 69543 147347 69646
rect 152940 70829 154305 70939
rect 152940 69647 153059 70829
rect 154183 69647 154305 70829
rect 152940 69544 154305 69647
rect 159857 70827 161222 70937
rect 159857 69645 159976 70827
rect 161100 69645 161222 70827
rect 159857 69542 161222 69645
rect 166822 70828 168187 70938
rect 166822 69646 166941 70828
rect 168065 69646 168187 70828
rect 166822 69543 168187 69646
rect 173780 70829 175145 70939
rect 173780 69647 173899 70829
rect 175023 69647 175145 70829
rect 173780 69544 175145 69647
rect 180585 70822 181950 70932
rect 180585 69640 180704 70822
rect 181828 69640 181950 70822
rect 180585 69537 181950 69640
rect 187550 70823 188915 70933
rect 187550 69641 187669 70823
rect 188793 69641 188915 70823
rect 187550 69538 188915 69641
rect 194508 70824 195873 70934
rect 194508 69642 194627 70824
rect 195751 69642 195873 70824
rect 194508 69539 195873 69642
rect 201428 70823 202793 70933
rect 201428 69641 201547 70823
rect 202671 69641 202793 70823
rect 201428 69538 202793 69641
rect 208393 70824 209758 70934
rect 208393 69642 208512 70824
rect 209636 69642 209758 70824
rect 208393 69539 209758 69642
rect 215351 70825 216716 70935
rect 215351 69643 215470 70825
rect 216594 69643 216716 70825
rect 215351 69540 216716 69643
rect 222268 70829 223633 70939
rect 222268 69647 222387 70829
rect 223511 69647 223633 70829
rect 222268 69544 223633 69647
rect 229233 70830 230598 70940
rect 229233 69648 229352 70830
rect 230476 69648 230598 70830
rect 229233 69545 230598 69648
rect 236191 70831 237556 70941
rect 236191 69649 236310 70831
rect 237434 69649 237556 70831
rect 236191 69546 237556 69649
rect 243108 70829 244473 70939
rect 243108 69647 243227 70829
rect 244351 69647 244473 70829
rect 243108 69544 244473 69647
rect 250073 70830 251438 70940
rect 250073 69648 250192 70830
rect 251316 69648 251438 70830
rect 250073 69545 251438 69648
rect 257031 70831 258396 70941
rect 257031 69649 257150 70831
rect 258274 69649 258396 70831
rect 257031 69546 258396 69649
rect 264171 70831 265536 70941
rect 264171 69649 264290 70831
rect 265414 69649 265536 70831
rect 264171 69546 265536 69649
rect 271129 70832 272494 70942
rect 271129 69650 271248 70832
rect 272372 69650 272494 70832
rect 271129 69547 272494 69650
rect 278265 70822 279630 70932
rect 278265 69640 278384 70822
rect 279508 69640 279630 70822
rect 278265 69537 279630 69640
rect 21000 64593 22365 64703
rect 21000 63411 21119 64593
rect 22243 63411 22365 64593
rect 21000 63308 22365 63411
rect 27958 64594 29323 64704
rect 27958 63412 28077 64594
rect 29201 63412 29323 64594
rect 27958 63309 29323 63412
rect 34878 64593 36243 64703
rect 34878 63411 34997 64593
rect 36121 63411 36243 64593
rect 34878 63308 36243 63411
rect 41843 64594 43208 64704
rect 41843 63412 41962 64594
rect 43086 63412 43208 64594
rect 41843 63309 43208 63412
rect 48801 64595 50166 64705
rect 48801 63413 48920 64595
rect 50044 63413 50166 64595
rect 48801 63310 50166 63413
rect 55718 64599 57083 64709
rect 55718 63417 55837 64599
rect 56961 63417 57083 64599
rect 55718 63314 57083 63417
rect 62683 64600 64048 64710
rect 62683 63418 62802 64600
rect 63926 63418 64048 64600
rect 62683 63315 64048 63418
rect 69641 64601 71006 64711
rect 69641 63419 69760 64601
rect 70884 63419 71006 64601
rect 69641 63316 71006 63419
rect 76558 64599 77923 64709
rect 76558 63417 76677 64599
rect 77801 63417 77923 64599
rect 76558 63314 77923 63417
rect 83523 64600 84888 64710
rect 83523 63418 83642 64600
rect 84766 63418 84888 64600
rect 83523 63315 84888 63418
rect 90481 64601 91846 64711
rect 90481 63419 90600 64601
rect 91724 63419 91846 64601
rect 90481 63316 91846 63419
rect 97299 64580 98664 64690
rect 97299 63398 97418 64580
rect 98542 63398 98664 64580
rect 97299 63295 98664 63398
rect 104264 64581 105629 64691
rect 104264 63399 104383 64581
rect 105507 63399 105629 64581
rect 104264 63296 105629 63399
rect 111222 64582 112587 64692
rect 111222 63400 111341 64582
rect 112465 63400 112587 64582
rect 111222 63297 112587 63400
rect 118142 64581 119507 64691
rect 118142 63399 118261 64581
rect 119385 63399 119507 64581
rect 118142 63296 119507 63399
rect 125107 64582 126472 64692
rect 125107 63400 125226 64582
rect 126350 63400 126472 64582
rect 125107 63297 126472 63400
rect 132065 64583 133430 64693
rect 132065 63401 132184 64583
rect 133308 63401 133430 64583
rect 132065 63298 133430 63401
rect 138982 64587 140347 64697
rect 138982 63405 139101 64587
rect 140225 63405 140347 64587
rect 138982 63302 140347 63405
rect 145947 64588 147312 64698
rect 145947 63406 146066 64588
rect 147190 63406 147312 64588
rect 145947 63303 147312 63406
rect 152905 64589 154270 64699
rect 152905 63407 153024 64589
rect 154148 63407 154270 64589
rect 152905 63304 154270 63407
rect 159822 64587 161187 64697
rect 159822 63405 159941 64587
rect 161065 63405 161187 64587
rect 159822 63302 161187 63405
rect 166787 64588 168152 64698
rect 166787 63406 166906 64588
rect 168030 63406 168152 64588
rect 166787 63303 168152 63406
rect 173745 64589 175110 64699
rect 173745 63407 173864 64589
rect 174988 63407 175110 64589
rect 173745 63304 175110 63407
rect 180550 64582 181915 64692
rect 180550 63400 180669 64582
rect 181793 63400 181915 64582
rect 180550 63297 181915 63400
rect 187515 64583 188880 64693
rect 187515 63401 187634 64583
rect 188758 63401 188880 64583
rect 187515 63298 188880 63401
rect 194473 64584 195838 64694
rect 194473 63402 194592 64584
rect 195716 63402 195838 64584
rect 194473 63299 195838 63402
rect 201393 64583 202758 64693
rect 201393 63401 201512 64583
rect 202636 63401 202758 64583
rect 201393 63298 202758 63401
rect 208358 64584 209723 64694
rect 208358 63402 208477 64584
rect 209601 63402 209723 64584
rect 208358 63299 209723 63402
rect 215316 64585 216681 64695
rect 215316 63403 215435 64585
rect 216559 63403 216681 64585
rect 215316 63300 216681 63403
rect 222233 64589 223598 64699
rect 222233 63407 222352 64589
rect 223476 63407 223598 64589
rect 222233 63304 223598 63407
rect 229198 64590 230563 64700
rect 229198 63408 229317 64590
rect 230441 63408 230563 64590
rect 229198 63305 230563 63408
rect 236156 64591 237521 64701
rect 236156 63409 236275 64591
rect 237399 63409 237521 64591
rect 236156 63306 237521 63409
rect 243073 64589 244438 64699
rect 243073 63407 243192 64589
rect 244316 63407 244438 64589
rect 243073 63304 244438 63407
rect 250038 64590 251403 64700
rect 250038 63408 250157 64590
rect 251281 63408 251403 64590
rect 250038 63305 251403 63408
rect 256996 64591 258361 64701
rect 256996 63409 257115 64591
rect 258239 63409 258361 64591
rect 256996 63306 258361 63409
rect 264136 64591 265501 64701
rect 264136 63409 264255 64591
rect 265379 63409 265501 64591
rect 264136 63306 265501 63409
rect 271094 64592 272459 64702
rect 271094 63410 271213 64592
rect 272337 63410 272459 64592
rect 271094 63307 272459 63410
rect 278230 64582 279595 64692
rect 278230 63400 278349 64582
rect 279473 63400 279595 64582
rect 278230 63297 279595 63400
rect 20965 58876 22330 58986
rect 20965 57694 21084 58876
rect 22208 57694 22330 58876
rect 20965 57591 22330 57694
rect 27923 58877 29288 58987
rect 27923 57695 28042 58877
rect 29166 57695 29288 58877
rect 27923 57592 29288 57695
rect 34843 58876 36208 58986
rect 34843 57694 34962 58876
rect 36086 57694 36208 58876
rect 34843 57591 36208 57694
rect 41808 58877 43173 58987
rect 41808 57695 41927 58877
rect 43051 57695 43173 58877
rect 41808 57592 43173 57695
rect 48766 58878 50131 58988
rect 48766 57696 48885 58878
rect 50009 57696 50131 58878
rect 48766 57593 50131 57696
rect 55683 58882 57048 58992
rect 55683 57700 55802 58882
rect 56926 57700 57048 58882
rect 55683 57597 57048 57700
rect 62648 58883 64013 58993
rect 62648 57701 62767 58883
rect 63891 57701 64013 58883
rect 62648 57598 64013 57701
rect 69606 58884 70971 58994
rect 69606 57702 69725 58884
rect 70849 57702 70971 58884
rect 69606 57599 70971 57702
rect 76523 58882 77888 58992
rect 76523 57700 76642 58882
rect 77766 57700 77888 58882
rect 76523 57597 77888 57700
rect 83488 58883 84853 58993
rect 83488 57701 83607 58883
rect 84731 57701 84853 58883
rect 83488 57598 84853 57701
rect 90446 58884 91811 58994
rect 90446 57702 90565 58884
rect 91689 57702 91811 58884
rect 90446 57599 91811 57702
rect 97264 58863 98629 58973
rect 97264 57681 97383 58863
rect 98507 57681 98629 58863
rect 97264 57578 98629 57681
rect 104229 58864 105594 58974
rect 104229 57682 104348 58864
rect 105472 57682 105594 58864
rect 104229 57579 105594 57682
rect 111187 58865 112552 58975
rect 111187 57683 111306 58865
rect 112430 57683 112552 58865
rect 111187 57580 112552 57683
rect 118107 58864 119472 58974
rect 118107 57682 118226 58864
rect 119350 57682 119472 58864
rect 118107 57579 119472 57682
rect 125072 58865 126437 58975
rect 125072 57683 125191 58865
rect 126315 57683 126437 58865
rect 125072 57580 126437 57683
rect 132030 58866 133395 58976
rect 132030 57684 132149 58866
rect 133273 57684 133395 58866
rect 132030 57581 133395 57684
rect 138947 58870 140312 58980
rect 138947 57688 139066 58870
rect 140190 57688 140312 58870
rect 138947 57585 140312 57688
rect 145912 58871 147277 58981
rect 145912 57689 146031 58871
rect 147155 57689 147277 58871
rect 145912 57586 147277 57689
rect 152870 58872 154235 58982
rect 152870 57690 152989 58872
rect 154113 57690 154235 58872
rect 152870 57587 154235 57690
rect 159787 58870 161152 58980
rect 159787 57688 159906 58870
rect 161030 57688 161152 58870
rect 159787 57585 161152 57688
rect 166752 58871 168117 58981
rect 166752 57689 166871 58871
rect 167995 57689 168117 58871
rect 166752 57586 168117 57689
rect 173710 58872 175075 58982
rect 173710 57690 173829 58872
rect 174953 57690 175075 58872
rect 173710 57587 175075 57690
rect 180515 58865 181880 58975
rect 180515 57683 180634 58865
rect 181758 57683 181880 58865
rect 180515 57580 181880 57683
rect 187480 58866 188845 58976
rect 187480 57684 187599 58866
rect 188723 57684 188845 58866
rect 187480 57581 188845 57684
rect 194438 58867 195803 58977
rect 194438 57685 194557 58867
rect 195681 57685 195803 58867
rect 194438 57582 195803 57685
rect 201358 58866 202723 58976
rect 201358 57684 201477 58866
rect 202601 57684 202723 58866
rect 201358 57581 202723 57684
rect 208323 58867 209688 58977
rect 208323 57685 208442 58867
rect 209566 57685 209688 58867
rect 208323 57582 209688 57685
rect 215281 58868 216646 58978
rect 215281 57686 215400 58868
rect 216524 57686 216646 58868
rect 215281 57583 216646 57686
rect 222198 58872 223563 58982
rect 222198 57690 222317 58872
rect 223441 57690 223563 58872
rect 222198 57587 223563 57690
rect 229163 58873 230528 58983
rect 229163 57691 229282 58873
rect 230406 57691 230528 58873
rect 229163 57588 230528 57691
rect 236121 58874 237486 58984
rect 236121 57692 236240 58874
rect 237364 57692 237486 58874
rect 236121 57589 237486 57692
rect 243038 58872 244403 58982
rect 243038 57690 243157 58872
rect 244281 57690 244403 58872
rect 243038 57587 244403 57690
rect 250003 58873 251368 58983
rect 250003 57691 250122 58873
rect 251246 57691 251368 58873
rect 250003 57588 251368 57691
rect 256961 58874 258326 58984
rect 256961 57692 257080 58874
rect 258204 57692 258326 58874
rect 256961 57589 258326 57692
rect 264101 58874 265466 58984
rect 264101 57692 264220 58874
rect 265344 57692 265466 58874
rect 264101 57589 265466 57692
rect 271059 58875 272424 58985
rect 271059 57693 271178 58875
rect 272302 57693 272424 58875
rect 271059 57590 272424 57693
rect 278195 58865 279560 58975
rect 278195 57683 278314 58865
rect 279438 57683 279560 58865
rect 278195 57580 279560 57683
rect 20896 52671 22261 52781
rect 20896 51489 21015 52671
rect 22139 51489 22261 52671
rect 20896 51386 22261 51489
rect 27854 52672 29219 52782
rect 27854 51490 27973 52672
rect 29097 51490 29219 52672
rect 27854 51387 29219 51490
rect 34774 52671 36139 52781
rect 34774 51489 34893 52671
rect 36017 51489 36139 52671
rect 34774 51386 36139 51489
rect 41739 52672 43104 52782
rect 41739 51490 41858 52672
rect 42982 51490 43104 52672
rect 41739 51387 43104 51490
rect 48697 52673 50062 52783
rect 48697 51491 48816 52673
rect 49940 51491 50062 52673
rect 48697 51388 50062 51491
rect 55614 52677 56979 52787
rect 55614 51495 55733 52677
rect 56857 51495 56979 52677
rect 55614 51392 56979 51495
rect 62579 52678 63944 52788
rect 62579 51496 62698 52678
rect 63822 51496 63944 52678
rect 62579 51393 63944 51496
rect 69537 52679 70902 52789
rect 69537 51497 69656 52679
rect 70780 51497 70902 52679
rect 69537 51394 70902 51497
rect 76454 52677 77819 52787
rect 76454 51495 76573 52677
rect 77697 51495 77819 52677
rect 76454 51392 77819 51495
rect 83419 52678 84784 52788
rect 83419 51496 83538 52678
rect 84662 51496 84784 52678
rect 83419 51393 84784 51496
rect 90377 52679 91742 52789
rect 90377 51497 90496 52679
rect 91620 51497 91742 52679
rect 90377 51394 91742 51497
rect 97195 52658 98560 52768
rect 97195 51476 97314 52658
rect 98438 51476 98560 52658
rect 97195 51373 98560 51476
rect 104160 52659 105525 52769
rect 104160 51477 104279 52659
rect 105403 51477 105525 52659
rect 104160 51374 105525 51477
rect 111118 52660 112483 52770
rect 111118 51478 111237 52660
rect 112361 51478 112483 52660
rect 111118 51375 112483 51478
rect 118038 52659 119403 52769
rect 118038 51477 118157 52659
rect 119281 51477 119403 52659
rect 118038 51374 119403 51477
rect 125003 52660 126368 52770
rect 125003 51478 125122 52660
rect 126246 51478 126368 52660
rect 125003 51375 126368 51478
rect 131961 52661 133326 52771
rect 131961 51479 132080 52661
rect 133204 51479 133326 52661
rect 131961 51376 133326 51479
rect 138878 52665 140243 52775
rect 138878 51483 138997 52665
rect 140121 51483 140243 52665
rect 138878 51380 140243 51483
rect 145843 52666 147208 52776
rect 145843 51484 145962 52666
rect 147086 51484 147208 52666
rect 145843 51381 147208 51484
rect 152801 52667 154166 52777
rect 152801 51485 152920 52667
rect 154044 51485 154166 52667
rect 152801 51382 154166 51485
rect 159718 52665 161083 52775
rect 159718 51483 159837 52665
rect 160961 51483 161083 52665
rect 159718 51380 161083 51483
rect 166683 52666 168048 52776
rect 166683 51484 166802 52666
rect 167926 51484 168048 52666
rect 166683 51381 168048 51484
rect 173641 52667 175006 52777
rect 173641 51485 173760 52667
rect 174884 51485 175006 52667
rect 173641 51382 175006 51485
rect 180446 52660 181811 52770
rect 180446 51478 180565 52660
rect 181689 51478 181811 52660
rect 180446 51375 181811 51478
rect 187411 52661 188776 52771
rect 187411 51479 187530 52661
rect 188654 51479 188776 52661
rect 187411 51376 188776 51479
rect 194369 52662 195734 52772
rect 194369 51480 194488 52662
rect 195612 51480 195734 52662
rect 194369 51377 195734 51480
rect 201289 52661 202654 52771
rect 201289 51479 201408 52661
rect 202532 51479 202654 52661
rect 201289 51376 202654 51479
rect 208254 52662 209619 52772
rect 208254 51480 208373 52662
rect 209497 51480 209619 52662
rect 208254 51377 209619 51480
rect 215212 52663 216577 52773
rect 215212 51481 215331 52663
rect 216455 51481 216577 52663
rect 215212 51378 216577 51481
rect 222129 52667 223494 52777
rect 222129 51485 222248 52667
rect 223372 51485 223494 52667
rect 222129 51382 223494 51485
rect 229094 52668 230459 52778
rect 229094 51486 229213 52668
rect 230337 51486 230459 52668
rect 229094 51383 230459 51486
rect 236052 52669 237417 52779
rect 236052 51487 236171 52669
rect 237295 51487 237417 52669
rect 236052 51384 237417 51487
rect 242969 52667 244334 52777
rect 242969 51485 243088 52667
rect 244212 51485 244334 52667
rect 242969 51382 244334 51485
rect 249934 52668 251299 52778
rect 249934 51486 250053 52668
rect 251177 51486 251299 52668
rect 249934 51383 251299 51486
rect 256892 52669 258257 52779
rect 256892 51487 257011 52669
rect 258135 51487 258257 52669
rect 256892 51384 258257 51487
rect 264032 52669 265397 52779
rect 264032 51487 264151 52669
rect 265275 51487 265397 52669
rect 264032 51384 265397 51487
rect 270990 52670 272355 52780
rect 270990 51488 271109 52670
rect 272233 51488 272355 52670
rect 270990 51385 272355 51488
rect 278126 52660 279491 52770
rect 278126 51478 278245 52660
rect 279369 51478 279491 52660
rect 278126 51375 279491 51478
rect 69249 44821 70614 44931
rect 69249 43639 69368 44821
rect 70492 43639 70614 44821
rect 69249 43536 70614 43639
rect 76166 44819 77531 44929
rect 76166 43637 76285 44819
rect 77409 43637 77531 44819
rect 76166 43534 77531 43637
rect 83131 44820 84496 44930
rect 83131 43638 83250 44820
rect 84374 43638 84496 44820
rect 83131 43535 84496 43638
rect 90089 44821 91454 44931
rect 90089 43639 90208 44821
rect 91332 43639 91454 44821
rect 90089 43536 91454 43639
rect 96907 44800 98272 44910
rect 96907 43618 97026 44800
rect 98150 43618 98272 44800
rect 96907 43515 98272 43618
rect 103872 44801 105237 44911
rect 103872 43619 103991 44801
rect 105115 43619 105237 44801
rect 103872 43516 105237 43619
rect 110830 44802 112195 44912
rect 110830 43620 110949 44802
rect 112073 43620 112195 44802
rect 110830 43517 112195 43620
rect 117750 44801 119115 44911
rect 117750 43619 117869 44801
rect 118993 43619 119115 44801
rect 117750 43516 119115 43619
rect 124715 44802 126080 44912
rect 124715 43620 124834 44802
rect 125958 43620 126080 44802
rect 124715 43517 126080 43620
rect 131673 44803 133038 44913
rect 131673 43621 131792 44803
rect 132916 43621 133038 44803
rect 131673 43518 133038 43621
rect 138590 44807 139955 44917
rect 138590 43625 138709 44807
rect 139833 43625 139955 44807
rect 138590 43522 139955 43625
rect 145555 44808 146920 44918
rect 145555 43626 145674 44808
rect 146798 43626 146920 44808
rect 145555 43523 146920 43626
rect 152513 44809 153878 44919
rect 152513 43627 152632 44809
rect 153756 43627 153878 44809
rect 152513 43524 153878 43627
rect 159430 44807 160795 44917
rect 159430 43625 159549 44807
rect 160673 43625 160795 44807
rect 159430 43522 160795 43625
rect 166395 44808 167760 44918
rect 166395 43626 166514 44808
rect 167638 43626 167760 44808
rect 166395 43523 167760 43626
rect 173353 44809 174718 44919
rect 173353 43627 173472 44809
rect 174596 43627 174718 44809
rect 173353 43524 174718 43627
rect 180158 44802 181523 44912
rect 180158 43620 180277 44802
rect 181401 43620 181523 44802
rect 180158 43517 181523 43620
rect 187123 44803 188488 44913
rect 187123 43621 187242 44803
rect 188366 43621 188488 44803
rect 187123 43518 188488 43621
rect 194081 44804 195446 44914
rect 194081 43622 194200 44804
rect 195324 43622 195446 44804
rect 194081 43519 195446 43622
rect 201001 44803 202366 44913
rect 201001 43621 201120 44803
rect 202244 43621 202366 44803
rect 201001 43518 202366 43621
rect 207966 44804 209331 44914
rect 207966 43622 208085 44804
rect 209209 43622 209331 44804
rect 207966 43519 209331 43622
rect 214924 44805 216289 44915
rect 214924 43623 215043 44805
rect 216167 43623 216289 44805
rect 214924 43520 216289 43623
rect 221841 44809 223206 44919
rect 221841 43627 221960 44809
rect 223084 43627 223206 44809
rect 221841 43524 223206 43627
rect 228806 44810 230171 44920
rect 228806 43628 228925 44810
rect 230049 43628 230171 44810
rect 228806 43525 230171 43628
rect 235764 44811 237129 44921
rect 235764 43629 235883 44811
rect 237007 43629 237129 44811
rect 235764 43526 237129 43629
rect 242681 44809 244046 44919
rect 242681 43627 242800 44809
rect 243924 43627 244046 44809
rect 242681 43524 244046 43627
rect 249646 44810 251011 44920
rect 249646 43628 249765 44810
rect 250889 43628 251011 44810
rect 249646 43525 251011 43628
rect 256604 44811 257969 44921
rect 256604 43629 256723 44811
rect 257847 43629 257969 44811
rect 256604 43526 257969 43629
rect 263744 44811 265109 44921
rect 263744 43629 263863 44811
rect 264987 43629 265109 44811
rect 263744 43526 265109 43629
rect 270702 44812 272067 44922
rect 270702 43630 270821 44812
rect 271945 43630 272067 44812
rect 270702 43527 272067 43630
rect 277838 44802 279203 44912
rect 277838 43620 277957 44802
rect 279081 43620 279203 44802
rect 277838 43517 279203 43620
rect 69249 38527 70614 38637
rect 69249 37345 69368 38527
rect 70492 37345 70614 38527
rect 69249 37242 70614 37345
rect 76166 38525 77531 38635
rect 76166 37343 76285 38525
rect 77409 37343 77531 38525
rect 76166 37240 77531 37343
rect 83131 38526 84496 38636
rect 83131 37344 83250 38526
rect 84374 37344 84496 38526
rect 83131 37241 84496 37344
rect 90089 38527 91454 38637
rect 90089 37345 90208 38527
rect 91332 37345 91454 38527
rect 90089 37242 91454 37345
rect 96907 38506 98272 38616
rect 96907 37324 97026 38506
rect 98150 37324 98272 38506
rect 96907 37221 98272 37324
rect 103872 38507 105237 38617
rect 103872 37325 103991 38507
rect 105115 37325 105237 38507
rect 103872 37222 105237 37325
rect 110830 38508 112195 38618
rect 110830 37326 110949 38508
rect 112073 37326 112195 38508
rect 110830 37223 112195 37326
rect 117750 38507 119115 38617
rect 117750 37325 117869 38507
rect 118993 37325 119115 38507
rect 117750 37222 119115 37325
rect 124715 38508 126080 38618
rect 124715 37326 124834 38508
rect 125958 37326 126080 38508
rect 124715 37223 126080 37326
rect 131673 38509 133038 38619
rect 131673 37327 131792 38509
rect 132916 37327 133038 38509
rect 131673 37224 133038 37327
rect 138590 38513 139955 38623
rect 138590 37331 138709 38513
rect 139833 37331 139955 38513
rect 138590 37228 139955 37331
rect 145555 38514 146920 38624
rect 145555 37332 145674 38514
rect 146798 37332 146920 38514
rect 145555 37229 146920 37332
rect 152513 38515 153878 38625
rect 152513 37333 152632 38515
rect 153756 37333 153878 38515
rect 152513 37230 153878 37333
rect 159430 38513 160795 38623
rect 159430 37331 159549 38513
rect 160673 37331 160795 38513
rect 159430 37228 160795 37331
rect 166395 38514 167760 38624
rect 166395 37332 166514 38514
rect 167638 37332 167760 38514
rect 166395 37229 167760 37332
rect 173353 38515 174718 38625
rect 173353 37333 173472 38515
rect 174596 37333 174718 38515
rect 173353 37230 174718 37333
rect 180158 38508 181523 38618
rect 180158 37326 180277 38508
rect 181401 37326 181523 38508
rect 180158 37223 181523 37326
rect 187123 38509 188488 38619
rect 187123 37327 187242 38509
rect 188366 37327 188488 38509
rect 187123 37224 188488 37327
rect 194081 38510 195446 38620
rect 194081 37328 194200 38510
rect 195324 37328 195446 38510
rect 194081 37225 195446 37328
rect 201001 38509 202366 38619
rect 201001 37327 201120 38509
rect 202244 37327 202366 38509
rect 201001 37224 202366 37327
rect 207966 38510 209331 38620
rect 207966 37328 208085 38510
rect 209209 37328 209331 38510
rect 207966 37225 209331 37328
rect 214924 38511 216289 38621
rect 214924 37329 215043 38511
rect 216167 37329 216289 38511
rect 214924 37226 216289 37329
rect 221841 38515 223206 38625
rect 221841 37333 221960 38515
rect 223084 37333 223206 38515
rect 221841 37230 223206 37333
rect 228806 38516 230171 38626
rect 228806 37334 228925 38516
rect 230049 37334 230171 38516
rect 228806 37231 230171 37334
rect 235764 38517 237129 38627
rect 235764 37335 235883 38517
rect 237007 37335 237129 38517
rect 235764 37232 237129 37335
rect 242681 38515 244046 38625
rect 242681 37333 242800 38515
rect 243924 37333 244046 38515
rect 242681 37230 244046 37333
rect 249646 38516 251011 38626
rect 249646 37334 249765 38516
rect 250889 37334 251011 38516
rect 249646 37231 251011 37334
rect 256604 38517 257969 38627
rect 256604 37335 256723 38517
rect 257847 37335 257969 38517
rect 256604 37232 257969 37335
rect 263744 38517 265109 38627
rect 263744 37335 263863 38517
rect 264987 37335 265109 38517
rect 263744 37232 265109 37335
rect 270702 38518 272067 38628
rect 270702 37336 270821 38518
rect 271945 37336 272067 38518
rect 270702 37233 272067 37336
rect 277838 38508 279203 38618
rect 277838 37326 277957 38508
rect 279081 37326 279203 38508
rect 277838 37223 279203 37326
rect 69249 32233 70614 32343
rect 69249 31051 69368 32233
rect 70492 31051 70614 32233
rect 69249 30948 70614 31051
rect 76166 32231 77531 32341
rect 76166 31049 76285 32231
rect 77409 31049 77531 32231
rect 76166 30946 77531 31049
rect 83131 32232 84496 32342
rect 83131 31050 83250 32232
rect 84374 31050 84496 32232
rect 83131 30947 84496 31050
rect 90089 32233 91454 32343
rect 90089 31051 90208 32233
rect 91332 31051 91454 32233
rect 90089 30948 91454 31051
rect 96907 32212 98272 32322
rect 96907 31030 97026 32212
rect 98150 31030 98272 32212
rect 96907 30927 98272 31030
rect 103872 32213 105237 32323
rect 103872 31031 103991 32213
rect 105115 31031 105237 32213
rect 103872 30928 105237 31031
rect 110830 32214 112195 32324
rect 110830 31032 110949 32214
rect 112073 31032 112195 32214
rect 110830 30929 112195 31032
rect 117750 32213 119115 32323
rect 117750 31031 117869 32213
rect 118993 31031 119115 32213
rect 117750 30928 119115 31031
rect 124715 32214 126080 32324
rect 124715 31032 124834 32214
rect 125958 31032 126080 32214
rect 124715 30929 126080 31032
rect 131673 32215 133038 32325
rect 131673 31033 131792 32215
rect 132916 31033 133038 32215
rect 131673 30930 133038 31033
rect 138590 32219 139955 32329
rect 138590 31037 138709 32219
rect 139833 31037 139955 32219
rect 138590 30934 139955 31037
rect 145555 32220 146920 32330
rect 145555 31038 145674 32220
rect 146798 31038 146920 32220
rect 145555 30935 146920 31038
rect 152513 32221 153878 32331
rect 152513 31039 152632 32221
rect 153756 31039 153878 32221
rect 152513 30936 153878 31039
rect 159430 32219 160795 32329
rect 159430 31037 159549 32219
rect 160673 31037 160795 32219
rect 159430 30934 160795 31037
rect 166395 32220 167760 32330
rect 166395 31038 166514 32220
rect 167638 31038 167760 32220
rect 166395 30935 167760 31038
rect 173353 32221 174718 32331
rect 173353 31039 173472 32221
rect 174596 31039 174718 32221
rect 173353 30936 174718 31039
rect 180158 32214 181523 32324
rect 180158 31032 180277 32214
rect 181401 31032 181523 32214
rect 180158 30929 181523 31032
rect 187123 32215 188488 32325
rect 187123 31033 187242 32215
rect 188366 31033 188488 32215
rect 187123 30930 188488 31033
rect 194081 32216 195446 32326
rect 194081 31034 194200 32216
rect 195324 31034 195446 32216
rect 194081 30931 195446 31034
rect 201001 32215 202366 32325
rect 201001 31033 201120 32215
rect 202244 31033 202366 32215
rect 201001 30930 202366 31033
rect 207966 32216 209331 32326
rect 207966 31034 208085 32216
rect 209209 31034 209331 32216
rect 207966 30931 209331 31034
rect 214924 32217 216289 32327
rect 214924 31035 215043 32217
rect 216167 31035 216289 32217
rect 214924 30932 216289 31035
rect 221841 32221 223206 32331
rect 221841 31039 221960 32221
rect 223084 31039 223206 32221
rect 221841 30936 223206 31039
rect 228806 32222 230171 32332
rect 228806 31040 228925 32222
rect 230049 31040 230171 32222
rect 228806 30937 230171 31040
rect 235764 32223 237129 32333
rect 235764 31041 235883 32223
rect 237007 31041 237129 32223
rect 235764 30938 237129 31041
rect 242681 32221 244046 32331
rect 242681 31039 242800 32221
rect 243924 31039 244046 32221
rect 242681 30936 244046 31039
rect 249646 32222 251011 32332
rect 249646 31040 249765 32222
rect 250889 31040 251011 32222
rect 249646 30937 251011 31040
rect 256604 32223 257969 32333
rect 256604 31041 256723 32223
rect 257847 31041 257969 32223
rect 256604 30938 257969 31041
rect 263744 32223 265109 32333
rect 263744 31041 263863 32223
rect 264987 31041 265109 32223
rect 263744 30938 265109 31041
rect 270702 32224 272067 32334
rect 270702 31042 270821 32224
rect 271945 31042 272067 32224
rect 270702 30939 272067 31042
rect 277838 32214 279203 32324
rect 277838 31032 277957 32214
rect 279081 31032 279203 32214
rect 277838 30929 279203 31032
rect 20624 21669 21989 21779
rect 20624 20487 20743 21669
rect 21867 20487 21989 21669
rect 20624 20384 21989 20487
rect 27582 21670 28947 21780
rect 27582 20488 27701 21670
rect 28825 20488 28947 21670
rect 27582 20385 28947 20488
rect 34502 21669 35867 21779
rect 34502 20487 34621 21669
rect 35745 20487 35867 21669
rect 34502 20384 35867 20487
rect 41467 21670 42832 21780
rect 41467 20488 41586 21670
rect 42710 20488 42832 21670
rect 41467 20385 42832 20488
rect 48425 21671 49790 21781
rect 48425 20489 48544 21671
rect 49668 20489 49790 21671
rect 48425 20386 49790 20489
rect 55342 21675 56707 21785
rect 55342 20493 55461 21675
rect 56585 20493 56707 21675
rect 55342 20390 56707 20493
rect 62307 21676 63672 21786
rect 62307 20494 62426 21676
rect 63550 20494 63672 21676
rect 62307 20391 63672 20494
rect 69265 21677 70630 21787
rect 69265 20495 69384 21677
rect 70508 20495 70630 21677
rect 69265 20392 70630 20495
rect 76182 21675 77547 21785
rect 76182 20493 76301 21675
rect 77425 20493 77547 21675
rect 76182 20390 77547 20493
rect 83147 21676 84512 21786
rect 83147 20494 83266 21676
rect 84390 20494 84512 21676
rect 83147 20391 84512 20494
rect 90105 21677 91470 21787
rect 90105 20495 90224 21677
rect 91348 20495 91470 21677
rect 90105 20392 91470 20495
rect 96923 21656 98288 21766
rect 96923 20474 97042 21656
rect 98166 20474 98288 21656
rect 96923 20371 98288 20474
rect 103888 21657 105253 21767
rect 103888 20475 104007 21657
rect 105131 20475 105253 21657
rect 103888 20372 105253 20475
rect 110846 21658 112211 21768
rect 110846 20476 110965 21658
rect 112089 20476 112211 21658
rect 110846 20373 112211 20476
rect 117766 21657 119131 21767
rect 117766 20475 117885 21657
rect 119009 20475 119131 21657
rect 117766 20372 119131 20475
rect 124731 21658 126096 21768
rect 124731 20476 124850 21658
rect 125974 20476 126096 21658
rect 124731 20373 126096 20476
rect 131689 21659 133054 21769
rect 131689 20477 131808 21659
rect 132932 20477 133054 21659
rect 131689 20374 133054 20477
rect 138606 21663 139971 21773
rect 138606 20481 138725 21663
rect 139849 20481 139971 21663
rect 138606 20378 139971 20481
rect 145571 21664 146936 21774
rect 145571 20482 145690 21664
rect 146814 20482 146936 21664
rect 145571 20379 146936 20482
rect 152529 21665 153894 21775
rect 152529 20483 152648 21665
rect 153772 20483 153894 21665
rect 152529 20380 153894 20483
rect 159446 21663 160811 21773
rect 159446 20481 159565 21663
rect 160689 20481 160811 21663
rect 159446 20378 160811 20481
rect 166411 21664 167776 21774
rect 166411 20482 166530 21664
rect 167654 20482 167776 21664
rect 166411 20379 167776 20482
rect 173369 21665 174734 21775
rect 173369 20483 173488 21665
rect 174612 20483 174734 21665
rect 173369 20380 174734 20483
rect 180174 21658 181539 21768
rect 180174 20476 180293 21658
rect 181417 20476 181539 21658
rect 180174 20373 181539 20476
rect 187139 21659 188504 21769
rect 187139 20477 187258 21659
rect 188382 20477 188504 21659
rect 187139 20374 188504 20477
rect 194097 21660 195462 21770
rect 194097 20478 194216 21660
rect 195340 20478 195462 21660
rect 194097 20375 195462 20478
rect 201017 21659 202382 21769
rect 201017 20477 201136 21659
rect 202260 20477 202382 21659
rect 201017 20374 202382 20477
rect 207982 21660 209347 21770
rect 207982 20478 208101 21660
rect 209225 20478 209347 21660
rect 207982 20375 209347 20478
rect 214940 21661 216305 21771
rect 214940 20479 215059 21661
rect 216183 20479 216305 21661
rect 214940 20376 216305 20479
rect 221857 21665 223222 21775
rect 221857 20483 221976 21665
rect 223100 20483 223222 21665
rect 221857 20380 223222 20483
rect 228822 21666 230187 21776
rect 228822 20484 228941 21666
rect 230065 20484 230187 21666
rect 228822 20381 230187 20484
rect 235780 21667 237145 21777
rect 235780 20485 235899 21667
rect 237023 20485 237145 21667
rect 235780 20382 237145 20485
rect 242697 21665 244062 21775
rect 242697 20483 242816 21665
rect 243940 20483 244062 21665
rect 242697 20380 244062 20483
rect 249662 21666 251027 21776
rect 249662 20484 249781 21666
rect 250905 20484 251027 21666
rect 249662 20381 251027 20484
rect 256620 21667 257985 21777
rect 256620 20485 256739 21667
rect 257863 20485 257985 21667
rect 256620 20382 257985 20485
rect 263760 21667 265125 21777
rect 263760 20485 263879 21667
rect 265003 20485 265125 21667
rect 263760 20382 265125 20485
rect 270718 21668 272083 21778
rect 270718 20486 270837 21668
rect 271961 20486 272083 21668
rect 270718 20383 272083 20486
rect 277854 21658 279219 21768
rect 277854 20476 277973 21658
rect 279097 20476 279219 21658
rect 277854 20373 279219 20476
rect 20608 15991 21973 16101
rect 20608 14809 20727 15991
rect 21851 14809 21973 15991
rect 20608 14706 21973 14809
rect 27566 15992 28931 16102
rect 27566 14810 27685 15992
rect 28809 14810 28931 15992
rect 27566 14707 28931 14810
rect 34486 15991 35851 16101
rect 34486 14809 34605 15991
rect 35729 14809 35851 15991
rect 34486 14706 35851 14809
rect 41451 15992 42816 16102
rect 41451 14810 41570 15992
rect 42694 14810 42816 15992
rect 41451 14707 42816 14810
rect 48409 15993 49774 16103
rect 48409 14811 48528 15993
rect 49652 14811 49774 15993
rect 48409 14708 49774 14811
rect 55326 15997 56691 16107
rect 55326 14815 55445 15997
rect 56569 14815 56691 15997
rect 55326 14712 56691 14815
rect 62291 15998 63656 16108
rect 62291 14816 62410 15998
rect 63534 14816 63656 15998
rect 62291 14713 63656 14816
rect 69249 15999 70614 16109
rect 69249 14817 69368 15999
rect 70492 14817 70614 15999
rect 69249 14714 70614 14817
rect 76166 15997 77531 16107
rect 76166 14815 76285 15997
rect 77409 14815 77531 15997
rect 76166 14712 77531 14815
rect 83131 15998 84496 16108
rect 83131 14816 83250 15998
rect 84374 14816 84496 15998
rect 83131 14713 84496 14816
rect 90089 15999 91454 16109
rect 90089 14817 90208 15999
rect 91332 14817 91454 15999
rect 90089 14714 91454 14817
rect 96907 15978 98272 16088
rect 96907 14796 97026 15978
rect 98150 14796 98272 15978
rect 96907 14693 98272 14796
rect 103872 15979 105237 16089
rect 103872 14797 103991 15979
rect 105115 14797 105237 15979
rect 103872 14694 105237 14797
rect 110830 15980 112195 16090
rect 110830 14798 110949 15980
rect 112073 14798 112195 15980
rect 110830 14695 112195 14798
rect 117750 15979 119115 16089
rect 117750 14797 117869 15979
rect 118993 14797 119115 15979
rect 117750 14694 119115 14797
rect 124715 15980 126080 16090
rect 124715 14798 124834 15980
rect 125958 14798 126080 15980
rect 124715 14695 126080 14798
rect 131673 15981 133038 16091
rect 131673 14799 131792 15981
rect 132916 14799 133038 15981
rect 131673 14696 133038 14799
rect 138590 15985 139955 16095
rect 138590 14803 138709 15985
rect 139833 14803 139955 15985
rect 138590 14700 139955 14803
rect 145555 15986 146920 16096
rect 145555 14804 145674 15986
rect 146798 14804 146920 15986
rect 145555 14701 146920 14804
rect 152513 15987 153878 16097
rect 152513 14805 152632 15987
rect 153756 14805 153878 15987
rect 152513 14702 153878 14805
rect 159430 15985 160795 16095
rect 159430 14803 159549 15985
rect 160673 14803 160795 15985
rect 159430 14700 160795 14803
rect 166395 15986 167760 16096
rect 166395 14804 166514 15986
rect 167638 14804 167760 15986
rect 166395 14701 167760 14804
rect 173353 15987 174718 16097
rect 173353 14805 173472 15987
rect 174596 14805 174718 15987
rect 173353 14702 174718 14805
rect 180158 15980 181523 16090
rect 180158 14798 180277 15980
rect 181401 14798 181523 15980
rect 180158 14695 181523 14798
rect 187123 15981 188488 16091
rect 187123 14799 187242 15981
rect 188366 14799 188488 15981
rect 187123 14696 188488 14799
rect 194081 15982 195446 16092
rect 194081 14800 194200 15982
rect 195324 14800 195446 15982
rect 194081 14697 195446 14800
rect 201001 15981 202366 16091
rect 201001 14799 201120 15981
rect 202244 14799 202366 15981
rect 201001 14696 202366 14799
rect 207966 15982 209331 16092
rect 207966 14800 208085 15982
rect 209209 14800 209331 15982
rect 207966 14697 209331 14800
rect 214924 15983 216289 16093
rect 214924 14801 215043 15983
rect 216167 14801 216289 15983
rect 214924 14698 216289 14801
rect 221841 15987 223206 16097
rect 221841 14805 221960 15987
rect 223084 14805 223206 15987
rect 221841 14702 223206 14805
rect 228806 15988 230171 16098
rect 228806 14806 228925 15988
rect 230049 14806 230171 15988
rect 228806 14703 230171 14806
rect 235764 15989 237129 16099
rect 235764 14807 235883 15989
rect 237007 14807 237129 15989
rect 235764 14704 237129 14807
rect 242681 15987 244046 16097
rect 242681 14805 242800 15987
rect 243924 14805 244046 15987
rect 242681 14702 244046 14805
rect 249646 15988 251011 16098
rect 249646 14806 249765 15988
rect 250889 14806 251011 15988
rect 249646 14703 251011 14806
rect 256604 15989 257969 16099
rect 256604 14807 256723 15989
rect 257847 14807 257969 15989
rect 256604 14704 257969 14807
rect 263744 15989 265109 16099
rect 263744 14807 263863 15989
rect 264987 14807 265109 15989
rect 263744 14704 265109 14807
rect 270702 15990 272067 16100
rect 270702 14808 270821 15990
rect 271945 14808 272067 15990
rect 270702 14705 272067 14808
rect 277838 15980 279203 16090
rect 277838 14798 277957 15980
rect 279081 14798 279203 15980
rect 277838 14695 279203 14798
rect 20608 8898 21973 9008
rect 20608 7716 20727 8898
rect 21851 7716 21973 8898
rect 20608 7613 21973 7716
rect 27566 8899 28931 9009
rect 27566 7717 27685 8899
rect 28809 7717 28931 8899
rect 27566 7614 28931 7717
rect 34486 8898 35851 9008
rect 34486 7716 34605 8898
rect 35729 7716 35851 8898
rect 34486 7613 35851 7716
rect 41451 8899 42816 9009
rect 41451 7717 41570 8899
rect 42694 7717 42816 8899
rect 41451 7614 42816 7717
rect 48409 8900 49774 9010
rect 48409 7718 48528 8900
rect 49652 7718 49774 8900
rect 48409 7615 49774 7718
rect 55326 8904 56691 9014
rect 55326 7722 55445 8904
rect 56569 7722 56691 8904
rect 55326 7619 56691 7722
rect 62291 8905 63656 9015
rect 62291 7723 62410 8905
rect 63534 7723 63656 8905
rect 62291 7620 63656 7723
rect 69249 8906 70614 9016
rect 69249 7724 69368 8906
rect 70492 7724 70614 8906
rect 69249 7621 70614 7724
rect 76166 8904 77531 9014
rect 76166 7722 76285 8904
rect 77409 7722 77531 8904
rect 76166 7619 77531 7722
rect 83131 8905 84496 9015
rect 83131 7723 83250 8905
rect 84374 7723 84496 8905
rect 83131 7620 84496 7723
rect 90089 8906 91454 9016
rect 90089 7724 90208 8906
rect 91332 7724 91454 8906
rect 90089 7621 91454 7724
rect 96907 8885 98272 8995
rect 96907 7703 97026 8885
rect 98150 7703 98272 8885
rect 96907 7600 98272 7703
rect 103872 8886 105237 8996
rect 103872 7704 103991 8886
rect 105115 7704 105237 8886
rect 103872 7601 105237 7704
rect 110830 8887 112195 8997
rect 110830 7705 110949 8887
rect 112073 7705 112195 8887
rect 110830 7602 112195 7705
rect 117750 8886 119115 8996
rect 117750 7704 117869 8886
rect 118993 7704 119115 8886
rect 117750 7601 119115 7704
rect 124715 8887 126080 8997
rect 124715 7705 124834 8887
rect 125958 7705 126080 8887
rect 124715 7602 126080 7705
rect 131673 8888 133038 8998
rect 131673 7706 131792 8888
rect 132916 7706 133038 8888
rect 131673 7603 133038 7706
rect 138590 8892 139955 9002
rect 138590 7710 138709 8892
rect 139833 7710 139955 8892
rect 138590 7607 139955 7710
rect 145555 8893 146920 9003
rect 145555 7711 145674 8893
rect 146798 7711 146920 8893
rect 145555 7608 146920 7711
rect 152513 8894 153878 9004
rect 152513 7712 152632 8894
rect 153756 7712 153878 8894
rect 152513 7609 153878 7712
rect 159430 8892 160795 9002
rect 159430 7710 159549 8892
rect 160673 7710 160795 8892
rect 159430 7607 160795 7710
rect 166395 8893 167760 9003
rect 166395 7711 166514 8893
rect 167638 7711 167760 8893
rect 166395 7608 167760 7711
rect 173353 8894 174718 9004
rect 173353 7712 173472 8894
rect 174596 7712 174718 8894
rect 173353 7609 174718 7712
rect 180158 8887 181523 8997
rect 180158 7705 180277 8887
rect 181401 7705 181523 8887
rect 180158 7602 181523 7705
rect 187123 8888 188488 8998
rect 187123 7706 187242 8888
rect 188366 7706 188488 8888
rect 187123 7603 188488 7706
rect 194081 8889 195446 8999
rect 194081 7707 194200 8889
rect 195324 7707 195446 8889
rect 194081 7604 195446 7707
rect 201001 8888 202366 8998
rect 201001 7706 201120 8888
rect 202244 7706 202366 8888
rect 201001 7603 202366 7706
rect 207966 8889 209331 8999
rect 207966 7707 208085 8889
rect 209209 7707 209331 8889
rect 207966 7604 209331 7707
rect 214924 8890 216289 9000
rect 214924 7708 215043 8890
rect 216167 7708 216289 8890
rect 214924 7605 216289 7708
rect 221841 8894 223206 9004
rect 221841 7712 221960 8894
rect 223084 7712 223206 8894
rect 221841 7609 223206 7712
rect 228806 8895 230171 9005
rect 228806 7713 228925 8895
rect 230049 7713 230171 8895
rect 228806 7610 230171 7713
rect 235764 8896 237129 9006
rect 235764 7714 235883 8896
rect 237007 7714 237129 8896
rect 235764 7611 237129 7714
rect 242681 8894 244046 9004
rect 242681 7712 242800 8894
rect 243924 7712 244046 8894
rect 242681 7609 244046 7712
rect 249646 8895 251011 9005
rect 249646 7713 249765 8895
rect 250889 7713 251011 8895
rect 249646 7610 251011 7713
rect 256604 8896 257969 9006
rect 256604 7714 256723 8896
rect 257847 7714 257969 8896
rect 256604 7611 257969 7714
rect 263744 8896 265109 9006
rect 263744 7714 263863 8896
rect 264987 7714 265109 8896
rect 263744 7611 265109 7714
rect 270702 8897 272067 9007
rect 270702 7715 270821 8897
rect 271945 7715 272067 8897
rect 270702 7612 272067 7715
rect 277838 8887 279203 8997
rect 277838 7705 277957 8887
rect 279081 7705 279203 8887
rect 277838 7602 279203 7705
<< nsubdiff >>
rect 26431 264775 26576 264790
rect 26431 264665 26446 264775
rect 26561 264665 26576 264775
rect 26431 264655 26576 264665
rect 23581 264447 23730 264462
rect 23581 264330 23597 264447
rect 23716 264330 23730 264447
rect 23581 264315 23730 264330
<< psubdiffcont >>
rect 69629 338866 70753 340048
rect 76546 338864 77670 340046
rect 83511 338865 84635 340047
rect 90469 338866 91593 340048
rect 97287 338845 98411 340027
rect 104252 338846 105376 340028
rect 111210 338847 112334 340029
rect 118130 338846 119254 340028
rect 125095 338847 126219 340029
rect 132053 338848 133177 340030
rect 138970 338852 140094 340034
rect 145935 338853 147059 340035
rect 152893 338854 154017 340036
rect 159810 338852 160934 340034
rect 166775 338853 167899 340035
rect 173733 338854 174857 340036
rect 180538 338847 181662 340029
rect 187503 338848 188627 340030
rect 194461 338849 195585 340031
rect 201381 338848 202505 340030
rect 208346 338849 209470 340031
rect 215304 338850 216428 340032
rect 69355 331736 70479 332918
rect 76272 331734 77396 332916
rect 83237 331735 84361 332917
rect 90195 331736 91319 332918
rect 97013 331715 98137 332897
rect 103978 331716 105102 332898
rect 110936 331717 112060 332899
rect 117856 331716 118980 332898
rect 124821 331717 125945 332899
rect 131779 331718 132903 332900
rect 138696 331722 139820 332904
rect 145661 331723 146785 332905
rect 152619 331724 153743 332906
rect 159536 331722 160660 332904
rect 166501 331723 167625 332905
rect 173459 331724 174583 332906
rect 180264 331717 181388 332899
rect 187229 331718 188353 332900
rect 194187 331719 195311 332901
rect 201107 331718 202231 332900
rect 208072 331719 209196 332901
rect 215030 331720 216154 332902
rect 69629 325408 70753 326590
rect 76546 325406 77670 326588
rect 83511 325407 84635 326589
rect 90469 325408 91593 326590
rect 97287 325387 98411 326569
rect 104252 325388 105376 326570
rect 111210 325389 112334 326571
rect 118130 325388 119254 326570
rect 125095 325389 126219 326571
rect 132053 325390 133177 326572
rect 138970 325394 140094 326576
rect 145935 325395 147059 326577
rect 152893 325396 154017 326578
rect 159810 325394 160934 326576
rect 166775 325395 167899 326577
rect 173733 325396 174857 326578
rect 180538 325389 181662 326571
rect 187503 325390 188627 326572
rect 194461 325391 195585 326573
rect 201381 325390 202505 326572
rect 208346 325391 209470 326573
rect 215304 325392 216428 326574
rect 69355 318278 70479 319460
rect 76272 318276 77396 319458
rect 83237 318277 84361 319459
rect 90195 318278 91319 319460
rect 97013 318257 98137 319439
rect 103978 318258 105102 319440
rect 110936 318259 112060 319441
rect 117856 318258 118980 319440
rect 124821 318259 125945 319441
rect 131779 318260 132903 319442
rect 138696 318264 139820 319446
rect 145661 318265 146785 319447
rect 152619 318266 153743 319448
rect 159536 318264 160660 319446
rect 166501 318265 167625 319447
rect 173459 318266 174583 319448
rect 180264 318259 181388 319441
rect 187229 318260 188353 319442
rect 194187 318261 195311 319443
rect 201107 318260 202231 319442
rect 208072 318261 209196 319443
rect 215030 318262 216154 319444
rect 20994 311139 22118 312321
rect 27952 311140 29076 312322
rect 34872 311139 35996 312321
rect 41837 311140 42961 312322
rect 48795 311141 49919 312323
rect 55712 311145 56836 312327
rect 62677 311146 63801 312328
rect 69635 311147 70759 312329
rect 76552 311145 77676 312327
rect 83517 311146 84641 312328
rect 90475 311147 91599 312329
rect 97293 311126 98417 312308
rect 104258 311127 105382 312309
rect 111216 311128 112340 312310
rect 118136 311127 119260 312309
rect 125101 311128 126225 312310
rect 132059 311129 133183 312311
rect 138976 311133 140100 312315
rect 145941 311134 147065 312316
rect 152899 311135 154023 312317
rect 159816 311133 160940 312315
rect 166781 311134 167905 312316
rect 173739 311135 174863 312317
rect 180544 311128 181668 312310
rect 187509 311129 188633 312311
rect 194467 311130 195591 312312
rect 201387 311129 202511 312311
rect 208352 311130 209476 312312
rect 215310 311131 216434 312313
rect 20720 304009 21844 305191
rect 27678 304010 28802 305192
rect 34598 304009 35722 305191
rect 41563 304010 42687 305192
rect 48521 304011 49645 305193
rect 55438 304015 56562 305197
rect 62403 304016 63527 305198
rect 69361 304017 70485 305199
rect 76278 304015 77402 305197
rect 83243 304016 84367 305198
rect 90201 304017 91325 305199
rect 97019 303996 98143 305178
rect 103984 303997 105108 305179
rect 110942 303998 112066 305180
rect 117862 303997 118986 305179
rect 124827 303998 125951 305180
rect 131785 303999 132909 305181
rect 138702 304003 139826 305185
rect 145667 304004 146791 305186
rect 152625 304005 153749 305187
rect 159542 304003 160666 305185
rect 166507 304004 167631 305186
rect 173465 304005 174589 305187
rect 180270 303998 181394 305180
rect 187235 303999 188359 305181
rect 194193 304000 195317 305182
rect 201113 303999 202237 305181
rect 208078 304000 209202 305182
rect 215036 304001 216160 305183
rect 21083 294780 22207 295962
rect 28041 294781 29165 295963
rect 34961 294780 36085 295962
rect 41926 294781 43050 295963
rect 48884 294782 50008 295964
rect 55801 294786 56925 295968
rect 62766 294787 63890 295969
rect 69724 294788 70848 295970
rect 76641 294786 77765 295968
rect 83606 294787 84730 295969
rect 90564 294788 91688 295970
rect 97382 294767 98506 295949
rect 104347 294768 105471 295950
rect 111305 294769 112429 295951
rect 118225 294768 119349 295950
rect 125190 294769 126314 295951
rect 132148 294770 133272 295952
rect 139065 294774 140189 295956
rect 146030 294775 147154 295957
rect 152988 294776 154112 295958
rect 159905 294774 161029 295956
rect 166870 294775 167994 295957
rect 173828 294776 174952 295958
rect 180633 294769 181757 295951
rect 187598 294770 188722 295952
rect 194556 294771 195680 295953
rect 201476 294770 202600 295952
rect 208441 294771 209565 295953
rect 215399 294772 216523 295954
rect 222316 294776 223440 295958
rect 229281 294777 230405 295959
rect 236239 294778 237363 295960
rect 243156 294776 244280 295958
rect 250121 294777 251245 295959
rect 257079 294778 258203 295960
rect 264219 294778 265343 295960
rect 271177 294779 272301 295961
rect 278313 294769 279437 295951
rect 20809 287650 21933 288832
rect 27767 287651 28891 288833
rect 34687 287650 35811 288832
rect 41652 287651 42776 288833
rect 48610 287652 49734 288834
rect 55527 287656 56651 288838
rect 62492 287657 63616 288839
rect 69450 287658 70574 288840
rect 76367 287656 77491 288838
rect 83332 287657 84456 288839
rect 90290 287658 91414 288840
rect 97108 287637 98232 288819
rect 104073 287638 105197 288820
rect 111031 287639 112155 288821
rect 117951 287638 119075 288820
rect 124916 287639 126040 288821
rect 131874 287640 132998 288822
rect 138791 287644 139915 288826
rect 145756 287645 146880 288827
rect 152714 287646 153838 288828
rect 159631 287644 160755 288826
rect 166596 287645 167720 288827
rect 173554 287646 174678 288828
rect 180359 287639 181483 288821
rect 187324 287640 188448 288822
rect 194282 287641 195406 288823
rect 201202 287640 202326 288822
rect 208167 287641 209291 288823
rect 215125 287642 216249 288824
rect 222042 287646 223166 288828
rect 229007 287647 230131 288829
rect 235965 287648 237089 288830
rect 242882 287646 244006 288828
rect 249847 287647 250971 288829
rect 256805 287648 257929 288830
rect 263945 287648 265069 288830
rect 270903 287649 272027 288831
rect 278039 287639 279163 288821
rect 20917 281237 22041 282419
rect 27875 281238 28999 282420
rect 34795 281237 35919 282419
rect 41760 281238 42884 282420
rect 48718 281239 49842 282421
rect 55635 281243 56759 282425
rect 62600 281244 63724 282426
rect 69558 281245 70682 282427
rect 76475 281243 77599 282425
rect 83440 281244 84564 282426
rect 90398 281245 91522 282427
rect 97216 281224 98340 282406
rect 104181 281225 105305 282407
rect 111139 281226 112263 282408
rect 118059 281225 119183 282407
rect 125024 281226 126148 282408
rect 131982 281227 133106 282409
rect 138899 281231 140023 282413
rect 145864 281232 146988 282414
rect 152822 281233 153946 282415
rect 159739 281231 160863 282413
rect 166704 281232 167828 282414
rect 173662 281233 174786 282415
rect 180467 281226 181591 282408
rect 187432 281227 188556 282409
rect 194390 281228 195514 282410
rect 201310 281227 202434 282409
rect 208275 281228 209399 282410
rect 215233 281229 216357 282411
rect 222150 281233 223274 282415
rect 229115 281234 230239 282416
rect 236073 281235 237197 282417
rect 242990 281233 244114 282415
rect 249955 281234 251079 282416
rect 256913 281235 258037 282417
rect 264053 281235 265177 282417
rect 271011 281236 272135 282418
rect 278147 281226 279271 282408
rect 69775 272380 70899 273562
rect 76692 272378 77816 273560
rect 83657 272379 84781 273561
rect 90615 272380 91739 273562
rect 97433 272359 98557 273541
rect 104398 272360 105522 273542
rect 111356 272361 112480 273543
rect 118276 272360 119400 273542
rect 125241 272361 126365 273543
rect 132199 272362 133323 273544
rect 139116 272366 140240 273548
rect 146081 272367 147205 273549
rect 153039 272368 154163 273550
rect 159956 272366 161080 273548
rect 166921 272367 168045 273549
rect 173879 272368 175003 273550
rect 180684 272361 181808 273543
rect 187649 272362 188773 273544
rect 194607 272363 195731 273545
rect 201527 272362 202651 273544
rect 208492 272363 209616 273545
rect 215450 272364 216574 273546
rect 222367 272368 223491 273550
rect 69501 265250 70625 266432
rect 76418 265248 77542 266430
rect 83383 265249 84507 266431
rect 90341 265250 91465 266432
rect 97159 265229 98283 266411
rect 104124 265230 105248 266412
rect 111082 265231 112206 266413
rect 118002 265230 119126 266412
rect 124967 265231 126091 266413
rect 131925 265232 133049 266414
rect 138842 265236 139966 266418
rect 145807 265237 146931 266419
rect 152765 265238 153889 266420
rect 159682 265236 160806 266418
rect 166647 265237 167771 266419
rect 173605 265238 174729 266420
rect 180410 265231 181534 266413
rect 187375 265232 188499 266414
rect 194333 265233 195457 266415
rect 201253 265232 202377 266414
rect 208218 265233 209342 266415
rect 215176 265234 216300 266416
rect 222093 265238 223217 266420
rect 69609 258837 70733 260019
rect 76526 258835 77650 260017
rect 83491 258836 84615 260018
rect 90449 258837 91573 260019
rect 97267 258816 98391 259998
rect 104232 258817 105356 259999
rect 111190 258818 112314 260000
rect 118110 258817 119234 259999
rect 125075 258818 126199 260000
rect 132033 258819 133157 260001
rect 138950 258823 140074 260005
rect 145915 258824 147039 260006
rect 152873 258825 153997 260007
rect 159790 258823 160914 260005
rect 166755 258824 167879 260006
rect 173713 258825 174837 260007
rect 180518 258818 181642 260000
rect 187483 258819 188607 260001
rect 194441 258820 195565 260002
rect 201361 258819 202485 260001
rect 208326 258820 209450 260002
rect 215284 258821 216408 260003
rect 222201 258825 223325 260007
rect 83688 248125 84812 249307
rect 90646 248126 91770 249308
rect 97464 248105 98588 249287
rect 104429 248106 105553 249288
rect 111387 248107 112511 249289
rect 118307 248106 119431 249288
rect 125272 248107 126396 249289
rect 132230 248108 133354 249290
rect 139147 248112 140271 249294
rect 146112 248113 147236 249295
rect 153070 248114 154194 249296
rect 159987 248112 161111 249294
rect 166952 248113 168076 249295
rect 173910 248114 175034 249296
rect 180715 248107 181839 249289
rect 187680 248108 188804 249290
rect 194638 248109 195762 249291
rect 201558 248108 202682 249290
rect 208523 248109 209647 249291
rect 215481 248110 216605 249292
rect 222398 248114 223522 249296
rect 83414 240995 84538 242177
rect 90372 240996 91496 242178
rect 97190 240975 98314 242157
rect 104155 240976 105279 242158
rect 111113 240977 112237 242159
rect 118033 240976 119157 242158
rect 124998 240977 126122 242159
rect 131956 240978 133080 242160
rect 138873 240982 139997 242164
rect 145838 240983 146962 242165
rect 152796 240984 153920 242166
rect 159713 240982 160837 242164
rect 166678 240983 167802 242165
rect 173636 240984 174760 242166
rect 180441 240977 181565 242159
rect 187406 240978 188530 242160
rect 194364 240979 195488 242161
rect 201284 240978 202408 242160
rect 208249 240979 209373 242161
rect 215207 240980 216331 242162
rect 222124 240984 223248 242166
rect 83522 234582 84646 235764
rect 90480 234583 91604 235765
rect 97298 234562 98422 235744
rect 104263 234563 105387 235745
rect 111221 234564 112345 235746
rect 118141 234563 119265 235745
rect 125106 234564 126230 235746
rect 132064 234565 133188 235747
rect 138981 234569 140105 235751
rect 145946 234570 147070 235752
rect 152904 234571 154028 235753
rect 159821 234569 160945 235751
rect 166786 234570 167910 235752
rect 173744 234571 174868 235753
rect 180549 234564 181673 235746
rect 187514 234565 188638 235747
rect 194472 234566 195596 235748
rect 201392 234565 202516 235747
rect 208357 234566 209481 235748
rect 215315 234567 216439 235749
rect 222232 234571 223356 235753
rect 49090 227854 50214 229036
rect 56007 227858 57131 229040
rect 62972 227859 64096 229041
rect 69930 227860 71054 229042
rect 76847 227858 77971 229040
rect 83812 227859 84936 229041
rect 90770 227860 91894 229042
rect 97588 227839 98712 229021
rect 104553 227840 105677 229022
rect 111511 227841 112635 229023
rect 118431 227840 119555 229022
rect 125396 227841 126520 229023
rect 132354 227842 133478 229024
rect 139271 227846 140395 229028
rect 146236 227847 147360 229029
rect 153194 227848 154318 229030
rect 160111 227846 161235 229028
rect 167076 227847 168200 229029
rect 174034 227848 175158 229030
rect 180839 227841 181963 229023
rect 187804 227842 188928 229024
rect 194762 227843 195886 229025
rect 201682 227842 202806 229024
rect 208647 227843 209771 229025
rect 215605 227844 216729 229026
rect 222522 227848 223646 229030
rect 229487 227849 230611 229031
rect 236445 227850 237569 229032
rect 243362 227848 244486 229030
rect 250327 227849 251451 229031
rect 257285 227850 258409 229032
rect 264425 227850 265549 229032
rect 271383 227851 272507 229033
rect 278519 227841 279643 229023
rect 49070 221992 50194 223174
rect 55987 221996 57111 223178
rect 62952 221997 64076 223179
rect 69910 221998 71034 223180
rect 76827 221996 77951 223178
rect 83792 221997 84916 223179
rect 90750 221998 91874 223180
rect 97568 221977 98692 223159
rect 104533 221978 105657 223160
rect 111491 221979 112615 223161
rect 118411 221978 119535 223160
rect 125376 221979 126500 223161
rect 132334 221980 133458 223162
rect 139251 221984 140375 223166
rect 146216 221985 147340 223167
rect 153174 221986 154298 223168
rect 160091 221984 161215 223166
rect 167056 221985 168180 223167
rect 174014 221986 175138 223168
rect 180819 221979 181943 223161
rect 187784 221980 188908 223162
rect 194742 221981 195866 223163
rect 201662 221980 202786 223162
rect 208627 221981 209751 223163
rect 215585 221982 216709 223164
rect 222502 221986 223626 223168
rect 229467 221987 230591 223169
rect 236425 221988 237549 223170
rect 243342 221986 244466 223168
rect 250307 221987 251431 223169
rect 257265 221988 258389 223170
rect 264405 221988 265529 223170
rect 271363 221989 272487 223171
rect 278499 221979 279623 223161
rect 21309 209927 22433 211109
rect 28267 209928 29391 211110
rect 35187 209927 36311 211109
rect 42152 209928 43276 211110
rect 49110 209929 50234 211111
rect 56027 209933 57151 211115
rect 62992 209934 64116 211116
rect 69950 209935 71074 211117
rect 76867 209933 77991 211115
rect 83832 209934 84956 211116
rect 90790 209935 91914 211117
rect 97608 209914 98732 211096
rect 104573 209915 105697 211097
rect 111531 209916 112655 211098
rect 118451 209915 119575 211097
rect 125416 209916 126540 211098
rect 132374 209917 133498 211099
rect 139291 209921 140415 211103
rect 146256 209922 147380 211104
rect 153214 209923 154338 211105
rect 160131 209921 161255 211103
rect 167096 209922 168220 211104
rect 174054 209923 175178 211105
rect 180859 209916 181983 211098
rect 187824 209917 188948 211099
rect 194782 209918 195906 211100
rect 201702 209917 202826 211099
rect 208667 209918 209791 211100
rect 215625 209919 216749 211101
rect 222542 209923 223666 211105
rect 229507 209924 230631 211106
rect 236465 209925 237589 211107
rect 243382 209923 244506 211105
rect 250347 209924 251471 211106
rect 257305 209925 258429 211107
rect 264445 209925 265569 211107
rect 271403 209926 272527 211108
rect 278539 209916 279663 211098
rect 21035 202797 22159 203979
rect 27993 202798 29117 203980
rect 34913 202797 36037 203979
rect 41878 202798 43002 203980
rect 48836 202799 49960 203981
rect 55753 202803 56877 203985
rect 62718 202804 63842 203986
rect 69676 202805 70800 203987
rect 76593 202803 77717 203985
rect 83558 202804 84682 203986
rect 90516 202805 91640 203987
rect 97334 202784 98458 203966
rect 104299 202785 105423 203967
rect 111257 202786 112381 203968
rect 118177 202785 119301 203967
rect 125142 202786 126266 203968
rect 132100 202787 133224 203969
rect 139017 202791 140141 203973
rect 145982 202792 147106 203974
rect 152940 202793 154064 203975
rect 159857 202791 160981 203973
rect 166822 202792 167946 203974
rect 173780 202793 174904 203975
rect 180585 202786 181709 203968
rect 187550 202787 188674 203969
rect 194508 202788 195632 203970
rect 201428 202787 202552 203969
rect 208393 202788 209517 203970
rect 215351 202789 216475 203971
rect 222268 202793 223392 203975
rect 229233 202794 230357 203976
rect 236191 202795 237315 203977
rect 243108 202793 244232 203975
rect 250073 202794 251197 203976
rect 257031 202795 258155 203977
rect 264171 202795 265295 203977
rect 271129 202796 272253 203978
rect 278265 202786 279389 203968
rect 21143 196384 22267 197566
rect 28101 196385 29225 197567
rect 35021 196384 36145 197566
rect 41986 196385 43110 197567
rect 48944 196386 50068 197568
rect 55861 196390 56985 197572
rect 62826 196391 63950 197573
rect 69784 196392 70908 197574
rect 76701 196390 77825 197572
rect 83666 196391 84790 197573
rect 90624 196392 91748 197574
rect 97442 196371 98566 197553
rect 104407 196372 105531 197554
rect 111365 196373 112489 197555
rect 118285 196372 119409 197554
rect 125250 196373 126374 197555
rect 132208 196374 133332 197556
rect 139125 196378 140249 197560
rect 146090 196379 147214 197561
rect 153048 196380 154172 197562
rect 159965 196378 161089 197560
rect 166930 196379 168054 197561
rect 173888 196380 175012 197562
rect 180693 196373 181817 197555
rect 187658 196374 188782 197556
rect 194616 196375 195740 197557
rect 201536 196374 202660 197556
rect 208501 196375 209625 197557
rect 215459 196376 216583 197558
rect 222376 196380 223500 197562
rect 229341 196381 230465 197563
rect 236299 196382 237423 197564
rect 243216 196380 244340 197562
rect 250181 196381 251305 197563
rect 257139 196382 258263 197564
rect 264279 196382 265403 197564
rect 271237 196383 272361 197565
rect 278373 196373 279497 197555
rect 76854 192040 77978 193222
rect 83819 192041 84943 193223
rect 90777 192042 91901 193224
rect 97595 192021 98719 193203
rect 104560 192022 105684 193204
rect 111518 192023 112642 193205
rect 118438 192022 119562 193204
rect 125403 192023 126527 193205
rect 132361 192024 133485 193206
rect 139278 192028 140402 193210
rect 146243 192029 147367 193211
rect 153201 192030 154325 193212
rect 160118 192028 161242 193210
rect 167083 192029 168207 193211
rect 174041 192030 175165 193212
rect 180846 192023 181970 193205
rect 187811 192024 188935 193206
rect 194769 192025 195893 193207
rect 201689 192024 202813 193206
rect 208654 192025 209778 193207
rect 215612 192026 216736 193208
rect 222529 192030 223653 193212
rect 229494 192031 230618 193213
rect 236452 192032 237576 193214
rect 243369 192030 244493 193212
rect 250334 192031 251458 193213
rect 257292 192032 258416 193214
rect 264432 192032 265556 193214
rect 271390 192033 272514 193215
rect 278526 192023 279650 193205
rect 76580 184910 77704 186092
rect 83545 184911 84669 186093
rect 90503 184912 91627 186094
rect 97321 184891 98445 186073
rect 104286 184892 105410 186074
rect 111244 184893 112368 186075
rect 118164 184892 119288 186074
rect 125129 184893 126253 186075
rect 132087 184894 133211 186076
rect 139004 184898 140128 186080
rect 145969 184899 147093 186081
rect 152927 184900 154051 186082
rect 159844 184898 160968 186080
rect 166809 184899 167933 186081
rect 173767 184900 174891 186082
rect 180572 184893 181696 186075
rect 187537 184894 188661 186076
rect 194495 184895 195619 186077
rect 201415 184894 202539 186076
rect 208380 184895 209504 186077
rect 215338 184896 216462 186078
rect 222255 184900 223379 186082
rect 229220 184901 230344 186083
rect 236178 184902 237302 186084
rect 243095 184900 244219 186082
rect 250060 184901 251184 186083
rect 257018 184902 258142 186084
rect 264158 184902 265282 186084
rect 271116 184903 272240 186085
rect 278252 184893 279376 186075
rect 76688 178497 77812 179679
rect 83653 178498 84777 179680
rect 90611 178499 91735 179681
rect 97429 178478 98553 179660
rect 104394 178479 105518 179661
rect 111352 178480 112476 179662
rect 118272 178479 119396 179661
rect 125237 178480 126361 179662
rect 132195 178481 133319 179663
rect 139112 178485 140236 179667
rect 146077 178486 147201 179668
rect 153035 178487 154159 179669
rect 159952 178485 161076 179667
rect 166917 178486 168041 179668
rect 173875 178487 174999 179669
rect 180680 178480 181804 179662
rect 187645 178481 188769 179663
rect 194603 178482 195727 179664
rect 201523 178481 202647 179663
rect 208488 178482 209612 179664
rect 215446 178483 216570 179665
rect 222363 178487 223487 179669
rect 229328 178488 230452 179670
rect 236286 178489 237410 179671
rect 243203 178487 244327 179669
rect 250168 178488 251292 179670
rect 257126 178489 258250 179671
rect 264266 178489 265390 179671
rect 271224 178490 272348 179672
rect 278360 178480 279484 179662
rect 48646 172579 49770 173761
rect 55563 172583 56687 173765
rect 62528 172584 63652 173766
rect 69486 172585 70610 173767
rect 76403 172583 77527 173765
rect 83368 172584 84492 173766
rect 90326 172585 91450 173767
rect 97144 172564 98268 173746
rect 104109 172565 105233 173747
rect 111067 172566 112191 173748
rect 117987 172565 119111 173747
rect 124952 172566 126076 173748
rect 131910 172567 133034 173749
rect 138827 172571 139951 173753
rect 145792 172572 146916 173754
rect 152750 172573 153874 173755
rect 159667 172571 160791 173753
rect 166632 172572 167756 173754
rect 173590 172573 174714 173755
rect 180395 172566 181519 173748
rect 187360 172567 188484 173749
rect 194318 172568 195442 173750
rect 201238 172567 202362 173749
rect 208203 172568 209327 173750
rect 215161 172569 216285 173751
rect 222078 172573 223202 173755
rect 229043 172574 230167 173756
rect 236001 172575 237125 173757
rect 242918 172573 244042 173755
rect 249883 172574 251007 173756
rect 256841 172575 257965 173757
rect 263981 172575 265105 173757
rect 270939 172576 272063 173758
rect 278075 172566 279199 173748
rect 48754 166166 49878 167348
rect 55671 166170 56795 167352
rect 62636 166171 63760 167353
rect 69594 166172 70718 167354
rect 76511 166170 77635 167352
rect 83476 166171 84600 167353
rect 90434 166172 91558 167354
rect 97252 166151 98376 167333
rect 104217 166152 105341 167334
rect 111175 166153 112299 167335
rect 118095 166152 119219 167334
rect 125060 166153 126184 167335
rect 132018 166154 133142 167336
rect 138935 166158 140059 167340
rect 145900 166159 147024 167341
rect 152858 166160 153982 167342
rect 159775 166158 160899 167340
rect 166740 166159 167864 167341
rect 173698 166160 174822 167342
rect 180503 166153 181627 167335
rect 187468 166154 188592 167336
rect 194426 166155 195550 167337
rect 201346 166154 202470 167336
rect 208311 166155 209435 167337
rect 215269 166156 216393 167338
rect 222186 166160 223310 167342
rect 229151 166161 230275 167343
rect 236109 166162 237233 167344
rect 243026 166160 244150 167342
rect 249991 166161 251115 167343
rect 256949 166162 258073 167344
rect 264089 166162 265213 167344
rect 271047 166163 272171 167345
rect 278183 166153 279307 167335
rect 21720 158825 22844 160007
rect 28678 158826 29802 160008
rect 35598 158825 36722 160007
rect 42563 158826 43687 160008
rect 49521 158827 50645 160009
rect 56438 158831 57562 160013
rect 63403 158832 64527 160014
rect 70361 158833 71485 160015
rect 77278 158831 78402 160013
rect 84243 158832 85367 160014
rect 91201 158833 92325 160015
rect 98019 158812 99143 159994
rect 104984 158813 106108 159995
rect 111942 158814 113066 159996
rect 118862 158813 119986 159995
rect 125827 158814 126951 159996
rect 132785 158815 133909 159997
rect 139702 158819 140826 160001
rect 146667 158820 147791 160002
rect 153625 158821 154749 160003
rect 160542 158819 161666 160001
rect 167507 158820 168631 160002
rect 174465 158821 175589 160003
rect 181270 158814 182394 159996
rect 188235 158815 189359 159997
rect 195193 158816 196317 159998
rect 202113 158815 203237 159997
rect 209078 158816 210202 159998
rect 216036 158817 217160 159999
rect 222953 158821 224077 160003
rect 229792 158816 230916 159998
rect 236757 158817 237881 159999
rect 243715 158818 244839 160000
rect 250632 158822 251756 160004
rect 257524 158805 258648 159987
rect 264489 158806 265613 159988
rect 271447 158807 272571 159989
rect 278364 158811 279488 159993
rect 22005 153992 23129 155174
rect 28963 153993 30087 155175
rect 35883 153992 37007 155174
rect 42848 153993 43972 155175
rect 49806 153994 50930 155176
rect 56723 153998 57847 155180
rect 63688 153999 64812 155181
rect 70646 154000 71770 155182
rect 77563 153998 78687 155180
rect 84528 153999 85652 155181
rect 91486 154000 92610 155182
rect 98304 153979 99428 155161
rect 105269 153980 106393 155162
rect 112227 153981 113351 155163
rect 119147 153980 120271 155162
rect 126112 153981 127236 155163
rect 133070 153982 134194 155164
rect 139987 153986 141111 155168
rect 146952 153987 148076 155169
rect 153910 153988 155034 155170
rect 160827 153986 161951 155168
rect 167792 153987 168916 155169
rect 174750 153988 175874 155170
rect 181555 153981 182679 155163
rect 188520 153982 189644 155164
rect 195478 153983 196602 155165
rect 202398 153982 203522 155164
rect 209363 153983 210487 155165
rect 216321 153984 217445 155166
rect 223238 153988 224362 155170
rect 230077 153983 231201 155165
rect 237042 153984 238166 155166
rect 244000 153985 245124 155167
rect 250917 153989 252041 155171
rect 257809 153972 258933 155154
rect 264774 153973 265898 155155
rect 271732 153974 272856 155156
rect 278649 153978 279773 155160
rect 22076 148732 23200 149914
rect 29034 148733 30158 149915
rect 35954 148732 37078 149914
rect 42919 148733 44043 149915
rect 49877 148734 51001 149916
rect 56794 148738 57918 149920
rect 63759 148739 64883 149921
rect 70717 148740 71841 149922
rect 77634 148738 78758 149920
rect 84599 148739 85723 149921
rect 91557 148740 92681 149922
rect 98375 148719 99499 149901
rect 105340 148720 106464 149902
rect 112298 148721 113422 149903
rect 119218 148720 120342 149902
rect 126183 148721 127307 149903
rect 133141 148722 134265 149904
rect 140058 148726 141182 149908
rect 147023 148727 148147 149909
rect 153981 148728 155105 149910
rect 160898 148726 162022 149908
rect 167863 148727 168987 149909
rect 174821 148728 175945 149910
rect 181626 148721 182750 149903
rect 188591 148722 189715 149904
rect 195549 148723 196673 149905
rect 202469 148722 203593 149904
rect 209434 148723 210558 149905
rect 216392 148724 217516 149906
rect 223309 148728 224433 149910
rect 230148 148723 231272 149905
rect 237113 148724 238237 149906
rect 244071 148725 245195 149907
rect 250988 148729 252112 149911
rect 257880 148712 259004 149894
rect 264845 148713 265969 149895
rect 271803 148714 272927 149896
rect 278720 148718 279844 149900
rect 22005 143258 23129 144440
rect 28963 143259 30087 144441
rect 35883 143258 37007 144440
rect 42848 143259 43972 144441
rect 49806 143260 50930 144442
rect 56723 143264 57847 144446
rect 63688 143265 64812 144447
rect 70646 143266 71770 144448
rect 77563 143264 78687 144446
rect 84528 143265 85652 144447
rect 91486 143266 92610 144448
rect 98304 143245 99428 144427
rect 105269 143246 106393 144428
rect 112227 143247 113351 144429
rect 119147 143246 120271 144428
rect 126112 143247 127236 144429
rect 133070 143248 134194 144430
rect 139987 143252 141111 144434
rect 146952 143253 148076 144435
rect 153910 143254 155034 144436
rect 160827 143252 161951 144434
rect 167792 143253 168916 144435
rect 174750 143254 175874 144436
rect 181555 143247 182679 144429
rect 188520 143248 189644 144430
rect 195478 143249 196602 144431
rect 202398 143248 203522 144430
rect 209363 143249 210487 144431
rect 216321 143250 217445 144432
rect 223238 143254 224362 144436
rect 22147 137146 23271 138328
rect 29105 137147 30229 138329
rect 36025 137146 37149 138328
rect 42990 137147 44114 138329
rect 49948 137148 51072 138330
rect 56865 137152 57989 138334
rect 63830 137153 64954 138335
rect 70788 137154 71912 138336
rect 77705 137152 78829 138334
rect 84670 137153 85794 138335
rect 91628 137154 92752 138336
rect 98446 137133 99570 138315
rect 105411 137134 106535 138316
rect 112369 137135 113493 138317
rect 119289 137134 120413 138316
rect 126254 137135 127378 138317
rect 133212 137136 134336 138318
rect 140129 137140 141253 138322
rect 147094 137141 148218 138323
rect 154052 137142 155176 138324
rect 160969 137140 162093 138322
rect 167934 137141 169058 138323
rect 174892 137142 176016 138324
rect 181697 137135 182821 138317
rect 188662 137136 189786 138318
rect 195620 137137 196744 138319
rect 202540 137136 203664 138318
rect 209505 137137 210629 138319
rect 216463 137138 217587 138320
rect 223380 137142 224504 138324
rect 21937 129272 23061 130454
rect 28895 129273 30019 130455
rect 35815 129272 36939 130454
rect 42780 129273 43904 130455
rect 49738 129274 50862 130456
rect 56655 129278 57779 130460
rect 63620 129279 64744 130461
rect 70578 129280 71702 130462
rect 77495 129278 78619 130460
rect 84460 129279 85584 130461
rect 91418 129280 92542 130462
rect 98236 129259 99360 130441
rect 105201 129260 106325 130442
rect 112159 129261 113283 130443
rect 119079 129260 120203 130442
rect 126044 129261 127168 130443
rect 133002 129262 134126 130444
rect 139919 129266 141043 130448
rect 146884 129267 148008 130449
rect 153842 129268 154966 130450
rect 160759 129266 161883 130448
rect 167724 129267 168848 130449
rect 174682 129268 175806 130450
rect 181487 129261 182611 130443
rect 188452 129262 189576 130444
rect 195410 129263 196534 130445
rect 202330 129262 203454 130444
rect 209295 129263 210419 130445
rect 216253 129264 217377 130446
rect 223170 129268 224294 130450
rect 21454 117956 22578 119138
rect 28412 117957 29536 119139
rect 35332 117956 36456 119138
rect 42297 117957 43421 119139
rect 49255 117958 50379 119140
rect 56172 117962 57296 119144
rect 63137 117963 64261 119145
rect 70095 117964 71219 119146
rect 77012 117962 78136 119144
rect 83977 117963 85101 119145
rect 90935 117964 92059 119146
rect 97753 117943 98877 119125
rect 104718 117944 105842 119126
rect 111676 117945 112800 119127
rect 118596 117944 119720 119126
rect 125561 117945 126685 119127
rect 132519 117946 133643 119128
rect 139436 117950 140560 119132
rect 146401 117951 147525 119133
rect 153359 117952 154483 119134
rect 160276 117950 161400 119132
rect 167241 117951 168365 119133
rect 174199 117952 175323 119134
rect 181004 117945 182128 119127
rect 187969 117946 189093 119128
rect 194927 117947 196051 119129
rect 201847 117946 202971 119128
rect 208812 117947 209936 119129
rect 215770 117948 216894 119130
rect 222687 117952 223811 119134
rect 229652 117953 230776 119135
rect 236610 117954 237734 119136
rect 243527 117952 244651 119134
rect 250492 117953 251616 119135
rect 257450 117954 258574 119136
rect 264590 117954 265714 119136
rect 271548 117955 272672 119137
rect 278684 117945 279808 119127
rect 21659 110004 22783 111186
rect 28617 110005 29741 111187
rect 35537 110004 36661 111186
rect 42502 110005 43626 111187
rect 49460 110006 50584 111188
rect 56377 110010 57501 111192
rect 63342 110011 64466 111193
rect 70300 110012 71424 111194
rect 77217 110010 78341 111192
rect 84182 110011 85306 111193
rect 91140 110012 92264 111194
rect 97958 109991 99082 111173
rect 104923 109992 106047 111174
rect 111881 109993 113005 111175
rect 118801 109992 119925 111174
rect 125766 109993 126890 111175
rect 132724 109994 133848 111176
rect 139641 109998 140765 111180
rect 146606 109999 147730 111181
rect 153564 110000 154688 111182
rect 160481 109998 161605 111180
rect 167446 109999 168570 111181
rect 174404 110000 175528 111182
rect 181209 109993 182333 111175
rect 188174 109994 189298 111176
rect 195132 109995 196256 111177
rect 202052 109994 203176 111176
rect 209017 109995 210141 111177
rect 215975 109996 217099 111178
rect 222892 110000 224016 111182
rect 229857 110001 230981 111183
rect 236815 110002 237939 111184
rect 243732 110000 244856 111182
rect 250697 110001 251821 111183
rect 257655 110002 258779 111184
rect 264795 110002 265919 111184
rect 271753 110003 272877 111185
rect 278889 109993 280013 111175
rect 21659 101778 22783 102960
rect 28617 101779 29741 102961
rect 35537 101778 36661 102960
rect 42502 101779 43626 102961
rect 49460 101780 50584 102962
rect 56377 101784 57501 102966
rect 63342 101785 64466 102967
rect 70300 101786 71424 102968
rect 77217 101784 78341 102966
rect 84182 101785 85306 102967
rect 91140 101786 92264 102968
rect 97958 101765 99082 102947
rect 104923 101766 106047 102948
rect 111881 101767 113005 102949
rect 118801 101766 119925 102948
rect 125766 101767 126890 102949
rect 132724 101768 133848 102950
rect 139641 101772 140765 102954
rect 146606 101773 147730 102955
rect 153564 101774 154688 102956
rect 160481 101772 161605 102954
rect 167446 101773 168570 102955
rect 174404 101774 175528 102956
rect 181209 101767 182333 102949
rect 188174 101768 189298 102950
rect 195132 101769 196256 102951
rect 202052 101768 203176 102950
rect 209017 101769 210141 102951
rect 215975 101770 217099 102952
rect 222892 101774 224016 102956
rect 229857 101775 230981 102957
rect 236815 101776 237939 102958
rect 243732 101774 244856 102956
rect 250697 101775 251821 102957
rect 257655 101776 258779 102958
rect 264795 101776 265919 102958
rect 271753 101777 272877 102959
rect 278889 101767 280013 102949
rect 21454 94374 22578 95556
rect 28412 94375 29536 95557
rect 35332 94374 36456 95556
rect 42297 94375 43421 95557
rect 49255 94376 50379 95558
rect 56172 94380 57296 95562
rect 63137 94381 64261 95563
rect 70095 94382 71219 95564
rect 77012 94380 78136 95562
rect 83977 94381 85101 95563
rect 90935 94382 92059 95564
rect 97753 94361 98877 95543
rect 104718 94362 105842 95544
rect 111676 94363 112800 95545
rect 118596 94362 119720 95544
rect 125561 94363 126685 95545
rect 132519 94364 133643 95546
rect 139436 94368 140560 95550
rect 146401 94369 147525 95551
rect 153359 94370 154483 95552
rect 160276 94368 161400 95550
rect 167241 94369 168365 95551
rect 174199 94370 175323 95552
rect 181004 94363 182128 95545
rect 187969 94364 189093 95546
rect 194927 94365 196051 95547
rect 201847 94364 202971 95546
rect 208812 94365 209936 95547
rect 215770 94366 216894 95548
rect 222687 94370 223811 95552
rect 229652 94371 230776 95553
rect 236610 94372 237734 95554
rect 243527 94370 244651 95552
rect 250492 94371 251616 95553
rect 257450 94372 258574 95554
rect 264590 94372 265714 95554
rect 271548 94373 272672 95555
rect 278684 94363 279808 95545
rect 21180 87244 22304 88426
rect 28138 87245 29262 88427
rect 35058 87244 36182 88426
rect 42023 87245 43147 88427
rect 48981 87246 50105 88428
rect 55898 87250 57022 88432
rect 62863 87251 63987 88433
rect 69821 87252 70945 88434
rect 76738 87250 77862 88432
rect 83703 87251 84827 88433
rect 90661 87252 91785 88434
rect 97479 87231 98603 88413
rect 104444 87232 105568 88414
rect 111402 87233 112526 88415
rect 118322 87232 119446 88414
rect 125287 87233 126411 88415
rect 132245 87234 133369 88416
rect 139162 87238 140286 88420
rect 146127 87239 147251 88421
rect 153085 87240 154209 88422
rect 160002 87238 161126 88420
rect 166967 87239 168091 88421
rect 173925 87240 175049 88422
rect 180730 87233 181854 88415
rect 187695 87234 188819 88416
rect 194653 87235 195777 88417
rect 201573 87234 202697 88416
rect 208538 87235 209662 88417
rect 215496 87236 216620 88418
rect 222413 87240 223537 88422
rect 229378 87241 230502 88423
rect 236336 87242 237460 88424
rect 243253 87240 244377 88422
rect 250218 87241 251342 88423
rect 257176 87242 258300 88424
rect 264316 87242 265440 88424
rect 271274 87243 272398 88425
rect 278410 87233 279534 88415
rect 21288 80831 22412 82013
rect 28246 80832 29370 82014
rect 35166 80831 36290 82013
rect 42131 80832 43255 82014
rect 49089 80833 50213 82015
rect 56006 80837 57130 82019
rect 62971 80838 64095 82020
rect 69929 80839 71053 82021
rect 76846 80837 77970 82019
rect 83811 80838 84935 82020
rect 90769 80839 91893 82021
rect 97587 80818 98711 82000
rect 104552 80819 105676 82001
rect 111510 80820 112634 82002
rect 118430 80819 119554 82001
rect 125395 80820 126519 82002
rect 132353 80821 133477 82003
rect 139270 80825 140394 82007
rect 146235 80826 147359 82008
rect 153193 80827 154317 82009
rect 160110 80825 161234 82007
rect 167075 80826 168199 82008
rect 174033 80827 175157 82009
rect 180838 80820 181962 82002
rect 187803 80821 188927 82003
rect 194761 80822 195885 82004
rect 201681 80821 202805 82003
rect 208646 80822 209770 82004
rect 215604 80823 216728 82005
rect 222521 80827 223645 82009
rect 229486 80828 230610 82010
rect 236444 80829 237568 82011
rect 243361 80827 244485 82009
rect 250326 80828 251450 82010
rect 257284 80829 258408 82011
rect 264424 80829 265548 82011
rect 271382 80830 272506 82012
rect 278518 80820 279642 82002
rect 21154 69651 22278 70833
rect 28112 69652 29236 70834
rect 35032 69651 36156 70833
rect 41997 69652 43121 70834
rect 48955 69653 50079 70835
rect 55872 69657 56996 70839
rect 62837 69658 63961 70840
rect 69795 69659 70919 70841
rect 76712 69657 77836 70839
rect 83677 69658 84801 70840
rect 90635 69659 91759 70841
rect 97453 69638 98577 70820
rect 104418 69639 105542 70821
rect 111376 69640 112500 70822
rect 118296 69639 119420 70821
rect 125261 69640 126385 70822
rect 132219 69641 133343 70823
rect 139136 69645 140260 70827
rect 146101 69646 147225 70828
rect 153059 69647 154183 70829
rect 159976 69645 161100 70827
rect 166941 69646 168065 70828
rect 173899 69647 175023 70829
rect 180704 69640 181828 70822
rect 187669 69641 188793 70823
rect 194627 69642 195751 70824
rect 201547 69641 202671 70823
rect 208512 69642 209636 70824
rect 215470 69643 216594 70825
rect 222387 69647 223511 70829
rect 229352 69648 230476 70830
rect 236310 69649 237434 70831
rect 243227 69647 244351 70829
rect 250192 69648 251316 70830
rect 257150 69649 258274 70831
rect 264290 69649 265414 70831
rect 271248 69650 272372 70832
rect 278384 69640 279508 70822
rect 21119 63411 22243 64593
rect 28077 63412 29201 64594
rect 34997 63411 36121 64593
rect 41962 63412 43086 64594
rect 48920 63413 50044 64595
rect 55837 63417 56961 64599
rect 62802 63418 63926 64600
rect 69760 63419 70884 64601
rect 76677 63417 77801 64599
rect 83642 63418 84766 64600
rect 90600 63419 91724 64601
rect 97418 63398 98542 64580
rect 104383 63399 105507 64581
rect 111341 63400 112465 64582
rect 118261 63399 119385 64581
rect 125226 63400 126350 64582
rect 132184 63401 133308 64583
rect 139101 63405 140225 64587
rect 146066 63406 147190 64588
rect 153024 63407 154148 64589
rect 159941 63405 161065 64587
rect 166906 63406 168030 64588
rect 173864 63407 174988 64589
rect 180669 63400 181793 64582
rect 187634 63401 188758 64583
rect 194592 63402 195716 64584
rect 201512 63401 202636 64583
rect 208477 63402 209601 64584
rect 215435 63403 216559 64585
rect 222352 63407 223476 64589
rect 229317 63408 230441 64590
rect 236275 63409 237399 64591
rect 243192 63407 244316 64589
rect 250157 63408 251281 64590
rect 257115 63409 258239 64591
rect 264255 63409 265379 64591
rect 271213 63410 272337 64592
rect 278349 63400 279473 64582
rect 21084 57694 22208 58876
rect 28042 57695 29166 58877
rect 34962 57694 36086 58876
rect 41927 57695 43051 58877
rect 48885 57696 50009 58878
rect 55802 57700 56926 58882
rect 62767 57701 63891 58883
rect 69725 57702 70849 58884
rect 76642 57700 77766 58882
rect 83607 57701 84731 58883
rect 90565 57702 91689 58884
rect 97383 57681 98507 58863
rect 104348 57682 105472 58864
rect 111306 57683 112430 58865
rect 118226 57682 119350 58864
rect 125191 57683 126315 58865
rect 132149 57684 133273 58866
rect 139066 57688 140190 58870
rect 146031 57689 147155 58871
rect 152989 57690 154113 58872
rect 159906 57688 161030 58870
rect 166871 57689 167995 58871
rect 173829 57690 174953 58872
rect 180634 57683 181758 58865
rect 187599 57684 188723 58866
rect 194557 57685 195681 58867
rect 201477 57684 202601 58866
rect 208442 57685 209566 58867
rect 215400 57686 216524 58868
rect 222317 57690 223441 58872
rect 229282 57691 230406 58873
rect 236240 57692 237364 58874
rect 243157 57690 244281 58872
rect 250122 57691 251246 58873
rect 257080 57692 258204 58874
rect 264220 57692 265344 58874
rect 271178 57693 272302 58875
rect 278314 57683 279438 58865
rect 21015 51489 22139 52671
rect 27973 51490 29097 52672
rect 34893 51489 36017 52671
rect 41858 51490 42982 52672
rect 48816 51491 49940 52673
rect 55733 51495 56857 52677
rect 62698 51496 63822 52678
rect 69656 51497 70780 52679
rect 76573 51495 77697 52677
rect 83538 51496 84662 52678
rect 90496 51497 91620 52679
rect 97314 51476 98438 52658
rect 104279 51477 105403 52659
rect 111237 51478 112361 52660
rect 118157 51477 119281 52659
rect 125122 51478 126246 52660
rect 132080 51479 133204 52661
rect 138997 51483 140121 52665
rect 145962 51484 147086 52666
rect 152920 51485 154044 52667
rect 159837 51483 160961 52665
rect 166802 51484 167926 52666
rect 173760 51485 174884 52667
rect 180565 51478 181689 52660
rect 187530 51479 188654 52661
rect 194488 51480 195612 52662
rect 201408 51479 202532 52661
rect 208373 51480 209497 52662
rect 215331 51481 216455 52663
rect 222248 51485 223372 52667
rect 229213 51486 230337 52668
rect 236171 51487 237295 52669
rect 243088 51485 244212 52667
rect 250053 51486 251177 52668
rect 257011 51487 258135 52669
rect 264151 51487 265275 52669
rect 271109 51488 272233 52670
rect 278245 51478 279369 52660
rect 69368 43639 70492 44821
rect 76285 43637 77409 44819
rect 83250 43638 84374 44820
rect 90208 43639 91332 44821
rect 97026 43618 98150 44800
rect 103991 43619 105115 44801
rect 110949 43620 112073 44802
rect 117869 43619 118993 44801
rect 124834 43620 125958 44802
rect 131792 43621 132916 44803
rect 138709 43625 139833 44807
rect 145674 43626 146798 44808
rect 152632 43627 153756 44809
rect 159549 43625 160673 44807
rect 166514 43626 167638 44808
rect 173472 43627 174596 44809
rect 180277 43620 181401 44802
rect 187242 43621 188366 44803
rect 194200 43622 195324 44804
rect 201120 43621 202244 44803
rect 208085 43622 209209 44804
rect 215043 43623 216167 44805
rect 221960 43627 223084 44809
rect 228925 43628 230049 44810
rect 235883 43629 237007 44811
rect 242800 43627 243924 44809
rect 249765 43628 250889 44810
rect 256723 43629 257847 44811
rect 263863 43629 264987 44811
rect 270821 43630 271945 44812
rect 277957 43620 279081 44802
rect 69368 37345 70492 38527
rect 76285 37343 77409 38525
rect 83250 37344 84374 38526
rect 90208 37345 91332 38527
rect 97026 37324 98150 38506
rect 103991 37325 105115 38507
rect 110949 37326 112073 38508
rect 117869 37325 118993 38507
rect 124834 37326 125958 38508
rect 131792 37327 132916 38509
rect 138709 37331 139833 38513
rect 145674 37332 146798 38514
rect 152632 37333 153756 38515
rect 159549 37331 160673 38513
rect 166514 37332 167638 38514
rect 173472 37333 174596 38515
rect 180277 37326 181401 38508
rect 187242 37327 188366 38509
rect 194200 37328 195324 38510
rect 201120 37327 202244 38509
rect 208085 37328 209209 38510
rect 215043 37329 216167 38511
rect 221960 37333 223084 38515
rect 228925 37334 230049 38516
rect 235883 37335 237007 38517
rect 242800 37333 243924 38515
rect 249765 37334 250889 38516
rect 256723 37335 257847 38517
rect 263863 37335 264987 38517
rect 270821 37336 271945 38518
rect 277957 37326 279081 38508
rect 69368 31051 70492 32233
rect 76285 31049 77409 32231
rect 83250 31050 84374 32232
rect 90208 31051 91332 32233
rect 97026 31030 98150 32212
rect 103991 31031 105115 32213
rect 110949 31032 112073 32214
rect 117869 31031 118993 32213
rect 124834 31032 125958 32214
rect 131792 31033 132916 32215
rect 138709 31037 139833 32219
rect 145674 31038 146798 32220
rect 152632 31039 153756 32221
rect 159549 31037 160673 32219
rect 166514 31038 167638 32220
rect 173472 31039 174596 32221
rect 180277 31032 181401 32214
rect 187242 31033 188366 32215
rect 194200 31034 195324 32216
rect 201120 31033 202244 32215
rect 208085 31034 209209 32216
rect 215043 31035 216167 32217
rect 221960 31039 223084 32221
rect 228925 31040 230049 32222
rect 235883 31041 237007 32223
rect 242800 31039 243924 32221
rect 249765 31040 250889 32222
rect 256723 31041 257847 32223
rect 263863 31041 264987 32223
rect 270821 31042 271945 32224
rect 277957 31032 279081 32214
rect 20743 20487 21867 21669
rect 27701 20488 28825 21670
rect 34621 20487 35745 21669
rect 41586 20488 42710 21670
rect 48544 20489 49668 21671
rect 55461 20493 56585 21675
rect 62426 20494 63550 21676
rect 69384 20495 70508 21677
rect 76301 20493 77425 21675
rect 83266 20494 84390 21676
rect 90224 20495 91348 21677
rect 97042 20474 98166 21656
rect 104007 20475 105131 21657
rect 110965 20476 112089 21658
rect 117885 20475 119009 21657
rect 124850 20476 125974 21658
rect 131808 20477 132932 21659
rect 138725 20481 139849 21663
rect 145690 20482 146814 21664
rect 152648 20483 153772 21665
rect 159565 20481 160689 21663
rect 166530 20482 167654 21664
rect 173488 20483 174612 21665
rect 180293 20476 181417 21658
rect 187258 20477 188382 21659
rect 194216 20478 195340 21660
rect 201136 20477 202260 21659
rect 208101 20478 209225 21660
rect 215059 20479 216183 21661
rect 221976 20483 223100 21665
rect 228941 20484 230065 21666
rect 235899 20485 237023 21667
rect 242816 20483 243940 21665
rect 249781 20484 250905 21666
rect 256739 20485 257863 21667
rect 263879 20485 265003 21667
rect 270837 20486 271961 21668
rect 277973 20476 279097 21658
rect 20727 14809 21851 15991
rect 27685 14810 28809 15992
rect 34605 14809 35729 15991
rect 41570 14810 42694 15992
rect 48528 14811 49652 15993
rect 55445 14815 56569 15997
rect 62410 14816 63534 15998
rect 69368 14817 70492 15999
rect 76285 14815 77409 15997
rect 83250 14816 84374 15998
rect 90208 14817 91332 15999
rect 97026 14796 98150 15978
rect 103991 14797 105115 15979
rect 110949 14798 112073 15980
rect 117869 14797 118993 15979
rect 124834 14798 125958 15980
rect 131792 14799 132916 15981
rect 138709 14803 139833 15985
rect 145674 14804 146798 15986
rect 152632 14805 153756 15987
rect 159549 14803 160673 15985
rect 166514 14804 167638 15986
rect 173472 14805 174596 15987
rect 180277 14798 181401 15980
rect 187242 14799 188366 15981
rect 194200 14800 195324 15982
rect 201120 14799 202244 15981
rect 208085 14800 209209 15982
rect 215043 14801 216167 15983
rect 221960 14805 223084 15987
rect 228925 14806 230049 15988
rect 235883 14807 237007 15989
rect 242800 14805 243924 15987
rect 249765 14806 250889 15988
rect 256723 14807 257847 15989
rect 263863 14807 264987 15989
rect 270821 14808 271945 15990
rect 277957 14798 279081 15980
rect 20727 7716 21851 8898
rect 27685 7717 28809 8899
rect 34605 7716 35729 8898
rect 41570 7717 42694 8899
rect 48528 7718 49652 8900
rect 55445 7722 56569 8904
rect 62410 7723 63534 8905
rect 69368 7724 70492 8906
rect 76285 7722 77409 8904
rect 83250 7723 84374 8905
rect 90208 7724 91332 8906
rect 97026 7703 98150 8885
rect 103991 7704 105115 8886
rect 110949 7705 112073 8887
rect 117869 7704 118993 8886
rect 124834 7705 125958 8887
rect 131792 7706 132916 8888
rect 138709 7710 139833 8892
rect 145674 7711 146798 8893
rect 152632 7712 153756 8894
rect 159549 7710 160673 8892
rect 166514 7711 167638 8893
rect 173472 7712 174596 8894
rect 180277 7705 181401 8887
rect 187242 7706 188366 8888
rect 194200 7707 195324 8889
rect 201120 7706 202244 8888
rect 208085 7707 209209 8889
rect 215043 7708 216167 8890
rect 221960 7712 223084 8894
rect 228925 7713 230049 8895
rect 235883 7714 237007 8896
rect 242800 7712 243924 8894
rect 249765 7713 250889 8895
rect 256723 7714 257847 8896
rect 263863 7714 264987 8896
rect 270821 7715 271945 8897
rect 277957 7705 279081 8887
<< nsubdiffcont >>
rect 26446 264665 26561 264775
rect 23597 264330 23716 264447
<< locali >>
rect 67252 340492 100486 340530
rect 102753 340517 141064 340530
rect 143513 340517 189653 340530
rect 102753 340495 189653 340517
rect 192003 340495 220030 340530
rect 102753 340492 220030 340495
rect 67252 340048 220030 340492
rect 67252 338866 69629 340048
rect 70753 340047 90469 340048
rect 70753 340046 83511 340047
rect 70753 338866 76546 340046
rect 67252 338864 76546 338866
rect 77670 338865 83511 340046
rect 84635 338866 90469 340047
rect 91593 340036 220030 340048
rect 91593 340035 152893 340036
rect 91593 340034 145935 340035
rect 91593 340030 138970 340034
rect 91593 340029 132053 340030
rect 91593 340028 111210 340029
rect 91593 340027 104252 340028
rect 91593 338866 97287 340027
rect 84635 338865 97287 338866
rect 77670 338864 97287 338865
rect 67252 338845 97287 338864
rect 98411 338846 104252 340027
rect 105376 338847 111210 340028
rect 112334 340028 125095 340029
rect 112334 338847 118130 340028
rect 105376 338846 118130 338847
rect 119254 338847 125095 340028
rect 126219 338848 132053 340029
rect 133177 338852 138970 340030
rect 140094 338853 145935 340034
rect 147059 338854 152893 340035
rect 154017 340035 173733 340036
rect 154017 340034 166775 340035
rect 154017 338854 159810 340034
rect 147059 338853 159810 338854
rect 140094 338852 159810 338853
rect 160934 339949 166775 340034
rect 160934 338852 164500 339949
rect 133177 338848 164500 338852
rect 126219 338847 164500 338848
rect 119254 338846 164500 338847
rect 98411 338845 164500 338846
rect 67252 338774 164500 338845
rect 165766 338853 166775 339949
rect 167899 338854 173733 340035
rect 174857 340032 220030 340036
rect 174857 340031 215304 340032
rect 174857 340030 194461 340031
rect 174857 340029 187503 340030
rect 174857 338854 180538 340029
rect 167899 338853 180538 338854
rect 165766 338847 180538 338853
rect 181662 338848 187503 340029
rect 188627 338849 194461 340030
rect 195585 340030 208346 340031
rect 195585 338849 201381 340030
rect 188627 338848 201381 338849
rect 202505 338849 208346 340030
rect 209470 338850 215304 340031
rect 216428 338850 220030 340032
rect 209470 338849 220030 338850
rect 202505 338848 220030 338849
rect 181662 338847 220030 338848
rect 165766 338774 220030 338847
rect 67252 338423 220030 338774
rect 100639 333400 102538 338423
rect 141388 333400 143287 338423
rect 189962 333400 191861 338423
rect 67252 332918 220030 333400
rect 67252 331736 69355 332918
rect 70479 332917 90195 332918
rect 70479 332916 83237 332917
rect 70479 331736 76272 332916
rect 67252 331734 76272 331736
rect 77396 331735 83237 332916
rect 84361 331736 90195 332917
rect 91319 332906 220030 332918
rect 91319 332905 152619 332906
rect 91319 332904 145661 332905
rect 91319 332900 138696 332904
rect 91319 332899 131779 332900
rect 91319 332898 110936 332899
rect 91319 332897 103978 332898
rect 91319 331736 97013 332897
rect 84361 331735 97013 331736
rect 77396 331734 97013 331735
rect 67252 331715 97013 331734
rect 98137 331716 103978 332897
rect 105102 331717 110936 332898
rect 112060 332898 124821 332899
rect 112060 331717 117856 332898
rect 105102 331716 117856 331717
rect 118980 331717 124821 332898
rect 125945 331718 131779 332899
rect 132903 331722 138696 332900
rect 139820 331723 145661 332904
rect 146785 331724 152619 332905
rect 153743 332905 173459 332906
rect 153743 332904 166501 332905
rect 153743 331724 159536 332904
rect 146785 331723 159536 331724
rect 139820 331722 159536 331723
rect 160660 332863 166501 332904
rect 160660 331722 164481 332863
rect 132903 331718 164481 331722
rect 125945 331717 164481 331718
rect 118980 331716 164481 331717
rect 98137 331715 164481 331716
rect 67252 331688 164481 331715
rect 165747 331723 166501 332863
rect 167625 331724 173459 332905
rect 174583 332902 220030 332906
rect 174583 332901 215030 332902
rect 174583 332900 194187 332901
rect 174583 332899 187229 332900
rect 174583 331724 180264 332899
rect 167625 331723 180264 331724
rect 165747 331717 180264 331723
rect 181388 331718 187229 332899
rect 188353 331719 194187 332900
rect 195311 332900 208072 332901
rect 195311 331719 201107 332900
rect 188353 331718 201107 331719
rect 202231 331719 208072 332900
rect 209196 331720 215030 332901
rect 216154 331720 220030 332902
rect 209196 331719 220030 331720
rect 202231 331718 220030 331719
rect 181388 331717 220030 331718
rect 165747 331688 220030 331717
rect 67252 331293 220030 331688
rect 100593 330649 102644 331293
rect 141388 330649 143422 331293
rect 100593 327072 102621 330649
rect 141394 327719 143422 330649
rect 141388 327072 143422 327719
rect 189886 330649 191921 331293
rect 189886 327072 191914 330649
rect 247445 329554 247576 329570
rect 247445 329454 247459 329554
rect 247560 329454 247576 329554
rect 247445 329439 247576 329454
rect 67252 326590 220030 327072
rect 67252 325408 69629 326590
rect 70753 326589 90469 326590
rect 70753 326588 83511 326589
rect 70753 325408 76546 326588
rect 67252 325406 76546 325408
rect 77670 325407 83511 326588
rect 84635 325408 90469 326589
rect 91593 326578 220030 326590
rect 91593 326577 152893 326578
rect 91593 326576 145935 326577
rect 91593 326572 138970 326576
rect 91593 326571 132053 326572
rect 91593 326570 111210 326571
rect 91593 326569 104252 326570
rect 91593 325408 97287 326569
rect 84635 325407 97287 325408
rect 77670 325406 97287 325407
rect 67252 325387 97287 325406
rect 98411 325388 104252 326569
rect 105376 325389 111210 326570
rect 112334 326570 125095 326571
rect 112334 325389 118130 326570
rect 105376 325388 118130 325389
rect 119254 325389 125095 326570
rect 126219 325390 132053 326571
rect 133177 325394 138970 326572
rect 140094 325395 145935 326576
rect 147059 325396 152893 326577
rect 154017 326577 173733 326578
rect 154017 326576 166775 326577
rect 154017 325396 159810 326576
rect 147059 325395 159810 325396
rect 140094 325394 159810 325395
rect 160934 326491 166775 326576
rect 160934 325394 164500 326491
rect 133177 325390 164500 325394
rect 126219 325389 164500 325390
rect 119254 325388 164500 325389
rect 98411 325387 164500 325388
rect 67252 325316 164500 325387
rect 165766 325395 166775 326491
rect 167899 325396 173733 326577
rect 174857 326574 220030 326578
rect 174857 326573 215304 326574
rect 174857 326572 194461 326573
rect 174857 326571 187503 326572
rect 174857 325396 180538 326571
rect 167899 325395 180538 325396
rect 165766 325389 180538 325395
rect 181662 325390 187503 326571
rect 188627 325391 194461 326572
rect 195585 326572 208346 326573
rect 195585 325391 201381 326572
rect 188627 325390 201381 325391
rect 202505 325391 208346 326572
rect 209470 325392 215304 326573
rect 216428 325392 220030 326574
rect 209470 325391 220030 325392
rect 202505 325390 220030 325391
rect 181662 325389 220030 325390
rect 165766 325316 220030 325389
rect 67252 324965 220030 325316
rect 100593 319942 102621 324965
rect 141388 319942 143422 324965
rect 189886 319942 191914 324965
rect 248420 324185 248457 324380
rect 248417 322901 248457 324185
rect 248907 323928 248944 324430
rect 248903 322951 248944 323928
rect 249397 323723 249434 324407
rect 248417 322751 248454 322901
rect 243780 322749 248454 322751
rect 243707 322706 248454 322749
rect 243707 322691 248438 322706
rect 67252 319460 220030 319942
rect 67252 318278 69355 319460
rect 70479 319459 90195 319460
rect 70479 319458 83237 319459
rect 70479 318278 76272 319458
rect 67252 318276 76272 318278
rect 77396 318277 83237 319458
rect 84361 318278 90195 319459
rect 91319 319448 220030 319460
rect 91319 319447 152619 319448
rect 91319 319446 145661 319447
rect 91319 319442 138696 319446
rect 91319 319441 131779 319442
rect 91319 319440 110936 319441
rect 91319 319439 103978 319440
rect 91319 318278 97013 319439
rect 84361 318277 97013 318278
rect 77396 318276 97013 318277
rect 67252 318257 97013 318276
rect 98137 318258 103978 319439
rect 105102 318259 110936 319440
rect 112060 319440 124821 319441
rect 112060 318259 117856 319440
rect 105102 318258 117856 318259
rect 118980 318259 124821 319440
rect 125945 318260 131779 319441
rect 132903 318264 138696 319442
rect 139820 318265 145661 319446
rect 146785 318266 152619 319447
rect 153743 319447 173459 319448
rect 153743 319446 166501 319447
rect 153743 318266 159536 319446
rect 146785 318265 159536 318266
rect 139820 318264 159536 318265
rect 160660 319405 166501 319446
rect 160660 318264 164481 319405
rect 132903 318260 164481 318264
rect 125945 318259 164481 318260
rect 118980 318258 164481 318259
rect 98137 318257 164481 318258
rect 67252 318230 164481 318257
rect 165747 318265 166501 319405
rect 167625 318266 173459 319447
rect 174583 319444 220030 319448
rect 174583 319443 215030 319444
rect 174583 319442 194187 319443
rect 174583 319441 187229 319442
rect 174583 318266 180264 319441
rect 167625 318265 180264 318266
rect 165747 318259 180264 318265
rect 181388 318260 187229 319441
rect 188353 318261 194187 319442
rect 195311 319442 208072 319443
rect 195311 318261 201107 319442
rect 188353 318260 201107 318261
rect 202231 318261 208072 319442
rect 209196 318262 215030 319443
rect 216154 318262 220030 319444
rect 209196 318261 220030 318262
rect 202231 318260 220030 318261
rect 181388 318259 220030 318260
rect 165747 318230 220030 318259
rect 67252 317835 220030 318230
rect 100593 317191 102644 317835
rect 141388 317191 143422 317835
rect 25883 316944 25997 316962
rect 25883 316894 25928 316944
rect 25978 316894 25997 316944
rect 25883 316882 25997 316894
rect 25892 316743 26006 316761
rect 25892 316693 25937 316743
rect 25987 316693 26006 316743
rect 25892 316681 26006 316693
rect 25877 316054 25991 316072
rect 25877 316004 25922 316054
rect 25972 316004 25991 316054
rect 25877 315992 25991 316004
rect 25883 315703 25997 315721
rect 25883 315653 25928 315703
rect 25978 315653 25997 315703
rect 25883 315641 25997 315653
rect 100593 313001 102621 317191
rect 141394 313182 143422 317191
rect 189886 317191 191921 317835
rect 100645 312811 102544 313001
rect 141394 312811 143293 313182
rect 189886 313114 191914 317191
rect 189968 312811 191867 313114
rect 17908 312798 30608 312811
rect 33967 312798 58547 312811
rect 61906 312798 220036 312811
rect 17908 312329 220036 312798
rect 17908 312328 69635 312329
rect 17908 312327 62677 312328
rect 17908 312323 55712 312327
rect 17908 312322 48795 312323
rect 17908 312321 27952 312322
rect 17908 311139 20994 312321
rect 22118 311140 27952 312321
rect 29076 312321 41837 312322
rect 29076 311140 34872 312321
rect 22118 311139 34872 311140
rect 35996 311140 41837 312321
rect 42961 311141 48795 312322
rect 49919 311145 55712 312323
rect 56836 311146 62677 312327
rect 63801 311147 69635 312328
rect 70759 312328 90475 312329
rect 70759 312327 83517 312328
rect 70759 311147 76552 312327
rect 63801 311146 76552 311147
rect 56836 311145 76552 311146
rect 77676 311146 83517 312327
rect 84641 311147 90475 312328
rect 91599 312317 220036 312329
rect 91599 312316 152899 312317
rect 91599 312315 145941 312316
rect 91599 312311 138976 312315
rect 91599 312310 132059 312311
rect 91599 312309 111216 312310
rect 91599 312308 104258 312309
rect 91599 311147 97293 312308
rect 84641 311146 97293 311147
rect 77676 311145 97293 311146
rect 49919 311141 97293 311145
rect 42961 311140 97293 311141
rect 35996 311139 97293 311140
rect 17908 311126 97293 311139
rect 98417 311127 104258 312308
rect 105382 311128 111216 312309
rect 112340 312309 125101 312310
rect 112340 311128 118136 312309
rect 105382 311127 118136 311128
rect 119260 311128 125101 312309
rect 126225 311129 132059 312310
rect 133183 311133 138976 312311
rect 140100 311134 145941 312315
rect 147065 311135 152899 312316
rect 154023 312316 173739 312317
rect 154023 312315 166781 312316
rect 154023 311135 159816 312315
rect 147065 311134 159816 311135
rect 140100 311133 159816 311134
rect 160940 312230 166781 312315
rect 160940 311133 164506 312230
rect 133183 311129 164506 311133
rect 126225 311128 164506 311129
rect 119260 311127 164506 311128
rect 98417 311126 164506 311127
rect 17908 311055 164506 311126
rect 165772 311134 166781 312230
rect 167905 311135 173739 312316
rect 174863 312313 220036 312317
rect 174863 312312 215310 312313
rect 174863 312311 194467 312312
rect 174863 312310 187509 312311
rect 174863 311135 180544 312310
rect 167905 311134 180544 311135
rect 165772 311128 180544 311134
rect 181668 311129 187509 312310
rect 188633 311130 194467 312311
rect 195591 312311 208352 312312
rect 195591 311130 201387 312311
rect 188633 311129 201387 311130
rect 202511 311130 208352 312311
rect 209476 311131 215310 312312
rect 216434 311131 220036 312313
rect 209476 311130 220036 311131
rect 202511 311129 220036 311130
rect 181668 311128 220036 311129
rect 165772 311055 220036 311128
rect 17908 310704 220036 311055
rect 30923 305681 32822 310704
rect 58769 305681 60668 310704
rect 100645 305681 102544 310704
rect 141394 305681 143293 310704
rect 189968 305681 191867 310704
rect 243707 306229 243802 322691
rect 248903 322469 248940 322951
rect 249397 322928 249436 323723
rect 249886 323493 249923 324432
rect 244003 322465 248940 322469
rect 243957 322449 248940 322465
rect 243957 322409 248935 322449
rect 243957 308695 244034 322409
rect 249399 322246 249436 322928
rect 249885 322953 249923 323493
rect 244260 322241 249440 322246
rect 244198 322186 249440 322241
rect 244198 311097 244284 322186
rect 244431 322041 244517 322052
rect 249885 322041 249922 322953
rect 244431 322014 249922 322041
rect 244431 321972 249919 322014
rect 244431 313581 244517 321972
rect 250376 321835 250413 324434
rect 244696 321819 250424 321835
rect 244655 321775 250424 321819
rect 244655 315946 244724 321775
rect 250970 321604 251007 324430
rect 244853 321527 251024 321604
rect 244853 318395 244939 321527
rect 244851 318388 244942 318395
rect 244851 318306 244859 318388
rect 244934 318306 244942 318388
rect 244851 318296 244942 318306
rect 245914 318392 246005 318400
rect 245914 318310 245922 318392
rect 245997 318310 246005 318392
rect 245914 318300 246005 318310
rect 244853 318184 244939 318296
rect 244645 315938 244736 315946
rect 244645 315856 244653 315938
rect 244728 315856 244736 315938
rect 244645 315846 244736 315856
rect 245820 315933 245911 315941
rect 245820 315851 245828 315933
rect 245903 315851 245911 315933
rect 244655 315798 244724 315846
rect 245820 315841 245911 315851
rect 244427 313573 244518 313581
rect 244427 313491 244435 313573
rect 244510 313491 244518 313573
rect 244427 313481 244518 313491
rect 245754 313549 245845 313557
rect 244431 313394 244517 313481
rect 245754 313467 245762 313549
rect 245837 313467 245845 313549
rect 245754 313457 245845 313467
rect 244195 311089 244286 311097
rect 244195 311007 244203 311089
rect 244278 311007 244286 311089
rect 244195 310997 244286 311007
rect 245669 311086 245760 311094
rect 245669 311004 245677 311086
rect 245752 311004 245760 311086
rect 244198 310965 244284 310997
rect 245669 310994 245760 311004
rect 245594 308710 245685 308718
rect 243953 308687 244044 308695
rect 243953 308605 243961 308687
rect 244036 308605 244044 308687
rect 245594 308628 245602 308710
rect 245677 308628 245685 308710
rect 245594 308618 245685 308628
rect 243953 308595 244044 308605
rect 243957 308459 244034 308595
rect 243708 306147 243716 306229
rect 243791 306147 243802 306229
rect 243708 306129 243802 306147
rect 245514 306235 245605 306243
rect 245514 306153 245522 306235
rect 245597 306153 245605 306235
rect 245514 306143 245605 306153
rect 243707 305917 243802 306129
rect 17908 305199 220036 305681
rect 17908 305198 69361 305199
rect 17908 305197 62403 305198
rect 17908 305193 55438 305197
rect 17908 305192 48521 305193
rect 17908 305191 27678 305192
rect 17908 304009 20720 305191
rect 21844 304010 27678 305191
rect 28802 305191 41563 305192
rect 28802 304010 34598 305191
rect 21844 304009 34598 304010
rect 35722 304010 41563 305191
rect 42687 304011 48521 305192
rect 49645 304015 55438 305193
rect 56562 304016 62403 305197
rect 63527 304017 69361 305198
rect 70485 305198 90201 305199
rect 70485 305197 83243 305198
rect 70485 304017 76278 305197
rect 63527 304016 76278 304017
rect 56562 304015 76278 304016
rect 77402 304016 83243 305197
rect 84367 304017 90201 305198
rect 91325 305187 220036 305199
rect 91325 305186 152625 305187
rect 91325 305185 145667 305186
rect 91325 305181 138702 305185
rect 91325 305180 131785 305181
rect 91325 305179 110942 305180
rect 91325 305178 103984 305179
rect 91325 304017 97019 305178
rect 84367 304016 97019 304017
rect 77402 304015 97019 304016
rect 49645 304011 97019 304015
rect 42687 304010 97019 304011
rect 35722 304009 97019 304010
rect 17908 303996 97019 304009
rect 98143 303997 103984 305178
rect 105108 303998 110942 305179
rect 112066 305179 124827 305180
rect 112066 303998 117862 305179
rect 105108 303997 117862 303998
rect 118986 303998 124827 305179
rect 125951 303999 131785 305180
rect 132909 304003 138702 305181
rect 139826 304004 145667 305185
rect 146791 304005 152625 305186
rect 153749 305186 173465 305187
rect 153749 305185 166507 305186
rect 153749 304005 159542 305185
rect 146791 304004 159542 304005
rect 139826 304003 159542 304004
rect 160666 305144 166507 305185
rect 160666 304003 164487 305144
rect 132909 303999 164487 304003
rect 125951 303998 164487 303999
rect 118986 303997 164487 303998
rect 98143 303996 164487 303997
rect 17908 303969 164487 303996
rect 165753 304004 166507 305144
rect 167631 304005 173465 305186
rect 174589 305183 220036 305187
rect 174589 305182 215036 305183
rect 174589 305181 194193 305182
rect 174589 305180 187235 305181
rect 174589 304005 180270 305180
rect 167631 304004 180270 304005
rect 165753 303998 180270 304004
rect 181394 303999 187235 305180
rect 188359 304000 194193 305181
rect 195317 305181 208078 305182
rect 195317 304000 201113 305181
rect 188359 303999 201113 304000
rect 202237 304000 208078 305181
rect 209202 304001 215036 305182
rect 216160 304001 220036 305183
rect 209202 304000 220036 304001
rect 202237 303999 220036 304000
rect 181394 303998 220036 303999
rect 165753 303969 220036 303998
rect 17908 303574 220036 303969
rect 30923 302753 32911 303574
rect 58769 302753 60786 303574
rect 100645 302753 102650 303574
rect 141394 302753 143412 303574
rect 30947 296598 32911 302753
rect 58822 296839 60786 302753
rect 31012 296452 32911 296598
rect 58858 296452 60757 296839
rect 100686 296667 102650 302753
rect 141448 296736 143412 302753
rect 189963 297099 191927 303574
rect 189963 296770 191956 297099
rect 100734 296452 102633 296667
rect 141483 296452 143382 296736
rect 190057 296452 191956 296770
rect 232340 296452 234239 297099
rect 267192 296452 269091 297099
rect 17997 296414 279970 296452
rect 17997 295970 281013 296414
rect 17997 295969 69724 295970
rect 17997 295968 62766 295969
rect 17997 295964 55801 295968
rect 17997 295963 48884 295964
rect 17997 295962 28041 295963
rect 17997 294780 21083 295962
rect 22207 294781 28041 295962
rect 29165 295962 41926 295963
rect 29165 294781 34961 295962
rect 22207 294780 34961 294781
rect 36085 294781 41926 295962
rect 43050 294782 48884 295963
rect 50008 294786 55801 295964
rect 56925 294787 62766 295968
rect 63890 294788 69724 295969
rect 70848 295969 90564 295970
rect 70848 295968 83606 295969
rect 70848 294788 76641 295968
rect 63890 294787 76641 294788
rect 56925 294786 76641 294787
rect 77765 294787 83606 295968
rect 84730 294788 90564 295969
rect 91688 295961 281013 295970
rect 91688 295960 271177 295961
rect 91688 295959 236239 295960
rect 91688 295958 229281 295959
rect 91688 295957 152988 295958
rect 91688 295956 146030 295957
rect 91688 295952 139065 295956
rect 91688 295951 132148 295952
rect 91688 295950 111305 295951
rect 91688 295949 104347 295950
rect 91688 294788 97382 295949
rect 84730 294787 97382 294788
rect 77765 294786 97382 294787
rect 50008 294782 97382 294786
rect 43050 294781 97382 294782
rect 36085 294780 97382 294781
rect 17997 294767 97382 294780
rect 98506 294768 104347 295949
rect 105471 294769 111305 295950
rect 112429 295950 125190 295951
rect 112429 294769 118225 295950
rect 105471 294768 118225 294769
rect 119349 294769 125190 295950
rect 126314 294770 132148 295951
rect 133272 294774 139065 295952
rect 140189 294775 146030 295956
rect 147154 294776 152988 295957
rect 154112 295957 173828 295958
rect 154112 295956 166870 295957
rect 154112 294776 159905 295956
rect 147154 294775 159905 294776
rect 140189 294774 159905 294775
rect 161029 295871 166870 295956
rect 161029 294774 164595 295871
rect 133272 294770 164595 294774
rect 126314 294769 164595 294770
rect 119349 294768 164595 294769
rect 98506 294767 164595 294768
rect 17997 294696 164595 294767
rect 165861 294775 166870 295871
rect 167994 294776 173828 295957
rect 174952 295954 222316 295958
rect 174952 295953 215399 295954
rect 174952 295952 194556 295953
rect 174952 295951 187598 295952
rect 174952 294776 180633 295951
rect 167994 294775 180633 294776
rect 165861 294769 180633 294775
rect 181757 294770 187598 295951
rect 188722 294771 194556 295952
rect 195680 295952 208441 295953
rect 195680 294771 201476 295952
rect 188722 294770 201476 294771
rect 202600 294771 208441 295952
rect 209565 294772 215399 295953
rect 216523 294776 222316 295954
rect 223440 294777 229281 295958
rect 230405 294778 236239 295959
rect 237363 295959 257079 295960
rect 237363 295958 250121 295959
rect 237363 294778 243156 295958
rect 230405 294777 243156 294778
rect 223440 294776 243156 294777
rect 244280 294777 250121 295958
rect 251245 294778 257079 295959
rect 258203 294778 264219 295960
rect 265343 294779 271177 295960
rect 272301 295951 281013 295961
rect 272301 294779 278313 295951
rect 265343 294778 278313 294779
rect 251245 294777 278313 294778
rect 244280 294776 278313 294777
rect 216523 294772 278313 294776
rect 209565 294771 278313 294772
rect 202600 294770 278313 294771
rect 181757 294769 278313 294770
rect 279437 294769 281013 295951
rect 165861 294696 281013 294769
rect 17997 294364 281013 294696
rect 17997 294345 279970 294364
rect 31012 289322 32911 294345
rect 58858 289322 60757 294345
rect 100734 289322 102633 294345
rect 141483 289322 143382 294345
rect 190057 289322 191956 294345
rect 232340 289322 234239 294345
rect 267192 289322 269091 294345
rect 17997 289284 279696 289322
rect 17997 288840 280739 289284
rect 17997 288839 69450 288840
rect 17997 288838 62492 288839
rect 17997 288834 55527 288838
rect 17997 288833 48610 288834
rect 17997 288832 27767 288833
rect 17997 287650 20809 288832
rect 21933 287651 27767 288832
rect 28891 288832 41652 288833
rect 28891 287651 34687 288832
rect 21933 287650 34687 287651
rect 35811 287651 41652 288832
rect 42776 287652 48610 288833
rect 49734 287656 55527 288834
rect 56651 287657 62492 288838
rect 63616 287658 69450 288839
rect 70574 288839 90290 288840
rect 70574 288838 83332 288839
rect 70574 287658 76367 288838
rect 63616 287657 76367 287658
rect 56651 287656 76367 287657
rect 77491 287657 83332 288838
rect 84456 287658 90290 288839
rect 91414 288831 280739 288840
rect 91414 288830 270903 288831
rect 91414 288829 235965 288830
rect 91414 288828 229007 288829
rect 91414 288827 152714 288828
rect 91414 288826 145756 288827
rect 91414 288822 138791 288826
rect 91414 288821 131874 288822
rect 91414 288820 111031 288821
rect 91414 288819 104073 288820
rect 91414 287658 97108 288819
rect 84456 287657 97108 287658
rect 77491 287656 97108 287657
rect 49734 287652 97108 287656
rect 42776 287651 97108 287652
rect 35811 287650 97108 287651
rect 17997 287637 97108 287650
rect 98232 287638 104073 288819
rect 105197 287639 111031 288820
rect 112155 288820 124916 288821
rect 112155 287639 117951 288820
rect 105197 287638 117951 287639
rect 119075 287639 124916 288820
rect 126040 287640 131874 288821
rect 132998 287644 138791 288822
rect 139915 287645 145756 288826
rect 146880 287646 152714 288827
rect 153838 288827 173554 288828
rect 153838 288826 166596 288827
rect 153838 287646 159631 288826
rect 146880 287645 159631 287646
rect 139915 287644 159631 287645
rect 160755 288785 166596 288826
rect 160755 287644 164576 288785
rect 132998 287640 164576 287644
rect 126040 287639 164576 287640
rect 119075 287638 164576 287639
rect 98232 287637 164576 287638
rect 17997 287610 164576 287637
rect 165842 287645 166596 288785
rect 167720 287646 173554 288827
rect 174678 288824 222042 288828
rect 174678 288823 215125 288824
rect 174678 288822 194282 288823
rect 174678 288821 187324 288822
rect 174678 287646 180359 288821
rect 167720 287645 180359 287646
rect 165842 287639 180359 287645
rect 181483 287640 187324 288821
rect 188448 287641 194282 288822
rect 195406 288822 208167 288823
rect 195406 287641 201202 288822
rect 188448 287640 201202 287641
rect 202326 287641 208167 288822
rect 209291 287642 215125 288823
rect 216249 287646 222042 288824
rect 223166 287647 229007 288828
rect 230131 287648 235965 288829
rect 237089 288829 256805 288830
rect 237089 288828 249847 288829
rect 237089 287648 242882 288828
rect 230131 287647 242882 287648
rect 223166 287646 242882 287647
rect 244006 287647 249847 288828
rect 250971 287648 256805 288829
rect 257929 287648 263945 288830
rect 265069 287649 270903 288830
rect 272027 288821 280739 288831
rect 272027 287649 278039 288821
rect 265069 287648 278039 287649
rect 250971 287647 278039 287648
rect 244006 287646 278039 287647
rect 216249 287642 278039 287646
rect 209291 287641 278039 287642
rect 202326 287640 278039 287641
rect 181483 287639 278039 287640
rect 279163 287639 280739 288821
rect 165842 287610 280739 287639
rect 17997 287234 280739 287610
rect 17997 287215 279696 287234
rect 31012 282909 32911 287215
rect 58858 282909 60757 287215
rect 100734 282909 102633 287215
rect 141483 282909 143382 287215
rect 190057 282909 191956 287215
rect 232340 282909 234239 287215
rect 267192 282909 269091 287215
rect 17997 282871 279804 282909
rect 17997 282427 280847 282871
rect 17997 282426 69558 282427
rect 17997 282425 62600 282426
rect 17997 282421 55635 282425
rect 17997 282420 48718 282421
rect 17997 282419 27875 282420
rect 17997 281237 20917 282419
rect 22041 281238 27875 282419
rect 28999 282419 41760 282420
rect 28999 281238 34795 282419
rect 22041 281237 34795 281238
rect 35919 281238 41760 282419
rect 42884 281239 48718 282420
rect 49842 281243 55635 282421
rect 56759 281244 62600 282425
rect 63724 281245 69558 282426
rect 70682 282426 90398 282427
rect 70682 282425 83440 282426
rect 70682 281245 76475 282425
rect 63724 281244 76475 281245
rect 56759 281243 76475 281244
rect 77599 281244 83440 282425
rect 84564 281245 90398 282426
rect 91522 282418 280847 282427
rect 91522 282417 271011 282418
rect 91522 282416 236073 282417
rect 91522 282415 229115 282416
rect 91522 282414 152822 282415
rect 91522 282413 145864 282414
rect 91522 282409 138899 282413
rect 91522 282408 131982 282409
rect 91522 282407 111139 282408
rect 91522 282406 104181 282407
rect 91522 281245 97216 282406
rect 84564 281244 97216 281245
rect 77599 281243 97216 281244
rect 49842 281239 97216 281243
rect 42884 281238 97216 281239
rect 35919 281237 97216 281238
rect 17997 281224 97216 281237
rect 98340 281225 104181 282406
rect 105305 281226 111139 282407
rect 112263 282407 125024 282408
rect 112263 281226 118059 282407
rect 105305 281225 118059 281226
rect 119183 281226 125024 282407
rect 126148 281227 131982 282408
rect 133106 281231 138899 282409
rect 140023 281232 145864 282413
rect 146988 281233 152822 282414
rect 153946 282414 173662 282415
rect 153946 282413 166704 282414
rect 153946 281233 159739 282413
rect 146988 281232 159739 281233
rect 140023 281231 159739 281232
rect 160863 282383 166704 282413
rect 160863 281231 164539 282383
rect 133106 281227 164539 281231
rect 126148 281226 164539 281227
rect 119183 281225 164539 281226
rect 98340 281224 164539 281225
rect 17997 281208 164539 281224
rect 165805 281232 166704 282383
rect 167828 281233 173662 282414
rect 174786 282411 222150 282415
rect 174786 282410 215233 282411
rect 174786 282409 194390 282410
rect 174786 282408 187432 282409
rect 174786 281233 180467 282408
rect 167828 281232 180467 281233
rect 165805 281226 180467 281232
rect 181591 281227 187432 282408
rect 188556 281228 194390 282409
rect 195514 282409 208275 282410
rect 195514 281228 201310 282409
rect 188556 281227 201310 281228
rect 202434 281228 208275 282409
rect 209399 281229 215233 282410
rect 216357 281233 222150 282411
rect 223274 281234 229115 282415
rect 230239 281235 236073 282416
rect 237197 282416 256913 282417
rect 237197 282415 249955 282416
rect 237197 281235 242990 282415
rect 230239 281234 242990 281235
rect 223274 281233 242990 281234
rect 244114 281234 249955 282415
rect 251079 281235 256913 282416
rect 258037 281235 264053 282417
rect 265177 281236 271011 282417
rect 272135 282408 280847 282418
rect 272135 281236 278147 282408
rect 265177 281235 278147 281236
rect 251079 281234 278147 281235
rect 244114 281233 278147 281234
rect 216357 281229 278147 281233
rect 209399 281228 278147 281229
rect 202434 281227 278147 281228
rect 181591 281226 278147 281227
rect 279271 281226 280847 282408
rect 165805 281208 280847 281226
rect 17997 280821 280847 281208
rect 17997 280802 279804 280821
rect 30688 280739 32778 280802
rect 58459 280781 60549 280802
rect 100327 274044 102704 280802
rect 141089 274044 143466 280802
rect 189461 274691 191838 280802
rect 231966 280229 234056 280802
rect 267079 280229 269169 280802
rect 189461 274044 192007 274691
rect 66323 273562 226094 274044
rect 66323 272380 69775 273562
rect 70899 273561 90615 273562
rect 70899 273560 83657 273561
rect 70899 272380 76692 273560
rect 66323 272378 76692 272380
rect 77816 272379 83657 273560
rect 84781 272380 90615 273561
rect 91739 273550 226094 273562
rect 91739 273549 153039 273550
rect 91739 273548 146081 273549
rect 91739 273544 139116 273548
rect 91739 273543 132199 273544
rect 91739 273542 111356 273543
rect 91739 273541 104398 273542
rect 91739 272380 97433 273541
rect 84781 272379 97433 272380
rect 77816 272378 97433 272379
rect 66323 272359 97433 272378
rect 98557 272360 104398 273541
rect 105522 272361 111356 273542
rect 112480 273542 125241 273543
rect 112480 272361 118276 273542
rect 105522 272360 118276 272361
rect 119400 272361 125241 273542
rect 126365 272362 132199 273543
rect 133323 272366 139116 273544
rect 140240 272367 146081 273548
rect 147205 272368 153039 273549
rect 154163 273549 173879 273550
rect 154163 273548 166921 273549
rect 154163 272368 159956 273548
rect 147205 272367 159956 272368
rect 140240 272366 159956 272367
rect 161080 273463 166921 273548
rect 161080 272366 164646 273463
rect 133323 272362 164646 272366
rect 126365 272361 164646 272362
rect 119400 272360 164646 272361
rect 98557 272359 164646 272360
rect 66323 272288 164646 272359
rect 165912 272367 166921 273463
rect 168045 272368 173879 273549
rect 175003 273546 222367 273550
rect 175003 273545 215450 273546
rect 175003 273544 194607 273545
rect 175003 273543 187649 273544
rect 175003 272368 180684 273543
rect 168045 272367 180684 272368
rect 165912 272361 180684 272367
rect 181808 272362 187649 273543
rect 188773 272363 194607 273544
rect 195731 273544 208492 273545
rect 195731 272363 201527 273544
rect 188773 272362 201527 272363
rect 202651 272363 208492 273544
rect 209616 272364 215450 273545
rect 216574 272368 222367 273546
rect 223491 272368 226094 273550
rect 216574 272364 226094 272368
rect 209616 272363 226094 272364
rect 202651 272362 226094 272363
rect 181808 272361 226094 272362
rect 165912 272288 226094 272361
rect 66323 271937 226094 272288
rect 29771 266041 30276 267017
rect 32451 266041 32956 267017
rect 35370 266058 35875 267034
rect 37561 266050 38066 267026
rect 39915 266067 40420 267043
rect 42432 266041 42937 267017
rect 44854 266041 45359 267017
rect 47097 266058 47602 267034
rect 49271 266041 49776 267017
rect 51291 265562 51784 267050
rect 53354 265587 53847 267075
rect 55794 265544 56287 267032
rect 58216 265570 58709 267058
rect 100785 266914 102684 271937
rect 141534 266914 143433 271937
rect 190108 266914 192007 271937
rect 66323 266432 226094 266914
rect 66323 265250 69501 266432
rect 70625 266431 90341 266432
rect 70625 266430 83383 266431
rect 70625 265250 76418 266430
rect 66323 265248 76418 265250
rect 77542 265249 83383 266430
rect 84507 265250 90341 266431
rect 91465 266420 226094 266432
rect 91465 266419 152765 266420
rect 91465 266418 145807 266419
rect 91465 266414 138842 266418
rect 91465 266413 131925 266414
rect 91465 266412 111082 266413
rect 91465 266411 104124 266412
rect 91465 265250 97159 266411
rect 84507 265249 97159 265250
rect 77542 265248 97159 265249
rect 66323 265229 97159 265248
rect 98283 265230 104124 266411
rect 105248 265231 111082 266412
rect 112206 266412 124967 266413
rect 112206 265231 118002 266412
rect 105248 265230 118002 265231
rect 119126 265231 124967 266412
rect 126091 265232 131925 266413
rect 133049 265236 138842 266414
rect 139966 265237 145807 266418
rect 146931 265238 152765 266419
rect 153889 266419 173605 266420
rect 153889 266418 166647 266419
rect 153889 265238 159682 266418
rect 146931 265237 159682 265238
rect 139966 265236 159682 265237
rect 160806 266377 166647 266418
rect 160806 265236 164627 266377
rect 133049 265232 164627 265236
rect 126091 265231 164627 265232
rect 119126 265230 164627 265231
rect 98283 265229 164627 265230
rect 66323 265202 164627 265229
rect 165893 265237 166647 266377
rect 167771 265238 173605 266419
rect 174729 266416 222093 266420
rect 174729 266415 215176 266416
rect 174729 266414 194333 266415
rect 174729 266413 187375 266414
rect 174729 265238 180410 266413
rect 167771 265237 180410 265238
rect 165893 265231 180410 265237
rect 181534 265232 187375 266413
rect 188499 265233 194333 266414
rect 195457 266414 208218 266415
rect 195457 265233 201253 266414
rect 188499 265232 201253 265233
rect 202377 265233 208218 266414
rect 209342 265234 215176 266415
rect 216300 265238 222093 266416
rect 223217 265238 226094 266420
rect 216300 265234 226094 265238
rect 209342 265233 226094 265234
rect 202377 265232 226094 265233
rect 181534 265231 226094 265232
rect 165893 265202 226094 265231
rect 66323 264807 226094 265202
rect 266009 265300 266147 265320
rect 266009 265202 266024 265300
rect 266126 265202 266147 265300
rect 266009 265179 266147 265202
rect 26436 264775 26571 264785
rect 26436 264665 26446 264775
rect 26561 264665 26571 264775
rect 26436 264660 26571 264665
rect 23581 264447 23730 264462
rect 23581 264330 23597 264447
rect 23716 264330 23730 264447
rect 23581 264315 23730 264330
rect 29735 263623 30347 264617
rect 32446 263589 33058 264583
rect 35412 263614 36024 264608
rect 37579 263580 38191 264574
rect 39823 263623 40435 264617
rect 42329 263623 42941 264617
rect 44870 263614 45482 264608
rect 47105 263606 47717 264600
rect 49255 263623 49867 264617
rect 26041 262939 28333 263156
rect 51473 263104 51966 264592
rect 53479 263130 53972 264618
rect 55850 263130 56343 264618
rect 58289 263121 58782 264609
rect 100785 260501 102684 264807
rect 141534 260501 143433 264807
rect 190108 260501 192007 264807
rect 265929 262942 266067 262962
rect 265929 262844 265944 262942
rect 266046 262844 266067 262942
rect 265929 262821 266067 262844
rect 66323 260019 226094 260501
rect 66323 258837 69609 260019
rect 70733 260018 90449 260019
rect 70733 260017 83491 260018
rect 70733 258837 76526 260017
rect 66323 258835 76526 258837
rect 77650 258836 83491 260017
rect 84615 258837 90449 260018
rect 91573 260007 226094 260019
rect 91573 260006 152873 260007
rect 91573 260005 145915 260006
rect 91573 260001 138950 260005
rect 91573 260000 132033 260001
rect 91573 259999 111190 260000
rect 91573 259998 104232 259999
rect 91573 258837 97267 259998
rect 84615 258836 97267 258837
rect 77650 258835 97267 258836
rect 66323 258816 97267 258835
rect 98391 258817 104232 259998
rect 105356 258818 111190 259999
rect 112314 259999 125075 260000
rect 112314 258818 118110 259999
rect 105356 258817 118110 258818
rect 119234 258818 125075 259999
rect 126199 258819 132033 260000
rect 133157 258823 138950 260001
rect 140074 258824 145915 260005
rect 147039 258825 152873 260006
rect 153997 260006 173713 260007
rect 153997 260005 166755 260006
rect 153997 258825 159790 260005
rect 147039 258824 159790 258825
rect 140074 258823 159790 258824
rect 160914 259975 166755 260005
rect 160914 258823 164590 259975
rect 133157 258819 164590 258823
rect 126199 258818 164590 258819
rect 119234 258817 164590 258818
rect 98391 258816 164590 258817
rect 66323 258800 164590 258816
rect 165856 258824 166755 259975
rect 167879 258825 173713 260006
rect 174837 260003 222201 260007
rect 174837 260002 215284 260003
rect 174837 260001 194441 260002
rect 174837 260000 187483 260001
rect 174837 258825 180518 260000
rect 167879 258824 180518 258825
rect 165856 258818 180518 258824
rect 181642 258819 187483 260000
rect 188607 258820 194441 260001
rect 195565 260001 208326 260002
rect 195565 258820 201361 260001
rect 188607 258819 201361 258820
rect 202485 258820 208326 260001
rect 209450 258821 215284 260002
rect 216408 258825 222201 260003
rect 223325 258825 226094 260007
rect 216408 258821 226094 258825
rect 209450 258820 226094 258821
rect 202485 258819 226094 258820
rect 181642 258818 226094 258819
rect 165856 258800 226094 258818
rect 66323 258394 226094 258800
rect 100447 257821 102801 258394
rect 141318 257821 143513 258394
rect 100748 250077 102801 257821
rect 141460 250096 143513 257821
rect 189592 250437 191978 258394
rect 100816 249790 102715 250077
rect 141565 249790 143464 250096
rect 189592 249790 192038 250437
rect 80519 249308 226125 249790
rect 80519 249307 90646 249308
rect 80519 248125 83688 249307
rect 84812 248126 90646 249307
rect 91770 249296 226125 249308
rect 91770 249295 153070 249296
rect 91770 249294 146112 249295
rect 91770 249290 139147 249294
rect 91770 249289 132230 249290
rect 91770 249288 111387 249289
rect 91770 249287 104429 249288
rect 91770 248126 97464 249287
rect 84812 248125 97464 248126
rect 80519 248105 97464 248125
rect 98588 248106 104429 249287
rect 105553 248107 111387 249288
rect 112511 249288 125272 249289
rect 112511 248107 118307 249288
rect 105553 248106 118307 248107
rect 119431 248107 125272 249288
rect 126396 248108 132230 249289
rect 133354 248112 139147 249290
rect 140271 248113 146112 249294
rect 147236 248114 153070 249295
rect 154194 249295 173910 249296
rect 154194 249294 166952 249295
rect 154194 248114 159987 249294
rect 147236 248113 159987 248114
rect 140271 248112 159987 248113
rect 161111 249209 166952 249294
rect 161111 248112 164677 249209
rect 133354 248108 164677 248112
rect 126396 248107 164677 248108
rect 119431 248106 164677 248107
rect 98588 248105 164677 248106
rect 80519 248034 164677 248105
rect 165943 248113 166952 249209
rect 168076 248114 173910 249295
rect 175034 249292 222398 249296
rect 175034 249291 215481 249292
rect 175034 249290 194638 249291
rect 175034 249289 187680 249290
rect 175034 248114 180715 249289
rect 168076 248113 180715 248114
rect 165943 248107 180715 248113
rect 181839 248108 187680 249289
rect 188804 248109 194638 249290
rect 195762 249290 208523 249291
rect 195762 248109 201558 249290
rect 188804 248108 201558 248109
rect 202682 248109 208523 249290
rect 209647 248110 215481 249291
rect 216605 248114 222398 249292
rect 223522 248114 226125 249296
rect 216605 248110 226125 248114
rect 209647 248109 226125 248110
rect 202682 248108 226125 248109
rect 181839 248107 226125 248108
rect 165943 248034 226125 248107
rect 80519 247683 226125 248034
rect 100816 242660 102715 247683
rect 141565 242660 143464 247683
rect 190139 242660 192038 247683
rect 80519 242178 226125 242660
rect 80519 242177 90372 242178
rect 80519 240995 83414 242177
rect 84538 240996 90372 242177
rect 91496 242166 226125 242178
rect 91496 242165 152796 242166
rect 91496 242164 145838 242165
rect 91496 242160 138873 242164
rect 91496 242159 131956 242160
rect 91496 242158 111113 242159
rect 91496 242157 104155 242158
rect 91496 240996 97190 242157
rect 84538 240995 97190 240996
rect 80519 240975 97190 240995
rect 98314 240976 104155 242157
rect 105279 240977 111113 242158
rect 112237 242158 124998 242159
rect 112237 240977 118033 242158
rect 105279 240976 118033 240977
rect 119157 240977 124998 242158
rect 126122 240978 131956 242159
rect 133080 240982 138873 242160
rect 139997 240983 145838 242164
rect 146962 240984 152796 242165
rect 153920 242165 173636 242166
rect 153920 242164 166678 242165
rect 153920 240984 159713 242164
rect 146962 240983 159713 240984
rect 139997 240982 159713 240983
rect 160837 242123 166678 242164
rect 160837 240982 164658 242123
rect 133080 240978 164658 240982
rect 126122 240977 164658 240978
rect 119157 240976 164658 240977
rect 98314 240975 164658 240976
rect 80519 240948 164658 240975
rect 165924 240983 166678 242123
rect 167802 240984 173636 242165
rect 174760 242162 222124 242166
rect 174760 242161 215207 242162
rect 174760 242160 194364 242161
rect 174760 242159 187406 242160
rect 174760 240984 180441 242159
rect 167802 240983 180441 240984
rect 165924 240977 180441 240983
rect 181565 240978 187406 242159
rect 188530 240979 194364 242160
rect 195488 242160 208249 242161
rect 195488 240979 201284 242160
rect 188530 240978 201284 240979
rect 202408 240979 208249 242160
rect 209373 240980 215207 242161
rect 216331 240984 222124 242162
rect 223248 240984 226125 242166
rect 216331 240980 226125 240984
rect 209373 240979 226125 240980
rect 202408 240978 226125 240979
rect 181565 240977 226125 240978
rect 165924 240948 226125 240977
rect 80519 240553 226125 240948
rect 63180 240219 63320 240238
rect 63180 240105 63189 240219
rect 63304 240105 63320 240219
rect 63180 240095 63320 240105
rect 63101 237883 63241 237902
rect 63101 237769 63110 237883
rect 63225 237769 63241 237883
rect 63101 237759 63241 237769
rect 100816 236247 102715 240553
rect 141565 236247 143464 240553
rect 190139 236247 192038 240553
rect 246845 237180 249936 237339
rect 247520 236863 247688 237180
rect 248653 236863 248821 237180
rect 246840 236704 249931 236863
rect 247520 236351 247688 236704
rect 248653 236351 248821 236704
rect 80519 235765 226125 236247
rect 246840 236192 249931 236351
rect 247520 235880 247688 236192
rect 248653 235880 248821 236192
rect 80519 235764 90480 235765
rect 63020 235399 63160 235418
rect 63020 235285 63029 235399
rect 63144 235285 63160 235399
rect 63020 235275 63160 235285
rect 80519 234582 83522 235764
rect 84646 234583 90480 235764
rect 91604 235753 226125 235765
rect 91604 235752 152904 235753
rect 91604 235751 145946 235752
rect 91604 235747 138981 235751
rect 91604 235746 132064 235747
rect 91604 235745 111221 235746
rect 91604 235744 104263 235745
rect 91604 234583 97298 235744
rect 84646 234582 97298 234583
rect 80519 234562 97298 234582
rect 98422 234563 104263 235744
rect 105387 234564 111221 235745
rect 112345 235745 125106 235746
rect 112345 234564 118141 235745
rect 105387 234563 118141 234564
rect 119265 234564 125106 235745
rect 126230 234565 132064 235746
rect 133188 234569 138981 235747
rect 140105 234570 145946 235751
rect 147070 234571 152904 235752
rect 154028 235752 173744 235753
rect 154028 235751 166786 235752
rect 154028 234571 159821 235751
rect 147070 234570 159821 234571
rect 140105 234569 159821 234570
rect 160945 235721 166786 235751
rect 160945 234569 164621 235721
rect 133188 234565 164621 234569
rect 126230 234564 164621 234565
rect 119265 234563 164621 234564
rect 98422 234562 164621 234563
rect 80519 234546 164621 234562
rect 165887 234570 166786 235721
rect 167910 234571 173744 235752
rect 174868 235749 222232 235753
rect 174868 235748 215315 235749
rect 174868 235747 194472 235748
rect 174868 235746 187514 235747
rect 174868 234571 180549 235746
rect 167910 234570 180549 234571
rect 165887 234564 180549 234570
rect 181673 234565 187514 235746
rect 188638 234566 194472 235747
rect 195596 235747 208357 235748
rect 195596 234566 201392 235747
rect 188638 234565 201392 234566
rect 202516 234566 208357 235747
rect 209481 234567 215315 235748
rect 216439 234571 222232 235749
rect 223356 234571 226125 235753
rect 246849 235721 249940 235880
rect 247520 235408 247688 235721
rect 248653 235408 248821 235721
rect 246863 235249 249954 235408
rect 216439 234567 226125 234571
rect 209481 234566 226125 234567
rect 202516 234565 226125 234566
rect 181673 234564 226125 234565
rect 165887 234546 226125 234564
rect 80519 234140 226125 234546
rect 100478 233567 102850 234140
rect 141349 233567 143486 234140
rect 63024 233192 63159 233203
rect 63024 233078 63033 233192
rect 63148 233078 63159 233192
rect 63024 233068 63159 233078
rect 100933 230190 102850 233567
rect 100940 229524 102839 230190
rect 141413 229545 143486 233567
rect 189617 233567 191774 234140
rect 141413 229524 143588 229545
rect 189617 229524 191690 233567
rect 46151 229501 58746 229524
rect 61078 229503 191690 229524
rect 192275 229503 232345 229524
rect 61078 229501 232345 229503
rect 46151 229496 232345 229501
rect 234575 229510 267314 229524
rect 269474 229510 280176 229524
rect 234575 229496 280176 229510
rect 46151 229486 280176 229496
rect 46151 229042 281219 229486
rect 46151 229041 69930 229042
rect 46151 229040 62972 229041
rect 46151 229036 56007 229040
rect 46151 227854 49090 229036
rect 50214 227858 56007 229036
rect 57131 227859 62972 229040
rect 64096 227860 69930 229041
rect 71054 229041 90770 229042
rect 71054 229040 83812 229041
rect 71054 227860 76847 229040
rect 64096 227859 76847 227860
rect 57131 227858 76847 227859
rect 77971 227859 83812 229040
rect 84936 227860 90770 229041
rect 91894 229033 281219 229042
rect 91894 229032 271383 229033
rect 91894 229031 236445 229032
rect 91894 229030 229487 229031
rect 91894 229029 153194 229030
rect 91894 229028 146236 229029
rect 91894 229024 139271 229028
rect 91894 229023 132354 229024
rect 91894 229022 111511 229023
rect 91894 229021 104553 229022
rect 91894 227860 97588 229021
rect 84936 227859 97588 227860
rect 77971 227858 97588 227859
rect 50214 227854 97588 227858
rect 46151 227839 97588 227854
rect 98712 227840 104553 229021
rect 105677 227841 111511 229022
rect 112635 229022 125396 229023
rect 112635 227841 118431 229022
rect 105677 227840 118431 227841
rect 119555 227841 125396 229022
rect 126520 227842 132354 229023
rect 133478 227846 139271 229024
rect 140395 227847 146236 229028
rect 147360 227848 153194 229029
rect 154318 229029 174034 229030
rect 154318 229028 167076 229029
rect 154318 227848 160111 229028
rect 147360 227847 160111 227848
rect 140395 227846 160111 227847
rect 161235 228943 167076 229028
rect 161235 227846 164801 228943
rect 133478 227842 164801 227846
rect 126520 227841 164801 227842
rect 119555 227840 164801 227841
rect 98712 227839 164801 227840
rect 46151 227768 164801 227839
rect 166067 227847 167076 228943
rect 168200 227848 174034 229029
rect 175158 229026 222522 229030
rect 175158 229025 215605 229026
rect 175158 229024 194762 229025
rect 175158 229023 187804 229024
rect 175158 227848 180839 229023
rect 168200 227847 180839 227848
rect 166067 227841 180839 227847
rect 181963 227842 187804 229023
rect 188928 227843 194762 229024
rect 195886 229024 208647 229025
rect 195886 227843 201682 229024
rect 188928 227842 201682 227843
rect 202806 227843 208647 229024
rect 209771 227844 215605 229025
rect 216729 227848 222522 229026
rect 223646 227849 229487 229030
rect 230611 227850 236445 229031
rect 237569 229031 257285 229032
rect 237569 229030 250327 229031
rect 237569 227850 243362 229030
rect 230611 227849 243362 227850
rect 223646 227848 243362 227849
rect 244486 227849 250327 229030
rect 251451 227850 257285 229031
rect 258409 227850 264425 229032
rect 265549 227851 271383 229032
rect 272507 229023 281219 229033
rect 272507 227851 278519 229023
rect 265549 227850 278519 227851
rect 251451 227849 278519 227850
rect 244486 227848 278519 227849
rect 216729 227844 278519 227848
rect 209771 227843 278519 227844
rect 202806 227842 278519 227843
rect 181963 227841 278519 227842
rect 279643 227841 281219 229023
rect 166067 227768 281219 227841
rect 46151 227436 281219 227768
rect 46151 227417 280176 227436
rect 59047 224776 60999 227417
rect 59044 223662 60999 224776
rect 100884 226887 102839 227417
rect 141689 226887 143654 227417
rect 100884 223662 102836 226887
rect 141702 224776 143654 226887
rect 141669 223662 143654 224776
rect 190179 226887 192162 227417
rect 190179 224776 192131 226887
rect 190179 223662 192142 224776
rect 232519 223662 234471 227417
rect 267372 223662 269324 227417
rect 46131 223624 280156 223662
rect 46131 223180 281199 223624
rect 46131 223179 69910 223180
rect 46131 223178 62952 223179
rect 46131 223174 55987 223178
rect 46131 221992 49070 223174
rect 50194 221996 55987 223174
rect 57111 221997 62952 223178
rect 64076 221998 69910 223179
rect 71034 223179 90750 223180
rect 71034 223178 83792 223179
rect 71034 221998 76827 223178
rect 64076 221997 76827 221998
rect 57111 221996 76827 221997
rect 77951 221997 83792 223178
rect 84916 221998 90750 223179
rect 91874 223171 281199 223180
rect 91874 223170 271363 223171
rect 91874 223169 236425 223170
rect 91874 223168 229467 223169
rect 91874 223167 153174 223168
rect 91874 223166 146216 223167
rect 91874 223162 139251 223166
rect 91874 223161 132334 223162
rect 91874 223160 111491 223161
rect 91874 223159 104533 223160
rect 91874 221998 97568 223159
rect 84916 221997 97568 221998
rect 77951 221996 97568 221997
rect 50194 221992 97568 221996
rect 46131 221977 97568 221992
rect 98692 221978 104533 223159
rect 105657 221979 111491 223160
rect 112615 223160 125376 223161
rect 112615 221979 118411 223160
rect 105657 221978 118411 221979
rect 119535 221979 125376 223160
rect 126500 221980 132334 223161
rect 133458 221984 139251 223162
rect 140375 221985 146216 223166
rect 147340 221986 153174 223167
rect 154298 223167 174014 223168
rect 154298 223166 167056 223167
rect 154298 221986 160091 223166
rect 147340 221985 160091 221986
rect 140375 221984 160091 221985
rect 161215 223081 167056 223166
rect 161215 221984 164781 223081
rect 133458 221980 164781 221984
rect 126500 221979 164781 221980
rect 119535 221978 164781 221979
rect 98692 221977 164781 221978
rect 46131 221906 164781 221977
rect 166047 221985 167056 223081
rect 168180 221986 174014 223167
rect 175138 223164 222502 223168
rect 175138 223163 215585 223164
rect 175138 223162 194742 223163
rect 175138 223161 187784 223162
rect 175138 221986 180819 223161
rect 168180 221985 180819 221986
rect 166047 221979 180819 221985
rect 181943 221980 187784 223161
rect 188908 221981 194742 223162
rect 195866 223162 208627 223163
rect 195866 221981 201662 223162
rect 188908 221980 201662 221981
rect 202786 221981 208627 223162
rect 209751 221982 215585 223163
rect 216709 221986 222502 223164
rect 223626 221987 229467 223168
rect 230591 221988 236425 223169
rect 237549 223169 257265 223170
rect 237549 223168 250307 223169
rect 237549 221988 243342 223168
rect 230591 221987 243342 221988
rect 223626 221986 243342 221987
rect 244466 221987 250307 223168
rect 251431 221988 257265 223169
rect 258389 221988 264405 223170
rect 265529 221989 271363 223170
rect 272487 223161 281199 223171
rect 272487 221989 278499 223161
rect 265529 221988 278499 221989
rect 251431 221987 278499 221988
rect 244466 221986 278499 221987
rect 216709 221982 278499 221986
rect 209751 221981 278499 221982
rect 202786 221980 278499 221981
rect 181943 221979 278499 221980
rect 279623 221979 281199 223161
rect 166047 221906 281199 221979
rect 46131 221574 281199 221906
rect 46131 221555 280156 221574
rect 59044 221025 60999 221555
rect 59047 212180 60999 221025
rect 100884 213295 102836 221555
rect 141669 221025 143654 221555
rect 100884 212669 102859 213295
rect 59084 211599 60983 212180
rect 100960 211599 102859 212669
rect 141702 212477 143654 221025
rect 190179 221025 192142 221555
rect 190179 213295 192131 221025
rect 190179 212674 192182 213295
rect 141709 211599 143608 212477
rect 190283 211599 192182 212674
rect 232519 212402 234471 221555
rect 267372 212458 269324 221555
rect 232566 211599 234465 212402
rect 267418 211599 269317 212458
rect 18223 211578 31024 211599
rect 33596 211578 280196 211599
rect 18223 211561 280196 211578
rect 18223 211117 281239 211561
rect 18223 211116 69950 211117
rect 18223 211115 62992 211116
rect 18223 211111 56027 211115
rect 18223 211110 49110 211111
rect 18223 211109 28267 211110
rect 18223 209927 21309 211109
rect 22433 209928 28267 211109
rect 29391 211109 42152 211110
rect 29391 209928 35187 211109
rect 22433 209927 35187 209928
rect 36311 209928 42152 211109
rect 43276 209929 49110 211110
rect 50234 209933 56027 211111
rect 57151 209934 62992 211115
rect 64116 209935 69950 211116
rect 71074 211116 90790 211117
rect 71074 211115 83832 211116
rect 71074 209935 76867 211115
rect 64116 209934 76867 209935
rect 57151 209933 76867 209934
rect 77991 209934 83832 211115
rect 84956 209935 90790 211116
rect 91914 211108 281239 211117
rect 91914 211107 271403 211108
rect 91914 211106 236465 211107
rect 91914 211105 229507 211106
rect 91914 211104 153214 211105
rect 91914 211103 146256 211104
rect 91914 211099 139291 211103
rect 91914 211098 132374 211099
rect 91914 211097 111531 211098
rect 91914 211096 104573 211097
rect 91914 209935 97608 211096
rect 84956 209934 97608 209935
rect 77991 209933 97608 209934
rect 50234 209929 97608 209933
rect 43276 209928 97608 209929
rect 36311 209927 97608 209928
rect 18223 209914 97608 209927
rect 98732 209915 104573 211096
rect 105697 209916 111531 211097
rect 112655 211097 125416 211098
rect 112655 209916 118451 211097
rect 105697 209915 118451 209916
rect 119575 209916 125416 211097
rect 126540 209917 132374 211098
rect 133498 209921 139291 211099
rect 140415 209922 146256 211103
rect 147380 209923 153214 211104
rect 154338 211104 174054 211105
rect 154338 211103 167096 211104
rect 154338 209923 160131 211103
rect 147380 209922 160131 209923
rect 140415 209921 160131 209922
rect 161255 211018 167096 211103
rect 161255 209921 164821 211018
rect 133498 209917 164821 209921
rect 126540 209916 164821 209917
rect 119575 209915 164821 209916
rect 98732 209914 164821 209915
rect 18223 209843 164821 209914
rect 166087 209922 167096 211018
rect 168220 209923 174054 211104
rect 175178 211101 222542 211105
rect 175178 211100 215625 211101
rect 175178 211099 194782 211100
rect 175178 211098 187824 211099
rect 175178 209923 180859 211098
rect 168220 209922 180859 209923
rect 166087 209916 180859 209922
rect 181983 209917 187824 211098
rect 188948 209918 194782 211099
rect 195906 211099 208667 211100
rect 195906 209918 201702 211099
rect 188948 209917 201702 209918
rect 202826 209918 208667 211099
rect 209791 209919 215625 211100
rect 216749 209923 222542 211101
rect 223666 209924 229507 211105
rect 230631 209925 236465 211106
rect 237589 211106 257305 211107
rect 237589 211105 250347 211106
rect 237589 209925 243382 211105
rect 230631 209924 243382 209925
rect 223666 209923 243382 209924
rect 244506 209924 250347 211105
rect 251471 209925 257305 211106
rect 258429 209925 264445 211107
rect 265569 209926 271403 211107
rect 272527 211098 281239 211108
rect 272527 209926 278539 211098
rect 265569 209925 278539 209926
rect 251471 209924 278539 209925
rect 244506 209923 278539 209924
rect 216749 209919 278539 209923
rect 209791 209918 278539 209919
rect 202826 209917 278539 209918
rect 181983 209916 278539 209917
rect 279663 209916 281239 211098
rect 166087 209843 281239 209916
rect 18223 209511 281239 209843
rect 18223 209492 280196 209511
rect 31238 204469 33137 209492
rect 59084 204469 60983 209492
rect 100960 204469 102859 209492
rect 141709 204469 143608 209492
rect 190283 204469 192182 209492
rect 232566 204469 234465 209492
rect 267418 204469 269317 209492
rect 18223 204431 279922 204469
rect 18223 203987 280965 204431
rect 18223 203986 69676 203987
rect 18223 203985 62718 203986
rect 18223 203981 55753 203985
rect 18223 203980 48836 203981
rect 18223 203979 27993 203980
rect 18223 202797 21035 203979
rect 22159 202798 27993 203979
rect 29117 203979 41878 203980
rect 29117 202798 34913 203979
rect 22159 202797 34913 202798
rect 36037 202798 41878 203979
rect 43002 202799 48836 203980
rect 49960 202803 55753 203981
rect 56877 202804 62718 203985
rect 63842 202805 69676 203986
rect 70800 203986 90516 203987
rect 70800 203985 83558 203986
rect 70800 202805 76593 203985
rect 63842 202804 76593 202805
rect 56877 202803 76593 202804
rect 77717 202804 83558 203985
rect 84682 202805 90516 203986
rect 91640 203978 280965 203987
rect 91640 203977 271129 203978
rect 91640 203976 236191 203977
rect 91640 203975 229233 203976
rect 91640 203974 152940 203975
rect 91640 203973 145982 203974
rect 91640 203969 139017 203973
rect 91640 203968 132100 203969
rect 91640 203967 111257 203968
rect 91640 203966 104299 203967
rect 91640 202805 97334 203966
rect 84682 202804 97334 202805
rect 77717 202803 97334 202804
rect 49960 202799 97334 202803
rect 43002 202798 97334 202799
rect 36037 202797 97334 202798
rect 18223 202784 97334 202797
rect 98458 202785 104299 203966
rect 105423 202786 111257 203967
rect 112381 203967 125142 203968
rect 112381 202786 118177 203967
rect 105423 202785 118177 202786
rect 119301 202786 125142 203967
rect 126266 202787 132100 203968
rect 133224 202791 139017 203969
rect 140141 202792 145982 203973
rect 147106 202793 152940 203974
rect 154064 203974 173780 203975
rect 154064 203973 166822 203974
rect 154064 202793 159857 203973
rect 147106 202792 159857 202793
rect 140141 202791 159857 202792
rect 160981 203932 166822 203973
rect 160981 202791 164802 203932
rect 133224 202787 164802 202791
rect 126266 202786 164802 202787
rect 119301 202785 164802 202786
rect 98458 202784 164802 202785
rect 18223 202757 164802 202784
rect 166068 202792 166822 203932
rect 167946 202793 173780 203974
rect 174904 203971 222268 203975
rect 174904 203970 215351 203971
rect 174904 203969 194508 203970
rect 174904 203968 187550 203969
rect 174904 202793 180585 203968
rect 167946 202792 180585 202793
rect 166068 202786 180585 202792
rect 181709 202787 187550 203968
rect 188674 202788 194508 203969
rect 195632 203969 208393 203970
rect 195632 202788 201428 203969
rect 188674 202787 201428 202788
rect 202552 202788 208393 203969
rect 209517 202789 215351 203970
rect 216475 202793 222268 203971
rect 223392 202794 229233 203975
rect 230357 202795 236191 203976
rect 237315 203976 257031 203977
rect 237315 203975 250073 203976
rect 237315 202795 243108 203975
rect 230357 202794 243108 202795
rect 223392 202793 243108 202794
rect 244232 202794 250073 203975
rect 251197 202795 257031 203976
rect 258155 202795 264171 203977
rect 265295 202796 271129 203977
rect 272253 203968 280965 203978
rect 272253 202796 278265 203968
rect 265295 202795 278265 202796
rect 251197 202794 278265 202795
rect 244232 202793 278265 202794
rect 216475 202789 278265 202793
rect 209517 202788 278265 202789
rect 202552 202787 278265 202788
rect 181709 202786 278265 202787
rect 279389 202786 280965 203968
rect 166068 202757 280965 202786
rect 18223 202381 280965 202757
rect 18223 202362 279922 202381
rect 31238 198056 33137 202362
rect 59084 198056 60983 202362
rect 100960 198056 102859 202362
rect 141709 198056 143608 202362
rect 190283 198056 192182 202362
rect 232566 198056 234465 202362
rect 267418 198056 269317 202362
rect 18223 198018 280030 198056
rect 18223 197574 281073 198018
rect 18223 197573 69784 197574
rect 18223 197572 62826 197573
rect 18223 197568 55861 197572
rect 18223 197567 48944 197568
rect 18223 197566 28101 197567
rect 18223 196384 21143 197566
rect 22267 196385 28101 197566
rect 29225 197566 41986 197567
rect 29225 196385 35021 197566
rect 22267 196384 35021 196385
rect 36145 196385 41986 197566
rect 43110 196386 48944 197567
rect 50068 196390 55861 197568
rect 56985 196391 62826 197572
rect 63950 196392 69784 197573
rect 70908 197573 90624 197574
rect 70908 197572 83666 197573
rect 70908 196392 76701 197572
rect 63950 196391 76701 196392
rect 56985 196390 76701 196391
rect 77825 196391 83666 197572
rect 84790 196392 90624 197573
rect 91748 197565 281073 197574
rect 91748 197564 271237 197565
rect 91748 197563 236299 197564
rect 91748 197562 229341 197563
rect 91748 197561 153048 197562
rect 91748 197560 146090 197561
rect 91748 197556 139125 197560
rect 91748 197555 132208 197556
rect 91748 197554 111365 197555
rect 91748 197553 104407 197554
rect 91748 196392 97442 197553
rect 84790 196391 97442 196392
rect 77825 196390 97442 196391
rect 50068 196386 97442 196390
rect 43110 196385 97442 196386
rect 36145 196384 97442 196385
rect 18223 196371 97442 196384
rect 98566 196372 104407 197553
rect 105531 196373 111365 197554
rect 112489 197554 125250 197555
rect 112489 196373 118285 197554
rect 105531 196372 118285 196373
rect 119409 196373 125250 197554
rect 126374 196374 132208 197555
rect 133332 196378 139125 197556
rect 140249 196379 146090 197560
rect 147214 196380 153048 197561
rect 154172 197561 173888 197562
rect 154172 197560 166930 197561
rect 154172 196380 159965 197560
rect 147214 196379 159965 196380
rect 140249 196378 159965 196379
rect 161089 197530 166930 197560
rect 161089 196378 164765 197530
rect 133332 196374 164765 196378
rect 126374 196373 164765 196374
rect 119409 196372 164765 196373
rect 98566 196371 164765 196372
rect 18223 196355 164765 196371
rect 166031 196379 166930 197530
rect 168054 196380 173888 197561
rect 175012 197558 222376 197562
rect 175012 197557 215459 197558
rect 175012 197556 194616 197557
rect 175012 197555 187658 197556
rect 175012 196380 180693 197555
rect 168054 196379 180693 196380
rect 166031 196373 180693 196379
rect 181817 196374 187658 197555
rect 188782 196375 194616 197556
rect 195740 197556 208501 197557
rect 195740 196375 201536 197556
rect 188782 196374 201536 196375
rect 202660 196375 208501 197556
rect 209625 196376 215459 197557
rect 216583 196380 222376 197558
rect 223500 196381 229341 197562
rect 230465 196382 236299 197563
rect 237423 197563 257139 197564
rect 237423 197562 250181 197563
rect 237423 196382 243216 197562
rect 230465 196381 243216 196382
rect 223500 196380 243216 196381
rect 244340 196381 250181 197562
rect 251305 196382 257139 197563
rect 258263 196382 264279 197564
rect 265403 196383 271237 197564
rect 272361 197555 281073 197565
rect 272361 196383 278373 197555
rect 265403 196382 278373 196383
rect 251305 196381 278373 196382
rect 244340 196380 278373 196381
rect 216583 196376 278373 196380
rect 209625 196375 278373 196376
rect 202660 196374 278373 196375
rect 181817 196373 278373 196374
rect 279497 196373 281073 197555
rect 166031 196355 281073 196373
rect 18223 195968 281073 196355
rect 18223 195949 280030 195968
rect 30914 195886 33004 195949
rect 58685 195928 60775 195949
rect 100622 194676 102712 195949
rect 141493 194676 143583 195949
rect 189828 194676 191918 195949
rect 232192 194676 234282 195949
rect 100622 193706 102846 194676
rect 141493 193706 143595 194676
rect 189828 193706 192169 194676
rect 232192 193706 234452 194676
rect 267305 193706 269395 195949
rect 73528 193668 280183 193706
rect 73528 193224 281226 193668
rect 73528 193223 90777 193224
rect 73528 193222 83819 193223
rect 73528 192040 76854 193222
rect 77978 192041 83819 193222
rect 84943 192042 90777 193223
rect 91901 193215 281226 193224
rect 91901 193214 271390 193215
rect 91901 193213 236452 193214
rect 91901 193212 229494 193213
rect 91901 193211 153201 193212
rect 91901 193210 146243 193211
rect 91901 193206 139278 193210
rect 91901 193205 132361 193206
rect 91901 193204 111518 193205
rect 91901 193203 104560 193204
rect 91901 192042 97595 193203
rect 84943 192041 97595 192042
rect 77978 192040 97595 192041
rect 73528 192021 97595 192040
rect 98719 192022 104560 193203
rect 105684 192023 111518 193204
rect 112642 193204 125403 193205
rect 112642 192023 118438 193204
rect 105684 192022 118438 192023
rect 119562 192023 125403 193204
rect 126527 192024 132361 193205
rect 133485 192028 139278 193206
rect 140402 192029 146243 193210
rect 147367 192030 153201 193211
rect 154325 193211 174041 193212
rect 154325 193210 167083 193211
rect 154325 192030 160118 193210
rect 147367 192029 160118 192030
rect 140402 192028 160118 192029
rect 161242 193125 167083 193210
rect 161242 192028 164808 193125
rect 133485 192024 164808 192028
rect 126527 192023 164808 192024
rect 119562 192022 164808 192023
rect 98719 192021 164808 192022
rect 73528 191950 164808 192021
rect 166074 192029 167083 193125
rect 168207 192030 174041 193211
rect 175165 193208 222529 193212
rect 175165 193207 215612 193208
rect 175165 193206 194769 193207
rect 175165 193205 187811 193206
rect 175165 192030 180846 193205
rect 168207 192029 180846 192030
rect 166074 192023 180846 192029
rect 181970 192024 187811 193205
rect 188935 192025 194769 193206
rect 195893 193206 208654 193207
rect 195893 192025 201689 193206
rect 188935 192024 201689 192025
rect 202813 192025 208654 193206
rect 209778 192026 215612 193207
rect 216736 192030 222529 193208
rect 223653 192031 229494 193212
rect 230618 192032 236452 193213
rect 237576 193213 257292 193214
rect 237576 193212 250334 193213
rect 237576 192032 243369 193212
rect 230618 192031 243369 192032
rect 223653 192030 243369 192031
rect 244493 192031 250334 193212
rect 251458 192032 257292 193213
rect 258416 192032 264432 193214
rect 265556 192033 271390 193214
rect 272514 193205 281226 193215
rect 272514 192033 278526 193205
rect 265556 192032 278526 192033
rect 251458 192031 278526 192032
rect 244493 192030 278526 192031
rect 216736 192026 278526 192030
rect 209778 192025 278526 192026
rect 202813 192024 278526 192025
rect 181970 192023 278526 192024
rect 279650 192023 281226 193205
rect 166074 191950 281226 192023
rect 73528 191618 281226 191950
rect 73528 191599 280183 191618
rect 100947 186576 102846 191599
rect 141696 186576 143595 191599
rect 190270 186576 192169 191599
rect 232553 186576 234452 191599
rect 267405 186576 269304 191599
rect 73528 186538 279909 186576
rect 61504 186500 61644 186521
rect 61504 186400 61518 186500
rect 61626 186400 61644 186500
rect 61504 186381 61644 186400
rect 73528 186094 280952 186538
rect 73528 186093 90503 186094
rect 73528 186092 83545 186093
rect 73528 184910 76580 186092
rect 77704 184911 83545 186092
rect 84669 184912 90503 186093
rect 91627 186085 280952 186094
rect 91627 186084 271116 186085
rect 91627 186083 236178 186084
rect 91627 186082 229220 186083
rect 91627 186081 152927 186082
rect 91627 186080 145969 186081
rect 91627 186076 139004 186080
rect 91627 186075 132087 186076
rect 91627 186074 111244 186075
rect 91627 186073 104286 186074
rect 91627 184912 97321 186073
rect 84669 184911 97321 184912
rect 77704 184910 97321 184911
rect 73528 184891 97321 184910
rect 98445 184892 104286 186073
rect 105410 184893 111244 186074
rect 112368 186074 125129 186075
rect 112368 184893 118164 186074
rect 105410 184892 118164 184893
rect 119288 184893 125129 186074
rect 126253 184894 132087 186075
rect 133211 184898 139004 186076
rect 140128 184899 145969 186080
rect 147093 184900 152927 186081
rect 154051 186081 173767 186082
rect 154051 186080 166809 186081
rect 154051 184900 159844 186080
rect 147093 184899 159844 184900
rect 140128 184898 159844 184899
rect 160968 186039 166809 186080
rect 160968 184898 164789 186039
rect 133211 184894 164789 184898
rect 126253 184893 164789 184894
rect 119288 184892 164789 184893
rect 98445 184891 164789 184892
rect 73528 184864 164789 184891
rect 166055 184899 166809 186039
rect 167933 184900 173767 186081
rect 174891 186078 222255 186082
rect 174891 186077 215338 186078
rect 174891 186076 194495 186077
rect 174891 186075 187537 186076
rect 174891 184900 180572 186075
rect 167933 184899 180572 184900
rect 166055 184893 180572 184899
rect 181696 184894 187537 186075
rect 188661 184895 194495 186076
rect 195619 186076 208380 186077
rect 195619 184895 201415 186076
rect 188661 184894 201415 184895
rect 202539 184895 208380 186076
rect 209504 184896 215338 186077
rect 216462 184900 222255 186078
rect 223379 184901 229220 186082
rect 230344 184902 236178 186083
rect 237302 186083 257018 186084
rect 237302 186082 250060 186083
rect 237302 184902 243095 186082
rect 230344 184901 243095 184902
rect 223379 184900 243095 184901
rect 244219 184901 250060 186082
rect 251184 184902 257018 186083
rect 258142 184902 264158 186084
rect 265282 184903 271116 186084
rect 272240 186075 280952 186085
rect 272240 184903 278252 186075
rect 265282 184902 278252 184903
rect 251184 184901 278252 184902
rect 244219 184900 278252 184901
rect 216462 184896 278252 184900
rect 209504 184895 278252 184896
rect 202539 184894 278252 184895
rect 181696 184893 278252 184894
rect 279376 184893 280952 186075
rect 166055 184864 280952 184893
rect 73528 184488 280952 184864
rect 73528 184469 279909 184488
rect 61424 184077 61564 184098
rect 61424 183977 61438 184077
rect 61546 183977 61564 184077
rect 61424 183958 61564 183977
rect 61345 181593 61485 181614
rect 61345 181493 61359 181593
rect 61467 181493 61485 181593
rect 61345 181474 61485 181493
rect 100947 180163 102846 184469
rect 141696 180163 143595 184469
rect 190270 180163 192169 184469
rect 232553 180163 234452 184469
rect 267405 180163 269304 184469
rect 73528 180125 280017 180163
rect 73528 179681 281060 180125
rect 73528 179680 90611 179681
rect 73528 179679 83653 179680
rect 73528 178497 76688 179679
rect 77812 178498 83653 179679
rect 84777 178499 90611 179680
rect 91735 179672 281060 179681
rect 91735 179671 271224 179672
rect 91735 179670 236286 179671
rect 91735 179669 229328 179670
rect 91735 179668 153035 179669
rect 91735 179667 146077 179668
rect 91735 179663 139112 179667
rect 91735 179662 132195 179663
rect 91735 179661 111352 179662
rect 91735 179660 104394 179661
rect 91735 178499 97429 179660
rect 84777 178498 97429 178499
rect 77812 178497 97429 178498
rect 73528 178478 97429 178497
rect 98553 178479 104394 179660
rect 105518 178480 111352 179661
rect 112476 179661 125237 179662
rect 112476 178480 118272 179661
rect 105518 178479 118272 178480
rect 119396 178480 125237 179661
rect 126361 178481 132195 179662
rect 133319 178485 139112 179663
rect 140236 178486 146077 179667
rect 147201 178487 153035 179668
rect 154159 179668 173875 179669
rect 154159 179667 166917 179668
rect 154159 178487 159952 179667
rect 147201 178486 159952 178487
rect 140236 178485 159952 178486
rect 161076 179637 166917 179667
rect 161076 178485 164752 179637
rect 133319 178481 164752 178485
rect 126361 178480 164752 178481
rect 119396 178479 164752 178480
rect 98553 178478 164752 178479
rect 73528 178462 164752 178478
rect 166018 178486 166917 179637
rect 168041 178487 173875 179668
rect 174999 179665 222363 179669
rect 174999 179664 215446 179665
rect 174999 179663 194603 179664
rect 174999 179662 187645 179663
rect 174999 178487 180680 179662
rect 168041 178486 180680 178487
rect 166018 178480 180680 178486
rect 181804 178481 187645 179662
rect 188769 178482 194603 179663
rect 195727 179663 208488 179664
rect 195727 178482 201523 179663
rect 188769 178481 201523 178482
rect 202647 178482 208488 179663
rect 209612 178483 215446 179664
rect 216570 178487 222363 179665
rect 223487 178488 229328 179669
rect 230452 178489 236286 179670
rect 237410 179670 257126 179671
rect 237410 179669 250168 179670
rect 237410 178489 243203 179669
rect 230452 178488 243203 178489
rect 223487 178487 243203 178488
rect 244327 178488 250168 179669
rect 251292 178489 257126 179670
rect 258250 178489 264266 179671
rect 265390 178490 271224 179671
rect 272348 179662 281060 179672
rect 272348 178490 278360 179662
rect 265390 178489 278360 178490
rect 251292 178488 278360 178489
rect 244327 178487 278360 178488
rect 216570 178483 278360 178487
rect 209612 178482 278360 178483
rect 202647 178481 278360 178482
rect 181804 178480 278360 178481
rect 279484 178480 281060 179662
rect 166018 178462 281060 178480
rect 73528 178075 281060 178462
rect 73528 178056 280017 178075
rect 100609 176358 102830 178056
rect 100674 174249 102830 176358
rect 141462 174249 143618 178056
rect 189815 176358 192042 178056
rect 189886 174249 192042 176358
rect 232171 176358 234269 178056
rect 267266 176358 269382 178056
rect 232171 175011 234265 176358
rect 267266 175011 269360 176358
rect 232171 174249 234275 175011
rect 267228 174249 269360 175011
rect 47149 174187 58627 174249
rect 61148 174211 279732 174249
rect 61148 174187 280775 174211
rect 47149 173767 280775 174187
rect 47149 173766 69486 173767
rect 47149 173765 62528 173766
rect 47149 173761 55563 173765
rect 47149 172579 48646 173761
rect 49770 172583 55563 173761
rect 56687 172584 62528 173765
rect 63652 172585 69486 173766
rect 70610 173766 90326 173767
rect 70610 173765 83368 173766
rect 70610 172585 76403 173765
rect 63652 172584 76403 172585
rect 56687 172583 76403 172584
rect 77527 172584 83368 173765
rect 84492 172585 90326 173766
rect 91450 173758 280775 173767
rect 91450 173757 270939 173758
rect 91450 173756 236001 173757
rect 91450 173755 229043 173756
rect 91450 173754 152750 173755
rect 91450 173753 145792 173754
rect 91450 173749 138827 173753
rect 91450 173748 131910 173749
rect 91450 173747 111067 173748
rect 91450 173746 104109 173747
rect 91450 172585 97144 173746
rect 84492 172584 97144 172585
rect 77527 172583 97144 172584
rect 49770 172579 97144 172583
rect 47149 172564 97144 172579
rect 98268 172565 104109 173746
rect 105233 172566 111067 173747
rect 112191 173747 124952 173748
rect 112191 172566 117987 173747
rect 105233 172565 117987 172566
rect 119111 172566 124952 173747
rect 126076 172567 131910 173748
rect 133034 172571 138827 173749
rect 139951 172572 145792 173753
rect 146916 172573 152750 173754
rect 153874 173754 173590 173755
rect 153874 173753 166632 173754
rect 153874 172573 159667 173753
rect 146916 172572 159667 172573
rect 139951 172571 159667 172572
rect 160791 173712 166632 173753
rect 160791 172571 164612 173712
rect 133034 172567 164612 172571
rect 126076 172566 164612 172567
rect 119111 172565 164612 172566
rect 98268 172564 164612 172565
rect 47149 172537 164612 172564
rect 165878 172572 166632 173712
rect 167756 172573 173590 173754
rect 174714 173751 222078 173755
rect 174714 173750 215161 173751
rect 174714 173749 194318 173750
rect 174714 173748 187360 173749
rect 174714 172573 180395 173748
rect 167756 172572 180395 172573
rect 165878 172566 180395 172572
rect 181519 172567 187360 173748
rect 188484 172568 194318 173749
rect 195442 173749 208203 173750
rect 195442 172568 201238 173749
rect 188484 172567 201238 172568
rect 202362 172568 208203 173749
rect 209327 172569 215161 173750
rect 216285 172573 222078 173751
rect 223202 172574 229043 173755
rect 230167 172575 236001 173756
rect 237125 173756 256841 173757
rect 237125 173755 249883 173756
rect 237125 172575 242918 173755
rect 230167 172574 242918 172575
rect 223202 172573 242918 172574
rect 244042 172574 249883 173755
rect 251007 172575 256841 173756
rect 257965 172575 263981 173757
rect 265105 172576 270939 173757
rect 272063 173748 280775 173758
rect 272063 172576 278075 173748
rect 265105 172575 278075 172576
rect 251007 172574 278075 172575
rect 244042 172573 278075 172574
rect 216285 172569 278075 172573
rect 209327 172568 278075 172569
rect 202362 172567 278075 172568
rect 181519 172566 278075 172567
rect 279199 172566 280775 173748
rect 165878 172537 280775 172566
rect 47149 172161 280775 172537
rect 47149 172142 279732 172161
rect 36481 170918 38491 171031
rect 36995 170522 37134 170918
rect 37814 170522 37953 170918
rect 36507 170409 38517 170522
rect 36995 170126 37134 170409
rect 37814 170126 37953 170409
rect 36509 170013 38519 170126
rect 36995 169779 37134 170013
rect 37814 169779 37953 170013
rect 36514 169666 38524 169779
rect 58894 167836 60793 172142
rect 100674 167836 102830 172142
rect 141462 167836 143618 172142
rect 189886 167836 192042 172142
rect 232171 167836 234275 172142
rect 267228 167836 269360 172142
rect 47149 167798 279840 167836
rect 47149 167354 280883 167798
rect 47149 167353 69594 167354
rect 47149 167352 62636 167353
rect 47149 167348 55671 167352
rect 47149 166166 48754 167348
rect 49878 166170 55671 167348
rect 56795 166171 62636 167352
rect 63760 166172 69594 167353
rect 70718 167353 90434 167354
rect 70718 167352 83476 167353
rect 70718 166172 76511 167352
rect 63760 166171 76511 166172
rect 56795 166170 76511 166171
rect 77635 166171 83476 167352
rect 84600 166172 90434 167353
rect 91558 167345 280883 167354
rect 91558 167344 271047 167345
rect 91558 167343 236109 167344
rect 91558 167342 229151 167343
rect 91558 167341 152858 167342
rect 91558 167340 145900 167341
rect 91558 167336 138935 167340
rect 91558 167335 132018 167336
rect 91558 167334 111175 167335
rect 91558 167333 104217 167334
rect 91558 166172 97252 167333
rect 84600 166171 97252 166172
rect 77635 166170 97252 166171
rect 49878 166166 97252 166170
rect 47149 166151 97252 166166
rect 98376 166152 104217 167333
rect 105341 166153 111175 167334
rect 112299 167334 125060 167335
rect 112299 166153 118095 167334
rect 105341 166152 118095 166153
rect 119219 166153 125060 167334
rect 126184 166154 132018 167335
rect 133142 166158 138935 167336
rect 140059 166159 145900 167340
rect 147024 166160 152858 167341
rect 153982 167341 173698 167342
rect 153982 167340 166740 167341
rect 153982 166160 159775 167340
rect 147024 166159 159775 166160
rect 140059 166158 159775 166159
rect 160899 167310 166740 167340
rect 160899 166158 164575 167310
rect 133142 166154 164575 166158
rect 126184 166153 164575 166154
rect 119219 166152 164575 166153
rect 98376 166151 164575 166152
rect 47149 166135 164575 166151
rect 165841 166159 166740 167310
rect 167864 166160 173698 167341
rect 174822 167338 222186 167342
rect 174822 167337 215269 167338
rect 174822 167336 194426 167337
rect 174822 167335 187468 167336
rect 174822 166160 180503 167335
rect 167864 166159 180503 166160
rect 165841 166153 180503 166159
rect 181627 166154 187468 167335
rect 188592 166155 194426 167336
rect 195550 167336 208311 167337
rect 195550 166155 201346 167336
rect 188592 166154 201346 166155
rect 202470 166155 208311 167336
rect 209435 166156 215269 167337
rect 216393 166160 222186 167338
rect 223310 166161 229151 167342
rect 230275 166162 236109 167343
rect 237233 167343 256949 167344
rect 237233 167342 249991 167343
rect 237233 166162 243026 167342
rect 230275 166161 243026 166162
rect 223310 166160 243026 166161
rect 244150 166161 249991 167342
rect 251115 166162 256949 167343
rect 258073 166162 264089 167344
rect 265213 166163 271047 167344
rect 272171 167335 280883 167345
rect 272171 166163 278183 167335
rect 265213 166162 278183 166163
rect 251115 166161 278183 166162
rect 244150 166160 278183 166161
rect 216393 166156 278183 166160
rect 209435 166155 278183 166156
rect 202470 166154 278183 166155
rect 181627 166153 278183 166154
rect 279307 166153 280883 167335
rect 165841 166135 280883 166153
rect 47149 165748 280883 166135
rect 47149 165729 279840 165748
rect 58495 165708 60585 165729
rect 100432 164985 102830 165729
rect 141303 164985 143618 165729
rect 189638 164985 192042 165729
rect 232002 164985 234265 165729
rect 267115 164985 269360 165729
rect 100674 160497 102830 164985
rect 141462 160497 143618 164985
rect 189886 160497 192042 164985
rect 225709 160546 226746 160583
rect 225709 160498 226764 160546
rect 232171 160498 234265 164985
rect 225709 160497 253730 160498
rect 18634 160488 143618 160497
rect 144252 160488 253730 160497
rect 18634 160049 253730 160488
rect 267266 160487 269360 164985
rect 18634 160015 164841 160049
rect 18634 160014 70361 160015
rect 18634 160013 63403 160014
rect 18634 160009 56438 160013
rect 18634 160008 49521 160009
rect 18634 160007 28678 160008
rect 18634 158825 21720 160007
rect 22844 158826 28678 160007
rect 29802 160007 42563 160008
rect 29802 158826 35598 160007
rect 22844 158825 35598 158826
rect 36722 158826 42563 160007
rect 43687 158827 49521 160008
rect 50645 158831 56438 160009
rect 57562 158832 63403 160013
rect 64527 158833 70361 160014
rect 71485 160014 91201 160015
rect 71485 160013 84243 160014
rect 71485 158833 77278 160013
rect 64527 158832 77278 158833
rect 57562 158831 77278 158832
rect 78402 158832 84243 160013
rect 85367 158833 91201 160014
rect 92325 160003 164841 160015
rect 92325 160002 153625 160003
rect 92325 160001 146667 160002
rect 92325 159997 139702 160001
rect 92325 159996 132785 159997
rect 92325 159995 111942 159996
rect 92325 159994 104984 159995
rect 92325 158833 98019 159994
rect 85367 158832 98019 158833
rect 78402 158831 98019 158832
rect 50645 158827 98019 158831
rect 43687 158826 98019 158827
rect 36722 158825 98019 158826
rect 18634 158812 98019 158825
rect 99143 158813 104984 159994
rect 106108 158814 111942 159995
rect 113066 159995 125827 159996
rect 113066 158814 118862 159995
rect 106108 158813 118862 158814
rect 119986 158814 125827 159995
rect 126951 158815 132785 159996
rect 133909 158819 139702 159997
rect 140826 158820 146667 160001
rect 147791 158821 153625 160002
rect 154749 160001 164841 160003
rect 154749 158821 160542 160001
rect 147791 158820 160542 158821
rect 140826 158819 160542 158820
rect 161666 158874 164841 160001
rect 166107 160004 253730 160049
rect 166107 160003 250632 160004
rect 166107 160002 174465 160003
rect 166107 158874 167507 160002
rect 161666 158820 167507 158874
rect 168631 158821 174465 160002
rect 175589 159999 222953 160003
rect 175589 159998 216036 159999
rect 175589 159997 195193 159998
rect 175589 159996 188235 159997
rect 175589 158821 181270 159996
rect 168631 158820 181270 158821
rect 161666 158819 181270 158820
rect 133909 158815 181270 158819
rect 126951 158814 181270 158815
rect 182394 158815 188235 159996
rect 189359 158816 195193 159997
rect 196317 159997 209078 159998
rect 196317 158816 202113 159997
rect 189359 158815 202113 158816
rect 203237 158816 209078 159997
rect 210202 158817 216036 159998
rect 217160 158821 222953 159999
rect 224077 160000 250632 160003
rect 224077 159999 243715 160000
rect 224077 159998 236757 159999
rect 224077 158821 229792 159998
rect 217160 158817 229792 158821
rect 210202 158816 229792 158817
rect 230916 158817 236757 159998
rect 237881 158818 243715 159999
rect 244839 158822 250632 160000
rect 251756 158822 253730 160004
rect 244839 158818 253730 158822
rect 237881 158817 253730 158818
rect 230916 158816 253730 158817
rect 203237 158815 253730 158816
rect 182394 158814 253730 158815
rect 119986 158813 253730 158814
rect 99143 158812 253730 158813
rect 18634 158394 253730 158812
rect 18634 158390 31100 158394
rect 31314 155664 33327 158394
rect 34165 158391 253730 158394
rect 253787 159993 281462 160487
rect 253787 159989 278364 159993
rect 253787 159988 271447 159989
rect 253787 159987 264489 159988
rect 253787 158805 257524 159987
rect 258648 158806 264489 159987
rect 265613 158807 271447 159988
rect 272571 158811 278364 159989
rect 279488 158811 281462 159993
rect 272571 158807 281462 158811
rect 265613 158806 281462 158807
rect 258648 158805 281462 158806
rect 34165 158390 226764 158391
rect 59124 158325 61394 158390
rect 101090 158325 103270 158390
rect 141462 158376 144019 158390
rect 141763 158325 144019 158376
rect 190340 158360 192593 158390
rect 225727 158361 226764 158390
rect 59124 155664 61137 158325
rect 101090 155664 103103 158325
rect 141763 155664 143776 158325
rect 190340 155664 192353 158360
rect 232171 155665 234265 158391
rect 253787 158380 281462 158805
rect 226055 155664 254015 155665
rect 18919 155654 254015 155664
rect 267266 155654 269360 158380
rect 18919 155209 281747 155654
rect 18919 155182 164822 155209
rect 18919 155181 70646 155182
rect 18919 155180 63688 155181
rect 18919 155176 56723 155180
rect 18919 155175 49806 155176
rect 18919 155174 28963 155175
rect 18919 153992 22005 155174
rect 23129 153993 28963 155174
rect 30087 155174 42848 155175
rect 30087 153993 35883 155174
rect 23129 153992 35883 153993
rect 37007 153993 42848 155174
rect 43972 153994 49806 155175
rect 50930 153998 56723 155176
rect 57847 153999 63688 155180
rect 64812 154000 70646 155181
rect 71770 155181 91486 155182
rect 71770 155180 84528 155181
rect 71770 154000 77563 155180
rect 64812 153999 77563 154000
rect 57847 153998 77563 153999
rect 78687 153999 84528 155180
rect 85652 154000 91486 155181
rect 92610 155170 164822 155182
rect 92610 155169 153910 155170
rect 92610 155168 146952 155169
rect 92610 155164 139987 155168
rect 92610 155163 133070 155164
rect 92610 155162 112227 155163
rect 92610 155161 105269 155162
rect 92610 154000 98304 155161
rect 85652 153999 98304 154000
rect 78687 153998 98304 153999
rect 50930 153994 98304 153998
rect 43972 153993 98304 153994
rect 37007 153992 98304 153993
rect 18919 153979 98304 153992
rect 99428 153980 105269 155161
rect 106393 153981 112227 155162
rect 113351 155162 126112 155163
rect 113351 153981 119147 155162
rect 106393 153980 119147 153981
rect 120271 153981 126112 155162
rect 127236 153982 133070 155163
rect 134194 153986 139987 155164
rect 141111 153987 146952 155168
rect 148076 153988 153910 155169
rect 155034 155168 164822 155170
rect 155034 153988 160827 155168
rect 148076 153987 160827 153988
rect 141111 153986 160827 153987
rect 161951 154034 164822 155168
rect 166088 155171 281747 155209
rect 166088 155170 250917 155171
rect 166088 155169 174750 155170
rect 166088 154034 167792 155169
rect 161951 153987 167792 154034
rect 168916 153988 174750 155169
rect 175874 155166 223238 155170
rect 175874 155165 216321 155166
rect 175874 155164 195478 155165
rect 175874 155163 188520 155164
rect 175874 153988 181555 155163
rect 168916 153987 181555 153988
rect 161951 153986 181555 153987
rect 134194 153982 181555 153986
rect 127236 153981 181555 153982
rect 182679 153982 188520 155163
rect 189644 153983 195478 155164
rect 196602 155164 209363 155165
rect 196602 153983 202398 155164
rect 189644 153982 202398 153983
rect 203522 153983 209363 155164
rect 210487 153984 216321 155165
rect 217445 153988 223238 155166
rect 224362 155167 250917 155170
rect 224362 155166 244000 155167
rect 224362 155165 237042 155166
rect 224362 153988 230077 155165
rect 217445 153984 230077 153988
rect 210487 153983 230077 153984
rect 231201 153984 237042 155165
rect 238166 153985 244000 155166
rect 245124 153989 250917 155167
rect 252041 155160 281747 155171
rect 252041 155156 278649 155160
rect 252041 155155 271732 155156
rect 252041 155154 264774 155155
rect 252041 153989 257809 155154
rect 245124 153985 257809 153989
rect 238166 153984 257809 153985
rect 231201 153983 257809 153984
rect 203522 153982 257809 153983
rect 182679 153981 257809 153982
rect 120271 153980 257809 153981
rect 99428 153979 257809 153980
rect 18919 153972 257809 153979
rect 258933 153973 264774 155154
rect 265898 153974 271732 155155
rect 272856 153978 278649 155156
rect 279773 153978 281747 155160
rect 272856 153974 281747 153978
rect 265898 153973 281747 153974
rect 258933 153972 281747 153973
rect 18919 153561 281747 153972
rect 18919 153557 33327 153561
rect 34450 153558 281747 153561
rect 34450 153557 226336 153558
rect 31314 150404 33327 153557
rect 59124 153492 61679 153557
rect 101090 153492 103555 153557
rect 141763 153492 144304 153557
rect 190340 153527 192878 153557
rect 59124 150404 61137 153492
rect 101090 150404 103103 153492
rect 141763 150404 143776 153492
rect 190340 150404 192353 153527
rect 232171 150405 234265 153558
rect 253787 153547 281747 153558
rect 226055 150404 254086 150405
rect 18990 150394 254086 150404
rect 267266 150394 269360 153547
rect 18990 149939 281818 150394
rect 18990 149922 164803 149939
rect 18990 149921 70717 149922
rect 18990 149920 63759 149921
rect 18990 149916 56794 149920
rect 18990 149915 49877 149916
rect 18990 149914 29034 149915
rect 18990 148732 22076 149914
rect 23200 148733 29034 149914
rect 30158 149914 42919 149915
rect 30158 148733 35954 149914
rect 23200 148732 35954 148733
rect 37078 148733 42919 149914
rect 44043 148734 49877 149915
rect 51001 148738 56794 149916
rect 57918 148739 63759 149920
rect 64883 148740 70717 149921
rect 71841 149921 91557 149922
rect 71841 149920 84599 149921
rect 71841 148740 77634 149920
rect 64883 148739 77634 148740
rect 57918 148738 77634 148739
rect 78758 148739 84599 149920
rect 85723 148740 91557 149921
rect 92681 149910 164803 149922
rect 92681 149909 153981 149910
rect 92681 149908 147023 149909
rect 92681 149904 140058 149908
rect 92681 149903 133141 149904
rect 92681 149902 112298 149903
rect 92681 149901 105340 149902
rect 92681 148740 98375 149901
rect 85723 148739 98375 148740
rect 78758 148738 98375 148739
rect 51001 148734 98375 148738
rect 44043 148733 98375 148734
rect 37078 148732 98375 148733
rect 18990 148719 98375 148732
rect 99499 148720 105340 149901
rect 106464 148721 112298 149902
rect 113422 149902 126183 149903
rect 113422 148721 119218 149902
rect 106464 148720 119218 148721
rect 120342 148721 126183 149902
rect 127307 148722 133141 149903
rect 134265 148726 140058 149904
rect 141182 148727 147023 149908
rect 148147 148728 153981 149909
rect 155105 149908 164803 149910
rect 155105 148728 160898 149908
rect 148147 148727 160898 148728
rect 141182 148726 160898 148727
rect 162022 148764 164803 149908
rect 166069 149911 281818 149939
rect 166069 149910 250988 149911
rect 166069 149909 174821 149910
rect 166069 148764 167863 149909
rect 162022 148727 167863 148764
rect 168987 148728 174821 149909
rect 175945 149906 223309 149910
rect 175945 149905 216392 149906
rect 175945 149904 195549 149905
rect 175945 149903 188591 149904
rect 175945 148728 181626 149903
rect 168987 148727 181626 148728
rect 162022 148726 181626 148727
rect 134265 148722 181626 148726
rect 127307 148721 181626 148722
rect 182750 148722 188591 149903
rect 189715 148723 195549 149904
rect 196673 149904 209434 149905
rect 196673 148723 202469 149904
rect 189715 148722 202469 148723
rect 203593 148723 209434 149904
rect 210558 148724 216392 149905
rect 217516 148728 223309 149906
rect 224433 149907 250988 149910
rect 224433 149906 244071 149907
rect 224433 149905 237113 149906
rect 224433 148728 230148 149905
rect 217516 148724 230148 148728
rect 210558 148723 230148 148724
rect 231272 148724 237113 149905
rect 238237 148725 244071 149906
rect 245195 148729 250988 149907
rect 252112 149900 281818 149911
rect 252112 149896 278720 149900
rect 252112 149895 271803 149896
rect 252112 149894 264845 149895
rect 252112 148729 257880 149894
rect 245195 148725 257880 148729
rect 238237 148724 257880 148725
rect 231272 148723 257880 148724
rect 203593 148722 257880 148723
rect 182750 148721 257880 148722
rect 120342 148720 257880 148721
rect 99499 148719 257880 148720
rect 18990 148712 257880 148719
rect 259004 148713 264845 149894
rect 265969 148714 271803 149895
rect 272927 148718 278720 149896
rect 279844 148718 281818 149900
rect 272927 148714 281818 148718
rect 265969 148713 281818 148714
rect 259004 148712 281818 148713
rect 18990 148301 281818 148712
rect 18990 148297 33327 148301
rect 34521 148298 281818 148301
rect 34521 148297 226407 148298
rect 31314 144930 33327 148297
rect 59124 148232 61750 148297
rect 101090 148232 103626 148297
rect 141763 148232 144375 148297
rect 190340 148267 192949 148297
rect 253787 148287 281818 148298
rect 59124 144930 61137 148232
rect 101090 144930 103103 148232
rect 141763 144930 143776 148232
rect 190340 144930 192353 148267
rect 18919 144448 226336 144930
rect 18919 144447 70646 144448
rect 18919 144446 63688 144447
rect 18919 144442 56723 144446
rect 18919 144441 49806 144442
rect 18919 144440 28963 144441
rect 18919 143258 22005 144440
rect 23129 143259 28963 144440
rect 30087 144440 42848 144441
rect 30087 143259 35883 144440
rect 23129 143258 35883 143259
rect 37007 143259 42848 144440
rect 43972 143260 49806 144441
rect 50930 143264 56723 144442
rect 57847 143265 63688 144446
rect 64812 143266 70646 144447
rect 71770 144447 91486 144448
rect 71770 144446 84528 144447
rect 71770 143266 77563 144446
rect 64812 143265 77563 143266
rect 57847 143264 77563 143265
rect 78687 143265 84528 144446
rect 85652 143266 91486 144447
rect 92610 144436 226336 144448
rect 92610 144435 153910 144436
rect 92610 144434 146952 144435
rect 92610 144430 139987 144434
rect 92610 144429 133070 144430
rect 92610 144428 112227 144429
rect 92610 144427 105269 144428
rect 92610 143266 98304 144427
rect 85652 143265 98304 143266
rect 78687 143264 98304 143265
rect 50930 143260 98304 143264
rect 43972 143259 98304 143260
rect 37007 143258 98304 143259
rect 18919 143245 98304 143258
rect 99428 143246 105269 144427
rect 106393 143247 112227 144428
rect 113351 144428 126112 144429
rect 113351 143247 119147 144428
rect 106393 143246 119147 143247
rect 120271 143247 126112 144428
rect 127236 143248 133070 144429
rect 134194 143252 139987 144430
rect 141111 143253 146952 144434
rect 148076 143254 153910 144435
rect 155034 144435 174750 144436
rect 155034 144434 167792 144435
rect 155034 143254 160827 144434
rect 148076 143253 160827 143254
rect 141111 143252 160827 143253
rect 161951 144387 167792 144434
rect 161951 143252 164785 144387
rect 134194 143248 164785 143252
rect 127236 143247 164785 143248
rect 120271 143246 164785 143247
rect 99428 143245 164785 143246
rect 18919 143212 164785 143245
rect 166051 143253 167792 144387
rect 168916 143254 174750 144435
rect 175874 144432 223238 144436
rect 175874 144431 216321 144432
rect 175874 144430 195478 144431
rect 175874 144429 188520 144430
rect 175874 143254 181555 144429
rect 168916 143253 181555 143254
rect 166051 143247 181555 143253
rect 182679 143248 188520 144429
rect 189644 143249 195478 144430
rect 196602 144430 209363 144431
rect 196602 143249 202398 144430
rect 189644 143248 202398 143249
rect 203522 143249 209363 144430
rect 210487 143250 216321 144431
rect 217445 143254 223238 144432
rect 224362 143254 226336 144436
rect 217445 143250 226336 143254
rect 210487 143249 226336 143250
rect 203522 143248 226336 143249
rect 182679 143247 226336 143248
rect 166051 143212 226336 143247
rect 18919 142827 226336 143212
rect 18919 142823 33327 142827
rect 34450 142823 226336 142827
rect 31314 138818 33327 142823
rect 59124 142758 61679 142823
rect 101090 142758 103555 142823
rect 141763 142758 144304 142823
rect 190340 142793 192878 142823
rect 59124 138818 61137 142758
rect 101090 138818 103103 142758
rect 141763 138818 143776 142758
rect 190340 138818 192353 142793
rect 268956 140387 269095 140414
rect 268956 140283 268969 140387
rect 269079 140283 269095 140387
rect 268956 140260 269095 140283
rect 19061 138336 226478 138818
rect 19061 138335 70788 138336
rect 19061 138334 63830 138335
rect 19061 138330 56865 138334
rect 19061 138329 49948 138330
rect 19061 138328 29105 138329
rect 19061 137146 22147 138328
rect 23271 137147 29105 138328
rect 30229 138328 42990 138329
rect 30229 137147 36025 138328
rect 23271 137146 36025 137147
rect 37149 137147 42990 138328
rect 44114 137148 49948 138329
rect 51072 137152 56865 138330
rect 57989 137153 63830 138334
rect 64954 137154 70788 138335
rect 71912 138335 91628 138336
rect 71912 138334 84670 138335
rect 71912 137154 77705 138334
rect 64954 137153 77705 137154
rect 57989 137152 77705 137153
rect 78829 137153 84670 138334
rect 85794 137154 91628 138335
rect 92752 138324 226478 138336
rect 92752 138323 154052 138324
rect 92752 138322 147094 138323
rect 92752 138318 140129 138322
rect 92752 138317 133212 138318
rect 92752 138316 112369 138317
rect 92752 138315 105411 138316
rect 92752 137154 98446 138315
rect 85794 137153 98446 137154
rect 78829 137152 98446 137153
rect 51072 137148 98446 137152
rect 44114 137147 98446 137148
rect 37149 137146 98446 137147
rect 19061 137133 98446 137146
rect 99570 137134 105411 138315
rect 106535 137135 112369 138316
rect 113493 138316 126254 138317
rect 113493 137135 119289 138316
rect 106535 137134 119289 137135
rect 120413 137135 126254 138316
rect 127378 137136 133212 138317
rect 134336 137140 140129 138318
rect 141253 137141 147094 138322
rect 148218 137142 154052 138323
rect 155176 138323 174892 138324
rect 155176 138322 167934 138323
rect 155176 137142 160969 138322
rect 148218 137141 160969 137142
rect 141253 137140 160969 137141
rect 162093 138197 167934 138322
rect 162093 137140 164785 138197
rect 134336 137136 164785 137140
rect 127378 137135 164785 137136
rect 120413 137134 164785 137135
rect 99570 137133 164785 137134
rect 19061 137022 164785 137133
rect 166051 137141 167934 138197
rect 169058 137142 174892 138323
rect 176016 138320 223380 138324
rect 176016 138319 216463 138320
rect 176016 138318 195620 138319
rect 176016 138317 188662 138318
rect 176016 137142 181697 138317
rect 169058 137141 181697 137142
rect 166051 137135 181697 137141
rect 182821 137136 188662 138317
rect 189786 137137 195620 138318
rect 196744 138318 209505 138319
rect 196744 137137 202540 138318
rect 189786 137136 202540 137137
rect 203664 137137 209505 138318
rect 210629 137138 216463 138319
rect 217587 137142 223380 138320
rect 224504 137142 226478 138324
rect 268877 137927 269017 137954
rect 268877 137823 268890 137927
rect 269000 137823 269017 137927
rect 268877 137800 269017 137823
rect 217587 137138 226478 137142
rect 210629 137137 226478 137138
rect 203664 137136 226478 137137
rect 182821 137135 226478 137136
rect 166051 137022 226478 137135
rect 19061 136715 226478 137022
rect 19061 136711 33327 136715
rect 34592 136711 226478 136715
rect 31314 130944 33327 136711
rect 59124 136646 61821 136711
rect 101090 136646 103697 136711
rect 141763 136646 144446 136711
rect 190340 136681 193020 136711
rect 59124 130944 61137 136646
rect 101090 130944 103103 136646
rect 141763 130944 143776 136646
rect 190340 130944 192353 136681
rect 18851 130462 226268 130944
rect 18851 130461 70578 130462
rect 18851 130460 63620 130461
rect 18851 130456 56655 130460
rect 18851 130455 49738 130456
rect 18851 130454 28895 130455
rect 18851 129272 21937 130454
rect 23061 129273 28895 130454
rect 30019 130454 42780 130455
rect 30019 129273 35815 130454
rect 23061 129272 35815 129273
rect 36939 129273 42780 130454
rect 43904 129274 49738 130455
rect 50862 129278 56655 130456
rect 57779 129279 63620 130460
rect 64744 129280 70578 130461
rect 71702 130461 91418 130462
rect 71702 130460 84460 130461
rect 71702 129280 77495 130460
rect 64744 129279 77495 129280
rect 57779 129278 77495 129279
rect 78619 129279 84460 130460
rect 85584 129280 91418 130461
rect 92542 130450 226268 130462
rect 92542 130449 153842 130450
rect 92542 130448 146884 130449
rect 92542 130444 139919 130448
rect 92542 130443 133002 130444
rect 92542 130442 112159 130443
rect 92542 130441 105201 130442
rect 92542 129280 98236 130441
rect 85584 129279 98236 129280
rect 78619 129278 98236 129279
rect 50862 129274 98236 129278
rect 43904 129273 98236 129274
rect 36939 129272 98236 129273
rect 18851 129259 98236 129272
rect 99360 129260 105201 130441
rect 106325 129261 112159 130442
rect 113283 130442 126044 130443
rect 113283 129261 119079 130442
rect 106325 129260 119079 129261
rect 120203 129261 126044 130442
rect 127168 129262 133002 130443
rect 134126 129266 139919 130444
rect 141043 129267 146884 130448
rect 148008 129268 153842 130449
rect 154966 130449 174682 130450
rect 154966 130448 167724 130449
rect 154966 129268 160759 130448
rect 148008 129267 160759 129268
rect 141043 129266 160759 129267
rect 161883 129267 167724 130448
rect 168848 129268 174682 130449
rect 175806 130446 223170 130450
rect 175806 130445 216253 130446
rect 175806 130444 195410 130445
rect 175806 130443 188452 130444
rect 175806 129268 181487 130443
rect 168848 129267 181487 129268
rect 161883 129266 181487 129267
rect 134126 129262 181487 129266
rect 127168 129261 181487 129262
rect 182611 129262 188452 130443
rect 189576 129263 195410 130444
rect 196534 130444 209295 130445
rect 196534 129263 202330 130444
rect 189576 129262 202330 129263
rect 203454 129263 209295 130444
rect 210419 129264 216253 130445
rect 217377 129268 223170 130446
rect 224294 129268 226268 130450
rect 217377 129264 226268 129268
rect 210419 129263 226268 129264
rect 203454 129262 226268 129263
rect 182611 129261 226268 129262
rect 120203 129260 226268 129261
rect 99360 129259 226268 129260
rect 18851 128841 226268 129259
rect 18851 128837 33327 128841
rect 34382 128837 226268 128841
rect 31314 119628 33327 128837
rect 59124 128772 61611 128837
rect 101090 128772 103487 128837
rect 141763 128772 144236 128837
rect 190340 128807 192810 128837
rect 59124 119628 61137 128772
rect 101090 119628 103103 128772
rect 141763 119628 143776 128772
rect 190340 119628 192353 128807
rect 18368 119590 280341 119628
rect 18368 119146 281384 119590
rect 18368 119145 70095 119146
rect 18368 119144 63137 119145
rect 18368 119140 56172 119144
rect 18368 119139 49255 119140
rect 18368 119138 28412 119139
rect 18368 117956 21454 119138
rect 22578 117957 28412 119138
rect 29536 119138 42297 119139
rect 29536 117957 35332 119138
rect 22578 117956 35332 117957
rect 36456 117957 42297 119138
rect 43421 117958 49255 119139
rect 50379 117962 56172 119140
rect 57296 117963 63137 119144
rect 64261 117964 70095 119145
rect 71219 119145 90935 119146
rect 71219 119144 83977 119145
rect 71219 117964 77012 119144
rect 64261 117963 77012 117964
rect 57296 117962 77012 117963
rect 78136 117963 83977 119144
rect 85101 117964 90935 119145
rect 92059 119137 281384 119146
rect 92059 119136 271548 119137
rect 92059 119135 236610 119136
rect 92059 119134 229652 119135
rect 92059 119133 153359 119134
rect 92059 119132 146401 119133
rect 92059 119128 139436 119132
rect 92059 119127 132519 119128
rect 92059 119126 111676 119127
rect 92059 119125 104718 119126
rect 92059 117964 97753 119125
rect 85101 117963 97753 117964
rect 78136 117962 97753 117963
rect 50379 117958 97753 117962
rect 43421 117957 97753 117958
rect 36456 117956 97753 117957
rect 18368 117943 97753 117956
rect 98877 117944 104718 119125
rect 105842 117945 111676 119126
rect 112800 119126 125561 119127
rect 112800 117945 118596 119126
rect 105842 117944 118596 117945
rect 119720 117945 125561 119126
rect 126685 117946 132519 119127
rect 133643 117950 139436 119128
rect 140560 117951 146401 119132
rect 147525 117952 153359 119133
rect 154483 119133 174199 119134
rect 154483 119132 167241 119133
rect 154483 117952 160276 119132
rect 147525 117951 160276 117952
rect 140560 117950 160276 117951
rect 161400 119093 167241 119132
rect 161400 117950 164793 119093
rect 133643 117946 164793 117950
rect 126685 117945 164793 117946
rect 119720 117944 164793 117945
rect 98877 117943 164793 117944
rect 18368 117918 164793 117943
rect 166059 117951 167241 119093
rect 168365 117952 174199 119133
rect 175323 119130 222687 119134
rect 175323 119129 215770 119130
rect 175323 119128 194927 119129
rect 175323 119127 187969 119128
rect 175323 117952 181004 119127
rect 168365 117951 181004 117952
rect 166059 117945 181004 117951
rect 182128 117946 187969 119127
rect 189093 117947 194927 119128
rect 196051 119128 208812 119129
rect 196051 117947 201847 119128
rect 189093 117946 201847 117947
rect 202971 117947 208812 119128
rect 209936 117948 215770 119129
rect 216894 117952 222687 119130
rect 223811 117953 229652 119134
rect 230776 117954 236610 119135
rect 237734 119135 257450 119136
rect 237734 119134 250492 119135
rect 237734 117954 243527 119134
rect 230776 117953 243527 117954
rect 223811 117952 243527 117953
rect 244651 117953 250492 119134
rect 251616 117954 257450 119135
rect 258574 117954 264590 119136
rect 265714 117955 271548 119136
rect 272672 119127 281384 119137
rect 272672 117955 278684 119127
rect 265714 117954 278684 117955
rect 251616 117953 278684 117954
rect 244651 117952 278684 117953
rect 216894 117948 278684 117952
rect 209936 117947 278684 117948
rect 202971 117946 278684 117947
rect 182128 117945 278684 117946
rect 279808 117945 281384 119127
rect 166059 117918 281384 117945
rect 18368 117540 281384 117918
rect 18368 117521 280341 117540
rect 31314 116424 33327 117521
rect 31383 111676 33282 116424
rect 59124 116136 61137 117521
rect 101090 116639 103103 117521
rect 141763 117070 143776 117521
rect 59229 111676 61128 116136
rect 101105 111676 103004 116639
rect 141854 111676 143753 117070
rect 190340 115921 192353 117521
rect 190428 111676 192327 115921
rect 232711 111676 234610 117521
rect 267563 111676 269462 117521
rect 18368 111638 280546 111676
rect 18368 111194 281589 111638
rect 18368 111193 70300 111194
rect 18368 111192 63342 111193
rect 18368 111188 56377 111192
rect 18368 111187 49460 111188
rect 18368 111186 28617 111187
rect 18368 110004 21659 111186
rect 22783 110005 28617 111186
rect 29741 111186 42502 111187
rect 29741 110005 35537 111186
rect 22783 110004 35537 110005
rect 36661 110005 42502 111186
rect 43626 110006 49460 111187
rect 50584 110010 56377 111188
rect 57501 110011 63342 111192
rect 64466 110012 70300 111193
rect 71424 111193 91140 111194
rect 71424 111192 84182 111193
rect 71424 110012 77217 111192
rect 64466 110011 77217 110012
rect 57501 110010 77217 110011
rect 78341 110011 84182 111192
rect 85306 110012 91140 111193
rect 92264 111185 281589 111194
rect 92264 111184 271753 111185
rect 92264 111183 236815 111184
rect 92264 111182 229857 111183
rect 92264 111181 153564 111182
rect 92264 111180 146606 111181
rect 92264 111176 139641 111180
rect 92264 111175 132724 111176
rect 92264 111174 111881 111175
rect 92264 111173 104923 111174
rect 92264 110012 97958 111173
rect 85306 110011 97958 110012
rect 78341 110010 97958 110011
rect 50584 110006 97958 110010
rect 43626 110005 97958 110006
rect 36661 110004 97958 110005
rect 18368 109991 97958 110004
rect 99082 109992 104923 111173
rect 106047 109993 111881 111174
rect 113005 111174 125766 111175
rect 113005 109993 118801 111174
rect 106047 109992 118801 109993
rect 119925 109993 125766 111174
rect 126890 109994 132724 111175
rect 133848 109998 139641 111176
rect 140765 109999 146606 111180
rect 147730 110000 153564 111181
rect 154688 111181 174404 111182
rect 154688 111180 167446 111181
rect 154688 110000 160481 111180
rect 147730 109999 160481 110000
rect 140765 109998 160481 109999
rect 161605 111166 167446 111180
rect 161605 109998 164902 111166
rect 133848 109994 164902 109998
rect 126890 109993 164902 109994
rect 119925 109992 164902 109993
rect 99082 109991 164902 109992
rect 166168 109999 167446 111166
rect 168570 110000 174404 111181
rect 175528 111178 222892 111182
rect 175528 111177 215975 111178
rect 175528 111176 195132 111177
rect 175528 111175 188174 111176
rect 175528 110000 181209 111175
rect 168570 109999 181209 110000
rect 166168 109993 181209 109999
rect 182333 109994 188174 111175
rect 189298 109995 195132 111176
rect 196256 111176 209017 111177
rect 196256 109995 202052 111176
rect 189298 109994 202052 109995
rect 203176 109995 209017 111176
rect 210141 109996 215975 111177
rect 217099 110000 222892 111178
rect 224016 110001 229857 111182
rect 230981 110002 236815 111183
rect 237939 111183 257655 111184
rect 237939 111182 250697 111183
rect 237939 110002 243732 111182
rect 230981 110001 243732 110002
rect 224016 110000 243732 110001
rect 244856 110001 250697 111182
rect 251821 110002 257655 111183
rect 258779 110002 264795 111184
rect 265919 110003 271753 111184
rect 272877 111175 281589 111185
rect 272877 110003 278889 111175
rect 265919 110002 278889 110003
rect 251821 110001 278889 110002
rect 244856 110000 278889 110001
rect 217099 109996 278889 110000
rect 210141 109995 278889 109996
rect 203176 109994 278889 109995
rect 182333 109993 278889 109994
rect 280013 109993 281589 111175
rect 166168 109991 281589 109993
rect 18368 109588 281589 109991
rect 18368 109569 280546 109588
rect 31383 103450 33282 109569
rect 59229 103450 61128 109569
rect 101105 103450 103004 109569
rect 141854 103450 143753 109569
rect 190428 103450 192327 109569
rect 232711 103450 234610 109569
rect 267563 103450 269462 109569
rect 18368 103412 280546 103450
rect 18368 102968 281589 103412
rect 18368 102967 70300 102968
rect 18368 102966 63342 102967
rect 18368 102962 56377 102966
rect 18368 102961 49460 102962
rect 18368 102960 28617 102961
rect 18368 101778 21659 102960
rect 22783 101779 28617 102960
rect 29741 102960 42502 102961
rect 29741 101779 35537 102960
rect 22783 101778 35537 101779
rect 36661 101779 42502 102960
rect 43626 101780 49460 102961
rect 50584 101784 56377 102962
rect 57501 101785 63342 102966
rect 64466 101786 70300 102967
rect 71424 102967 91140 102968
rect 71424 102966 84182 102967
rect 71424 101786 77217 102966
rect 64466 101785 77217 101786
rect 57501 101784 77217 101785
rect 78341 101785 84182 102966
rect 85306 101786 91140 102967
rect 92264 102964 281589 102968
rect 92264 102956 165003 102964
rect 92264 102955 153564 102956
rect 92264 102954 146606 102955
rect 92264 102950 139641 102954
rect 92264 102949 132724 102950
rect 92264 102948 111881 102949
rect 92264 102947 104923 102948
rect 92264 101786 97958 102947
rect 85306 101785 97958 101786
rect 78341 101784 97958 101785
rect 50584 101780 97958 101784
rect 43626 101779 97958 101780
rect 36661 101778 97958 101779
rect 18368 101765 97958 101778
rect 99082 101766 104923 102947
rect 106047 101767 111881 102948
rect 113005 102948 125766 102949
rect 113005 101767 118801 102948
rect 106047 101766 118801 101767
rect 119925 101767 125766 102948
rect 126890 101768 132724 102949
rect 133848 101772 139641 102950
rect 140765 101773 146606 102954
rect 147730 101774 153564 102955
rect 154688 102954 165003 102956
rect 154688 101774 160481 102954
rect 147730 101773 160481 101774
rect 140765 101772 160481 101773
rect 161605 101789 165003 102954
rect 166269 102959 281589 102964
rect 166269 102958 271753 102959
rect 166269 102957 236815 102958
rect 166269 102956 229857 102957
rect 166269 102955 174404 102956
rect 166269 101789 167446 102955
rect 161605 101773 167446 101789
rect 168570 101774 174404 102955
rect 175528 102952 222892 102956
rect 175528 102951 215975 102952
rect 175528 102950 195132 102951
rect 175528 102949 188174 102950
rect 175528 101774 181209 102949
rect 168570 101773 181209 101774
rect 161605 101772 181209 101773
rect 133848 101768 181209 101772
rect 126890 101767 181209 101768
rect 182333 101768 188174 102949
rect 189298 101769 195132 102950
rect 196256 102950 209017 102951
rect 196256 101769 202052 102950
rect 189298 101768 202052 101769
rect 203176 101769 209017 102950
rect 210141 101770 215975 102951
rect 217099 101774 222892 102952
rect 224016 101775 229857 102956
rect 230981 101776 236815 102957
rect 237939 102957 257655 102958
rect 237939 102956 250697 102957
rect 237939 101776 243732 102956
rect 230981 101775 243732 101776
rect 224016 101774 243732 101775
rect 244856 101775 250697 102956
rect 251821 101776 257655 102957
rect 258779 101776 264795 102958
rect 265919 101777 271753 102958
rect 272877 102949 281589 102959
rect 272877 101777 278889 102949
rect 265919 101776 278889 101777
rect 251821 101775 278889 101776
rect 244856 101774 278889 101775
rect 217099 101770 278889 101774
rect 210141 101769 278889 101770
rect 203176 101768 278889 101769
rect 182333 101767 278889 101768
rect 280013 101767 281589 102949
rect 119925 101766 281589 101767
rect 99082 101765 281589 101766
rect 18368 101362 281589 101765
rect 18368 101343 280546 101362
rect 31383 96046 33282 101343
rect 59229 96046 61128 101343
rect 101105 96046 103004 101343
rect 141854 96046 143753 101343
rect 190428 96046 192327 101343
rect 232711 96046 234610 101343
rect 267563 96046 269462 101343
rect 18368 96008 280341 96046
rect 18368 95564 281384 96008
rect 18368 95563 70095 95564
rect 18368 95562 63137 95563
rect 18368 95558 56172 95562
rect 18368 95557 49255 95558
rect 18368 95556 28412 95557
rect 18368 94374 21454 95556
rect 22578 94375 28412 95556
rect 29536 95556 42297 95557
rect 29536 94375 35332 95556
rect 22578 94374 35332 94375
rect 36456 94375 42297 95556
rect 43421 94376 49255 95557
rect 50379 94380 56172 95558
rect 57296 94381 63137 95562
rect 64261 94382 70095 95563
rect 71219 95563 90935 95564
rect 71219 95562 83977 95563
rect 71219 94382 77012 95562
rect 64261 94381 77012 94382
rect 57296 94380 77012 94381
rect 78136 94381 83977 95562
rect 85101 94382 90935 95563
rect 92059 95555 281384 95564
rect 92059 95554 271548 95555
rect 92059 95553 236610 95554
rect 92059 95552 229652 95553
rect 92059 95551 153359 95552
rect 92059 95550 146401 95551
rect 92059 95546 139436 95550
rect 92059 95545 132519 95546
rect 92059 95544 111676 95545
rect 92059 95543 104718 95544
rect 92059 94382 97753 95543
rect 85101 94381 97753 94382
rect 78136 94380 97753 94381
rect 50379 94376 97753 94380
rect 43421 94375 97753 94376
rect 36456 94374 97753 94375
rect 18368 94361 97753 94374
rect 98877 94362 104718 95543
rect 105842 94363 111676 95544
rect 112800 95544 125561 95545
rect 112800 94363 118596 95544
rect 105842 94362 118596 94363
rect 119720 94363 125561 95544
rect 126685 94364 132519 95545
rect 133643 94368 139436 95546
rect 140560 94369 146401 95550
rect 147525 94370 153359 95551
rect 154483 95551 174199 95552
rect 154483 95550 167241 95551
rect 154483 94370 160276 95550
rect 147525 94369 160276 94370
rect 140560 94368 160276 94369
rect 161400 95465 167241 95550
rect 161400 94368 164966 95465
rect 133643 94364 164966 94368
rect 126685 94363 164966 94364
rect 119720 94362 164966 94363
rect 98877 94361 164966 94362
rect 18368 94290 164966 94361
rect 166232 94369 167241 95465
rect 168365 94370 174199 95551
rect 175323 95548 222687 95552
rect 175323 95547 215770 95548
rect 175323 95546 194927 95547
rect 175323 95545 187969 95546
rect 175323 94370 181004 95545
rect 168365 94369 181004 94370
rect 166232 94363 181004 94369
rect 182128 94364 187969 95545
rect 189093 94365 194927 95546
rect 196051 95546 208812 95547
rect 196051 94365 201847 95546
rect 189093 94364 201847 94365
rect 202971 94365 208812 95546
rect 209936 94366 215770 95547
rect 216894 94370 222687 95548
rect 223811 94371 229652 95552
rect 230776 94372 236610 95553
rect 237734 95553 257450 95554
rect 237734 95552 250492 95553
rect 237734 94372 243527 95552
rect 230776 94371 243527 94372
rect 223811 94370 243527 94371
rect 244651 94371 250492 95552
rect 251616 94372 257450 95553
rect 258574 94372 264590 95554
rect 265714 94373 271548 95554
rect 272672 95545 281384 95555
rect 272672 94373 278684 95545
rect 265714 94372 278684 94373
rect 251616 94371 278684 94372
rect 244651 94370 278684 94371
rect 216894 94366 278684 94370
rect 209936 94365 278684 94366
rect 202971 94364 278684 94365
rect 182128 94363 278684 94364
rect 279808 94363 281384 95545
rect 166232 94290 281384 94363
rect 18368 93958 281384 94290
rect 18368 93939 280341 93958
rect 31383 88916 33282 93939
rect 59229 88916 61128 93939
rect 101105 88916 103004 93939
rect 141854 88916 143753 93939
rect 190428 88916 192327 93939
rect 232711 88916 234610 93939
rect 267563 88916 269462 93939
rect 18368 88878 280067 88916
rect 18368 88434 281110 88878
rect 18368 88433 69821 88434
rect 18368 88432 62863 88433
rect 18368 88428 55898 88432
rect 18368 88427 48981 88428
rect 18368 88426 28138 88427
rect 18368 87244 21180 88426
rect 22304 87245 28138 88426
rect 29262 88426 42023 88427
rect 29262 87245 35058 88426
rect 22304 87244 35058 87245
rect 36182 87245 42023 88426
rect 43147 87246 48981 88427
rect 50105 87250 55898 88428
rect 57022 87251 62863 88432
rect 63987 87252 69821 88433
rect 70945 88433 90661 88434
rect 70945 88432 83703 88433
rect 70945 87252 76738 88432
rect 63987 87251 76738 87252
rect 57022 87250 76738 87251
rect 77862 87251 83703 88432
rect 84827 87252 90661 88433
rect 91785 88425 281110 88434
rect 91785 88424 271274 88425
rect 91785 88423 236336 88424
rect 91785 88422 229378 88423
rect 91785 88421 153085 88422
rect 91785 88420 146127 88421
rect 91785 88416 139162 88420
rect 91785 88415 132245 88416
rect 91785 88414 111402 88415
rect 91785 88413 104444 88414
rect 91785 87252 97479 88413
rect 84827 87251 97479 87252
rect 77862 87250 97479 87251
rect 50105 87246 97479 87250
rect 43147 87245 97479 87246
rect 36182 87244 97479 87245
rect 18368 87231 97479 87244
rect 98603 87232 104444 88413
rect 105568 87233 111402 88414
rect 112526 88414 125287 88415
rect 112526 87233 118322 88414
rect 105568 87232 118322 87233
rect 119446 87233 125287 88414
rect 126411 87234 132245 88415
rect 133369 87238 139162 88416
rect 140286 87239 146127 88420
rect 147251 87240 153085 88421
rect 154209 88421 173925 88422
rect 154209 88420 166967 88421
rect 154209 87240 160002 88420
rect 147251 87239 160002 87240
rect 140286 87238 160002 87239
rect 161126 88379 166967 88420
rect 161126 87238 164947 88379
rect 133369 87234 164947 87238
rect 126411 87233 164947 87234
rect 119446 87232 164947 87233
rect 98603 87231 164947 87232
rect 18368 87204 164947 87231
rect 166213 87239 166967 88379
rect 168091 87240 173925 88421
rect 175049 88418 222413 88422
rect 175049 88417 215496 88418
rect 175049 88416 194653 88417
rect 175049 88415 187695 88416
rect 175049 87240 180730 88415
rect 168091 87239 180730 87240
rect 166213 87233 180730 87239
rect 181854 87234 187695 88415
rect 188819 87235 194653 88416
rect 195777 88416 208538 88417
rect 195777 87235 201573 88416
rect 188819 87234 201573 87235
rect 202697 87235 208538 88416
rect 209662 87236 215496 88417
rect 216620 87240 222413 88418
rect 223537 87241 229378 88422
rect 230502 87242 236336 88423
rect 237460 88423 257176 88424
rect 237460 88422 250218 88423
rect 237460 87242 243253 88422
rect 230502 87241 243253 87242
rect 223537 87240 243253 87241
rect 244377 87241 250218 88422
rect 251342 87242 257176 88423
rect 258300 87242 264316 88424
rect 265440 87243 271274 88424
rect 272398 88415 281110 88425
rect 272398 87243 278410 88415
rect 265440 87242 278410 87243
rect 251342 87241 278410 87242
rect 244377 87240 278410 87241
rect 216620 87236 278410 87240
rect 209662 87235 278410 87236
rect 202697 87234 278410 87235
rect 181854 87233 278410 87234
rect 279534 87233 281110 88415
rect 166213 87204 281110 87233
rect 18368 86828 281110 87204
rect 18368 86809 280067 86828
rect 31383 82503 33282 86809
rect 59229 82503 61128 86809
rect 101105 82503 103004 86809
rect 141854 82503 143753 86809
rect 190428 82503 192327 86809
rect 232711 82503 234610 86809
rect 267563 82503 269462 86809
rect 18368 82465 280175 82503
rect 18368 82021 281218 82465
rect 18368 82020 69929 82021
rect 18368 82019 62971 82020
rect 18368 82015 56006 82019
rect 18368 82014 49089 82015
rect 18368 82013 28246 82014
rect 18368 80831 21288 82013
rect 22412 80832 28246 82013
rect 29370 82013 42131 82014
rect 29370 80832 35166 82013
rect 22412 80831 35166 80832
rect 36290 80832 42131 82013
rect 43255 80833 49089 82014
rect 50213 80837 56006 82015
rect 57130 80838 62971 82019
rect 64095 80839 69929 82020
rect 71053 82020 90769 82021
rect 71053 82019 83811 82020
rect 71053 80839 76846 82019
rect 64095 80838 76846 80839
rect 57130 80837 76846 80838
rect 77970 80838 83811 82019
rect 84935 80839 90769 82020
rect 91893 82012 281218 82021
rect 91893 82011 271382 82012
rect 91893 82010 236444 82011
rect 91893 82009 229486 82010
rect 91893 82008 153193 82009
rect 91893 82007 146235 82008
rect 91893 82003 139270 82007
rect 91893 82002 132353 82003
rect 91893 82001 111510 82002
rect 91893 82000 104552 82001
rect 91893 80839 97587 82000
rect 84935 80838 97587 80839
rect 77970 80837 97587 80838
rect 50213 80833 97587 80837
rect 43255 80832 97587 80833
rect 36290 80831 97587 80832
rect 18368 80818 97587 80831
rect 98711 80819 104552 82000
rect 105676 80820 111510 82001
rect 112634 82001 125395 82002
rect 112634 80820 118430 82001
rect 105676 80819 118430 80820
rect 119554 80820 125395 82001
rect 126519 80821 132353 82002
rect 133477 80825 139270 82003
rect 140394 80826 146235 82007
rect 147359 80827 153193 82008
rect 154317 82008 174033 82009
rect 154317 82007 167075 82008
rect 154317 80827 160110 82007
rect 147359 80826 160110 80827
rect 140394 80825 160110 80826
rect 161234 81977 167075 82007
rect 161234 80825 164910 81977
rect 133477 80821 164910 80825
rect 126519 80820 164910 80821
rect 119554 80819 164910 80820
rect 98711 80818 164910 80819
rect 18368 80802 164910 80818
rect 166176 80826 167075 81977
rect 168199 80827 174033 82008
rect 175157 82005 222521 82009
rect 175157 82004 215604 82005
rect 175157 82003 194761 82004
rect 175157 82002 187803 82003
rect 175157 80827 180838 82002
rect 168199 80826 180838 80827
rect 166176 80820 180838 80826
rect 181962 80821 187803 82002
rect 188927 80822 194761 82003
rect 195885 82003 208646 82004
rect 195885 80822 201681 82003
rect 188927 80821 201681 80822
rect 202805 80822 208646 82003
rect 209770 80823 215604 82004
rect 216728 80827 222521 82005
rect 223645 80828 229486 82009
rect 230610 80829 236444 82010
rect 237568 82010 257284 82011
rect 237568 82009 250326 82010
rect 237568 80829 243361 82009
rect 230610 80828 243361 80829
rect 223645 80827 243361 80828
rect 244485 80828 250326 82009
rect 251450 80829 257284 82010
rect 258408 80829 264424 82011
rect 265548 80830 271382 82011
rect 272506 82002 281218 82012
rect 272506 80830 278518 82002
rect 265548 80829 278518 80830
rect 251450 80828 278518 80829
rect 244485 80827 278518 80828
rect 216728 80823 278518 80827
rect 209770 80822 278518 80823
rect 202805 80821 278518 80822
rect 181962 80820 278518 80821
rect 279642 80820 281218 82002
rect 166176 80802 281218 80820
rect 18368 80415 281218 80802
rect 18368 80396 280175 80415
rect 31059 71323 33149 80396
rect 58830 71584 60920 80396
rect 100767 71584 102857 80396
rect 58830 71323 60994 71584
rect 100767 71323 102870 71584
rect 141638 71323 143728 80396
rect 189973 71584 192063 80396
rect 232337 71584 234427 80396
rect 267450 71584 269540 80396
rect 189973 71323 192193 71584
rect 232337 71323 234476 71584
rect 267429 71323 269540 71584
rect 18234 71285 280041 71323
rect 18234 70841 281084 71285
rect 18234 70840 69795 70841
rect 18234 70839 62837 70840
rect 18234 70835 55872 70839
rect 18234 70834 48955 70835
rect 18234 70833 28112 70834
rect 18234 69651 21154 70833
rect 22278 69652 28112 70833
rect 29236 70833 41997 70834
rect 29236 69652 35032 70833
rect 22278 69651 35032 69652
rect 36156 69652 41997 70833
rect 43121 69653 48955 70834
rect 50079 69657 55872 70835
rect 56996 69658 62837 70839
rect 63961 69659 69795 70840
rect 70919 70840 90635 70841
rect 70919 70839 83677 70840
rect 70919 69659 76712 70839
rect 63961 69658 76712 69659
rect 56996 69657 76712 69658
rect 77836 69658 83677 70839
rect 84801 69659 90635 70840
rect 91759 70832 281084 70841
rect 91759 70831 271248 70832
rect 91759 70830 236310 70831
rect 91759 70829 229352 70830
rect 91759 70828 153059 70829
rect 91759 70827 146101 70828
rect 91759 70823 139136 70827
rect 91759 70822 132219 70823
rect 91759 70821 111376 70822
rect 91759 70820 104418 70821
rect 91759 69659 97453 70820
rect 84801 69658 97453 69659
rect 77836 69657 97453 69658
rect 50079 69653 97453 69657
rect 43121 69652 97453 69653
rect 36156 69651 97453 69652
rect 18234 69638 97453 69651
rect 98577 69639 104418 70820
rect 105542 69640 111376 70821
rect 112500 70821 125261 70822
rect 112500 69640 118296 70821
rect 105542 69639 118296 69640
rect 119420 69640 125261 70821
rect 126385 69641 132219 70822
rect 133343 69645 139136 70823
rect 140260 69646 146101 70827
rect 147225 69647 153059 70828
rect 154183 70828 173899 70829
rect 154183 70827 166941 70828
rect 154183 69647 159976 70827
rect 147225 69646 159976 69647
rect 140260 69645 159976 69646
rect 161100 70727 166941 70827
rect 161100 69645 164892 70727
rect 133343 69641 164892 69645
rect 126385 69640 164892 69641
rect 119420 69639 164892 69640
rect 98577 69638 164892 69639
rect 18234 69552 164892 69638
rect 166158 69646 166941 70727
rect 168065 69647 173899 70828
rect 175023 70825 222387 70829
rect 175023 70824 215470 70825
rect 175023 70823 194627 70824
rect 175023 70822 187669 70823
rect 175023 69647 180704 70822
rect 168065 69646 180704 69647
rect 166158 69640 180704 69646
rect 181828 69641 187669 70822
rect 188793 69642 194627 70823
rect 195751 70823 208512 70824
rect 195751 69642 201547 70823
rect 188793 69641 201547 69642
rect 202671 69642 208512 70823
rect 209636 69643 215470 70824
rect 216594 69647 222387 70825
rect 223511 69648 229352 70829
rect 230476 69649 236310 70830
rect 237434 70830 257150 70831
rect 237434 70829 250192 70830
rect 237434 69649 243227 70829
rect 230476 69648 243227 69649
rect 223511 69647 243227 69648
rect 244351 69648 250192 70829
rect 251316 69649 257150 70830
rect 258274 69649 264290 70831
rect 265414 69650 271248 70831
rect 272372 70822 281084 70832
rect 272372 69650 278384 70822
rect 265414 69649 278384 69650
rect 251316 69648 278384 69649
rect 244351 69647 278384 69648
rect 216594 69643 278384 69647
rect 209636 69642 278384 69643
rect 202671 69641 278384 69642
rect 181828 69640 278384 69641
rect 279508 69640 281084 70822
rect 166158 69552 281084 69640
rect 18234 69235 281084 69552
rect 18234 69216 280041 69235
rect 31059 65083 33149 69216
rect 58830 65344 60920 69216
rect 58830 65083 60959 65344
rect 100767 65083 102857 69216
rect 141638 65083 143728 69216
rect 189973 65344 192063 69216
rect 232337 65344 234427 69216
rect 267450 65344 269540 69216
rect 189973 65083 192158 65344
rect 232337 65083 234441 65344
rect 267394 65083 269540 65344
rect 18199 65045 280006 65083
rect 18199 64732 281049 65045
rect 18199 64601 164818 64732
rect 18199 64600 69760 64601
rect 18199 64599 62802 64600
rect 18199 64595 55837 64599
rect 18199 64594 48920 64595
rect 18199 64593 28077 64594
rect 18199 63411 21119 64593
rect 22243 63412 28077 64593
rect 29201 64593 41962 64594
rect 29201 63412 34997 64593
rect 22243 63411 34997 63412
rect 36121 63412 41962 64593
rect 43086 63413 48920 64594
rect 50044 63417 55837 64595
rect 56961 63418 62802 64599
rect 63926 63419 69760 64600
rect 70884 64600 90600 64601
rect 70884 64599 83642 64600
rect 70884 63419 76677 64599
rect 63926 63418 76677 63419
rect 56961 63417 76677 63418
rect 77801 63418 83642 64599
rect 84766 63419 90600 64600
rect 91724 64589 164818 64601
rect 91724 64588 153024 64589
rect 91724 64587 146066 64588
rect 91724 64583 139101 64587
rect 91724 64582 132184 64583
rect 91724 64581 111341 64582
rect 91724 64580 104383 64581
rect 91724 63419 97418 64580
rect 84766 63418 97418 63419
rect 77801 63417 97418 63418
rect 50044 63413 97418 63417
rect 43086 63412 97418 63413
rect 36121 63411 97418 63412
rect 18199 63398 97418 63411
rect 98542 63399 104383 64580
rect 105507 63400 111341 64581
rect 112465 64581 125226 64582
rect 112465 63400 118261 64581
rect 105507 63399 118261 63400
rect 119385 63400 125226 64581
rect 126350 63401 132184 64582
rect 133308 63405 139101 64583
rect 140225 63406 146066 64587
rect 147190 63407 153024 64588
rect 154148 64587 164818 64589
rect 154148 63407 159941 64587
rect 147190 63406 159941 63407
rect 140225 63405 159941 63406
rect 161065 63557 164818 64587
rect 166084 64592 281049 64732
rect 166084 64591 271213 64592
rect 166084 64590 236275 64591
rect 166084 64589 229317 64590
rect 166084 64588 173864 64589
rect 166084 63557 166906 64588
rect 161065 63406 166906 63557
rect 168030 63407 173864 64588
rect 174988 64585 222352 64589
rect 174988 64584 215435 64585
rect 174988 64583 194592 64584
rect 174988 64582 187634 64583
rect 174988 63407 180669 64582
rect 168030 63406 180669 63407
rect 161065 63405 180669 63406
rect 133308 63401 180669 63405
rect 126350 63400 180669 63401
rect 181793 63401 187634 64582
rect 188758 63402 194592 64583
rect 195716 64583 208477 64584
rect 195716 63402 201512 64583
rect 188758 63401 201512 63402
rect 202636 63402 208477 64583
rect 209601 63403 215435 64584
rect 216559 63407 222352 64585
rect 223476 63408 229317 64589
rect 230441 63409 236275 64590
rect 237399 64590 257115 64591
rect 237399 64589 250157 64590
rect 237399 63409 243192 64589
rect 230441 63408 243192 63409
rect 223476 63407 243192 63408
rect 244316 63408 250157 64589
rect 251281 63409 257115 64590
rect 258239 63409 264255 64591
rect 265379 63410 271213 64591
rect 272337 64582 281049 64592
rect 272337 63410 278349 64582
rect 265379 63409 278349 63410
rect 251281 63408 278349 63409
rect 244316 63407 278349 63408
rect 216559 63403 278349 63407
rect 209601 63402 278349 63403
rect 202636 63401 278349 63402
rect 181793 63400 278349 63401
rect 279473 63400 281049 64582
rect 119385 63399 281049 63400
rect 98542 63398 281049 63399
rect 18199 62995 281049 63398
rect 18199 62976 280006 62995
rect 31059 59366 33149 62976
rect 58830 59627 60920 62976
rect 58830 59366 60924 59627
rect 100767 59366 102857 62976
rect 141638 59366 143728 62976
rect 189973 59627 192063 62976
rect 189973 59366 192123 59627
rect 232337 59366 234427 62976
rect 267450 59627 269540 62976
rect 267359 59366 269540 59627
rect 18164 59328 279971 59366
rect 18164 58904 281014 59328
rect 18164 58884 164855 58904
rect 18164 58883 69725 58884
rect 18164 58882 62767 58883
rect 18164 58878 55802 58882
rect 18164 58877 48885 58878
rect 18164 58876 28042 58877
rect 18164 57694 21084 58876
rect 22208 57695 28042 58876
rect 29166 58876 41927 58877
rect 29166 57695 34962 58876
rect 22208 57694 34962 57695
rect 36086 57695 41927 58876
rect 43051 57696 48885 58877
rect 50009 57700 55802 58878
rect 56926 57701 62767 58882
rect 63891 57702 69725 58883
rect 70849 58883 90565 58884
rect 70849 58882 83607 58883
rect 70849 57702 76642 58882
rect 63891 57701 76642 57702
rect 56926 57700 76642 57701
rect 77766 57701 83607 58882
rect 84731 57702 90565 58883
rect 91689 58872 164855 58884
rect 91689 58871 152989 58872
rect 91689 58870 146031 58871
rect 91689 58866 139066 58870
rect 91689 58865 132149 58866
rect 91689 58864 111306 58865
rect 91689 58863 104348 58864
rect 91689 57702 97383 58863
rect 84731 57701 97383 57702
rect 77766 57700 97383 57701
rect 50009 57696 97383 57700
rect 43051 57695 97383 57696
rect 36086 57694 97383 57695
rect 18164 57681 97383 57694
rect 98507 57682 104348 58863
rect 105472 57683 111306 58864
rect 112430 58864 125191 58865
rect 112430 57683 118226 58864
rect 105472 57682 118226 57683
rect 119350 57683 125191 58864
rect 126315 57684 132149 58865
rect 133273 57688 139066 58866
rect 140190 57689 146031 58870
rect 147155 57690 152989 58871
rect 154113 58870 164855 58872
rect 154113 57690 159906 58870
rect 147155 57689 159906 57690
rect 140190 57688 159906 57689
rect 161030 57729 164855 58870
rect 166121 58875 281014 58904
rect 166121 58874 271178 58875
rect 166121 58873 236240 58874
rect 166121 58872 229282 58873
rect 166121 58871 173829 58872
rect 166121 57729 166871 58871
rect 161030 57689 166871 57729
rect 167995 57690 173829 58871
rect 174953 58868 222317 58872
rect 174953 58867 215400 58868
rect 174953 58866 194557 58867
rect 174953 58865 187599 58866
rect 174953 57690 180634 58865
rect 167995 57689 180634 57690
rect 161030 57688 180634 57689
rect 133273 57684 180634 57688
rect 126315 57683 180634 57684
rect 181758 57684 187599 58865
rect 188723 57685 194557 58866
rect 195681 58866 208442 58867
rect 195681 57685 201477 58866
rect 188723 57684 201477 57685
rect 202601 57685 208442 58866
rect 209566 57686 215400 58867
rect 216524 57690 222317 58868
rect 223441 57691 229282 58872
rect 230406 57692 236240 58873
rect 237364 58873 257080 58874
rect 237364 58872 250122 58873
rect 237364 57692 243157 58872
rect 230406 57691 243157 57692
rect 223441 57690 243157 57691
rect 244281 57691 250122 58872
rect 251246 57692 257080 58873
rect 258204 57692 264220 58874
rect 265344 57693 271178 58874
rect 272302 58865 281014 58875
rect 272302 57693 278314 58865
rect 265344 57692 278314 57693
rect 251246 57691 278314 57692
rect 244281 57690 278314 57691
rect 216524 57686 278314 57690
rect 209566 57685 278314 57686
rect 202601 57684 278314 57685
rect 181758 57683 278314 57684
rect 279438 57683 281014 58865
rect 119350 57682 281014 57683
rect 98507 57681 281014 57682
rect 18164 57278 281014 57681
rect 18164 57259 279971 57278
rect 31059 53161 33149 57259
rect 58830 53161 60920 57259
rect 100767 53161 102857 57259
rect 141638 53422 143728 57259
rect 141581 53161 143728 53422
rect 189973 53161 192063 57259
rect 232337 53161 234427 57259
rect 267450 53422 269540 57259
rect 267290 53161 269540 53422
rect 18095 53123 279902 53161
rect 18095 52817 280945 53123
rect 18095 52679 164929 52817
rect 18095 52678 69656 52679
rect 18095 52677 62698 52678
rect 18095 52673 55733 52677
rect 18095 52672 48816 52673
rect 18095 52671 27973 52672
rect 18095 51489 21015 52671
rect 22139 51490 27973 52671
rect 29097 52671 41858 52672
rect 29097 51490 34893 52671
rect 22139 51489 34893 51490
rect 36017 51490 41858 52671
rect 42982 51491 48816 52672
rect 49940 51495 55733 52673
rect 56857 51496 62698 52677
rect 63822 51497 69656 52678
rect 70780 52678 90496 52679
rect 70780 52677 83538 52678
rect 70780 51497 76573 52677
rect 63822 51496 76573 51497
rect 56857 51495 76573 51496
rect 77697 51496 83538 52677
rect 84662 51497 90496 52678
rect 91620 52667 164929 52679
rect 91620 52666 152920 52667
rect 91620 52665 145962 52666
rect 91620 52661 138997 52665
rect 91620 52660 132080 52661
rect 91620 52659 111237 52660
rect 91620 52658 104279 52659
rect 91620 51497 97314 52658
rect 84662 51496 97314 51497
rect 77697 51495 97314 51496
rect 49940 51491 97314 51495
rect 42982 51490 97314 51491
rect 36017 51489 97314 51490
rect 18095 51476 97314 51489
rect 98438 51477 104279 52658
rect 105403 51478 111237 52659
rect 112361 52659 125122 52660
rect 112361 51478 118157 52659
rect 105403 51477 118157 51478
rect 119281 51478 125122 52659
rect 126246 51479 132080 52660
rect 133204 51483 138997 52661
rect 140121 51484 145962 52665
rect 147086 51485 152920 52666
rect 154044 52665 164929 52667
rect 154044 51485 159837 52665
rect 147086 51484 159837 51485
rect 140121 51483 159837 51484
rect 160961 51642 164929 52665
rect 166195 52670 280945 52817
rect 166195 52669 271109 52670
rect 166195 52668 236171 52669
rect 166195 52667 229213 52668
rect 166195 52666 173760 52667
rect 166195 51642 166802 52666
rect 160961 51484 166802 51642
rect 167926 51485 173760 52666
rect 174884 52663 222248 52667
rect 174884 52662 215331 52663
rect 174884 52661 194488 52662
rect 174884 52660 187530 52661
rect 174884 51485 180565 52660
rect 167926 51484 180565 51485
rect 160961 51483 180565 51484
rect 133204 51479 180565 51483
rect 126246 51478 180565 51479
rect 181689 51479 187530 52660
rect 188654 51480 194488 52661
rect 195612 52661 208373 52662
rect 195612 51480 201408 52661
rect 188654 51479 201408 51480
rect 202532 51480 208373 52661
rect 209497 51481 215331 52662
rect 216455 51485 222248 52663
rect 223372 51486 229213 52667
rect 230337 51487 236171 52668
rect 237295 52668 257011 52669
rect 237295 52667 250053 52668
rect 237295 51487 243088 52667
rect 230337 51486 243088 51487
rect 223372 51485 243088 51486
rect 244212 51486 250053 52667
rect 251177 51487 257011 52668
rect 258135 51487 264151 52669
rect 265275 51488 271109 52669
rect 272233 52660 280945 52670
rect 272233 51488 278245 52660
rect 265275 51487 278245 51488
rect 251177 51486 278245 51487
rect 244212 51485 278245 51486
rect 216455 51481 278245 51485
rect 209497 51480 278245 51481
rect 202532 51479 278245 51480
rect 181689 51478 278245 51479
rect 279369 51478 280945 52660
rect 119281 51477 280945 51478
rect 98438 51476 280945 51477
rect 18095 51073 280945 51476
rect 18095 51054 279902 51073
rect 100312 46276 102598 51054
rect 100312 45303 102638 46276
rect 141218 45303 143504 51054
rect 189692 45476 191978 51054
rect 189685 45303 191978 45476
rect 231872 45303 234143 51054
rect 266830 45303 269345 51054
rect 66199 45300 100228 45303
rect 100312 45300 279614 45303
rect 66199 45265 279614 45300
rect 66199 44959 280657 45265
rect 27245 44887 27349 44898
rect 27245 44794 27254 44887
rect 27342 44794 27349 44887
rect 27245 44788 27349 44794
rect 66199 44821 164641 44959
rect 36700 43332 37109 44326
rect 38160 43332 38569 44370
rect 39718 43332 40127 44397
rect 41748 43332 42157 44370
rect 43387 43332 43796 44353
rect 36700 42847 43796 43332
rect 66199 43639 69368 44821
rect 70492 44820 90208 44821
rect 70492 44819 83250 44820
rect 70492 43639 76285 44819
rect 66199 43637 76285 43639
rect 77409 43638 83250 44819
rect 84374 43639 90208 44820
rect 91332 44809 164641 44821
rect 91332 44808 152632 44809
rect 91332 44807 145674 44808
rect 91332 44803 138709 44807
rect 91332 44802 131792 44803
rect 91332 44801 110949 44802
rect 91332 44800 103991 44801
rect 91332 43639 97026 44800
rect 84374 43638 97026 43639
rect 77409 43637 97026 43638
rect 66199 43618 97026 43637
rect 98150 43619 103991 44800
rect 105115 43620 110949 44801
rect 112073 44801 124834 44802
rect 112073 43620 117869 44801
rect 105115 43619 117869 43620
rect 118993 43620 124834 44801
rect 125958 43621 131792 44802
rect 132916 43625 138709 44803
rect 139833 43626 145674 44807
rect 146798 43627 152632 44808
rect 153756 44807 164641 44809
rect 153756 43627 159549 44807
rect 146798 43626 159549 43627
rect 139833 43625 159549 43626
rect 160673 43784 164641 44807
rect 165907 44812 280657 44959
rect 165907 44811 270821 44812
rect 165907 44810 235883 44811
rect 165907 44809 228925 44810
rect 165907 44808 173472 44809
rect 165907 43784 166514 44808
rect 160673 43626 166514 43784
rect 167638 43627 173472 44808
rect 174596 44805 221960 44809
rect 174596 44804 215043 44805
rect 174596 44803 194200 44804
rect 174596 44802 187242 44803
rect 174596 43627 180277 44802
rect 167638 43626 180277 43627
rect 160673 43625 180277 43626
rect 132916 43621 180277 43625
rect 125958 43620 180277 43621
rect 181401 43621 187242 44802
rect 188366 43622 194200 44803
rect 195324 44803 208085 44804
rect 195324 43622 201120 44803
rect 188366 43621 201120 43622
rect 202244 43622 208085 44803
rect 209209 43623 215043 44804
rect 216167 43627 221960 44805
rect 223084 43628 228925 44809
rect 230049 43629 235883 44810
rect 237007 44810 256723 44811
rect 237007 44809 249765 44810
rect 237007 43629 242800 44809
rect 230049 43628 242800 43629
rect 223084 43627 242800 43628
rect 243924 43628 249765 44809
rect 250889 43629 256723 44810
rect 257847 43629 263863 44811
rect 264987 43630 270821 44811
rect 271945 44802 280657 44812
rect 271945 43630 277957 44802
rect 264987 43629 277957 43630
rect 250889 43628 277957 43629
rect 243924 43627 277957 43628
rect 216167 43623 277957 43627
rect 209209 43622 277957 43623
rect 202244 43621 277957 43622
rect 181401 43620 277957 43621
rect 279081 43620 280657 44802
rect 118993 43619 280657 43620
rect 98150 43618 280657 43619
rect 66199 43215 280657 43618
rect 66199 43196 279614 43215
rect 36700 41468 37109 42847
rect 38160 41512 38569 42847
rect 39718 41539 40127 42847
rect 41748 41512 42157 42847
rect 43387 41495 43796 42847
rect 100312 39818 102638 43196
rect 100312 39009 102642 39818
rect 141218 39009 143504 43196
rect 189615 42901 191978 43196
rect 189692 39182 191978 42901
rect 189685 39009 191978 39182
rect 231872 39009 234143 43196
rect 266830 39009 269345 43196
rect 66199 39006 100228 39009
rect 100312 39006 279614 39009
rect 66199 38971 279614 39006
rect 66199 38665 280657 38971
rect 66199 38527 164641 38665
rect 66199 37345 69368 38527
rect 70492 38526 90208 38527
rect 70492 38525 83250 38526
rect 70492 37345 76285 38525
rect 66199 37343 76285 37345
rect 77409 37344 83250 38525
rect 84374 37345 90208 38526
rect 91332 38515 164641 38527
rect 91332 38514 152632 38515
rect 91332 38513 145674 38514
rect 91332 38509 138709 38513
rect 91332 38508 131792 38509
rect 91332 38507 110949 38508
rect 91332 38506 103991 38507
rect 91332 37345 97026 38506
rect 84374 37344 97026 37345
rect 77409 37343 97026 37344
rect 66199 37324 97026 37343
rect 98150 37325 103991 38506
rect 105115 37326 110949 38507
rect 112073 38507 124834 38508
rect 112073 37326 117869 38507
rect 105115 37325 117869 37326
rect 118993 37326 124834 38507
rect 125958 37327 131792 38508
rect 132916 37331 138709 38509
rect 139833 37332 145674 38513
rect 146798 37333 152632 38514
rect 153756 38513 164641 38515
rect 153756 37333 159549 38513
rect 146798 37332 159549 37333
rect 139833 37331 159549 37332
rect 160673 37490 164641 38513
rect 165907 38518 280657 38665
rect 165907 38517 270821 38518
rect 165907 38516 235883 38517
rect 165907 38515 228925 38516
rect 165907 38514 173472 38515
rect 165907 37490 166514 38514
rect 160673 37332 166514 37490
rect 167638 37333 173472 38514
rect 174596 38511 221960 38515
rect 174596 38510 215043 38511
rect 174596 38509 194200 38510
rect 174596 38508 187242 38509
rect 174596 37333 180277 38508
rect 167638 37332 180277 37333
rect 160673 37331 180277 37332
rect 132916 37327 180277 37331
rect 125958 37326 180277 37327
rect 181401 37327 187242 38508
rect 188366 37328 194200 38509
rect 195324 38509 208085 38510
rect 195324 37328 201120 38509
rect 188366 37327 201120 37328
rect 202244 37328 208085 38509
rect 209209 37329 215043 38510
rect 216167 37333 221960 38511
rect 223084 37334 228925 38515
rect 230049 37335 235883 38516
rect 237007 38516 256723 38517
rect 237007 38515 249765 38516
rect 237007 37335 242800 38515
rect 230049 37334 242800 37335
rect 223084 37333 242800 37334
rect 243924 37334 249765 38515
rect 250889 37335 256723 38516
rect 257847 37335 263863 38517
rect 264987 37336 270821 38517
rect 271945 38508 280657 38518
rect 271945 37336 277957 38508
rect 264987 37335 277957 37336
rect 250889 37334 277957 37335
rect 243924 37333 277957 37334
rect 216167 37329 277957 37333
rect 209209 37328 277957 37329
rect 202244 37327 277957 37328
rect 181401 37326 277957 37327
rect 279081 37326 280657 38508
rect 118993 37325 280657 37326
rect 98150 37324 280657 37325
rect 66199 36921 280657 37324
rect 66199 36902 279614 36921
rect 100312 32715 102642 36902
rect 141218 32715 143504 36902
rect 189615 36607 191978 36902
rect 189692 32888 191978 36607
rect 189685 32715 191978 32888
rect 231872 32715 234143 36902
rect 266830 32715 269345 36902
rect 66199 32712 100228 32715
rect 100312 32712 279614 32715
rect 66199 32677 279614 32712
rect 66199 32371 280657 32677
rect 66199 32233 164641 32371
rect 66199 31051 69368 32233
rect 70492 32232 90208 32233
rect 70492 32231 83250 32232
rect 70492 31051 76285 32231
rect 66199 31049 76285 31051
rect 77409 31050 83250 32231
rect 84374 31051 90208 32232
rect 91332 32221 164641 32233
rect 91332 32220 152632 32221
rect 91332 32219 145674 32220
rect 91332 32215 138709 32219
rect 91332 32214 131792 32215
rect 91332 32213 110949 32214
rect 91332 32212 103991 32213
rect 91332 31051 97026 32212
rect 84374 31050 97026 31051
rect 77409 31049 97026 31050
rect 66199 31030 97026 31049
rect 98150 31031 103991 32212
rect 105115 31032 110949 32213
rect 112073 32213 124834 32214
rect 112073 31032 117869 32213
rect 105115 31031 117869 31032
rect 118993 31032 124834 32213
rect 125958 31033 131792 32214
rect 132916 31037 138709 32215
rect 139833 31038 145674 32219
rect 146798 31039 152632 32220
rect 153756 32219 164641 32221
rect 153756 31039 159549 32219
rect 146798 31038 159549 31039
rect 139833 31037 159549 31038
rect 160673 31196 164641 32219
rect 165907 32224 280657 32371
rect 165907 32223 270821 32224
rect 165907 32222 235883 32223
rect 165907 32221 228925 32222
rect 165907 32220 173472 32221
rect 165907 31196 166514 32220
rect 160673 31038 166514 31196
rect 167638 31039 173472 32220
rect 174596 32217 221960 32221
rect 174596 32216 215043 32217
rect 174596 32215 194200 32216
rect 174596 32214 187242 32215
rect 174596 31039 180277 32214
rect 167638 31038 180277 31039
rect 160673 31037 180277 31038
rect 132916 31033 180277 31037
rect 125958 31032 180277 31033
rect 181401 31033 187242 32214
rect 188366 31034 194200 32215
rect 195324 32215 208085 32216
rect 195324 31034 201120 32215
rect 188366 31033 201120 31034
rect 202244 31034 208085 32215
rect 209209 31035 215043 32216
rect 216167 31039 221960 32217
rect 223084 31040 228925 32221
rect 230049 31041 235883 32222
rect 237007 32222 256723 32223
rect 237007 32221 249765 32222
rect 237007 31041 242800 32221
rect 230049 31040 242800 31041
rect 223084 31039 242800 31040
rect 243924 31040 249765 32221
rect 250889 31041 256723 32222
rect 257847 31041 263863 32223
rect 264987 31042 270821 32223
rect 271945 32214 280657 32224
rect 271945 31042 277957 32214
rect 264987 31041 277957 31042
rect 250889 31040 277957 31041
rect 243924 31039 277957 31040
rect 216167 31035 277957 31039
rect 209209 31034 277957 31035
rect 202244 31033 277957 31034
rect 181401 31032 277957 31033
rect 279081 31032 280657 32214
rect 118993 31031 280657 31032
rect 98150 31030 280657 31031
rect 66199 30627 280657 31030
rect 66199 30608 279614 30627
rect 17823 22151 30545 22159
rect 34439 22151 58495 22159
rect 17823 22136 58495 22151
rect 60871 22156 100244 22159
rect 100312 22156 102598 30608
rect 141218 22159 143504 30608
rect 189615 30313 191978 30608
rect 189692 22159 191978 30313
rect 231872 22332 234143 30608
rect 231872 22159 234155 22332
rect 266830 22159 269345 30608
rect 102620 22156 279630 22159
rect 60871 22136 279630 22156
rect 17823 22121 279630 22136
rect 17823 21815 280673 22121
rect 17823 21677 164657 21815
rect 17823 21676 69384 21677
rect 17823 21675 62426 21676
rect 17823 21671 55461 21675
rect 17823 21670 48544 21671
rect 17823 21669 27701 21670
rect 17823 20487 20743 21669
rect 21867 20488 27701 21669
rect 28825 21669 41586 21670
rect 28825 20488 34621 21669
rect 21867 20487 34621 20488
rect 35745 20488 41586 21669
rect 42710 20489 48544 21670
rect 49668 20493 55461 21671
rect 56585 20494 62426 21675
rect 63550 20495 69384 21676
rect 70508 21676 90224 21677
rect 70508 21675 83266 21676
rect 70508 20495 76301 21675
rect 63550 20494 76301 20495
rect 56585 20493 76301 20494
rect 77425 20494 83266 21675
rect 84390 20495 90224 21676
rect 91348 21665 164657 21677
rect 91348 21664 152648 21665
rect 91348 21663 145690 21664
rect 91348 21659 138725 21663
rect 91348 21658 131808 21659
rect 91348 21657 110965 21658
rect 91348 21656 104007 21657
rect 91348 20495 97042 21656
rect 84390 20494 97042 20495
rect 77425 20493 97042 20494
rect 49668 20489 97042 20493
rect 42710 20488 97042 20489
rect 35745 20487 97042 20488
rect 17823 20474 97042 20487
rect 98166 20475 104007 21656
rect 105131 20476 110965 21657
rect 112089 21657 124850 21658
rect 112089 20476 117885 21657
rect 105131 20475 117885 20476
rect 119009 20476 124850 21657
rect 125974 20477 131808 21658
rect 132932 20481 138725 21659
rect 139849 20482 145690 21663
rect 146814 20483 152648 21664
rect 153772 21663 164657 21665
rect 153772 20483 159565 21663
rect 146814 20482 159565 20483
rect 139849 20481 159565 20482
rect 160689 20640 164657 21663
rect 165923 21668 280673 21815
rect 165923 21667 270837 21668
rect 165923 21666 235899 21667
rect 165923 21665 228941 21666
rect 165923 21664 173488 21665
rect 165923 20640 166530 21664
rect 160689 20482 166530 20640
rect 167654 20483 173488 21664
rect 174612 21661 221976 21665
rect 174612 21660 215059 21661
rect 174612 21659 194216 21660
rect 174612 21658 187258 21659
rect 174612 20483 180293 21658
rect 167654 20482 180293 20483
rect 160689 20481 180293 20482
rect 132932 20477 180293 20481
rect 125974 20476 180293 20477
rect 181417 20477 187258 21658
rect 188382 20478 194216 21659
rect 195340 21659 208101 21660
rect 195340 20478 201136 21659
rect 188382 20477 201136 20478
rect 202260 20478 208101 21659
rect 209225 20479 215059 21660
rect 216183 20483 221976 21661
rect 223100 20484 228941 21665
rect 230065 20485 235899 21666
rect 237023 21666 256739 21667
rect 237023 21665 249781 21666
rect 237023 20485 242816 21665
rect 230065 20484 242816 20485
rect 223100 20483 242816 20484
rect 243940 20484 249781 21665
rect 250905 20485 256739 21666
rect 257863 20485 263879 21667
rect 265003 20486 270837 21667
rect 271961 21658 280673 21668
rect 271961 20486 277973 21658
rect 265003 20485 277973 20486
rect 250905 20484 277973 20485
rect 243940 20483 277973 20484
rect 216183 20479 277973 20483
rect 209225 20478 277973 20479
rect 202260 20477 277973 20478
rect 181417 20476 277973 20477
rect 279097 20476 280673 21658
rect 119009 20475 280673 20476
rect 98166 20474 280673 20475
rect 17823 20071 280673 20474
rect 17823 20052 279630 20071
rect 30633 16654 32837 20052
rect 30633 16481 32861 16654
rect 58459 16481 60770 20052
rect 100312 19359 102598 20052
rect 141218 19404 143504 20052
rect 100414 16481 102573 19359
rect 141287 16481 143446 19404
rect 189631 16481 191790 20052
rect 231962 16654 234121 20052
rect 231962 16481 234139 16654
rect 266893 16481 269285 20052
rect 17807 16443 279614 16481
rect 17807 16137 280657 16443
rect 17807 15999 164641 16137
rect 17807 15998 69368 15999
rect 17807 15997 62410 15998
rect 17807 15993 55445 15997
rect 17807 15992 48528 15993
rect 17807 15991 27685 15992
rect 17807 14809 20727 15991
rect 21851 14810 27685 15991
rect 28809 15991 41570 15992
rect 28809 14810 34605 15991
rect 21851 14809 34605 14810
rect 35729 14810 41570 15991
rect 42694 14811 48528 15992
rect 49652 14815 55445 15993
rect 56569 14816 62410 15997
rect 63534 14817 69368 15998
rect 70492 15998 90208 15999
rect 70492 15997 83250 15998
rect 70492 14817 76285 15997
rect 63534 14816 76285 14817
rect 56569 14815 76285 14816
rect 77409 14816 83250 15997
rect 84374 14817 90208 15998
rect 91332 15987 164641 15999
rect 91332 15986 152632 15987
rect 91332 15985 145674 15986
rect 91332 15981 138709 15985
rect 91332 15980 131792 15981
rect 91332 15979 110949 15980
rect 91332 15978 103991 15979
rect 91332 14817 97026 15978
rect 84374 14816 97026 14817
rect 77409 14815 97026 14816
rect 49652 14811 97026 14815
rect 42694 14810 97026 14811
rect 35729 14809 97026 14810
rect 17807 14796 97026 14809
rect 98150 14797 103991 15978
rect 105115 14798 110949 15979
rect 112073 15979 124834 15980
rect 112073 14798 117869 15979
rect 105115 14797 117869 14798
rect 118993 14798 124834 15979
rect 125958 14799 131792 15980
rect 132916 14803 138709 15981
rect 139833 14804 145674 15985
rect 146798 14805 152632 15986
rect 153756 15985 164641 15987
rect 153756 14805 159549 15985
rect 146798 14804 159549 14805
rect 139833 14803 159549 14804
rect 160673 14962 164641 15985
rect 165907 15990 280657 16137
rect 165907 15989 270821 15990
rect 165907 15988 235883 15989
rect 165907 15987 228925 15988
rect 165907 15986 173472 15987
rect 165907 14962 166514 15986
rect 160673 14804 166514 14962
rect 167638 14805 173472 15986
rect 174596 15983 221960 15987
rect 174596 15982 215043 15983
rect 174596 15981 194200 15982
rect 174596 15980 187242 15981
rect 174596 14805 180277 15980
rect 167638 14804 180277 14805
rect 160673 14803 180277 14804
rect 132916 14799 180277 14803
rect 125958 14798 180277 14799
rect 181401 14799 187242 15980
rect 188366 14800 194200 15981
rect 195324 15981 208085 15982
rect 195324 14800 201120 15981
rect 188366 14799 201120 14800
rect 202244 14800 208085 15981
rect 209209 14801 215043 15982
rect 216167 14805 221960 15983
rect 223084 14806 228925 15987
rect 230049 14807 235883 15988
rect 237007 15988 256723 15989
rect 237007 15987 249765 15988
rect 237007 14807 242800 15987
rect 230049 14806 242800 14807
rect 223084 14805 242800 14806
rect 243924 14806 249765 15987
rect 250889 14807 256723 15988
rect 257847 14807 263863 15989
rect 264987 14808 270821 15989
rect 271945 15980 280657 15990
rect 271945 14808 277957 15980
rect 264987 14807 277957 14808
rect 250889 14806 277957 14807
rect 243924 14805 277957 14806
rect 216167 14801 277957 14805
rect 209209 14800 277957 14801
rect 202244 14799 277957 14800
rect 181401 14798 277957 14799
rect 279081 14798 280657 15980
rect 118993 14797 280657 14798
rect 98150 14796 280657 14797
rect 17807 14393 280657 14796
rect 17807 14374 279614 14393
rect 30633 9561 32837 14374
rect 30633 9388 32861 9561
rect 58459 9388 60770 14374
rect 100414 9388 102573 14374
rect 141287 9388 143446 14374
rect 189631 9388 191790 14374
rect 231962 9561 234121 14374
rect 231962 9388 234139 9561
rect 266893 9388 269285 14374
rect 17807 9350 279614 9388
rect 17807 9044 280657 9350
rect 17807 8906 164641 9044
rect 17807 8905 69368 8906
rect 17807 8904 62410 8905
rect 17807 8900 55445 8904
rect 17807 8899 48528 8900
rect 17807 8898 27685 8899
rect 17807 7716 20727 8898
rect 21851 7717 27685 8898
rect 28809 8898 41570 8899
rect 28809 7717 34605 8898
rect 21851 7716 34605 7717
rect 35729 7717 41570 8898
rect 42694 7718 48528 8899
rect 49652 7722 55445 8900
rect 56569 7723 62410 8904
rect 63534 7724 69368 8905
rect 70492 8905 90208 8906
rect 70492 8904 83250 8905
rect 70492 7724 76285 8904
rect 63534 7723 76285 7724
rect 56569 7722 76285 7723
rect 77409 7723 83250 8904
rect 84374 7724 90208 8905
rect 91332 8894 164641 8906
rect 91332 8893 152632 8894
rect 91332 8892 145674 8893
rect 91332 8888 138709 8892
rect 91332 8887 131792 8888
rect 91332 8886 110949 8887
rect 91332 8885 103991 8886
rect 91332 7724 97026 8885
rect 84374 7723 97026 7724
rect 77409 7722 97026 7723
rect 49652 7718 97026 7722
rect 42694 7717 97026 7718
rect 35729 7716 97026 7717
rect 17807 7703 97026 7716
rect 98150 7704 103991 8885
rect 105115 7705 110949 8886
rect 112073 8886 124834 8887
rect 112073 7705 117869 8886
rect 105115 7704 117869 7705
rect 118993 7705 124834 8886
rect 125958 7706 131792 8887
rect 132916 7710 138709 8888
rect 139833 7711 145674 8892
rect 146798 7712 152632 8893
rect 153756 8892 164641 8894
rect 153756 7712 159549 8892
rect 146798 7711 159549 7712
rect 139833 7710 159549 7711
rect 160673 7869 164641 8892
rect 165907 8897 280657 9044
rect 165907 8896 270821 8897
rect 165907 8895 235883 8896
rect 165907 8894 228925 8895
rect 165907 8893 173472 8894
rect 165907 7869 166514 8893
rect 160673 7711 166514 7869
rect 167638 7712 173472 8893
rect 174596 8890 221960 8894
rect 174596 8889 215043 8890
rect 174596 8888 194200 8889
rect 174596 8887 187242 8888
rect 174596 7712 180277 8887
rect 167638 7711 180277 7712
rect 160673 7710 180277 7711
rect 132916 7706 180277 7710
rect 125958 7705 180277 7706
rect 181401 7706 187242 8887
rect 188366 7707 194200 8888
rect 195324 8888 208085 8889
rect 195324 7707 201120 8888
rect 188366 7706 201120 7707
rect 202244 7707 208085 8888
rect 209209 7708 215043 8889
rect 216167 7712 221960 8890
rect 223084 7713 228925 8894
rect 230049 7714 235883 8895
rect 237007 8895 256723 8896
rect 237007 8894 249765 8895
rect 237007 7714 242800 8894
rect 230049 7713 242800 7714
rect 223084 7712 242800 7713
rect 243924 7713 249765 8894
rect 250889 7714 256723 8895
rect 257847 7714 263863 8896
rect 264987 7715 270821 8896
rect 271945 8887 280657 8897
rect 271945 7715 277957 8887
rect 264987 7714 277957 7715
rect 250889 7713 277957 7714
rect 243924 7712 277957 7713
rect 216167 7708 277957 7712
rect 209209 7707 277957 7708
rect 202244 7706 277957 7707
rect 181401 7705 277957 7706
rect 279081 7705 280657 8887
rect 118993 7704 280657 7705
rect 98150 7703 280657 7704
rect 17807 7300 280657 7703
rect 17807 7281 279614 7300
<< viali >>
rect 164500 338774 165766 339949
rect 164481 331688 165747 332863
rect 247701 329822 247772 329890
rect 247459 329454 247560 329554
rect 164500 325316 165766 326491
rect 164481 318230 165747 319405
rect 25928 316894 25978 316944
rect 25937 316693 25987 316743
rect 25922 316004 25972 316054
rect 25928 315653 25978 315703
rect 164506 311055 165772 312230
rect 244859 318306 244934 318388
rect 245922 318310 245997 318392
rect 244653 315856 244728 315938
rect 245828 315851 245903 315933
rect 244435 313491 244510 313573
rect 245762 313467 245837 313549
rect 244203 311007 244278 311089
rect 245677 311004 245752 311086
rect 243961 308605 244036 308687
rect 245602 308628 245677 308710
rect 243716 306147 243791 306229
rect 245522 306153 245597 306235
rect 164487 303969 165753 305144
rect 164595 294696 165861 295871
rect 164576 287610 165842 288785
rect 164539 281208 165805 282383
rect 164646 272288 165912 273463
rect 164627 265202 165893 266377
rect 266024 265202 266126 265300
rect 26446 264665 26561 264775
rect 23597 264330 23716 264447
rect 265944 262844 266046 262942
rect 265865 260359 265967 260457
rect 164590 258800 165856 259975
rect 164677 248034 165943 249209
rect 164658 240948 165924 242123
rect 242684 240947 242756 241013
rect 63189 240105 63304 240219
rect 63110 237769 63225 237883
rect 63029 235285 63144 235399
rect 164621 234546 165887 235721
rect 63033 233078 63148 233192
rect 164801 227768 166067 228943
rect 164781 221906 166047 223081
rect 164821 209843 166087 211018
rect 164802 202757 166068 203932
rect 164765 196355 166031 197530
rect 164808 191950 166074 193125
rect 61518 186400 61626 186500
rect 164789 184864 166055 186039
rect 61438 183977 61546 184077
rect 61359 181493 61467 181593
rect 61360 179342 61468 179442
rect 164752 178462 166018 179637
rect 164612 172537 165878 173712
rect 164575 166135 165841 167310
rect 164841 158874 166107 160049
rect 164822 154034 166088 155209
rect 164803 148764 166069 149939
rect 164785 143212 166051 144387
rect 269050 142679 269160 142783
rect 268969 140283 269079 140387
rect 164785 137022 166051 138197
rect 268890 137823 269000 137927
rect 164793 117918 166059 119093
rect 164902 109991 166168 111166
rect 165003 101789 166269 102964
rect 164966 94290 166232 95465
rect 164947 87204 166213 88379
rect 164910 80802 166176 81977
rect 164892 69552 166158 70727
rect 164818 63557 166084 64732
rect 164855 57729 166121 58904
rect 164929 51642 166195 52817
rect 27254 44794 27342 44887
rect 164641 43784 165907 44959
rect 164641 37490 165907 38665
rect 164641 31196 165907 32371
rect 164657 20640 165923 21815
rect 164641 14962 165907 16137
rect 164641 7869 165907 9044
<< metal1 >>
rect 164427 339949 165848 340032
rect 164427 338774 164500 339949
rect 165766 338774 165848 339949
rect 164427 338683 165848 338774
rect 164408 332863 165829 332946
rect 164408 331688 164481 332863
rect 165747 331688 165829 332863
rect 164408 331597 165829 331688
rect 247694 329890 247780 329899
rect 247694 329822 247701 329890
rect 247772 329822 247780 329890
rect 247694 329815 247780 329822
rect 247445 329554 247576 329570
rect 247445 329454 247459 329554
rect 247560 329454 247576 329554
rect 247445 329439 247576 329454
rect 164427 326491 165848 326574
rect 164427 325316 164500 326491
rect 165766 325316 165848 326491
rect 164427 325225 165848 325316
rect 164408 319405 165829 319488
rect 164408 318230 164481 319405
rect 165747 318230 165829 319405
rect 244825 318392 246016 318414
rect 244825 318388 245922 318392
rect 244825 318306 244859 318388
rect 244934 318310 245922 318388
rect 245997 318310 246016 318392
rect 244934 318306 246016 318310
rect 244825 318282 246016 318306
rect 164408 318139 165829 318230
rect 25918 316944 25988 316954
rect 25918 316894 25928 316944
rect 25978 316894 25988 316944
rect 25918 316884 25988 316894
rect 25927 316743 25997 316753
rect 25927 316693 25937 316743
rect 25987 316693 25997 316743
rect 25927 316683 25997 316693
rect 25912 316054 25982 316064
rect 25912 316004 25922 316054
rect 25972 316004 25982 316054
rect 25912 315994 25982 316004
rect 244622 315938 245929 315985
rect 244622 315856 244653 315938
rect 244728 315933 245929 315938
rect 244728 315856 245828 315933
rect 244622 315851 245828 315856
rect 245903 315851 245929 315933
rect 244622 315815 245929 315851
rect 25918 315703 25988 315713
rect 25918 315653 25928 315703
rect 25978 315653 25988 315703
rect 25918 315643 25988 315653
rect 244395 313573 245853 313599
rect 244395 313491 244435 313573
rect 244510 313549 245853 313573
rect 244510 313491 245762 313549
rect 244395 313467 245762 313491
rect 245837 313467 245853 313549
rect 244395 313434 245853 313467
rect 164433 312230 165854 312313
rect 164433 311055 164506 312230
rect 165772 311055 165854 312230
rect 164433 310964 165854 311055
rect 244145 311089 245782 311155
rect 244145 311007 244203 311089
rect 244278 311086 245782 311089
rect 244278 311007 245677 311086
rect 244145 311004 245677 311007
rect 245752 311004 245782 311086
rect 244145 310972 245782 311004
rect 243931 308710 245701 308760
rect 243931 308687 245602 308710
rect 243931 308605 243961 308687
rect 244036 308628 245602 308687
rect 245677 308628 245701 308710
rect 244036 308605 245701 308628
rect 243931 308542 245701 308605
rect 243681 306235 245612 306299
rect 243681 306229 245522 306235
rect 243681 306147 243716 306229
rect 243791 306153 245522 306229
rect 245597 306153 245612 306235
rect 243791 306147 245612 306153
rect 243681 306085 245612 306147
rect 164414 305144 165835 305227
rect 164414 303969 164487 305144
rect 165753 303969 165835 305144
rect 164414 303878 165835 303969
rect 164522 295871 165943 295954
rect 164522 294696 164595 295871
rect 165861 294696 165943 295871
rect 164522 294605 165943 294696
rect 164503 288785 165924 288868
rect 164503 287610 164576 288785
rect 165842 287610 165924 288785
rect 164503 287519 165924 287610
rect 164466 282383 165887 282466
rect 164466 281208 164539 282383
rect 165805 281208 165887 282383
rect 164466 281117 165887 281208
rect 164573 273463 165994 273546
rect 164573 272288 164646 273463
rect 165912 272288 165994 273463
rect 164573 272197 165994 272288
rect 164554 266377 165975 266460
rect 164554 265202 164627 266377
rect 165893 265202 165975 266377
rect 164554 265111 165975 265202
rect 266017 265300 266133 265309
rect 266017 265202 266024 265300
rect 266126 265202 266133 265300
rect 266017 265191 266133 265202
rect 26436 264775 26571 264785
rect 26436 264665 26446 264775
rect 26561 264665 26571 264775
rect 26436 264660 26571 264665
rect 23581 264447 23730 264462
rect 23581 264330 23597 264447
rect 23716 264330 23730 264447
rect 23581 264315 23730 264330
rect 265937 262942 266053 262951
rect 265937 262844 265944 262942
rect 266046 262844 266053 262942
rect 265937 262833 266053 262844
rect 265858 260457 265974 260466
rect 265858 260359 265865 260457
rect 265967 260359 265974 260457
rect 265858 260348 265974 260359
rect 164517 259975 165938 260058
rect 164517 258800 164590 259975
rect 165856 258800 165938 259975
rect 164517 258709 165938 258800
rect 164604 249209 166025 249292
rect 164604 248034 164677 249209
rect 165943 248034 166025 249209
rect 164604 247943 166025 248034
rect 164585 242123 166006 242206
rect 164585 240948 164658 242123
rect 165924 240948 166006 242123
rect 164585 240857 166006 240948
rect 242679 241013 242763 241022
rect 242679 240947 242684 241013
rect 242756 240947 242763 241013
rect 242679 240939 242763 240947
rect 63180 240219 63315 240230
rect 63180 240105 63189 240219
rect 63304 240105 63315 240219
rect 63180 240095 63315 240105
rect 63101 237883 63236 237894
rect 63101 237769 63110 237883
rect 63225 237769 63236 237883
rect 63101 237759 63236 237769
rect 164548 235721 165969 235804
rect 63020 235399 63155 235410
rect 63020 235285 63029 235399
rect 63144 235285 63155 235399
rect 63020 235275 63155 235285
rect 164548 234546 164621 235721
rect 165887 234546 165969 235721
rect 164548 234455 165969 234546
rect 63024 233192 63159 233203
rect 63024 233078 63033 233192
rect 63148 233078 63159 233192
rect 63024 233068 63159 233078
rect 164728 228943 166149 229026
rect 164728 227768 164801 228943
rect 166067 227768 166149 228943
rect 164728 227677 166149 227768
rect 164708 223081 166129 223164
rect 164708 221906 164781 223081
rect 166047 221906 166129 223081
rect 164708 221815 166129 221906
rect 164748 211018 166169 211101
rect 164748 209843 164821 211018
rect 166087 209843 166169 211018
rect 164748 209752 166169 209843
rect 164729 203932 166150 204015
rect 164729 202757 164802 203932
rect 166068 202757 166150 203932
rect 164729 202666 166150 202757
rect 164692 197530 166113 197613
rect 164692 196355 164765 197530
rect 166031 196355 166113 197530
rect 164692 196264 166113 196355
rect 164735 193125 166156 193208
rect 164735 191950 164808 193125
rect 166074 191950 166156 193125
rect 164735 191859 166156 191950
rect 61507 186500 61636 186511
rect 61507 186400 61518 186500
rect 61626 186400 61636 186500
rect 61507 186389 61636 186400
rect 164716 186039 166137 186122
rect 164716 184864 164789 186039
rect 166055 184864 166137 186039
rect 164716 184773 166137 184864
rect 61427 184077 61556 184088
rect 61427 183977 61438 184077
rect 61546 183977 61556 184077
rect 61427 183966 61556 183977
rect 61348 181593 61477 181604
rect 61348 181493 61359 181593
rect 61467 181493 61477 181593
rect 61348 181482 61477 181493
rect 164679 179637 166100 179720
rect 61349 179442 61478 179453
rect 61349 179342 61360 179442
rect 61468 179342 61478 179442
rect 61349 179331 61478 179342
rect 164679 178462 164752 179637
rect 166018 178462 166100 179637
rect 164679 178371 166100 178462
rect 164539 173712 165960 173795
rect 164539 172537 164612 173712
rect 165878 172537 165960 173712
rect 164539 172446 165960 172537
rect 164502 167310 165923 167393
rect 164502 166135 164575 167310
rect 165841 166135 165923 167310
rect 164502 166044 165923 166135
rect 164768 160049 166189 160132
rect 164768 158874 164841 160049
rect 166107 158874 166189 160049
rect 164768 158783 166189 158874
rect 164749 155209 166170 155292
rect 164749 154034 164822 155209
rect 166088 154034 166170 155209
rect 164749 153943 166170 154034
rect 164730 149939 166151 150022
rect 164730 148764 164803 149939
rect 166069 148764 166151 149939
rect 164730 148673 166151 148764
rect 164712 144387 166133 144470
rect 164712 143212 164785 144387
rect 166051 143212 166133 144387
rect 164712 143121 166133 143212
rect 269038 142783 269176 142796
rect 269038 142679 269050 142783
rect 269160 142679 269176 142783
rect 269038 142667 269176 142679
rect 268957 140387 269095 140400
rect 268957 140283 268969 140387
rect 269079 140283 269095 140387
rect 268957 140271 269095 140283
rect 164712 138197 166133 138280
rect 164712 137022 164785 138197
rect 166051 137022 166133 138197
rect 268878 137927 269016 137940
rect 268878 137823 268890 137927
rect 269000 137823 269016 137927
rect 268878 137811 269016 137823
rect 164712 136931 166133 137022
rect 164720 119093 166141 119176
rect 164720 117918 164793 119093
rect 166059 117918 166141 119093
rect 164720 117827 166141 117918
rect 164829 111166 166250 111249
rect 164829 109991 164902 111166
rect 166168 109991 166250 111166
rect 164829 109900 166250 109991
rect 164930 102964 166351 103047
rect 164930 101789 165003 102964
rect 166269 101789 166351 102964
rect 164930 101698 166351 101789
rect 164893 95465 166314 95548
rect 164893 94290 164966 95465
rect 166232 94290 166314 95465
rect 164893 94199 166314 94290
rect 164874 88379 166295 88462
rect 164874 87204 164947 88379
rect 166213 87204 166295 88379
rect 164874 87113 166295 87204
rect 164837 81977 166258 82060
rect 164837 80802 164910 81977
rect 166176 80802 166258 81977
rect 164837 80711 166258 80802
rect 164819 70727 166240 70810
rect 164819 69552 164892 70727
rect 166158 69552 166240 70727
rect 164819 69461 166240 69552
rect 164745 64732 166166 64815
rect 164745 63557 164818 64732
rect 166084 63557 166166 64732
rect 164745 63466 166166 63557
rect 164782 58904 166203 58987
rect 164782 57729 164855 58904
rect 166121 57729 166203 58904
rect 164782 57638 166203 57729
rect 164856 52817 166277 52900
rect 164856 51642 164929 52817
rect 166195 51642 166277 52817
rect 164856 51551 166277 51642
rect 164568 44959 165989 45042
rect 26613 44887 27349 44921
rect 26613 44794 27254 44887
rect 27342 44794 27349 44887
rect 26613 44778 27349 44794
rect 26616 44748 26821 44778
rect 26618 40297 26821 44748
rect 164568 43784 164641 44959
rect 165907 43784 165989 44959
rect 164568 43693 165989 43784
rect 26618 40296 30982 40297
rect 26618 40291 32860 40296
rect 26618 40290 37181 40291
rect 26618 40115 40438 40290
rect 27767 40114 40438 40115
rect 32817 40109 40438 40114
rect 36074 40108 40438 40109
rect 164568 38665 165989 38748
rect 164568 37490 164641 38665
rect 165907 37490 165989 38665
rect 164568 37399 165989 37490
rect 164568 32371 165989 32454
rect 164568 31196 164641 32371
rect 165907 31196 165989 32371
rect 164568 31105 165989 31196
rect 164584 21815 166005 21898
rect 164584 20640 164657 21815
rect 165923 20640 166005 21815
rect 164584 20549 166005 20640
rect 164517 16137 166098 16247
rect 164517 14962 164641 16137
rect 165907 14962 166098 16137
rect 164517 14797 166098 14962
rect 164568 9044 165989 9127
rect 164568 7869 164641 9044
rect 165907 7869 165989 9044
rect 164568 7778 165989 7869
<< via1 >>
rect 164500 338774 165766 339949
rect 164481 331688 165747 332863
rect 247701 329822 247772 329890
rect 247459 329454 247560 329554
rect 164500 325316 165766 326491
rect 164481 318230 165747 319405
rect 25928 316894 25978 316944
rect 25937 316693 25987 316743
rect 25922 316004 25972 316054
rect 25928 315653 25978 315703
rect 164506 311055 165772 312230
rect 164487 303969 165753 305144
rect 164595 294696 165861 295871
rect 164576 287610 165842 288785
rect 164539 281208 165805 282383
rect 164646 272288 165912 273463
rect 164627 265202 165893 266377
rect 266024 265202 266126 265300
rect 26446 264665 26561 264775
rect 23597 264330 23716 264447
rect 265944 262844 266046 262942
rect 265865 260359 265967 260457
rect 164590 258800 165856 259975
rect 164677 248034 165943 249209
rect 164658 240948 165924 242123
rect 242684 240947 242756 241013
rect 63189 240105 63304 240219
rect 63110 237769 63225 237883
rect 63029 235285 63144 235399
rect 164621 234546 165887 235721
rect 63033 233078 63148 233192
rect 164801 227768 166067 228943
rect 164781 221906 166047 223081
rect 164821 209843 166087 211018
rect 164802 202757 166068 203932
rect 164765 196355 166031 197530
rect 164808 191950 166074 193125
rect 61518 186400 61626 186500
rect 164789 184864 166055 186039
rect 61438 183977 61546 184077
rect 61359 181493 61467 181593
rect 61360 179342 61468 179442
rect 164752 178462 166018 179637
rect 164612 172537 165878 173712
rect 164575 166135 165841 167310
rect 164841 158874 166107 160049
rect 164822 154034 166088 155209
rect 164803 148764 166069 149939
rect 164785 143212 166051 144387
rect 269050 142679 269160 142783
rect 268969 140283 269079 140387
rect 164785 137022 166051 138197
rect 268890 137823 269000 137927
rect 164793 117918 166059 119093
rect 164902 109991 166168 111166
rect 165003 101789 166269 102964
rect 164966 94290 166232 95465
rect 164947 87204 166213 88379
rect 164910 80802 166176 81977
rect 164892 69552 166158 70727
rect 164818 63557 166084 64732
rect 164855 57729 166121 58904
rect 164929 51642 166195 52817
rect 164641 43784 165907 44959
rect 164641 37490 165907 38665
rect 164641 31196 165907 32371
rect 164657 20640 165923 21815
rect 164641 14962 165907 16137
rect 164641 7869 165907 9044
<< metal2 >>
rect 164427 339949 165848 340032
rect 164427 338774 164500 339949
rect 165766 338774 165848 339949
rect 164427 338683 165848 338774
rect 164408 332863 165829 332946
rect 164408 331688 164481 332863
rect 165747 331688 165829 332863
rect 164408 331597 165829 331688
rect 247049 329859 247236 330039
rect 247694 329890 247780 329899
rect 247694 329822 247701 329890
rect 247772 329822 247780 329890
rect 247694 329815 247780 329822
rect 247445 329554 247576 329570
rect 247445 329454 247459 329554
rect 247560 329454 247576 329554
rect 247445 329439 247576 329454
rect 164427 326491 165848 326574
rect 164427 325316 164500 326491
rect 165766 325316 165848 326491
rect 164427 325225 165848 325316
rect 164408 319405 165829 319488
rect 164408 318230 164481 319405
rect 165747 318230 165829 319405
rect 164408 318139 165829 318230
rect 25918 316944 25988 316954
rect 25918 316894 25928 316944
rect 25978 316894 25988 316944
rect 25918 316884 25988 316894
rect 25927 316743 25997 316753
rect 25927 316693 25937 316743
rect 25987 316693 25997 316743
rect 25927 316683 25997 316693
rect 25912 316054 25982 316064
rect 25912 316004 25922 316054
rect 25972 316004 25982 316054
rect 25912 315994 25982 316004
rect 25918 315703 25988 315713
rect 25918 315653 25928 315703
rect 25978 315653 25988 315703
rect 25918 315643 25988 315653
rect 164433 312230 165854 312313
rect 164433 311055 164506 312230
rect 165772 311055 165854 312230
rect 164433 310964 165854 311055
rect 164414 305144 165835 305227
rect 164414 303969 164487 305144
rect 165753 303969 165835 305144
rect 164414 303878 165835 303969
rect 164522 295871 165943 295954
rect 164522 294696 164595 295871
rect 165861 294696 165943 295871
rect 164522 294605 165943 294696
rect 164503 288785 165924 288868
rect 164503 287610 164576 288785
rect 165842 287610 165924 288785
rect 164503 287519 165924 287610
rect 164466 282383 165887 282466
rect 164466 281208 164539 282383
rect 165805 281208 165887 282383
rect 164466 281117 165887 281208
rect 164573 273463 165994 273546
rect 164573 272288 164646 273463
rect 165912 272288 165994 273463
rect 164573 272197 165994 272288
rect 164554 266377 165975 266460
rect 164554 265202 164627 266377
rect 165893 265202 165975 266377
rect 164554 265111 165975 265202
rect 266017 265300 266133 265309
rect 266017 265202 266024 265300
rect 266126 265202 266133 265300
rect 266017 265191 266133 265202
rect 26436 264775 26571 264785
rect 26436 264665 26446 264775
rect 26561 264665 26571 264775
rect 26436 264660 26571 264665
rect 23581 264447 23730 264462
rect 23581 264330 23597 264447
rect 23716 264330 23730 264447
rect 23581 264315 23730 264330
rect 265937 262942 266053 262951
rect 265937 262844 265944 262942
rect 266046 262844 266053 262942
rect 265937 262833 266053 262844
rect 265858 260457 265974 260466
rect 265858 260359 265865 260457
rect 265967 260359 265974 260457
rect 265858 260348 265974 260359
rect 164517 259975 165938 260058
rect 164517 258800 164590 259975
rect 165856 258800 165938 259975
rect 164517 258709 165938 258800
rect 164604 249209 166025 249292
rect 164604 248034 164677 249209
rect 165943 248034 166025 249209
rect 164604 247943 166025 248034
rect 164585 242123 166006 242206
rect 164585 240948 164658 242123
rect 165924 240948 166006 242123
rect 164585 240857 166006 240948
rect 242679 241013 242763 241022
rect 242679 240947 242684 241013
rect 242756 240947 242763 241013
rect 242679 240939 242763 240947
rect 63180 240219 63315 240230
rect 63180 240105 63189 240219
rect 63304 240105 63315 240219
rect 63180 240095 63315 240105
rect 63101 237883 63236 237894
rect 63101 237769 63110 237883
rect 63225 237769 63236 237883
rect 63101 237759 63236 237769
rect 164548 235721 165969 235804
rect 63020 235399 63155 235410
rect 63020 235285 63029 235399
rect 63144 235285 63155 235399
rect 63020 235275 63155 235285
rect 164548 234546 164621 235721
rect 165887 234546 165969 235721
rect 164548 234455 165969 234546
rect 63024 233192 63159 233203
rect 63024 233078 63033 233192
rect 63148 233078 63159 233192
rect 63024 233068 63159 233078
rect 164728 228943 166149 229026
rect 164728 227768 164801 228943
rect 166067 227768 166149 228943
rect 164728 227677 166149 227768
rect 164708 223081 166129 223164
rect 164708 221906 164781 223081
rect 166047 221906 166129 223081
rect 164708 221815 166129 221906
rect 164748 211018 166169 211101
rect 164748 209843 164821 211018
rect 166087 209843 166169 211018
rect 164748 209752 166169 209843
rect 164729 203932 166150 204015
rect 164729 202757 164802 203932
rect 166068 202757 166150 203932
rect 164729 202666 166150 202757
rect 164692 197530 166113 197613
rect 164692 196355 164765 197530
rect 166031 196355 166113 197530
rect 164692 196264 166113 196355
rect 164735 193125 166156 193208
rect 164735 191950 164808 193125
rect 166074 191950 166156 193125
rect 164735 191859 166156 191950
rect 61507 186500 61636 186511
rect 61507 186400 61518 186500
rect 61626 186400 61636 186500
rect 61507 186389 61636 186400
rect 164716 186039 166137 186122
rect 164716 184864 164789 186039
rect 166055 184864 166137 186039
rect 164716 184773 166137 184864
rect 61427 184077 61556 184088
rect 61427 183977 61438 184077
rect 61546 183977 61556 184077
rect 61427 183966 61556 183977
rect 61348 181593 61477 181604
rect 61348 181493 61359 181593
rect 61467 181493 61477 181593
rect 61348 181482 61477 181493
rect 164679 179637 166100 179720
rect 61349 179442 61478 179453
rect 61349 179342 61360 179442
rect 61468 179342 61478 179442
rect 61349 179331 61478 179342
rect 164679 178462 164752 179637
rect 166018 178462 166100 179637
rect 164679 178371 166100 178462
rect 164539 173712 165960 173795
rect 164539 172537 164612 173712
rect 165878 172537 165960 173712
rect 164539 172446 165960 172537
rect 164502 167310 165923 167393
rect 164502 166135 164575 167310
rect 165841 166135 165923 167310
rect 164502 166044 165923 166135
rect 164768 160049 166189 160132
rect 164768 158874 164841 160049
rect 166107 158874 166189 160049
rect 164768 158783 166189 158874
rect 164749 155209 166170 155292
rect 164749 154034 164822 155209
rect 166088 154034 166170 155209
rect 164749 153943 166170 154034
rect 164730 149939 166151 150022
rect 164730 148764 164803 149939
rect 166069 148764 166151 149939
rect 164730 148673 166151 148764
rect 164712 144387 166133 144470
rect 164712 143212 164785 144387
rect 166051 143212 166133 144387
rect 164712 143121 166133 143212
rect 269038 142783 269176 142796
rect 269038 142679 269050 142783
rect 269160 142679 269176 142783
rect 269038 142667 269176 142679
rect 268957 140387 269095 140400
rect 268957 140283 268969 140387
rect 269079 140283 269095 140387
rect 268957 140271 269095 140283
rect 164712 138197 166133 138280
rect 164712 137022 164785 138197
rect 166051 137022 166133 138197
rect 268878 137927 269016 137940
rect 268878 137823 268890 137927
rect 269000 137823 269016 137927
rect 268878 137811 269016 137823
rect 164712 136931 166133 137022
rect 164720 119093 166141 119176
rect 164720 117918 164793 119093
rect 166059 117918 166141 119093
rect 164720 117827 166141 117918
rect 164829 111166 166250 111249
rect 164829 109991 164902 111166
rect 166168 109991 166250 111166
rect 164829 109900 166250 109991
rect 164930 102964 166351 103047
rect 164930 101789 165003 102964
rect 166269 101789 166351 102964
rect 164930 101698 166351 101789
rect 164893 95465 166314 95548
rect 164893 94290 164966 95465
rect 166232 94290 166314 95465
rect 164893 94199 166314 94290
rect 164874 88379 166295 88462
rect 164874 87204 164947 88379
rect 166213 87204 166295 88379
rect 164874 87113 166295 87204
rect 164837 81977 166258 82060
rect 164837 80802 164910 81977
rect 166176 80802 166258 81977
rect 164837 80711 166258 80802
rect 164819 70727 166240 70810
rect 164819 69552 164892 70727
rect 166158 69552 166240 70727
rect 164819 69461 166240 69552
rect 164745 64732 166166 64815
rect 164745 63557 164818 64732
rect 166084 63557 166166 64732
rect 164745 63466 166166 63557
rect 164782 58904 166203 58987
rect 164782 57729 164855 58904
rect 166121 57729 166203 58904
rect 164782 57638 166203 57729
rect 164856 52817 166277 52900
rect 164856 51642 164929 52817
rect 166195 51642 166277 52817
rect 164856 51551 166277 51642
rect 164568 44959 165989 45042
rect 164568 43784 164641 44959
rect 165907 43784 165989 44959
rect 164568 43693 165989 43784
rect 164568 38665 165989 38748
rect 164568 37490 164641 38665
rect 165907 37490 165989 38665
rect 164568 37399 165989 37490
rect 164568 32371 165989 32454
rect 164568 31196 164641 32371
rect 165907 31196 165989 32371
rect 164568 31105 165989 31196
rect 164584 21815 166005 21898
rect 164584 20640 164657 21815
rect 165923 20640 166005 21815
rect 164584 20549 166005 20640
rect 164517 16137 166098 16247
rect 164517 14962 164641 16137
rect 165907 14962 166098 16137
rect 164517 14797 166098 14962
rect 164568 9044 165989 9127
rect 164568 7869 164641 9044
rect 165907 7869 165989 9044
rect 164568 7778 165989 7869
rect 262 -400 318 240
rect 853 -400 909 240
rect 1444 -400 1500 240
rect 2035 -400 2091 240
rect 2626 -400 2682 240
rect 3217 -400 3273 240
rect 3808 -400 3864 240
rect 4399 -400 4455 240
rect 4990 -400 5046 240
rect 5581 -400 5637 240
rect 6172 -400 6228 240
rect 6763 -400 6819 240
rect 7354 -400 7410 240
rect 7945 -400 8001 240
rect 8536 -400 8592 240
rect 9127 -400 9183 240
rect 9718 -400 9774 240
rect 10309 -400 10365 240
rect 10900 -400 10956 240
rect 11491 -400 11547 240
rect 12082 -400 12138 240
rect 12673 -400 12729 240
rect 13264 -400 13320 240
rect 13855 -400 13911 240
rect 14446 -400 14502 240
rect 15037 -400 15093 240
rect 15628 -400 15684 240
rect 16219 -400 16275 240
rect 16810 -400 16866 240
rect 17401 -400 17457 240
rect 17992 -400 18048 240
rect 18583 -400 18639 240
rect 19174 -400 19230 240
rect 19765 -400 19821 240
rect 20356 -400 20412 240
rect 20947 -400 21003 240
rect 21538 -400 21594 240
rect 22129 -400 22185 240
rect 22720 -400 22776 240
rect 23311 -400 23367 240
rect 23902 -400 23958 240
rect 24493 -400 24549 240
rect 25084 -400 25140 240
rect 25675 -400 25731 240
rect 26266 -400 26322 240
rect 26857 -400 26913 240
rect 27448 -400 27504 240
rect 28039 -400 28095 240
rect 28630 -400 28686 240
rect 29221 -400 29277 240
rect 29812 -400 29868 240
rect 30403 -400 30459 240
rect 30994 -400 31050 240
rect 31585 -400 31641 240
rect 32176 -400 32232 240
rect 32767 -400 32823 240
rect 33358 -400 33414 240
rect 33949 -400 34005 240
rect 34540 -400 34596 240
rect 35131 -400 35187 240
rect 35722 -400 35778 240
rect 36313 -400 36369 240
rect 36904 -400 36960 240
rect 37495 -400 37551 240
rect 38086 -400 38142 240
rect 38677 -400 38733 240
rect 39268 -400 39324 240
rect 39859 -400 39915 240
rect 40450 -400 40506 240
rect 41041 -400 41097 240
rect 41632 -400 41688 240
rect 42223 -400 42279 240
rect 42814 -400 42870 240
rect 43405 -400 43461 240
rect 43996 -400 44052 240
rect 44587 -400 44643 240
rect 45178 -400 45234 240
rect 45769 -400 45825 240
rect 46360 -400 46416 240
rect 46951 -400 47007 240
rect 47542 -400 47598 240
rect 48133 -400 48189 240
rect 48724 -400 48780 240
rect 49315 -400 49371 240
rect 49906 -400 49962 240
rect 50497 -400 50553 240
rect 51088 -400 51144 240
rect 51679 -400 51735 240
rect 52270 -400 52326 240
rect 52861 -400 52917 240
rect 53452 -400 53508 240
rect 54043 -400 54099 240
rect 54634 -400 54690 240
rect 55225 -400 55281 240
rect 55816 -400 55872 240
rect 56407 -400 56463 240
rect 56998 -400 57054 240
rect 57589 -400 57645 240
rect 58180 -400 58236 240
rect 58771 -400 58827 240
rect 59362 -400 59418 240
rect 59953 -400 60009 240
rect 60544 -400 60600 240
rect 61135 -400 61191 240
rect 61726 -400 61782 240
rect 62317 -400 62373 240
rect 62908 -400 62964 240
rect 63499 -400 63555 240
rect 64090 -400 64146 240
rect 64681 -400 64737 240
rect 65272 -400 65328 240
rect 65863 -400 65919 240
rect 66454 -400 66510 240
rect 67045 -400 67101 240
rect 67636 -400 67692 240
rect 68227 -400 68283 240
rect 68818 -400 68874 240
rect 69409 -400 69465 240
rect 70000 -400 70056 240
rect 70591 -400 70647 240
rect 71182 -400 71238 240
rect 71773 -400 71829 240
rect 72364 -400 72420 240
rect 72955 -400 73011 240
rect 73546 -400 73602 240
rect 74137 -400 74193 240
rect 74728 -400 74784 240
rect 75319 -400 75375 240
rect 75910 -400 75966 240
rect 76501 -400 76557 240
rect 77092 -400 77148 240
rect 77683 -400 77739 240
rect 78274 -400 78330 240
rect 78865 -400 78921 240
rect 79456 -400 79512 240
rect 80047 -400 80103 240
rect 80638 -400 80694 240
rect 81229 -400 81285 240
rect 81820 -400 81876 240
rect 82411 -400 82467 240
rect 83002 -400 83058 240
rect 83593 -400 83649 240
rect 84184 -400 84240 240
rect 84775 -400 84831 240
rect 85366 -400 85422 240
rect 85957 -400 86013 240
rect 86548 -400 86604 240
rect 87139 -400 87195 240
rect 87730 -400 87786 240
rect 88321 -400 88377 240
rect 88912 -400 88968 240
rect 89503 -400 89559 240
rect 90094 -400 90150 240
rect 90685 -400 90741 240
rect 91276 -400 91332 240
rect 91867 -400 91923 240
rect 92458 -400 92514 240
rect 93049 -400 93105 240
rect 93640 -400 93696 240
rect 94231 -400 94287 240
rect 94822 -400 94878 240
rect 95413 -400 95469 240
rect 96004 -400 96060 240
rect 96595 -400 96651 240
rect 97186 -400 97242 240
rect 97777 -400 97833 240
rect 98368 -400 98424 240
rect 98959 -400 99015 240
rect 99550 -400 99606 240
rect 100141 -400 100197 240
rect 100732 -400 100788 240
rect 101323 -400 101379 240
rect 101914 -400 101970 240
rect 102505 -400 102561 240
rect 103096 -400 103152 240
rect 103687 -400 103743 240
rect 104278 -400 104334 240
rect 104869 -400 104925 240
rect 105460 -400 105516 240
rect 106051 -400 106107 240
rect 106642 -400 106698 240
rect 107233 -400 107289 240
rect 107824 -400 107880 240
rect 108415 -400 108471 240
rect 109006 -400 109062 240
rect 109597 -400 109653 240
rect 110188 -400 110244 240
rect 110779 -400 110835 240
rect 111370 -400 111426 240
rect 111961 -400 112017 240
rect 112552 -400 112608 240
rect 113143 -400 113199 240
rect 113734 -400 113790 240
rect 114325 -400 114381 240
rect 114916 -400 114972 240
rect 115507 -400 115563 240
rect 116098 -400 116154 240
rect 116689 -400 116745 240
rect 117280 -400 117336 240
rect 117871 -400 117927 240
rect 118462 -400 118518 240
rect 119053 -400 119109 240
rect 119644 -400 119700 240
rect 120235 -400 120291 240
rect 120826 -400 120882 240
rect 121417 -400 121473 240
rect 122008 -400 122064 240
rect 122599 -400 122655 240
rect 123190 -400 123246 240
rect 123781 -400 123837 240
rect 124372 -400 124428 240
rect 124963 -400 125019 240
rect 125554 -400 125610 240
rect 126145 -400 126201 240
rect 126736 -400 126792 240
rect 127327 -400 127383 240
rect 127918 -400 127974 240
rect 128509 -400 128565 240
rect 129100 -400 129156 240
rect 129691 -400 129747 240
rect 130282 -400 130338 240
rect 130873 -400 130929 240
rect 131464 -400 131520 240
rect 132055 -400 132111 240
rect 132646 -400 132702 240
rect 133237 -400 133293 240
rect 133828 -400 133884 240
rect 134419 -400 134475 240
rect 135010 -400 135066 240
rect 135601 -400 135657 240
rect 136192 -400 136248 240
rect 136783 -400 136839 240
rect 137374 -400 137430 240
rect 137965 -400 138021 240
rect 138556 -400 138612 240
rect 139147 -400 139203 240
rect 139738 -400 139794 240
rect 140329 -400 140385 240
rect 140920 -400 140976 240
rect 141511 -400 141567 240
rect 142102 -400 142158 240
rect 142693 -400 142749 240
rect 143284 -400 143340 240
rect 143875 -400 143931 240
rect 144466 -400 144522 240
rect 145057 -400 145113 240
rect 145648 -400 145704 240
rect 146239 -400 146295 240
rect 146830 -400 146886 240
rect 147421 -400 147477 240
rect 148012 -400 148068 240
rect 148603 -400 148659 240
rect 149194 -400 149250 240
rect 149785 -400 149841 240
rect 150376 -400 150432 240
rect 150967 -400 151023 240
rect 151558 -400 151614 240
rect 152149 -400 152205 240
rect 152740 -400 152796 240
rect 153331 -400 153387 240
rect 153922 -400 153978 240
rect 154513 -400 154569 240
rect 155104 -400 155160 240
rect 155695 -400 155751 240
rect 156286 -400 156342 240
rect 156877 -400 156933 240
rect 157468 -400 157524 240
rect 158059 -400 158115 240
rect 158650 -400 158706 240
rect 159241 -400 159297 240
rect 159832 -400 159888 240
rect 160423 -400 160479 240
rect 161014 -400 161070 240
rect 161605 -400 161661 240
rect 162196 -400 162252 240
rect 162787 -400 162843 240
rect 163378 -400 163434 240
rect 163969 -400 164025 240
rect 164560 -400 164616 240
rect 165151 -400 165207 240
rect 165742 -400 165798 240
rect 166333 -400 166389 240
rect 166924 -400 166980 240
rect 167515 -400 167571 240
rect 168106 -400 168162 240
rect 168697 -400 168753 240
rect 169288 -400 169344 240
rect 169879 -400 169935 240
rect 170470 -400 170526 240
rect 171061 -400 171117 240
rect 171652 -400 171708 240
rect 172243 -400 172299 240
rect 172834 -400 172890 240
rect 173425 -400 173481 240
rect 174016 -400 174072 240
rect 174607 -400 174663 240
rect 175198 -400 175254 240
rect 175789 -400 175845 240
rect 176380 -400 176436 240
rect 176971 -400 177027 240
rect 177562 -400 177618 240
rect 178153 -400 178209 240
rect 178744 -400 178800 240
rect 179335 -400 179391 240
rect 179926 -400 179982 240
rect 180517 -400 180573 240
rect 181108 -400 181164 240
rect 181699 -400 181755 240
rect 182290 -400 182346 240
rect 182881 -400 182937 240
rect 183472 -400 183528 240
rect 184063 -400 184119 240
rect 184654 -400 184710 240
rect 185245 -400 185301 240
rect 185836 -400 185892 240
rect 186427 -400 186483 240
rect 187018 -400 187074 240
rect 187609 -400 187665 240
rect 188200 -400 188256 240
rect 188791 -400 188847 240
rect 189382 -400 189438 240
rect 189973 -400 190029 240
rect 190564 -400 190620 240
rect 191155 -400 191211 240
rect 191746 -400 191802 240
rect 192337 -400 192393 240
rect 192928 -400 192984 240
rect 193519 -400 193575 240
rect 194110 -400 194166 240
rect 194701 -400 194757 240
rect 195292 -400 195348 240
rect 195883 -400 195939 240
rect 196474 -400 196530 240
rect 197065 -400 197121 240
rect 197656 -400 197712 240
rect 198247 -400 198303 240
rect 198838 -400 198894 240
rect 199429 -400 199485 240
rect 200020 -400 200076 240
rect 200611 -400 200667 240
rect 201202 -400 201258 240
rect 201793 -400 201849 240
rect 202384 -400 202440 240
rect 202975 -400 203031 240
rect 203566 -400 203622 240
rect 204157 -400 204213 240
rect 204748 -400 204804 240
rect 205339 -400 205395 240
rect 205930 -400 205986 240
rect 206521 -400 206577 240
rect 207112 -400 207168 240
rect 207703 -400 207759 240
rect 208294 -400 208350 240
rect 208885 -400 208941 240
rect 209476 -400 209532 240
rect 210067 -400 210123 240
rect 210658 -400 210714 240
rect 211249 -400 211305 240
rect 211840 -400 211896 240
rect 212431 -400 212487 240
rect 213022 -400 213078 240
rect 213613 -400 213669 240
rect 214204 -400 214260 240
rect 214795 -400 214851 240
rect 215386 -400 215442 240
rect 215977 -400 216033 240
rect 216568 -400 216624 240
rect 217159 -400 217215 240
rect 217750 -400 217806 240
rect 218341 -400 218397 240
rect 218932 -400 218988 240
rect 219523 -400 219579 240
rect 220114 -400 220170 240
rect 220705 -400 220761 240
rect 221296 -400 221352 240
rect 221887 -400 221943 240
rect 222478 -400 222534 240
rect 223069 -400 223125 240
rect 223660 -400 223716 240
rect 224251 -400 224307 240
rect 224842 -400 224898 240
rect 225433 -400 225489 240
rect 226024 -400 226080 240
rect 226615 -400 226671 240
rect 227206 -400 227262 240
rect 227797 -400 227853 240
rect 228388 -400 228444 240
rect 228979 -400 229035 240
rect 229570 -400 229626 240
rect 230161 -400 230217 240
rect 230752 -400 230808 240
rect 231343 -400 231399 240
rect 231934 -400 231990 240
rect 232525 -400 232581 240
rect 233116 -400 233172 240
rect 233707 -400 233763 240
rect 234298 -400 234354 240
rect 234889 -400 234945 240
rect 235480 -400 235536 240
rect 236071 -400 236127 240
rect 236662 -400 236718 240
rect 237253 -400 237309 240
rect 237844 -400 237900 240
rect 238435 -400 238491 240
rect 239026 -400 239082 240
rect 239617 -400 239673 240
rect 240208 -400 240264 240
rect 240799 -400 240855 240
rect 241390 -400 241446 240
rect 241981 -400 242037 240
rect 242572 -400 242628 240
rect 243163 -400 243219 240
rect 243754 -400 243810 240
rect 244345 -400 244401 240
rect 244936 -400 244992 240
rect 245527 -400 245583 240
rect 246118 -400 246174 240
rect 246709 -400 246765 240
rect 247300 -400 247356 240
rect 247891 -400 247947 240
rect 248482 -400 248538 240
rect 249073 -400 249129 240
rect 249664 -400 249720 240
rect 250255 -400 250311 240
rect 250846 -400 250902 240
rect 251437 -400 251493 240
rect 252028 -400 252084 240
rect 252619 -400 252675 240
rect 253210 -400 253266 240
rect 253801 -400 253857 240
rect 254392 -400 254448 240
rect 254983 -400 255039 240
rect 255574 -400 255630 240
rect 256165 -400 256221 240
rect 256756 -400 256812 240
rect 257347 -400 257403 240
rect 257938 -400 257994 240
rect 258529 -400 258585 240
rect 259120 -400 259176 240
rect 259711 -400 259767 240
rect 260302 -400 260358 240
rect 260893 -400 260949 240
rect 261484 -400 261540 240
rect 262075 -400 262131 240
rect 262666 -400 262722 240
rect 263257 -400 263313 240
rect 263848 -400 263904 240
rect 264439 -400 264495 240
rect 265030 -400 265086 240
rect 265621 -400 265677 240
rect 266212 -400 266268 240
rect 266803 -400 266859 240
rect 267394 -400 267450 240
rect 267985 -400 268041 240
rect 268576 -400 268632 240
rect 269167 -400 269223 240
rect 269758 -400 269814 240
rect 270349 -400 270405 240
rect 270940 -400 270996 240
rect 271531 -400 271587 240
rect 272122 -400 272178 240
rect 272713 -400 272769 240
rect 273304 -400 273360 240
rect 273895 -400 273951 240
rect 274486 -400 274542 240
rect 275077 -400 275133 240
rect 275668 -400 275724 240
rect 276259 -400 276315 240
rect 276850 -400 276906 240
rect 277441 -400 277497 240
rect 278032 -400 278088 240
rect 278623 -400 278679 240
rect 279214 -400 279270 240
rect 279805 -400 279861 240
rect 280396 -400 280452 240
rect 280987 -400 281043 240
rect 281578 -400 281634 240
rect 282169 -400 282225 240
rect 282760 -400 282816 240
rect 283351 -400 283407 240
rect 283942 -400 283998 240
rect 284533 -400 284589 240
rect 285124 -400 285180 240
rect 285715 -400 285771 240
rect 286306 -400 286362 240
rect 286897 -400 286953 240
rect 287488 -400 287544 240
rect 288079 -400 288135 240
rect 288670 -400 288726 240
rect 289261 -400 289317 240
rect 289852 -400 289908 240
rect 290443 -400 290499 240
rect 291034 -400 291090 240
rect 291625 -400 291681 240
<< via2 >>
rect 164500 338774 165766 339949
rect 164481 331688 165747 332863
rect 247701 329822 247772 329890
rect 247459 329454 247560 329554
rect 164500 325316 165766 326491
rect 164481 318230 165747 319405
rect 25928 316894 25978 316944
rect 25937 316693 25987 316743
rect 25922 316004 25972 316054
rect 25928 315653 25978 315703
rect 164506 311055 165772 312230
rect 164487 303969 165753 305144
rect 164595 294696 165861 295871
rect 164576 287610 165842 288785
rect 164539 281208 165805 282383
rect 164646 272288 165912 273463
rect 164627 265202 165893 266377
rect 266024 265202 266126 265300
rect 26446 264665 26561 264775
rect 265944 262844 266046 262942
rect 265865 260359 265967 260457
rect 164590 258800 165856 259975
rect 164677 248034 165943 249209
rect 164658 240948 165924 242123
rect 242684 240947 242756 241013
rect 63189 240105 63304 240219
rect 63110 237769 63225 237883
rect 63029 235285 63144 235399
rect 164621 234546 165887 235721
rect 63033 233078 63148 233192
rect 164801 227768 166067 228943
rect 164781 221906 166047 223081
rect 164821 209843 166087 211018
rect 164802 202757 166068 203932
rect 164765 196355 166031 197530
rect 164808 191950 166074 193125
rect 61518 186400 61626 186500
rect 164789 184864 166055 186039
rect 61438 183977 61546 184077
rect 61359 181493 61467 181593
rect 61360 179342 61468 179442
rect 164752 178462 166018 179637
rect 164612 172537 165878 173712
rect 164575 166135 165841 167310
rect 164841 158874 166107 160049
rect 164822 154034 166088 155209
rect 164803 148764 166069 149939
rect 164785 143212 166051 144387
rect 269050 142679 269160 142783
rect 268969 140283 269079 140387
rect 164785 137022 166051 138197
rect 268890 137823 269000 137927
rect 164793 117918 166059 119093
rect 164902 109991 166168 111166
rect 165003 101789 166269 102964
rect 164966 94290 166232 95465
rect 164947 87204 166213 88379
rect 164910 80802 166176 81977
rect 164892 69552 166158 70727
rect 164818 63557 166084 64732
rect 164855 57729 166121 58904
rect 164929 51642 166195 52817
rect 164641 43784 165907 44959
rect 164641 37490 165907 38665
rect 164641 31196 165907 32371
rect 164657 20640 165923 21815
rect 164641 14962 165907 16137
rect 164641 7869 165907 9044
<< metal3 >>
rect 8097 351150 10597 352400
rect 34097 351150 36597 352400
rect 60097 351150 62597 352400
rect 82797 351150 85297 352400
rect 85447 351150 86547 352400
rect 86697 351150 87797 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 111297 351150 112397 352400
rect 112547 351150 113647 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 162147 351150 163247 352400
rect 163397 351150 164497 352400
rect 164647 351150 167147 352400
rect 206697 351150 209197 352400
rect 232697 351150 235197 352400
rect 255297 351170 257697 352400
rect 260297 351170 262697 352400
rect 8376 349233 10412 351150
rect 34331 349233 36367 351150
rect 60339 349338 62375 351150
rect 82963 349244 84999 351150
rect 88168 349208 90204 351150
rect 108814 349155 110850 351150
rect 114054 349155 116090 351150
rect 159668 349191 161704 351150
rect 164874 349155 166910 351150
rect 206890 349311 208926 351150
rect 232866 349389 234902 351150
rect 255440 349320 257476 351170
rect 260451 349303 262487 351170
rect 283297 351150 285797 352400
rect 283588 349206 285624 351150
rect -400 342364 850 342621
rect -400 340471 4906 342364
rect 291150 341209 292400 341492
rect -400 340121 850 340471
rect 164427 339949 165848 340032
rect 164427 338774 164500 339949
rect 165766 338774 165848 339949
rect 287117 339172 292400 341209
rect 291150 338992 292400 339172
rect 164427 338683 165848 338774
rect 164408 332863 165829 332946
rect 164408 331688 164481 332863
rect 165747 331688 165829 332863
rect 164408 331597 165829 331688
rect 247049 330028 247236 330039
rect 247049 330027 247778 330028
rect 247049 330024 247782 330027
rect 247049 329881 247062 330024
rect 247219 329940 247782 330024
rect 247219 329881 247236 329940
rect 247049 329859 247236 329881
rect 247681 329890 247782 329940
rect 247681 329822 247701 329890
rect 247772 329822 247782 329890
rect 247681 329815 247782 329822
rect 247445 329554 247576 329570
rect 247445 329454 247459 329554
rect 247560 329454 247576 329554
rect 247445 329439 247576 329454
rect 164427 326491 165848 326574
rect 164427 325316 164500 326491
rect 165766 325316 165848 326491
rect 164427 325225 165848 325316
rect -400 324049 830 324321
rect -400 322156 4976 324049
rect -400 321921 830 322156
rect 291170 322092 292400 322292
rect 287015 320055 292400 322092
rect 291170 319892 292400 320055
rect 164408 319405 165829 319488
rect -400 319125 830 319321
rect -400 317232 4906 319125
rect 164408 318230 164481 319405
rect 165747 318230 165829 319405
rect 164408 318139 165829 318230
rect -400 316921 830 317232
rect 291170 317127 292400 317292
rect 25918 316944 25997 316959
rect 25918 316943 25928 316944
rect 25918 316893 25927 316943
rect 25978 316893 25997 316944
rect 25918 316882 25997 316893
rect 25927 316743 26006 316758
rect 25927 316742 25937 316743
rect 25927 316692 25936 316742
rect 25987 316692 26006 316743
rect 25927 316681 26006 316692
rect 25912 316054 25991 316069
rect 25912 316053 25922 316054
rect 25912 316003 25921 316053
rect 25972 316003 25991 316054
rect 25912 315992 25991 316003
rect 25918 315703 25997 315718
rect 25918 315702 25928 315703
rect 25918 315652 25927 315702
rect 25978 315652 25997 315703
rect 25918 315641 25997 315652
rect 287114 315090 292400 317127
rect 291170 314892 292400 315090
rect 164433 312230 165854 312313
rect 164433 311055 164506 312230
rect 165772 311055 165854 312230
rect 164433 310964 165854 311055
rect 164414 305144 165835 305227
rect 164414 303969 164487 305144
rect 165753 303969 165835 305144
rect 164414 303878 165835 303969
rect 164522 295871 165943 295954
rect 164522 294696 164595 295871
rect 165861 294696 165943 295871
rect 291760 294736 292400 294792
rect 164522 294605 165943 294696
rect 291760 294145 292400 294201
rect 291760 293554 292400 293610
rect 291760 292963 292400 293019
rect 287531 292428 291858 292545
rect 287531 292372 292400 292428
rect 287531 292267 291858 292372
rect 287523 291837 291850 291977
rect 287523 291781 292400 291837
rect 287523 291699 291850 291781
rect 164503 288785 165924 288868
rect 164503 287610 164576 288785
rect 165842 287610 165924 288785
rect 164503 287519 165924 287610
rect 164466 282383 165887 282466
rect -400 281893 830 282121
rect -400 280000 4941 281893
rect 164466 281208 164539 282383
rect 165805 281208 165887 282383
rect 164466 281117 165887 281208
rect -400 279721 830 280000
rect 273285 277424 287287 277475
rect 291170 277424 292400 277681
rect -400 276863 830 277121
rect 273285 276989 292400 277424
rect -400 274970 4906 276863
rect 273285 275847 273813 276989
rect 275123 275847 292400 276989
rect 273285 275531 292400 275847
rect 273285 275503 287287 275531
rect 291170 275281 292400 275531
rect -400 274721 830 274970
rect 164573 273463 165994 273546
rect 164573 272288 164646 273463
rect 165912 272288 165994 273463
rect 291170 272430 292400 272681
rect 164573 272197 165994 272288
rect 286997 270537 292400 272430
rect 291170 270281 292400 270537
rect 164554 266377 165975 266460
rect 164554 265202 164627 266377
rect 165893 265202 165975 266377
rect 164554 265111 165975 265202
rect 266017 265300 266133 265309
rect 266017 265202 266024 265300
rect 266126 265202 266133 265300
rect 266017 265191 266133 265202
rect 26436 264775 26571 264785
rect 26436 264665 26446 264775
rect 26561 264665 26571 264775
rect 26436 264660 26571 264665
rect 265937 262942 266053 262951
rect 265937 262844 265944 262942
rect 266046 262844 266053 262942
rect 265937 262833 266053 262844
rect 265858 260457 265974 260466
rect 265858 260359 265865 260457
rect 265967 260359 265974 260457
rect 265858 260348 265974 260359
rect 164517 259975 165938 260058
rect 164517 258800 164590 259975
rect 165856 258800 165938 259975
rect 164517 258709 165938 258800
rect 176 255821 1564 255918
rect -400 255765 1564 255821
rect 176 255663 1564 255765
rect 190 255230 1578 255336
rect -400 255174 1578 255230
rect 190 255081 1578 255174
rect -400 254583 240 254639
rect -400 253992 240 254048
rect -400 253401 240 253457
rect -400 252810 240 252866
rect 291760 250025 292400 250081
rect 291760 249434 292400 249490
rect 164604 249209 166025 249292
rect 164604 248034 164677 249209
rect 165943 248034 166025 249209
rect 291760 248843 292400 248899
rect 291760 248252 292400 248308
rect 164604 247943 166025 248034
rect 291760 247661 292400 247717
rect 291760 247070 292400 247126
rect 164585 242123 166006 242206
rect 164585 240948 164658 242123
rect 165924 240948 166006 242123
rect 164585 240857 166006 240948
rect 242679 241013 242763 241022
rect 242679 240947 242684 241013
rect 242756 240947 242763 241013
rect 242679 240939 242763 240947
rect 63180 240219 63315 240230
rect 63180 240105 63189 240219
rect 63304 240105 63315 240219
rect 63180 240095 63315 240105
rect 63101 237883 63236 237894
rect 63101 237769 63110 237883
rect 63225 237769 63236 237883
rect 63101 237759 63236 237769
rect 164548 235721 165969 235804
rect 63020 235399 63155 235410
rect 63020 235285 63029 235399
rect 63144 235285 63155 235399
rect 63020 235275 63155 235285
rect 164548 234546 164621 235721
rect 165887 234546 165969 235721
rect 164548 234455 165969 234546
rect 153 234210 1541 234292
rect -400 234154 1541 234210
rect 153 234037 1541 234154
rect 176 233619 1564 233734
rect -400 233563 1564 233619
rect 176 233479 1564 233563
rect 63024 233192 63159 233203
rect 63024 233078 63033 233192
rect 63148 233078 63159 233192
rect 63024 233068 63159 233078
rect -400 232972 240 233028
rect -400 232381 240 232437
rect -400 231790 240 231846
rect -400 231199 240 231255
rect 164728 228943 166149 229026
rect 164728 227768 164801 228943
rect 166067 227768 166149 228943
rect 291760 227814 292400 227870
rect 164728 227677 166149 227768
rect 291760 227223 292400 227279
rect 291760 226632 292400 226688
rect 291760 226041 292400 226097
rect 291760 225450 292400 225506
rect 291760 224859 292400 224915
rect 164708 223081 166129 223164
rect 164708 221906 164781 223081
rect 166047 221906 166129 223081
rect 164708 221815 166129 221906
rect 171 212599 1559 212727
rect -400 212543 1559 212599
rect 171 212472 1559 212543
rect 175 212008 1563 212112
rect -400 211952 1563 212008
rect 175 211857 1563 211952
rect -400 211361 240 211417
rect 164748 211018 166169 211101
rect -400 210770 240 210826
rect -400 210179 240 210235
rect 164748 209843 164821 211018
rect 166087 209843 166169 211018
rect 164748 209752 166169 209843
rect -400 209588 240 209644
rect 291760 205603 292400 205659
rect 291760 205012 292400 205068
rect 291760 204421 292400 204477
rect 164729 203932 166150 204015
rect 164729 202757 164802 203932
rect 166068 202757 166150 203932
rect 291760 203830 292400 203886
rect 291760 203239 292400 203295
rect 164729 202666 166150 202757
rect 291760 202648 292400 202704
rect 164692 197530 166113 197613
rect 164692 196355 164765 197530
rect 166031 196355 166113 197530
rect 164692 196264 166113 196355
rect 164735 193125 166156 193208
rect 164735 191950 164808 193125
rect 166074 191950 166156 193125
rect 164735 191859 166156 191950
rect 185 190988 1573 191097
rect -400 190932 1573 190988
rect 185 190842 1573 190932
rect 204 190397 1592 190525
rect -400 190341 1592 190397
rect 204 190270 1592 190341
rect -400 189750 240 189806
rect -400 189159 240 189215
rect -400 188568 240 188624
rect -400 187977 240 188033
rect 61507 186500 61636 186511
rect 61507 186400 61518 186500
rect 61626 186400 61636 186500
rect 61507 186389 61636 186400
rect 164716 186039 166137 186122
rect 164716 184864 164789 186039
rect 166055 184864 166137 186039
rect 164716 184773 166137 184864
rect 61427 184077 61556 184088
rect 61427 183977 61438 184077
rect 61546 183977 61556 184077
rect 61427 183966 61556 183977
rect 291760 182392 292400 182448
rect 291760 181801 292400 181857
rect 61348 181593 61477 181604
rect 61348 181493 61359 181593
rect 61467 181493 61477 181593
rect 61348 181482 61477 181493
rect 291760 181210 292400 181266
rect 291760 180619 292400 180675
rect 291760 180028 292400 180084
rect 164679 179637 166100 179720
rect 61349 179442 61478 179453
rect 61349 179342 61360 179442
rect 61468 179342 61478 179442
rect 61349 179331 61478 179342
rect 164679 178462 164752 179637
rect 166018 178462 166100 179637
rect 291760 179437 292400 179493
rect 164679 178371 166100 178462
rect 164539 173712 165960 173795
rect 164539 172537 164612 173712
rect 165878 172537 165960 173712
rect 164539 172446 165960 172537
rect 181 169377 1569 169509
rect -400 169321 1569 169377
rect 181 169254 1569 169321
rect 199 168786 1587 168886
rect -400 168730 1587 168786
rect 199 168631 1587 168730
rect -400 168139 240 168195
rect -400 167548 240 167604
rect 164502 167310 165923 167393
rect -400 166957 240 167013
rect -400 166366 240 166422
rect 164502 166135 164575 167310
rect 165841 166135 165923 167310
rect 164502 166044 165923 166135
rect 164768 160049 166189 160132
rect 164768 158874 164841 160049
rect 166107 158874 166189 160049
rect 291760 159781 292400 159837
rect 291760 159190 292400 159246
rect 164768 158783 166189 158874
rect 291760 158599 292400 158655
rect 291760 158008 292400 158064
rect 291760 157417 292400 157473
rect 291760 156826 292400 156882
rect 164749 155209 166170 155292
rect 164749 154034 164822 155209
rect 166088 154034 166170 155209
rect 164749 153943 166170 154034
rect 164730 149939 166151 150022
rect 164730 148764 164803 149939
rect 166069 148764 166151 149939
rect 164730 148673 166151 148764
rect 190 147766 1578 147897
rect -400 147710 1578 147766
rect 190 147642 1578 147710
rect 218 147175 1606 147320
rect -400 147119 1606 147175
rect 218 147065 1606 147119
rect -400 146528 240 146584
rect -400 145937 240 145993
rect -400 145346 240 145402
rect -400 144755 240 144811
rect 164712 144387 166133 144470
rect 164712 143212 164785 144387
rect 166051 143212 166133 144387
rect 164712 143121 166133 143212
rect 269038 142783 269176 142796
rect 269038 142679 269050 142783
rect 269160 142679 269176 142783
rect 269038 142667 269176 142679
rect 268957 140387 269095 140400
rect 268957 140283 268969 140387
rect 269079 140283 269095 140387
rect 268957 140271 269095 140283
rect 164712 138197 166133 138280
rect 164712 137022 164785 138197
rect 166051 137022 166133 138197
rect 268878 137927 269016 137940
rect 268878 137823 268890 137927
rect 269000 137823 269016 137927
rect 268878 137811 269016 137823
rect 291760 137570 292400 137626
rect 164712 136931 166133 137022
rect 291760 136979 292400 137035
rect 291760 136388 292400 136444
rect 291760 135797 292400 135853
rect 291760 135206 292400 135262
rect 291760 134615 292400 134671
rect 195 126255 1583 126392
rect -400 126199 1583 126255
rect 195 126137 1583 126199
rect 204 125664 1592 125824
rect -400 125608 1592 125664
rect 204 125569 1592 125608
rect -400 125017 240 125073
rect -400 124426 240 124482
rect -400 123835 240 123891
rect -400 123244 240 123300
rect 164720 119093 166141 119176
rect 164720 117918 164793 119093
rect 166059 117918 166141 119093
rect 164720 117827 166141 117918
rect 291170 117615 292400 120015
rect 291170 112615 292400 115015
rect 164829 111166 166250 111249
rect 164829 109991 164902 111166
rect 166168 109991 166250 111166
rect 164829 109900 166250 109991
rect -400 109532 830 109844
rect -400 107639 4916 109532
rect -400 107444 830 107639
rect -400 104575 830 104844
rect -400 102682 4916 104575
rect 164930 102964 166351 103047
rect -400 102444 830 102682
rect 164930 101789 165003 102964
rect 166269 101789 166351 102964
rect 164930 101698 166351 101789
rect 291170 95715 292400 98115
rect 164893 95465 166314 95548
rect 164893 94290 164966 95465
rect 166232 94290 166314 95465
rect 164893 94199 166314 94290
rect 291170 90715 292400 93115
rect -400 88533 830 88844
rect -400 86640 4920 88533
rect 164874 88379 166295 88462
rect 164874 87204 164947 88379
rect 166213 87204 166295 88379
rect 164874 87113 166295 87204
rect -400 86444 830 86640
rect -400 83589 830 83844
rect -400 81696 4990 83589
rect 164837 81977 166258 82060
rect -400 81444 830 81696
rect 164837 80802 164910 81977
rect 166176 80802 166258 81977
rect 164837 80711 166258 80802
rect 280813 75549 287932 75721
rect 291170 75549 292400 75815
rect 280813 75451 292400 75549
rect 280813 73748 281123 75451
rect 282980 73748 292400 75451
rect 280813 73656 292400 73748
rect 280813 73516 287932 73656
rect 291170 73415 292400 73656
rect 164819 70727 166240 70810
rect 164819 69552 164892 70727
rect 166158 69552 166240 70727
rect 291170 70535 292400 70815
rect 164819 69461 166240 69552
rect 287095 68642 292400 70535
rect 291170 68415 292400 68642
rect 164745 64732 166166 64815
rect 164745 63557 164818 64732
rect 166084 63557 166166 64732
rect 164745 63466 166166 63557
rect 181 62444 1569 62587
rect -400 62388 1569 62444
rect 181 62332 1569 62388
rect 199 61853 1587 62001
rect -400 61797 1587 61853
rect 199 61746 1587 61797
rect -400 61206 240 61262
rect -400 60615 240 60671
rect -400 60024 240 60080
rect -400 59433 240 59489
rect 164782 58904 166203 58987
rect 164782 57729 164855 58904
rect 166121 57729 166203 58904
rect 164782 57638 166203 57729
rect 164856 52817 166277 52900
rect 164856 51642 164929 52817
rect 166195 51642 166277 52817
rect 164856 51551 166277 51642
rect 291760 47559 292400 47615
rect 291760 46968 292400 47024
rect 291760 46377 292400 46433
rect 291760 45786 292400 45842
rect 164568 44959 165989 45042
rect 164568 43784 164641 44959
rect 165907 43784 165989 44959
rect 164568 43693 165989 43784
rect 195 40833 1583 41003
rect -400 40777 1583 40833
rect 195 40748 1583 40777
rect 204 40242 1592 40399
rect -400 40186 1592 40242
rect 204 40144 1592 40186
rect -400 39595 240 39651
rect -400 39004 240 39060
rect 164568 38665 165989 38748
rect -400 38413 240 38469
rect -400 37822 240 37878
rect 164568 37490 164641 38665
rect 165907 37490 165989 38665
rect 164568 37399 165989 37490
rect 164568 32371 165989 32454
rect 164568 31196 164641 32371
rect 165907 31196 165989 32371
rect 164568 31105 165989 31196
rect 39779 30775 40392 30778
rect 39734 30146 40392 30775
rect 39734 30143 40347 30146
rect 39831 30099 40271 30143
rect 39831 29869 39950 30099
rect 40206 29869 40271 30099
rect 39831 29839 40271 29869
rect 291760 25230 292400 25286
rect 291760 24639 292400 24695
rect 291760 24048 292400 24104
rect 291760 23457 292400 23513
rect 164584 21815 166005 21898
rect 164584 20640 164657 21815
rect 165923 20640 166005 21815
rect 164584 20549 166005 20640
rect 199 19222 1587 19359
rect -400 19166 1587 19222
rect 199 19104 1587 19166
rect 195 18631 1583 18746
rect -400 18575 1583 18631
rect 195 18491 1583 18575
rect -400 17984 240 18040
rect -400 17393 240 17449
rect -400 16802 240 16858
rect -400 16211 240 16267
rect 164517 16137 166098 16247
rect 164517 14962 164641 16137
rect 165907 14962 166098 16137
rect 164517 14797 166098 14962
rect 291760 12001 292400 12057
rect 291760 11410 292400 11466
rect 291760 10819 292400 10875
rect 291760 10228 292400 10284
rect 291760 9637 292400 9693
rect 164568 9044 165989 9127
rect 291760 9046 292400 9102
rect 195 8511 1583 8651
rect -400 8455 1583 8511
rect 195 8396 1583 8455
rect 213 7920 1601 8041
rect -400 7864 1601 7920
rect 213 7786 1601 7864
rect 164568 7869 164641 9044
rect 165907 7869 165989 9044
rect 291760 8455 292400 8511
rect 164568 7778 165989 7869
rect 291760 7864 292400 7920
rect -400 7273 240 7329
rect 291760 7273 292400 7329
rect -400 6682 240 6738
rect 291760 6682 292400 6738
rect -400 6091 240 6147
rect 291760 6091 292400 6147
rect -400 5500 240 5556
rect 291760 5500 292400 5556
rect -400 4909 240 4965
rect 291760 4909 292400 4965
rect -400 4318 240 4374
rect 291760 4318 292400 4374
rect -400 3727 240 3783
rect 291760 3727 292400 3783
rect -400 3136 240 3192
rect 291760 3136 292400 3192
rect -400 2545 240 2601
rect 291760 2545 292400 2601
rect -400 1954 240 2010
rect 291760 1954 292400 2010
rect -400 1363 240 1419
rect 291760 1363 292400 1419
rect -400 772 240 828
rect 291760 772 292400 828
<< via3 >>
rect 164500 338774 165766 339949
rect 243932 337228 243984 337283
rect 243852 334765 243904 334815
rect 164481 331688 165747 332863
rect 247062 329881 247219 330024
rect 247459 329454 247560 329554
rect 164500 325316 165766 326491
rect 164481 318230 165747 319405
rect 245761 318620 245811 318670
rect 25927 316894 25928 316943
rect 25928 316894 25978 316943
rect 25927 316893 25978 316894
rect 25936 316693 25937 316742
rect 25937 316693 25987 316742
rect 25936 316692 25987 316693
rect 25921 316292 25972 316342
rect 245682 316154 245732 316204
rect 25921 316004 25922 316053
rect 25922 316004 25972 316053
rect 25921 316003 25972 316004
rect 25927 315653 25928 315702
rect 25928 315653 25978 315702
rect 25927 315652 25978 315653
rect 245602 313769 245652 313819
rect 164506 311055 165772 312230
rect 245523 311303 245573 311353
rect 245443 308917 245493 308967
rect 245363 306451 245413 306501
rect 164487 303969 165753 305144
rect 164595 294696 165861 295871
rect 164576 287610 165842 288785
rect 164539 281208 165805 282383
rect 273813 275847 275123 276989
rect 164646 272288 165912 273463
rect 164627 265202 165893 266377
rect 266024 265202 266126 265300
rect 26446 264665 26561 264775
rect 265944 262844 266046 262942
rect 265865 260359 265967 260457
rect 164590 258800 165856 259975
rect 164677 248034 165943 249209
rect 164658 240948 165924 242123
rect 242684 240947 242756 241013
rect 63189 240105 63304 240219
rect 63110 237769 63225 237883
rect 63029 235285 63144 235399
rect 164621 234546 165887 235721
rect 63033 233078 63148 233192
rect 164801 227768 166067 228943
rect 164781 221906 166047 223081
rect 164821 209843 166087 211018
rect 164802 202757 166068 203932
rect 164765 196355 166031 197530
rect 164808 191950 166074 193125
rect 61518 186400 61626 186500
rect 164789 184864 166055 186039
rect 61438 183977 61546 184077
rect 61359 181493 61467 181593
rect 61360 179342 61468 179442
rect 164752 178462 166018 179637
rect 164612 172537 165878 173712
rect 164575 166135 165841 167310
rect 164841 158874 166107 160049
rect 164822 154034 166088 155209
rect 164803 148764 166069 149939
rect 164785 143212 166051 144387
rect 269050 142679 269160 142783
rect 268969 140283 269079 140387
rect 164785 137022 166051 138197
rect 268890 137823 269000 137927
rect 164793 117918 166059 119093
rect 164902 109991 166168 111166
rect 165003 101789 166269 102964
rect 164966 94290 166232 95465
rect 164947 87204 166213 88379
rect 164910 80802 166176 81977
rect 281123 73748 282980 75451
rect 164892 69552 166158 70727
rect 164818 63557 166084 64732
rect 164855 57729 166121 58904
rect 164929 51642 166195 52817
rect 164641 43784 165907 44959
rect 164641 37490 165907 38665
rect 164641 31196 165907 32371
rect 39950 29869 40206 30099
rect 164657 20640 165923 21815
rect 164641 14962 165907 16137
rect 164641 7869 165907 9044
<< metal4 >>
rect 82797 351150 85297 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 164647 351150 167147 352400
rect 82963 349244 84999 351150
rect 88168 349208 90204 351150
rect 108814 349155 110850 351150
rect 114054 349155 116090 351150
rect 159668 349191 161704 351150
rect 164874 349155 166910 351150
rect 164359 341807 166659 342174
rect 164270 341177 166659 341807
rect 163899 339949 166659 341177
rect 163899 338774 164500 339949
rect 165766 338774 166659 339949
rect 163899 337301 166659 338774
rect 241132 337306 243344 338090
rect 243555 337802 243747 337814
rect 243555 337682 243571 337802
rect 243704 337737 243747 337802
rect 243704 337682 244231 337737
rect 243555 337669 244231 337682
rect 243555 337668 243747 337669
rect 163899 333969 166665 337301
rect 163791 332863 166665 333969
rect 163791 331688 164481 332863
rect 165747 331688 166665 332863
rect 163791 331547 166665 331688
rect 28402 331370 28612 331410
rect 28402 331218 28429 331370
rect 28585 331218 28612 331370
rect 28402 330731 28612 331218
rect 28977 331369 29187 331403
rect 28977 331217 29002 331369
rect 29158 331217 29187 331369
rect 28977 330724 29187 331217
rect 163789 330649 166665 331547
rect 164365 328716 166665 330649
rect 164359 328349 166665 328716
rect 164270 327719 166665 328349
rect 163899 326491 166665 327719
rect 163899 325316 164500 326491
rect 165766 325316 166665 326491
rect 163899 320511 166665 325316
rect 163791 319405 166665 320511
rect 163791 318230 164481 319405
rect 165747 318230 166665 319405
rect 163791 318089 166665 318230
rect 163789 317191 166665 318089
rect 24667 316962 25534 316964
rect 24667 316943 25997 316962
rect 24667 316893 25927 316943
rect 25978 316893 25997 316943
rect 24667 316882 25997 316893
rect 24667 316761 25534 316882
rect 24667 316742 26006 316761
rect 24667 316692 25936 316742
rect 25987 316692 26006 316742
rect 24667 316681 26006 316692
rect 24667 316438 25534 316681
rect 24670 316361 25532 316438
rect 24670 316342 25991 316361
rect 24670 316292 25921 316342
rect 25972 316292 25991 316342
rect 24670 316281 25991 316292
rect 24670 316072 25532 316281
rect 24670 316053 25991 316072
rect 24670 316003 25921 316053
rect 25972 316003 25991 316053
rect 24670 315992 25991 316003
rect 24670 315721 25532 315992
rect 24670 315702 25997 315721
rect 24670 315652 25927 315702
rect 25978 315652 25997 315702
rect 24670 315641 25997 315652
rect 24670 301000 25532 315641
rect 164365 314088 166665 317191
rect 164276 313458 166665 314088
rect 163905 312230 166665 313458
rect 163905 311055 164506 312230
rect 165772 311055 166665 312230
rect 163905 306250 166665 311055
rect 163797 305144 166665 306250
rect 163797 303969 164487 305144
rect 165753 303969 166665 305144
rect 163797 303828 166665 303969
rect 163795 302921 166665 303828
rect 163905 302753 166665 302921
rect 164365 301000 166665 302753
rect 241132 337283 244009 337306
rect 241132 337228 243932 337283
rect 243984 337228 244009 337283
rect 241132 337208 244009 337228
rect 241132 334841 243344 337208
rect 243506 335283 244150 335311
rect 243506 335143 243515 335283
rect 243666 335143 244150 335283
rect 243506 335128 244150 335143
rect 241132 334815 243924 334841
rect 241132 334765 243852 334815
rect 243904 334765 243924 334815
rect 241132 334737 243924 334765
rect 241132 329591 243344 334737
rect 247049 330024 247236 330039
rect 247049 329881 247062 330024
rect 247219 329881 247236 330024
rect 247049 329859 247236 329881
rect 241132 329554 247591 329591
rect 241132 329454 247459 329554
rect 247560 329454 247591 329554
rect 241132 329410 247591 329454
rect 241132 327660 243344 329410
rect 241132 327511 247307 327660
rect 241132 325878 243344 327511
rect 241132 325729 247285 325878
rect 241132 324107 243344 325729
rect 241132 323958 247312 324107
rect 241132 318705 243344 323958
rect 245408 319188 245640 319191
rect 245408 319175 246066 319188
rect 245408 319023 245432 319175
rect 245588 319023 246066 319175
rect 245408 319013 246066 319023
rect 245408 319001 245640 319013
rect 241132 318670 245856 318705
rect 241132 318620 245761 318670
rect 245811 318620 245856 318670
rect 241132 318570 245856 318620
rect 241132 316244 243344 318570
rect 245385 316705 245617 316713
rect 245385 316692 245985 316705
rect 245385 316540 245417 316692
rect 245576 316540 245985 316692
rect 245385 316529 245985 316540
rect 245385 316523 245617 316529
rect 241132 316204 245768 316244
rect 241132 316154 245682 316204
rect 245732 316154 245768 316204
rect 241132 316109 245768 316154
rect 241132 313866 243344 316109
rect 245501 314300 245547 314305
rect 245501 314291 245902 314300
rect 245207 314266 245902 314291
rect 245207 314132 245226 314266
rect 245364 314132 245902 314266
rect 245207 314114 245902 314132
rect 245501 314107 245902 314114
rect 245501 314093 245547 314107
rect 241132 313819 245684 313866
rect 241132 313769 245602 313819
rect 245652 313769 245684 313819
rect 241132 313740 245684 313769
rect 241132 311381 243344 313740
rect 245128 311854 245825 311890
rect 245128 311699 245151 311854
rect 245319 311699 245825 311854
rect 245128 311676 245825 311699
rect 241132 311353 245610 311381
rect 241132 311303 245523 311353
rect 245573 311303 245610 311353
rect 241132 311275 245610 311303
rect 241132 308994 243344 311275
rect 245072 309456 245751 309488
rect 245072 309309 245095 309456
rect 245251 309309 245751 309456
rect 245072 309282 245751 309309
rect 241132 308967 245508 308994
rect 241132 308917 245443 308967
rect 245493 308917 245508 308967
rect 241132 308897 245508 308917
rect 241132 306523 243344 308897
rect 244991 307058 245669 307089
rect 244991 306904 245010 307058
rect 245165 306904 245669 307058
rect 244991 306887 245669 306904
rect 241132 306501 245439 306523
rect 241132 306451 245363 306501
rect 245413 306451 245439 306501
rect 241132 306426 245439 306451
rect 241132 301000 243344 306426
rect 11000 299000 280000 301000
rect 164365 297099 166665 299000
rect 163994 295871 166665 297099
rect 163994 294696 164595 295871
rect 165861 294696 166665 295871
rect 163994 289891 166665 294696
rect 163886 288785 166665 289891
rect 163886 287610 164576 288785
rect 165842 287610 166665 288785
rect 163886 287469 166665 287610
rect 163884 286562 166665 287469
rect 163994 282383 166665 286562
rect 163994 281208 164539 282383
rect 165805 282016 166665 282383
rect 165805 281208 166759 282016
rect 163994 281056 166759 281208
rect 163992 280229 166759 281056
rect 164356 274691 166759 280229
rect 273495 276989 275423 277344
rect 273495 275847 273813 276989
rect 275123 275847 275423 276989
rect 273495 275548 275423 275847
rect 164045 273463 166759 274691
rect 164045 272288 164646 273463
rect 165912 272547 166759 273463
rect 165912 272524 166735 272547
rect 165912 272288 166716 272524
rect 164045 267483 166716 272288
rect 28721 266590 28859 267193
rect 26420 266258 28859 266590
rect 28721 265891 28859 266258
rect 163937 266377 166716 267483
rect 163937 265202 164627 266377
rect 165893 265202 166716 266377
rect 229932 266148 234831 266175
rect 229932 266001 230173 266148
rect 230330 266144 234831 266148
rect 230330 266001 230413 266144
rect 229932 265997 230413 266001
rect 230570 266142 234831 266144
rect 230570 265997 230649 266142
rect 229932 265995 230649 265997
rect 230806 266139 234831 266142
rect 230806 265995 230895 266139
rect 229932 265992 230895 265995
rect 231052 265992 234831 266139
rect 229932 265953 234831 265992
rect 266660 265320 267646 266008
rect 163937 265061 166716 265202
rect 266009 265300 267646 265320
rect 266009 265202 266024 265300
rect 266126 265202 267646 265300
rect 266009 265179 267646 265202
rect 26424 264775 26589 264812
rect 26424 264665 26446 264775
rect 26561 264665 26589 264775
rect 26424 264625 26589 264665
rect 28636 263423 28777 264812
rect 163935 264154 166716 265061
rect 18465 263165 20622 263265
rect 18465 262910 21722 263165
rect 18465 257000 20622 262910
rect 164045 259975 166716 264154
rect 230106 263775 234757 263808
rect 230106 263772 230409 263775
rect 230106 263625 230168 263772
rect 230325 263628 230409 263772
rect 230566 263771 234757 263775
rect 230566 263628 230645 263771
rect 230325 263625 230645 263628
rect 230106 263624 230645 263625
rect 230802 263624 230878 263771
rect 231035 263624 234757 263771
rect 230106 263599 234757 263624
rect 266660 262962 267646 265179
rect 265929 262942 267646 262962
rect 265929 262844 265944 262942
rect 266046 262844 267646 262942
rect 265929 262821 267646 262844
rect 229767 261289 233522 261293
rect 229767 261269 234677 261289
rect 229767 261267 230426 261269
rect 229767 261120 230199 261267
rect 230356 261122 230426 261267
rect 230583 261122 230643 261269
rect 230800 261267 234677 261269
rect 230800 261122 230862 261267
rect 230356 261120 230862 261122
rect 231019 261120 234677 261267
rect 229767 261115 234677 261120
rect 230922 261111 234677 261115
rect 266660 260481 267646 262821
rect 265847 260457 267646 260481
rect 265847 260359 265865 260457
rect 265967 260359 267646 260457
rect 265847 260332 267646 260359
rect 164045 258800 164590 259975
rect 165856 259608 166716 259975
rect 165856 258800 166810 259608
rect 164045 258648 166810 258800
rect 164043 257821 166810 258648
rect 164365 257000 166810 257821
rect 266660 257000 267646 260332
rect 10000 256982 62683 257000
rect 70642 256982 275000 257000
rect 10000 255000 275000 256982
rect 164365 250449 166665 255000
rect 164365 250437 166790 250449
rect 164076 249209 166790 250437
rect 164076 248034 164677 249209
rect 165943 248293 166790 249209
rect 165943 248270 166766 248293
rect 165943 248034 166747 248270
rect 164076 243229 166747 248034
rect 163968 242123 166747 243229
rect 242644 242302 242798 242305
rect 27160 241019 32004 241039
rect 27160 241014 27403 241019
rect 27160 240838 27170 241014
rect 27341 240843 27403 241014
rect 27574 240843 32004 241019
rect 27341 240838 32004 240843
rect 27160 240822 32004 240838
rect 63989 240238 65695 241256
rect 163968 240948 164658 242123
rect 165924 240948 166747 242123
rect 242643 242271 242798 242302
rect 242643 242153 242652 242271
rect 242787 242153 242798 242271
rect 242643 242101 242798 242153
rect 242643 241983 242654 242101
rect 242789 241983 242798 242101
rect 242643 241939 242798 241983
rect 242643 241821 242651 241939
rect 242786 241821 242798 241939
rect 242643 241798 242798 241821
rect 242643 241713 242792 241798
rect 163968 240807 166747 240948
rect 242644 241013 242792 241713
rect 242644 240947 242684 241013
rect 242756 240947 242792 241013
rect 242644 240939 242792 240947
rect 63180 240219 65695 240238
rect 63180 240105 63189 240219
rect 63304 240105 65695 240219
rect 63180 240095 65695 240105
rect 27092 238592 31936 238610
rect 27092 238416 27144 238592
rect 27315 238416 27403 238592
rect 27574 238416 31936 238592
rect 27092 238393 31936 238416
rect 63989 237902 65695 240095
rect 163966 239900 166747 240807
rect 63101 237883 65695 237902
rect 63101 237769 63110 237883
rect 63225 237769 65695 237883
rect 63101 237759 65695 237769
rect 27013 236134 31857 236153
rect 27013 235958 27109 236134
rect 27280 236130 31857 236134
rect 27280 235958 27376 236130
rect 27013 235954 27376 235958
rect 27547 235954 31857 236130
rect 27013 235936 31857 235954
rect 63989 235418 65695 237759
rect 63020 235399 65695 235418
rect 63020 235285 63029 235399
rect 63144 235285 65695 235399
rect 63020 235275 65695 235285
rect 27013 233961 31857 233976
rect 27013 233785 27061 233961
rect 27232 233785 27346 233961
rect 27517 233785 31857 233961
rect 27013 233759 31857 233785
rect 63989 233211 65695 235275
rect 164076 235721 166747 239900
rect 164076 234546 164621 235721
rect 165887 235354 166747 235721
rect 165887 234546 166841 235354
rect 164076 234394 166841 234546
rect 164074 233567 166841 234394
rect 63024 233192 65695 233211
rect 63024 233078 63033 233192
rect 63148 233078 65695 233192
rect 63024 233068 65695 233078
rect 63989 232000 65695 233068
rect 164365 233402 166841 233567
rect 164365 232000 166665 233402
rect 243457 232000 243989 234641
rect 246008 232000 246540 234632
rect 251025 232000 251514 235394
rect 11000 230004 276000 232000
rect 11000 230000 58746 230004
rect 61078 230000 267314 230004
rect 269474 230000 276000 230004
rect 141157 229989 144509 230000
rect 164200 228943 166666 230000
rect 231612 229991 234962 230000
rect 164200 227768 164801 228943
rect 166067 227768 166666 228943
rect 164200 227671 166666 227768
rect 164200 226887 166717 227671
rect 36596 225511 36738 225709
rect 36596 225389 36608 225511
rect 36727 225389 36738 225511
rect 36596 225326 36738 225389
rect 36596 225204 36610 225326
rect 36729 225204 36738 225326
rect 36596 225144 36738 225204
rect 36596 225022 36608 225144
rect 36727 225022 36738 225144
rect 36596 223492 36738 225022
rect 164365 224776 166665 226887
rect 164180 223081 166665 224776
rect 37934 221852 38078 222960
rect 36774 221726 38078 221852
rect 164180 221906 164781 223081
rect 166047 221906 166665 223081
rect 164180 221809 166665 221906
rect 36774 221670 38069 221726
rect 36784 220934 36926 221670
rect 37207 220934 37398 221670
rect 37707 220934 37849 221670
rect 164180 221025 166697 221809
rect 36784 220743 37849 220934
rect 36784 220000 36926 220743
rect 37207 220000 37398 220743
rect 37707 220000 37849 220743
rect 164365 220000 166665 221025
rect 10000 218000 275000 220000
rect 164365 213295 166665 218000
rect 164220 212168 166665 213295
rect 164220 211018 166686 212168
rect 164220 209843 164821 211018
rect 166087 209843 166686 211018
rect 164220 209746 166686 209843
rect 164220 208839 166737 209746
rect 164220 205038 166665 208839
rect 164112 203932 166665 205038
rect 164112 202757 164802 203932
rect 166068 202757 166665 203932
rect 164112 202616 166665 202757
rect 164110 201709 166665 202616
rect 164220 197530 166665 201709
rect 164220 196355 164765 197530
rect 166031 196355 166665 197530
rect 164220 196203 166665 196355
rect 164218 194676 166665 196203
rect 164207 194275 166665 194676
rect 164207 193125 166673 194275
rect 164207 191950 164808 193125
rect 166074 191950 166673 193125
rect 164207 191853 166673 191950
rect 164207 190946 166724 191853
rect 27587 187275 30331 187301
rect 27587 187145 27672 187275
rect 27843 187271 30331 187275
rect 27843 187145 27936 187271
rect 27587 187141 27936 187145
rect 28107 187141 28236 187271
rect 28407 187141 30331 187271
rect 164207 187145 166665 190946
rect 27587 187109 30331 187141
rect 62513 186521 64054 186993
rect 61504 186500 64054 186521
rect 61504 186400 61518 186500
rect 61626 186400 64054 186500
rect 61504 186381 64054 186400
rect 27501 184893 30245 184918
rect 27501 184763 27728 184893
rect 27899 184888 28223 184893
rect 27899 184763 27987 184888
rect 27501 184758 27987 184763
rect 28158 184763 28223 184888
rect 28394 184763 30245 184893
rect 28158 184758 30245 184763
rect 27501 184726 30245 184758
rect 62513 184098 64054 186381
rect 164099 186039 166665 187145
rect 164099 184864 164789 186039
rect 166055 184864 166665 186039
rect 164099 184723 166665 184864
rect 61424 184077 64054 184098
rect 61424 183977 61438 184077
rect 61546 183977 64054 184077
rect 61424 183958 64054 183977
rect 27427 182427 30171 182461
rect 27427 182297 27751 182427
rect 27922 182297 27982 182427
rect 28153 182297 28227 182427
rect 28398 182297 30171 182427
rect 27427 182269 30171 182297
rect 62513 181614 64054 183958
rect 164097 183816 166665 184723
rect 61345 181593 64054 181614
rect 61345 181493 61359 181593
rect 61467 181493 64054 181593
rect 61345 181474 64054 181493
rect 27431 180169 30175 180208
rect 27431 180039 27723 180169
rect 27894 180039 27959 180169
rect 28130 180039 28209 180169
rect 28380 180039 30175 180169
rect 27431 180016 30175 180039
rect 62513 179463 64054 181474
rect 61336 179442 64054 179463
rect 61336 179342 61360 179442
rect 61468 179342 64054 179442
rect 61336 179323 64054 179342
rect 35548 171266 35763 171272
rect 35547 171142 38630 171266
rect 27897 170817 32147 170839
rect 35548 170825 35763 171142
rect 27897 170816 28218 170817
rect 27897 170624 27924 170816
rect 28106 170625 28218 170816
rect 28400 170625 32147 170817
rect 28106 170624 32147 170625
rect 27897 170608 32147 170624
rect 32734 169146 33021 169470
rect 32579 165000 33270 169146
rect 62513 165000 64054 179323
rect 164207 179637 166665 183816
rect 164207 178462 164752 179637
rect 166018 178462 166665 179637
rect 164207 178310 166665 178462
rect 164205 176358 166665 178310
rect 164365 175011 166665 176358
rect 164030 174818 166665 175011
rect 163922 173712 166665 174818
rect 163922 172537 164612 173712
rect 165878 172537 166665 173712
rect 163922 172396 166665 172537
rect 163920 171489 166665 172396
rect 164030 167310 166665 171489
rect 164030 166135 164575 167310
rect 165841 166135 166665 167310
rect 164030 165983 166665 166135
rect 164028 165000 166665 165983
rect 11000 163000 276000 165000
rect 164365 160826 166665 163000
rect 164148 160049 167097 160826
rect 164148 158874 164841 160049
rect 166107 158874 167097 160049
rect 164148 158644 167097 158874
rect 164148 158070 167148 158644
rect 164365 155993 166665 158070
rect 164365 155209 167382 155993
rect 164365 154034 164822 155209
rect 166088 154034 167382 155209
rect 164365 153811 167382 154034
rect 164365 153237 167433 153811
rect 164365 150733 166665 153237
rect 164365 149939 167453 150733
rect 164365 148764 164803 149939
rect 166069 148764 167453 149939
rect 164365 148551 167453 148764
rect 164365 147977 167504 148551
rect 164365 145259 166665 147977
rect 164365 144387 167382 145259
rect 164365 143212 164785 144387
rect 166051 143212 167382 144387
rect 232782 143586 237864 143606
rect 232782 143583 234136 143586
rect 232782 143377 233504 143583
rect 233720 143377 233803 143583
rect 234019 143380 234136 143583
rect 234352 143583 237864 143586
rect 234352 143380 234419 143583
rect 234019 143377 234419 143380
rect 234635 143377 237864 143583
rect 232782 143365 237864 143377
rect 234498 143364 237864 143365
rect 164365 143077 167382 143212
rect 164365 142503 167433 143077
rect 270847 142813 272858 143119
rect 269026 142783 272858 142813
rect 269026 142679 269050 142783
rect 269160 142679 272858 142783
rect 269026 142654 272858 142679
rect 164365 139147 166665 142503
rect 234416 141214 237782 141216
rect 233039 141204 237782 141214
rect 233039 140998 233595 141204
rect 233811 141201 237782 141204
rect 233811 141198 234187 141201
rect 233811 140998 233915 141198
rect 233039 140992 233915 140998
rect 234131 140995 234187 141198
rect 234403 141198 237782 141201
rect 234403 140995 234462 141198
rect 234131 140992 234462 140995
rect 234678 140992 237782 141198
rect 233039 140974 237782 140992
rect 233039 140973 235327 140974
rect 270847 140419 272858 142654
rect 270754 140414 272858 140419
rect 268956 140387 272858 140414
rect 268956 140283 268969 140387
rect 269079 140283 272858 140387
rect 268956 140260 272858 140283
rect 270754 140258 272858 140260
rect 164365 138197 167524 139147
rect 234336 138761 237702 138762
rect 233130 138747 237702 138761
rect 233130 138744 234158 138747
rect 233130 138538 233536 138744
rect 233752 138538 233854 138744
rect 234070 138541 234158 138744
rect 234374 138541 234435 138747
rect 234651 138541 237702 138747
rect 234070 138538 237702 138541
rect 233130 138520 237702 138538
rect 164365 137022 164785 138197
rect 166051 137022 167524 138197
rect 270847 137976 272858 140258
rect 270706 137954 272858 137976
rect 268877 137927 272858 137954
rect 268877 137823 268890 137927
rect 269000 137823 272858 137927
rect 268877 137800 272858 137823
rect 270706 137789 272858 137800
rect 164365 136965 167524 137022
rect 164365 136391 167575 136965
rect 164365 131451 166665 136391
rect 164365 129091 167314 131451
rect 244745 130625 247049 130643
rect 244745 130459 244789 130625
rect 244953 130623 247049 130625
rect 244953 130459 244999 130623
rect 244745 130457 244999 130459
rect 245163 130457 247049 130623
rect 244745 130429 247049 130457
rect 164365 128188 167365 129091
rect 164365 127000 166665 128188
rect 248303 127000 248716 129374
rect 270847 127000 272858 137789
rect 12000 125000 277000 127000
rect 164365 120197 166665 125000
rect 164365 119093 166831 120197
rect 164365 117918 164793 119093
rect 166059 117918 166831 119093
rect 164365 117775 166831 117918
rect 164365 116868 166882 117775
rect 164365 112245 166665 116868
rect 164365 111166 167036 112245
rect 164365 109991 164902 111166
rect 166168 109991 167036 111166
rect 164365 109823 167036 109991
rect 164365 108916 167087 109823
rect 164365 104019 166665 108916
rect 164365 102964 167036 104019
rect 164365 101789 165003 102964
rect 166269 101789 167036 102964
rect 164365 101597 167036 101789
rect 164365 100690 167087 101597
rect 164365 96615 166665 100690
rect 164365 95465 166831 96615
rect 164365 94290 164966 95465
rect 166232 94290 166831 95465
rect 164365 94193 166831 94290
rect 164365 93286 166882 94193
rect 164365 89485 166665 93286
rect 164257 88379 166665 89485
rect 164257 87204 164947 88379
rect 166213 87204 166665 88379
rect 164257 87063 166665 87204
rect 164255 86156 166665 87063
rect 164365 81977 166665 86156
rect 164365 80802 164910 81977
rect 166176 80802 166665 81977
rect 164365 80650 166665 80802
rect 164363 75873 166716 80650
rect 7143 75808 242368 75873
rect 253842 75808 279373 75823
rect 7143 75789 279373 75808
rect 7143 75451 283186 75789
rect 7143 73748 281123 75451
rect 282980 73748 283186 75451
rect 7143 73486 283186 73748
rect 7143 73379 242368 73486
rect 247695 73413 283186 73486
rect 278502 73408 283186 73413
rect 164363 71584 166716 73379
rect 164231 70727 166716 71584
rect 164231 69552 164892 70727
rect 166158 69552 166716 70727
rect 164231 69470 166716 69552
rect 164229 69372 166716 69470
rect 164229 68908 166665 69372
rect 164365 65344 166665 68908
rect 164196 64732 166665 65344
rect 164196 63557 164818 64732
rect 166084 63557 166665 64732
rect 164196 63230 166665 63557
rect 164194 62668 166665 63230
rect 164365 59627 166665 62668
rect 164161 58904 166665 59627
rect 164161 57729 164855 58904
rect 166121 57729 166665 58904
rect 164161 57513 166665 57729
rect 164159 56951 166665 57513
rect 164365 53422 166665 56951
rect 164092 52817 166665 53422
rect 164092 51642 164929 52817
rect 166195 51642 166665 52817
rect 164092 51308 166665 51642
rect 164090 50746 166665 51308
rect 164365 45727 166665 50746
rect 24119 45664 27392 45667
rect 24119 45662 24978 45664
rect 24119 45659 24694 45662
rect 24119 45655 24430 45659
rect 24119 45531 24178 45655
rect 24302 45535 24430 45655
rect 24554 45538 24694 45659
rect 24818 45540 24978 45662
rect 25102 45659 27392 45664
rect 25102 45540 25207 45659
rect 24818 45538 25207 45540
rect 24554 45535 25207 45538
rect 25331 45657 27392 45659
rect 25331 45535 25464 45657
rect 24302 45533 25464 45535
rect 25588 45653 27392 45657
rect 25588 45533 25709 45653
rect 24302 45531 25709 45533
rect 24119 45529 25709 45531
rect 25833 45529 27392 45653
rect 24119 45514 27392 45529
rect 164349 45476 166665 45727
rect 163804 44959 166977 45476
rect 163804 43784 164641 44959
rect 165907 43784 166977 44959
rect 163804 43450 166977 43784
rect 163802 43049 166977 43450
rect 164349 42901 166665 43049
rect 164365 39433 166665 42901
rect 164349 39182 166665 39433
rect 163804 38665 166977 39182
rect 163804 37490 164641 38665
rect 165907 37490 166977 38665
rect 163804 37156 166977 37490
rect 163802 36755 166977 37156
rect 164349 36607 166665 36755
rect 164365 33139 166665 36607
rect 164349 32888 166665 33139
rect 163804 32371 166977 32888
rect 163804 31196 164641 32371
rect 165907 31196 166977 32371
rect 163804 30862 166977 31196
rect 163802 30461 166977 30862
rect 164349 30313 166665 30461
rect 39396 30099 40707 30135
rect 39396 29869 39950 30099
rect 40206 29869 40707 30099
rect 39396 28000 40707 29869
rect 46028 28000 48233 28003
rect 164365 28000 166665 30313
rect 11000 26000 276000 28000
rect 164365 22332 166665 26000
rect 163820 21815 166993 22332
rect 163820 20640 164657 21815
rect 165923 20640 166993 21815
rect 163820 20306 166993 20640
rect 163818 19905 166993 20306
rect 164365 16654 166665 19905
rect 163804 16137 166977 16654
rect 163804 14962 164641 16137
rect 165907 14962 166977 16137
rect 163804 14628 166977 14962
rect 163802 14227 166977 14628
rect 164365 9561 166665 14227
rect 163804 9044 166977 9561
rect 163804 7869 164641 9044
rect 165907 7869 166977 9044
rect 163804 7535 166977 7869
rect 163802 7134 166977 7535
rect 164365 6011 166665 7134
<< via4 >>
rect 243571 337682 243704 337802
rect 28429 331218 28585 331370
rect 29002 331217 29158 331369
rect 243515 335143 243666 335283
rect 247062 329881 247219 330024
rect 245432 319023 245588 319175
rect 245417 316540 245576 316692
rect 245226 314132 245364 314266
rect 245151 311699 245319 311854
rect 245095 309309 245251 309456
rect 245010 306904 245165 307058
rect 273813 275847 275123 276989
rect 22917 266518 23059 266651
rect 23442 266522 23582 266657
rect 230173 266001 230330 266148
rect 230413 265997 230570 266144
rect 230649 265995 230806 266142
rect 230895 265992 231052 266139
rect 230168 263625 230325 263772
rect 230409 263628 230566 263775
rect 230645 263624 230802 263771
rect 230878 263624 231035 263771
rect 230199 261120 230356 261267
rect 230426 261122 230583 261269
rect 230643 261122 230800 261269
rect 230862 261120 231019 261267
rect 27170 240838 27341 241014
rect 27403 240843 27574 241019
rect 242652 242153 242787 242271
rect 242654 241983 242789 242101
rect 242651 241821 242786 241939
rect 27144 238416 27315 238592
rect 27403 238416 27574 238592
rect 27109 235958 27280 236134
rect 27376 235954 27547 236130
rect 27061 233785 27232 233961
rect 27346 233785 27517 233961
rect 36608 225389 36727 225511
rect 36610 225204 36729 225326
rect 36608 225022 36727 225144
rect 27672 187145 27843 187275
rect 27936 187141 28107 187271
rect 28236 187141 28407 187271
rect 27728 184763 27899 184893
rect 27987 184758 28158 184888
rect 28223 184763 28394 184893
rect 27751 182297 27922 182427
rect 27982 182297 28153 182427
rect 28227 182297 28398 182427
rect 27723 180039 27894 180169
rect 27959 180039 28130 180169
rect 28209 180039 28380 180169
rect 27924 170624 28106 170816
rect 28218 170625 28400 170817
rect 233504 143377 233720 143583
rect 233803 143377 234019 143583
rect 234136 143380 234352 143586
rect 234419 143377 234635 143583
rect 233595 140998 233811 141204
rect 233915 140992 234131 141198
rect 234187 140995 234403 141201
rect 234462 140992 234678 141198
rect 233536 138538 233752 138744
rect 233854 138538 234070 138744
rect 234158 138541 234374 138747
rect 234435 138541 234651 138747
rect 244789 130459 244953 130625
rect 244999 130457 245163 130623
rect 24178 45531 24302 45655
rect 24430 45535 24554 45659
rect 24694 45538 24818 45662
rect 24978 45540 25102 45664
rect 25207 45535 25331 45659
rect 25464 45533 25588 45657
rect 25709 45529 25833 45653
<< metal5 >>
rect 82797 351150 85297 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 164647 351150 167147 352400
rect 82963 349244 84999 351150
rect 88168 349208 90204 351150
rect 108814 349155 110850 351150
rect 114054 349155 116090 351150
rect 159668 349191 161704 351150
rect 164874 349155 166910 351150
rect 10000 341000 279000 343000
rect 28333 331370 29338 341000
rect 100337 340994 103311 341000
rect 140522 340966 144447 341000
rect 156586 340685 160000 341000
rect 189353 340946 193169 341000
rect 156557 337000 160000 340685
rect 238022 337829 240372 341000
rect 238022 337802 243719 337829
rect 238022 337682 243571 337802
rect 243704 337682 243719 337802
rect 238022 337655 243719 337682
rect 156557 333969 159446 337000
rect 156478 332036 159446 333969
rect 28333 331218 28429 331370
rect 28585 331369 29338 331370
rect 28585 331218 29002 331369
rect 28333 331217 29002 331218
rect 29158 331217 29338 331369
rect 28333 331175 29338 331217
rect 156419 330649 159446 332036
rect 238022 335302 240372 337655
rect 238022 335283 243683 335302
rect 238022 335143 243515 335283
rect 243666 335143 243683 335283
rect 238022 335126 243683 335143
rect 157052 328716 159393 330649
rect 157046 328349 159393 328716
rect 156957 327719 159393 328349
rect 156586 327227 159393 327719
rect 156557 323816 159393 327227
rect 238022 330054 240372 335126
rect 238022 330024 247243 330054
rect 238022 329881 247062 330024
rect 247219 329881 247243 330024
rect 238022 329844 247243 329881
rect 156557 320511 159446 323816
rect 156478 318578 159446 320511
rect 156419 317191 159446 318578
rect 238022 319187 240372 329844
rect 238022 319175 245605 319187
rect 238022 319023 245432 319175
rect 245588 319023 245605 319175
rect 238022 319008 245605 319023
rect 157052 314088 159393 317191
rect 156963 313458 159393 314088
rect 156592 312966 159393 313458
rect 156563 309555 159393 312966
rect 238022 316709 240372 319008
rect 238022 316692 245596 316709
rect 238022 316540 245417 316692
rect 245576 316540 245596 316692
rect 238022 316527 245596 316540
rect 238022 314287 240372 316527
rect 238022 314286 245208 314287
rect 238022 314266 245383 314286
rect 238022 314132 245226 314266
rect 245364 314132 245383 314266
rect 238022 314115 245383 314132
rect 238022 311881 240372 314115
rect 238022 311854 245369 311881
rect 238022 311699 245151 311854
rect 245319 311699 245369 311854
rect 238022 311676 245369 311699
rect 156563 306250 159452 309555
rect 156484 304317 159452 306250
rect 238022 309474 240372 311676
rect 238022 309456 245265 309474
rect 238022 309309 245095 309456
rect 245251 309309 245265 309456
rect 238022 309295 245265 309309
rect 238022 307081 240372 309295
rect 238022 307058 245191 307081
rect 238022 306904 245010 307058
rect 245165 306904 245191 307058
rect 238022 306879 245191 306904
rect 238022 306014 240372 306879
rect 156425 302921 159452 304317
rect 156592 302753 159452 302921
rect 157052 297099 159393 302753
rect 156681 296607 159393 297099
rect 156652 293196 159393 296607
rect 156652 289891 159541 293196
rect 156573 287958 159541 289891
rect 156514 286562 159541 287958
rect 156681 286108 159541 286562
rect 156681 281545 159393 286108
rect 156622 281056 159393 281545
rect 156622 280229 159389 281056
rect 157010 277890 159389 280229
rect 255736 277912 260234 277918
rect 255736 277906 272994 277912
rect 255736 277890 275442 277906
rect 9908 276989 275442 277890
rect 9908 275847 273813 276989
rect 275123 275847 275442 276989
rect 9908 275136 275442 275847
rect 9908 275109 272994 275136
rect 9908 274976 260234 275109
rect 9908 274941 256191 274976
rect 9908 274937 14729 274941
rect 17925 274937 256191 274941
rect 22523 267082 24124 274937
rect 157010 274691 159444 274937
rect 156732 274199 159444 274691
rect 156703 270788 159444 274199
rect 156703 267483 159592 270788
rect 22903 266651 23075 267082
rect 22903 266518 22917 266651
rect 23059 266518 23075 266651
rect 22903 266505 23075 266518
rect 23424 266657 23603 267082
rect 23424 266522 23442 266657
rect 23582 266522 23603 266657
rect 22903 266504 23070 266505
rect 23424 266499 23603 266522
rect 156624 265550 159592 267483
rect 156565 264154 159592 265550
rect 156732 263700 159592 264154
rect 229206 266148 231073 274937
rect 229206 266001 230173 266148
rect 230330 266144 231073 266148
rect 230330 266001 230413 266144
rect 229206 265997 230413 266001
rect 230570 266142 231073 266144
rect 230570 265997 230649 266142
rect 229206 265995 230649 265997
rect 230806 266139 231073 266142
rect 230806 265995 230895 266139
rect 229206 265992 230895 265995
rect 231052 265992 231073 266139
rect 229206 263775 231073 265992
rect 229206 263772 230409 263775
rect 156732 259137 159444 263700
rect 229206 263625 230168 263772
rect 230325 263628 230409 263772
rect 230566 263771 231073 263775
rect 230566 263628 230645 263771
rect 230325 263625 230645 263628
rect 229206 263624 230645 263625
rect 230802 263624 230878 263771
rect 231035 263624 231073 263771
rect 229206 261269 231073 263624
rect 229206 261267 230426 261269
rect 229206 261120 230199 261267
rect 230356 261122 230426 261267
rect 230583 261122 230643 261269
rect 230800 261267 231073 261269
rect 230800 261122 230862 261267
rect 230356 261120 230862 261122
rect 231019 261120 231073 261267
rect 229206 260070 231073 261120
rect 156673 258648 159444 259137
rect 156673 257821 159440 258648
rect 157052 256386 159440 257821
rect 157052 253620 159393 256386
rect 156887 250449 159424 253620
rect 156887 250437 159475 250449
rect 156763 249945 159475 250437
rect 156734 246534 159475 249945
rect 122960 245000 130971 245011
rect 156734 245000 159623 246534
rect 9000 243072 274000 245000
rect 9000 243000 226843 243072
rect 234785 243000 239793 243072
rect 26157 241019 27614 243000
rect 122960 242990 130971 243000
rect 156655 241296 159623 243000
rect 242462 242271 243000 243072
rect 247735 243000 274000 243072
rect 242462 242153 242652 242271
rect 242787 242153 243000 242271
rect 242462 242101 243000 242153
rect 242462 241983 242654 242101
rect 242789 241983 243000 242101
rect 242462 241939 243000 241983
rect 242462 241821 242651 241939
rect 242786 241821 243000 241939
rect 242462 241804 243000 241821
rect 26157 241014 27403 241019
rect 26157 240838 27170 241014
rect 27341 240843 27403 241014
rect 27574 240843 27614 241019
rect 27341 240838 27614 240843
rect 26157 238592 27614 240838
rect 156596 239900 159623 241296
rect 26157 238416 27144 238592
rect 27315 238416 27403 238592
rect 27574 238416 27614 238592
rect 26157 236134 27614 238416
rect 26157 235958 27109 236134
rect 27280 236130 27614 236134
rect 27280 235958 27376 236130
rect 26157 235954 27376 235958
rect 27547 235954 27614 236130
rect 26157 233961 27614 235954
rect 156763 239446 159623 239900
rect 156763 234883 159475 239446
rect 26157 233785 27061 233961
rect 27232 233785 27346 233961
rect 27517 233785 27614 233961
rect 26157 233383 27614 233785
rect 156704 234394 159475 234883
rect 156704 233567 159471 234394
rect 157052 233402 159471 233567
rect 157052 230638 159393 233402
rect 156887 230093 159393 230638
rect 156887 229679 159394 230093
rect 156858 227000 159445 229679
rect 10000 225511 275000 227000
rect 10000 225389 36608 225511
rect 36727 225389 275000 225511
rect 10000 225326 275000 225389
rect 10000 225204 36610 225326
rect 36729 225204 275000 225326
rect 10000 225144 275000 225204
rect 10000 225022 36608 225144
rect 36727 225022 275000 225144
rect 10000 225000 275000 225022
rect 157052 224776 159393 225000
rect 156867 223817 159393 224776
rect 156838 221025 159425 223817
rect 157052 213295 159393 221025
rect 156907 212168 159393 213295
rect 156907 211754 159414 212168
rect 156878 205038 159465 211754
rect 156799 203105 159465 205038
rect 156740 202843 159465 203105
rect 156740 201709 159393 202843
rect 156907 196692 159393 201709
rect 156848 194275 159393 196692
rect 156848 193861 159401 194275
rect 156848 193531 159452 193861
rect 27342 187275 28458 187920
rect 27342 187145 27672 187275
rect 27843 187271 28458 187275
rect 27843 187145 27936 187271
rect 27342 187141 27936 187145
rect 28107 187141 28236 187271
rect 28407 187141 28458 187271
rect 156865 187145 159452 193531
rect 27342 184893 28458 187141
rect 156786 185212 159452 187145
rect 27342 184763 27728 184893
rect 27899 184888 28223 184893
rect 27899 184763 27987 184888
rect 27342 184758 27987 184763
rect 28158 184763 28223 184888
rect 28394 184763 28458 184893
rect 28158 184758 28458 184763
rect 27342 182427 28458 184758
rect 156727 184950 159452 185212
rect 156727 183816 159393 184950
rect 27342 182297 27751 182427
rect 27922 182297 27982 182427
rect 28153 182297 28227 182427
rect 28398 182297 28458 182427
rect 27342 180169 28458 182297
rect 27342 180039 27723 180169
rect 27894 180039 27959 180169
rect 28130 180039 28209 180169
rect 28380 180039 28458 180169
rect 27342 177000 28458 180039
rect 156894 178799 159393 183816
rect 156835 177000 159393 178799
rect 12000 175016 277000 177000
rect 12000 175000 58627 175016
rect 61148 175000 277000 175016
rect 27364 171169 28450 175000
rect 156688 174818 159393 175000
rect 156609 172885 159393 174818
rect 156550 171489 159393 172885
rect 27362 170817 28452 171169
rect 27362 170816 28218 170817
rect 27362 170624 27924 170816
rect 28106 170625 28218 170816
rect 28400 170625 28452 170817
rect 28106 170624 28452 170625
rect 27362 170528 28452 170624
rect 156717 166472 159393 171489
rect 156658 164985 159393 166472
rect 157052 160826 159393 164985
rect 156835 158070 159825 160826
rect 157052 155993 159393 158070
rect 157052 153237 160110 155993
rect 157052 150733 159393 153237
rect 157052 147977 160181 150733
rect 157052 145259 159393 147977
rect 157052 142503 160110 145259
rect 232121 143586 234728 144087
rect 232121 143583 234136 143586
rect 232121 143377 233504 143583
rect 233720 143377 233803 143583
rect 234019 143380 234136 143583
rect 234352 143583 234728 143586
rect 234352 143380 234419 143583
rect 234019 143377 234419 143380
rect 234635 143377 234728 143583
rect 157052 139147 159393 142503
rect 232121 141204 234728 143377
rect 232121 140998 233595 141204
rect 233811 141201 234728 141204
rect 233811 141198 234187 141201
rect 233811 140998 233915 141198
rect 232121 140992 233915 140998
rect 234131 140995 234187 141198
rect 234403 141198 234728 141201
rect 234403 140995 234462 141198
rect 234131 140992 234462 140995
rect 234678 140992 234728 141198
rect 157052 136391 160252 139147
rect 232121 138747 234728 140992
rect 232121 138744 234158 138747
rect 232121 138538 233536 138744
rect 233752 138538 233854 138744
rect 234070 138541 234158 138744
rect 234374 138541 234435 138747
rect 234651 138541 234728 138747
rect 234070 138538 234728 138541
rect 157052 135000 159393 136391
rect 232121 135000 234728 138538
rect 11000 133000 276000 135000
rect 157052 131451 159393 133000
rect 157052 128209 160042 131451
rect 244660 130625 245186 133000
rect 244660 130459 244789 130625
rect 244953 130623 245186 130625
rect 244953 130459 244999 130623
rect 244660 130457 244999 130459
rect 245163 130457 245186 130623
rect 244660 130410 245186 130457
rect 157052 128188 160040 128209
rect 157052 120197 159393 128188
rect 157052 116893 159559 120197
rect 157052 116868 159557 116893
rect 157052 112245 159393 116868
rect 157052 108941 159764 112245
rect 157052 108916 159762 108941
rect 157052 104019 159393 108916
rect 157052 100715 159764 104019
rect 157052 100690 159762 100715
rect 157052 96615 159393 100690
rect 157052 93311 159559 96615
rect 157052 93286 159557 93311
rect 157052 89485 159393 93286
rect 156944 87552 159393 89485
rect 156885 86156 159393 87552
rect 157052 81139 159393 86156
rect 156993 79768 159393 81139
rect 156993 71584 159391 79768
rect 156918 70211 159391 71584
rect 156918 69959 159393 70211
rect 156859 68908 159393 69959
rect 157052 65344 159393 68908
rect 156883 63719 159393 65344
rect 156824 62668 159393 63719
rect 157052 59627 159393 62668
rect 156848 58002 159393 59627
rect 156789 56951 159393 58002
rect 157052 53422 159393 56951
rect 156779 51797 159393 53422
rect 156720 50746 159393 51797
rect 157052 50000 159393 50746
rect 11000 48000 276000 50000
rect 22603 45664 25872 48000
rect 157052 45727 159393 48000
rect 22603 45662 24978 45664
rect 22603 45659 24694 45662
rect 22603 45655 24430 45659
rect 22603 45531 24178 45655
rect 24302 45535 24430 45655
rect 24554 45538 24694 45659
rect 24818 45540 24978 45662
rect 25102 45659 25872 45664
rect 25102 45540 25207 45659
rect 24818 45538 25207 45540
rect 24554 45535 25207 45538
rect 25331 45657 25872 45659
rect 25331 45535 25464 45657
rect 24302 45533 25464 45535
rect 25588 45653 25872 45657
rect 25588 45533 25709 45653
rect 24302 45531 25709 45533
rect 22603 45529 25709 45531
rect 25833 45529 25872 45653
rect 22603 44698 25872 45529
rect 157036 45476 159393 45727
rect 156491 43939 159705 45476
rect 156432 43049 159705 43939
rect 157036 42901 159393 43049
rect 157052 39433 159393 42901
rect 157036 39182 159393 39433
rect 156491 37645 159705 39182
rect 156432 36755 159705 37645
rect 157036 36607 159393 36755
rect 157052 33139 159393 36607
rect 157036 32888 159393 33139
rect 156491 31351 159705 32888
rect 156432 30461 159705 31351
rect 157036 30313 159393 30461
rect 157052 22332 159393 30313
rect 156507 20795 159721 22332
rect 156448 19905 159721 20795
rect 157052 16654 159393 19905
rect 156491 15117 159705 16654
rect 156432 14227 159705 15117
rect 157052 9561 159393 14227
rect 156491 8024 159705 9561
rect 156432 7134 159705 8024
rect 157052 6011 159393 7134
<< comment >>
rect -50 352000 292050 352050
rect -50 0 0 352000
rect 292000 0 292050 352000
rect -50 -50 292050 0
use filter  filter_1
timestamp 1640983258
transform 1 0 38025 0 1 41313
box -1800 -11005 6240 390
use divbuf  divbuf_19
timestamp 1641017053
transform 1 0 27511 0 1 45357
box -460 -1085 31200 495
use pd  pd_5
timestamp 1644268929
transform 1 0 38673 0 1 170517
box -215 -855 1685 810
use divider  divider_3
timestamp 1644268929
transform 1 0 31863 0 1 169542
box -490 -235 4690 2150
use divider  divider_0
timestamp 1644268929
transform 1 0 246803 0 1 129340
box -490 -235 4690 2150
use divbuf  divbuf_25
timestamp 1641017053
transform 1 0 237817 0 1 138431
box -460 -1085 31200 495
use divbuf  divbuf_24
timestamp 1641017053
transform 1 0 237896 0 1 140897
box -460 -1085 31200 495
use divbuf  divbuf_23
timestamp 1641017053
transform 1 0 237976 0 1 143283
box -460 -1085 31200 495
use divbuf  divbuf_18
timestamp 1641017053
transform 1 0 30445 0 1 186973
box -460 -1085 31200 495
use divbuf  divbuf_17
timestamp 1641017053
transform 1 0 30365 0 1 184587
box -460 -1085 31200 495
use divbuf  divbuf_16
timestamp 1641017053
transform 1 0 30286 0 1 182121
box -460 -1085 31200 495
use divbuf  divbuf_15
timestamp 1641017053
transform 1 0 30286 0 1 179927
box -460 -1085 31200 495
use pd  pd_4
timestamp 1644268929
transform 1 0 36668 0 1 222858
box -215 -855 1685 810
use cp  cp_0
timestamp 1640911461
transform 1 0 21911 0 1 264642
box -415 -1715 4690 2035
use divbuf  divbuf_14
timestamp 1641017053
transform 1 0 31964 0 1 233669
box -460 -1085 31200 495
use divbuf  divbuf_13
timestamp 1641017053
transform 1 0 31964 0 1 235863
box -460 -1085 31200 495
use divbuf  divbuf_12
timestamp 1641017053
transform 1 0 32043 0 1 238329
box -460 -1085 31200 495
use divbuf  divbuf_11
timestamp 1641017053
transform 1 0 32123 0 1 240715
box -460 -1085 31200 495
use divbuf  divbuf_8
timestamp 1641017053
transform 1 0 28673 0 1 263178
box -460 -1085 31200 495
use ro_complete  ro_complete_0
timestamp 1644268929
transform 1 0 242309 0 1 239846
box -348 -5690 4661 1440
use divider  divider_1
timestamp 1644268929
transform 1 0 250269 0 1 235475
box -490 -235 4690 2150
use divbuf  divbuf_21
timestamp 1641017053
transform 1 0 234867 0 1 263433
box -460 -1085 31200 495
use divbuf  divbuf_20
timestamp 1641017053
transform 1 0 234788 0 1 260967
box -460 -1085 31200 495
use divbuf  divbuf_10
timestamp 1641017053
transform 1 0 28832 0 1 268030
box -460 -1085 31200 495
use divbuf  divbuf_9
timestamp 1641017053
transform 1 0 28752 0 1 265644
box -460 -1085 31200 495
use divbuf  divbuf_22
timestamp 1641017053
transform 1 0 234947 0 1 265819
box -460 -1085 31200 495
use divbuf  divbuf_7
timestamp 1641017053
transform 1 0 245779 0 1 306691
box -460 -1085 31200 495
use divbuf  divbuf_6
timestamp 1641017053
transform 1 0 245858 0 1 309157
box -460 -1085 31200 495
use divbuf  divbuf_5
timestamp 1641017053
transform 1 0 245938 0 1 311543
box -460 -1085 31200 495
use pll_full  pll_full_1
timestamp 1644268929
transform 1 0 31292 0 1 318138
box -5794 -2690 26430 12835
use ro_complete  ro_complete_1
timestamp 1644268929
transform 1 0 247313 0 1 328719
box -348 -5690 4661 1440
use divbuf  divbuf_2
timestamp 1641017053
transform 1 0 246097 0 1 316394
box -460 -1085 31200 495
use divbuf  divbuf_4
timestamp 1641017053
transform 1 0 246017 0 1 314009
box -460 -1085 31200 495
use divbuf  divbuf_1
timestamp 1641017053
transform 1 0 246176 0 1 318860
box -460 -1085 31200 495
use divbuf  divbuf_0
timestamp 1641017053
transform 1 0 244268 0 1 335005
box -460 -1085 31200 495
use divbuf  divbuf_3
timestamp 1641017053
transform 1 0 244347 0 1 337471
box -460 -1085 31200 495
<< labels >>
flabel metal3 s 291760 134615 292400 134671 0 FreeSans 560 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -400 190932 240 190988 0 FreeSans 560 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -400 169321 240 169377 0 FreeSans 560 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -400 147710 240 147766 0 FreeSans 560 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -400 126199 240 126255 0 FreeSans 560 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -400 62388 240 62444 0 FreeSans 560 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -400 40777 240 40833 0 FreeSans 560 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -400 19166 240 19222 0 FreeSans 560 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -400 8455 240 8511 0 FreeSans 560 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 291760 156826 292400 156882 0 FreeSans 560 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 291760 179437 292400 179493 0 FreeSans 560 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 291760 202648 292400 202704 0 FreeSans 560 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 291760 224859 292400 224915 0 FreeSans 560 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 291760 247070 292400 247126 0 FreeSans 560 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 291760 291781 292400 291837 0 FreeSans 560 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -400 255765 240 255821 0 FreeSans 560 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -400 234154 240 234210 0 FreeSans 560 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -400 212543 240 212599 0 FreeSans 560 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 291760 135206 292400 135262 0 FreeSans 560 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -400 190341 240 190397 0 FreeSans 560 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -400 168730 240 168786 0 FreeSans 560 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -400 147119 240 147175 0 FreeSans 560 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -400 125608 240 125664 0 FreeSans 560 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -400 61797 240 61853 0 FreeSans 560 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -400 40186 240 40242 0 FreeSans 560 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -400 18575 240 18631 0 FreeSans 560 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -400 7864 240 7920 0 FreeSans 560 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 291760 157417 292400 157473 0 FreeSans 560 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 291760 180028 292400 180084 0 FreeSans 560 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 291760 203239 292400 203295 0 FreeSans 560 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 291760 225450 292400 225506 0 FreeSans 560 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 291760 247661 292400 247717 0 FreeSans 560 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 291760 292372 292400 292428 0 FreeSans 560 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -400 255174 240 255230 0 FreeSans 560 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -400 233563 240 233619 0 FreeSans 560 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -400 211952 240 212008 0 FreeSans 560 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 291150 338992 292400 341492 0 FreeSans 560 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 340121 850 342621 0 FreeSans 560 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 283297 351150 285797 352400 0 FreeSans 960 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 232697 351150 235197 352400 0 FreeSans 960 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 206697 351150 209197 352400 0 FreeSans 960 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 164647 351150 167147 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 8097 351150 10597 352400 0 FreeSans 960 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 159497 351150 161997 352400 0 FreeSans 960 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 163397 351150 164497 352400 0 FreeSans 960 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 162147 351150 163247 352400 0 FreeSans 960 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 291760 1363 292400 1419 0 FreeSans 560 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 291760 204421 292400 204477 0 FreeSans 560 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 291760 226632 292400 226688 0 FreeSans 560 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 291760 248843 292400 248899 0 FreeSans 560 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 291760 293554 292400 293610 0 FreeSans 560 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -400 253992 240 254048 0 FreeSans 560 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -400 232381 240 232437 0 FreeSans 560 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -400 210770 240 210826 0 FreeSans 560 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -400 189159 240 189215 0 FreeSans 560 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -400 167548 240 167604 0 FreeSans 560 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -400 145937 240 145993 0 FreeSans 560 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 291760 3727 292400 3783 0 FreeSans 560 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -400 124426 240 124482 0 FreeSans 560 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -400 60615 240 60671 0 FreeSans 560 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -400 39004 240 39060 0 FreeSans 560 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -400 17393 240 17449 0 FreeSans 560 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -400 6682 240 6738 0 FreeSans 560 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -400 4318 240 4374 0 FreeSans 560 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -400 1954 240 2010 0 FreeSans 560 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 291760 6091 292400 6147 0 FreeSans 560 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 291760 8455 292400 8511 0 FreeSans 560 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 291760 10819 292400 10875 0 FreeSans 560 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 291760 24048 292400 24104 0 FreeSans 560 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 291760 46377 292400 46433 0 FreeSans 560 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 291760 136388 292400 136444 0 FreeSans 560 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 291760 158599 292400 158655 0 FreeSans 560 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 291760 181210 292400 181266 0 FreeSans 560 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 291760 772 292400 828 0 FreeSans 560 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 291760 203830 292400 203886 0 FreeSans 560 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 291760 226041 292400 226097 0 FreeSans 560 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 291760 248252 292400 248308 0 FreeSans 560 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 291760 292963 292400 293019 0 FreeSans 560 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -400 254583 240 254639 0 FreeSans 560 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -400 232972 240 233028 0 FreeSans 560 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -400 211361 240 211417 0 FreeSans 560 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -400 189750 240 189806 0 FreeSans 560 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -400 168139 240 168195 0 FreeSans 560 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -400 146528 240 146584 0 FreeSans 560 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 291760 3136 292400 3192 0 FreeSans 560 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -400 125017 240 125073 0 FreeSans 560 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -400 61206 240 61262 0 FreeSans 560 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -400 39595 240 39651 0 FreeSans 560 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -400 17984 240 18040 0 FreeSans 560 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -400 7273 240 7329 0 FreeSans 560 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -400 4909 240 4965 0 FreeSans 560 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -400 2545 240 2601 0 FreeSans 560 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 291760 5500 292400 5556 0 FreeSans 560 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 291760 7864 292400 7920 0 FreeSans 560 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 291760 10228 292400 10284 0 FreeSans 560 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 291760 23457 292400 23513 0 FreeSans 560 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 291760 45786 292400 45842 0 FreeSans 560 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 291760 135797 292400 135853 0 FreeSans 560 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 291760 158008 292400 158064 0 FreeSans 560 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 291760 180619 292400 180675 0 FreeSans 560 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 291760 2545 292400 2601 0 FreeSans 560 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 291760 205603 292400 205659 0 FreeSans 560 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 291760 227814 292400 227870 0 FreeSans 560 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 291760 250025 292400 250081 0 FreeSans 560 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 291760 294736 292400 294792 0 FreeSans 560 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -400 252810 240 252866 0 FreeSans 560 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -400 231199 240 231255 0 FreeSans 560 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -400 209588 240 209644 0 FreeSans 560 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -400 187977 240 188033 0 FreeSans 560 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -400 166366 240 166422 0 FreeSans 560 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -400 144755 240 144811 0 FreeSans 560 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 291760 4909 292400 4965 0 FreeSans 560 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -400 123244 240 123300 0 FreeSans 560 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -400 59433 240 59489 0 FreeSans 560 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -400 37822 240 37878 0 FreeSans 560 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -400 16211 240 16267 0 FreeSans 560 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -400 5500 240 5556 0 FreeSans 560 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -400 3136 240 3192 0 FreeSans 560 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -400 772 240 828 0 FreeSans 560 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 291760 7273 292400 7329 0 FreeSans 560 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 291760 9637 292400 9693 0 FreeSans 560 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 291760 12001 292400 12057 0 FreeSans 560 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 291760 25230 292400 25286 0 FreeSans 560 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 291760 47559 292400 47615 0 FreeSans 560 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 291760 137570 292400 137626 0 FreeSans 560 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 291760 159781 292400 159837 0 FreeSans 560 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 291760 182392 292400 182448 0 FreeSans 560 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 291760 1954 292400 2010 0 FreeSans 560 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 291760 205012 292400 205068 0 FreeSans 560 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 291760 227223 292400 227279 0 FreeSans 560 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 291760 249434 292400 249490 0 FreeSans 560 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 291760 294145 292400 294201 0 FreeSans 560 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -400 253401 240 253457 0 FreeSans 560 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -400 231790 240 231846 0 FreeSans 560 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -400 210179 240 210235 0 FreeSans 560 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -400 188568 240 188624 0 FreeSans 560 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -400 166957 240 167013 0 FreeSans 560 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -400 145346 240 145402 0 FreeSans 560 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 291760 4318 292400 4374 0 FreeSans 560 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -400 123835 240 123891 0 FreeSans 560 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -400 60024 240 60080 0 FreeSans 560 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -400 38413 240 38469 0 FreeSans 560 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -400 16802 240 16858 0 FreeSans 560 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -400 6091 240 6147 0 FreeSans 560 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -400 3727 240 3783 0 FreeSans 560 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -400 1363 240 1419 0 FreeSans 560 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 291760 6682 292400 6738 0 FreeSans 560 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 291760 9046 292400 9102 0 FreeSans 560 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 291760 11410 292400 11466 0 FreeSans 560 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 291760 24639 292400 24695 0 FreeSans 560 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 291760 46968 292400 47024 0 FreeSans 560 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 291760 136979 292400 137035 0 FreeSans 560 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 291760 159190 292400 159246 0 FreeSans 560 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 291760 181801 292400 181857 0 FreeSans 560 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 62908 -400 62964 240 0 FreeSans 560 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 240208 -400 240264 240 0 FreeSans 560 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 241981 -400 242037 240 0 FreeSans 560 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 243754 -400 243810 240 0 FreeSans 560 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 245527 -400 245583 240 0 FreeSans 560 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 247300 -400 247356 240 0 FreeSans 560 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 249073 -400 249129 240 0 FreeSans 560 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 250846 -400 250902 240 0 FreeSans 560 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 252619 -400 252675 240 0 FreeSans 560 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 254392 -400 254448 240 0 FreeSans 560 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 256165 -400 256221 240 0 FreeSans 560 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 80638 -400 80694 240 0 FreeSans 560 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 257938 -400 257994 240 0 FreeSans 560 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 259711 -400 259767 240 0 FreeSans 560 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 261484 -400 261540 240 0 FreeSans 560 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 263257 -400 263313 240 0 FreeSans 560 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 265030 -400 265086 240 0 FreeSans 560 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 266803 -400 266859 240 0 FreeSans 560 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 268576 -400 268632 240 0 FreeSans 560 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 270349 -400 270405 240 0 FreeSans 560 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 272122 -400 272178 240 0 FreeSans 560 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 273895 -400 273951 240 0 FreeSans 560 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 82411 -400 82467 240 0 FreeSans 560 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 275668 -400 275724 240 0 FreeSans 560 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 277441 -400 277497 240 0 FreeSans 560 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 279214 -400 279270 240 0 FreeSans 560 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 280987 -400 281043 240 0 FreeSans 560 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 282760 -400 282816 240 0 FreeSans 560 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 284533 -400 284589 240 0 FreeSans 560 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 286306 -400 286362 240 0 FreeSans 560 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 288079 -400 288135 240 0 FreeSans 560 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 84184 -400 84240 240 0 FreeSans 560 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 85957 -400 86013 240 0 FreeSans 560 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 87730 -400 87786 240 0 FreeSans 560 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 89503 -400 89559 240 0 FreeSans 560 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 91276 -400 91332 240 0 FreeSans 560 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 93049 -400 93105 240 0 FreeSans 560 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 94822 -400 94878 240 0 FreeSans 560 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 96595 -400 96651 240 0 FreeSans 560 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 64681 -400 64737 240 0 FreeSans 560 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 98368 -400 98424 240 0 FreeSans 560 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 100141 -400 100197 240 0 FreeSans 560 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 101914 -400 101970 240 0 FreeSans 560 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 103687 -400 103743 240 0 FreeSans 560 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 105460 -400 105516 240 0 FreeSans 560 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 107233 -400 107289 240 0 FreeSans 560 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 109006 -400 109062 240 0 FreeSans 560 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 110779 -400 110835 240 0 FreeSans 560 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 112552 -400 112608 240 0 FreeSans 560 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 114325 -400 114381 240 0 FreeSans 560 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 66454 -400 66510 240 0 FreeSans 560 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 116098 -400 116154 240 0 FreeSans 560 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 117871 -400 117927 240 0 FreeSans 560 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 119644 -400 119700 240 0 FreeSans 560 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 121417 -400 121473 240 0 FreeSans 560 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 123190 -400 123246 240 0 FreeSans 560 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 124963 -400 125019 240 0 FreeSans 560 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 126736 -400 126792 240 0 FreeSans 560 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 128509 -400 128565 240 0 FreeSans 560 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 130282 -400 130338 240 0 FreeSans 560 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 132055 -400 132111 240 0 FreeSans 560 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 68227 -400 68283 240 0 FreeSans 560 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 133828 -400 133884 240 0 FreeSans 560 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 135601 -400 135657 240 0 FreeSans 560 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 137374 -400 137430 240 0 FreeSans 560 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 139147 -400 139203 240 0 FreeSans 560 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 140920 -400 140976 240 0 FreeSans 560 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 142693 -400 142749 240 0 FreeSans 560 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 144466 -400 144522 240 0 FreeSans 560 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 146239 -400 146295 240 0 FreeSans 560 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 148012 -400 148068 240 0 FreeSans 560 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 149785 -400 149841 240 0 FreeSans 560 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 70000 -400 70056 240 0 FreeSans 560 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 151558 -400 151614 240 0 FreeSans 560 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 153331 -400 153387 240 0 FreeSans 560 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 155104 -400 155160 240 0 FreeSans 560 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 156877 -400 156933 240 0 FreeSans 560 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 158650 -400 158706 240 0 FreeSans 560 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 160423 -400 160479 240 0 FreeSans 560 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 162196 -400 162252 240 0 FreeSans 560 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 163969 -400 164025 240 0 FreeSans 560 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 165742 -400 165798 240 0 FreeSans 560 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 167515 -400 167571 240 0 FreeSans 560 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 71773 -400 71829 240 0 FreeSans 560 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 169288 -400 169344 240 0 FreeSans 560 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 171061 -400 171117 240 0 FreeSans 560 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 172834 -400 172890 240 0 FreeSans 560 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 174607 -400 174663 240 0 FreeSans 560 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 176380 -400 176436 240 0 FreeSans 560 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 178153 -400 178209 240 0 FreeSans 560 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 179926 -400 179982 240 0 FreeSans 560 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 181699 -400 181755 240 0 FreeSans 560 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 183472 -400 183528 240 0 FreeSans 560 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 185245 -400 185301 240 0 FreeSans 560 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 73546 -400 73602 240 0 FreeSans 560 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 187018 -400 187074 240 0 FreeSans 560 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 188791 -400 188847 240 0 FreeSans 560 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 190564 -400 190620 240 0 FreeSans 560 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 192337 -400 192393 240 0 FreeSans 560 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 194110 -400 194166 240 0 FreeSans 560 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 195883 -400 195939 240 0 FreeSans 560 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 197656 -400 197712 240 0 FreeSans 560 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 199429 -400 199485 240 0 FreeSans 560 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 201202 -400 201258 240 0 FreeSans 560 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 202975 -400 203031 240 0 FreeSans 560 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 75319 -400 75375 240 0 FreeSans 560 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 204748 -400 204804 240 0 FreeSans 560 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 206521 -400 206577 240 0 FreeSans 560 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 208294 -400 208350 240 0 FreeSans 560 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 210067 -400 210123 240 0 FreeSans 560 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 211840 -400 211896 240 0 FreeSans 560 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 213613 -400 213669 240 0 FreeSans 560 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 215386 -400 215442 240 0 FreeSans 560 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 217159 -400 217215 240 0 FreeSans 560 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 218932 -400 218988 240 0 FreeSans 560 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 220705 -400 220761 240 0 FreeSans 560 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 77092 -400 77148 240 0 FreeSans 560 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 222478 -400 222534 240 0 FreeSans 560 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 224251 -400 224307 240 0 FreeSans 560 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 226024 -400 226080 240 0 FreeSans 560 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 227797 -400 227853 240 0 FreeSans 560 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 229570 -400 229626 240 0 FreeSans 560 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 231343 -400 231399 240 0 FreeSans 560 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 233116 -400 233172 240 0 FreeSans 560 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 234889 -400 234945 240 0 FreeSans 560 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 236662 -400 236718 240 0 FreeSans 560 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 238435 -400 238491 240 0 FreeSans 560 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 78865 -400 78921 240 0 FreeSans 560 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 63499 -400 63555 240 0 FreeSans 560 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 240799 -400 240855 240 0 FreeSans 560 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 242572 -400 242628 240 0 FreeSans 560 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 244345 -400 244401 240 0 FreeSans 560 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 246118 -400 246174 240 0 FreeSans 560 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 247891 -400 247947 240 0 FreeSans 560 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 249664 -400 249720 240 0 FreeSans 560 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 251437 -400 251493 240 0 FreeSans 560 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 253210 -400 253266 240 0 FreeSans 560 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 254983 -400 255039 240 0 FreeSans 560 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 256756 -400 256812 240 0 FreeSans 560 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 81229 -400 81285 240 0 FreeSans 560 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 258529 -400 258585 240 0 FreeSans 560 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 260302 -400 260358 240 0 FreeSans 560 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 262075 -400 262131 240 0 FreeSans 560 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 263848 -400 263904 240 0 FreeSans 560 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 265621 -400 265677 240 0 FreeSans 560 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 267394 -400 267450 240 0 FreeSans 560 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 269167 -400 269223 240 0 FreeSans 560 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 270940 -400 270996 240 0 FreeSans 560 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 272713 -400 272769 240 0 FreeSans 560 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 274486 -400 274542 240 0 FreeSans 560 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 83002 -400 83058 240 0 FreeSans 560 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 276259 -400 276315 240 0 FreeSans 560 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 278032 -400 278088 240 0 FreeSans 560 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 279805 -400 279861 240 0 FreeSans 560 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 281578 -400 281634 240 0 FreeSans 560 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 283351 -400 283407 240 0 FreeSans 560 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 285124 -400 285180 240 0 FreeSans 560 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 286897 -400 286953 240 0 FreeSans 560 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 288670 -400 288726 240 0 FreeSans 560 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 84775 -400 84831 240 0 FreeSans 560 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 86548 -400 86604 240 0 FreeSans 560 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 88321 -400 88377 240 0 FreeSans 560 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 90094 -400 90150 240 0 FreeSans 560 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 91867 -400 91923 240 0 FreeSans 560 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 93640 -400 93696 240 0 FreeSans 560 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 95413 -400 95469 240 0 FreeSans 560 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 97186 -400 97242 240 0 FreeSans 560 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 65272 -400 65328 240 0 FreeSans 560 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 98959 -400 99015 240 0 FreeSans 560 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 100732 -400 100788 240 0 FreeSans 560 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 102505 -400 102561 240 0 FreeSans 560 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 104278 -400 104334 240 0 FreeSans 560 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 106051 -400 106107 240 0 FreeSans 560 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 107824 -400 107880 240 0 FreeSans 560 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 109597 -400 109653 240 0 FreeSans 560 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 111370 -400 111426 240 0 FreeSans 560 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 113143 -400 113199 240 0 FreeSans 560 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 114916 -400 114972 240 0 FreeSans 560 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 67045 -400 67101 240 0 FreeSans 560 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 116689 -400 116745 240 0 FreeSans 560 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 118462 -400 118518 240 0 FreeSans 560 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 120235 -400 120291 240 0 FreeSans 560 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 122008 -400 122064 240 0 FreeSans 560 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 123781 -400 123837 240 0 FreeSans 560 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 125554 -400 125610 240 0 FreeSans 560 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 127327 -400 127383 240 0 FreeSans 560 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 129100 -400 129156 240 0 FreeSans 560 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 130873 -400 130929 240 0 FreeSans 560 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 132646 -400 132702 240 0 FreeSans 560 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 68818 -400 68874 240 0 FreeSans 560 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 134419 -400 134475 240 0 FreeSans 560 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 136192 -400 136248 240 0 FreeSans 560 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 137965 -400 138021 240 0 FreeSans 560 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 139738 -400 139794 240 0 FreeSans 560 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 141511 -400 141567 240 0 FreeSans 560 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 143284 -400 143340 240 0 FreeSans 560 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 145057 -400 145113 240 0 FreeSans 560 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 146830 -400 146886 240 0 FreeSans 560 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 148603 -400 148659 240 0 FreeSans 560 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 150376 -400 150432 240 0 FreeSans 560 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 70591 -400 70647 240 0 FreeSans 560 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 152149 -400 152205 240 0 FreeSans 560 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 153922 -400 153978 240 0 FreeSans 560 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 155695 -400 155751 240 0 FreeSans 560 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 157468 -400 157524 240 0 FreeSans 560 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 159241 -400 159297 240 0 FreeSans 560 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 161014 -400 161070 240 0 FreeSans 560 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 162787 -400 162843 240 0 FreeSans 560 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 164560 -400 164616 240 0 FreeSans 560 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 166333 -400 166389 240 0 FreeSans 560 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 168106 -400 168162 240 0 FreeSans 560 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 72364 -400 72420 240 0 FreeSans 560 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 169879 -400 169935 240 0 FreeSans 560 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 171652 -400 171708 240 0 FreeSans 560 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 173425 -400 173481 240 0 FreeSans 560 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 175198 -400 175254 240 0 FreeSans 560 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 176971 -400 177027 240 0 FreeSans 560 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 178744 -400 178800 240 0 FreeSans 560 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 180517 -400 180573 240 0 FreeSans 560 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 182290 -400 182346 240 0 FreeSans 560 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 184063 -400 184119 240 0 FreeSans 560 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 185836 -400 185892 240 0 FreeSans 560 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 74137 -400 74193 240 0 FreeSans 560 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 187609 -400 187665 240 0 FreeSans 560 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 189382 -400 189438 240 0 FreeSans 560 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 191155 -400 191211 240 0 FreeSans 560 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 192928 -400 192984 240 0 FreeSans 560 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 194701 -400 194757 240 0 FreeSans 560 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 196474 -400 196530 240 0 FreeSans 560 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 198247 -400 198303 240 0 FreeSans 560 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 200020 -400 200076 240 0 FreeSans 560 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 201793 -400 201849 240 0 FreeSans 560 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 203566 -400 203622 240 0 FreeSans 560 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 75910 -400 75966 240 0 FreeSans 560 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 205339 -400 205395 240 0 FreeSans 560 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 207112 -400 207168 240 0 FreeSans 560 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 208885 -400 208941 240 0 FreeSans 560 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 210658 -400 210714 240 0 FreeSans 560 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 212431 -400 212487 240 0 FreeSans 560 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 214204 -400 214260 240 0 FreeSans 560 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 215977 -400 216033 240 0 FreeSans 560 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 217750 -400 217806 240 0 FreeSans 560 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 219523 -400 219579 240 0 FreeSans 560 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 221296 -400 221352 240 0 FreeSans 560 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 77683 -400 77739 240 0 FreeSans 560 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 223069 -400 223125 240 0 FreeSans 560 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 224842 -400 224898 240 0 FreeSans 560 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 226615 -400 226671 240 0 FreeSans 560 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 228388 -400 228444 240 0 FreeSans 560 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 230161 -400 230217 240 0 FreeSans 560 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 231934 -400 231990 240 0 FreeSans 560 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 233707 -400 233763 240 0 FreeSans 560 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 235480 -400 235536 240 0 FreeSans 560 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 237253 -400 237309 240 0 FreeSans 560 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 239026 -400 239082 240 0 FreeSans 560 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 79456 -400 79512 240 0 FreeSans 560 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 64090 -400 64146 240 0 FreeSans 560 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 241390 -400 241446 240 0 FreeSans 560 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 243163 -400 243219 240 0 FreeSans 560 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 244936 -400 244992 240 0 FreeSans 560 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 246709 -400 246765 240 0 FreeSans 560 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 248482 -400 248538 240 0 FreeSans 560 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 250255 -400 250311 240 0 FreeSans 560 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 252028 -400 252084 240 0 FreeSans 560 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 253801 -400 253857 240 0 FreeSans 560 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 255574 -400 255630 240 0 FreeSans 560 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 257347 -400 257403 240 0 FreeSans 560 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 81820 -400 81876 240 0 FreeSans 560 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 259120 -400 259176 240 0 FreeSans 560 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 260893 -400 260949 240 0 FreeSans 560 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 262666 -400 262722 240 0 FreeSans 560 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 264439 -400 264495 240 0 FreeSans 560 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 266212 -400 266268 240 0 FreeSans 560 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 267985 -400 268041 240 0 FreeSans 560 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 269758 -400 269814 240 0 FreeSans 560 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 271531 -400 271587 240 0 FreeSans 560 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 273304 -400 273360 240 0 FreeSans 560 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 275077 -400 275133 240 0 FreeSans 560 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 83593 -400 83649 240 0 FreeSans 560 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 276850 -400 276906 240 0 FreeSans 560 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 278623 -400 278679 240 0 FreeSans 560 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 280396 -400 280452 240 0 FreeSans 560 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 282169 -400 282225 240 0 FreeSans 560 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 283942 -400 283998 240 0 FreeSans 560 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 285715 -400 285771 240 0 FreeSans 560 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 287488 -400 287544 240 0 FreeSans 560 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 289261 -400 289317 240 0 FreeSans 560 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 85366 -400 85422 240 0 FreeSans 560 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 87139 -400 87195 240 0 FreeSans 560 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 88912 -400 88968 240 0 FreeSans 560 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 90685 -400 90741 240 0 FreeSans 560 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 92458 -400 92514 240 0 FreeSans 560 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 94231 -400 94287 240 0 FreeSans 560 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 96004 -400 96060 240 0 FreeSans 560 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 97777 -400 97833 240 0 FreeSans 560 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 65863 -400 65919 240 0 FreeSans 560 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 99550 -400 99606 240 0 FreeSans 560 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 101323 -400 101379 240 0 FreeSans 560 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 103096 -400 103152 240 0 FreeSans 560 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 104869 -400 104925 240 0 FreeSans 560 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 106642 -400 106698 240 0 FreeSans 560 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 108415 -400 108471 240 0 FreeSans 560 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 110188 -400 110244 240 0 FreeSans 560 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 111961 -400 112017 240 0 FreeSans 560 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 113734 -400 113790 240 0 FreeSans 560 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 115507 -400 115563 240 0 FreeSans 560 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 67636 -400 67692 240 0 FreeSans 560 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 117280 -400 117336 240 0 FreeSans 560 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 119053 -400 119109 240 0 FreeSans 560 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 120826 -400 120882 240 0 FreeSans 560 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 122599 -400 122655 240 0 FreeSans 560 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 124372 -400 124428 240 0 FreeSans 560 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 126145 -400 126201 240 0 FreeSans 560 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 127918 -400 127974 240 0 FreeSans 560 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 129691 -400 129747 240 0 FreeSans 560 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 131464 -400 131520 240 0 FreeSans 560 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 133237 -400 133293 240 0 FreeSans 560 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 69409 -400 69465 240 0 FreeSans 560 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 135010 -400 135066 240 0 FreeSans 560 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 136783 -400 136839 240 0 FreeSans 560 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 138556 -400 138612 240 0 FreeSans 560 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 140329 -400 140385 240 0 FreeSans 560 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 142102 -400 142158 240 0 FreeSans 560 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 143875 -400 143931 240 0 FreeSans 560 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 145648 -400 145704 240 0 FreeSans 560 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 147421 -400 147477 240 0 FreeSans 560 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 149194 -400 149250 240 0 FreeSans 560 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 150967 -400 151023 240 0 FreeSans 560 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 71182 -400 71238 240 0 FreeSans 560 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 152740 -400 152796 240 0 FreeSans 560 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 154513 -400 154569 240 0 FreeSans 560 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 156286 -400 156342 240 0 FreeSans 560 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 158059 -400 158115 240 0 FreeSans 560 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 159832 -400 159888 240 0 FreeSans 560 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 161605 -400 161661 240 0 FreeSans 560 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 163378 -400 163434 240 0 FreeSans 560 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 165151 -400 165207 240 0 FreeSans 560 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 166924 -400 166980 240 0 FreeSans 560 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 168697 -400 168753 240 0 FreeSans 560 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 72955 -400 73011 240 0 FreeSans 560 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 170470 -400 170526 240 0 FreeSans 560 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 172243 -400 172299 240 0 FreeSans 560 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 174016 -400 174072 240 0 FreeSans 560 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 175789 -400 175845 240 0 FreeSans 560 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 177562 -400 177618 240 0 FreeSans 560 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 179335 -400 179391 240 0 FreeSans 560 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 181108 -400 181164 240 0 FreeSans 560 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 182881 -400 182937 240 0 FreeSans 560 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 184654 -400 184710 240 0 FreeSans 560 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 186427 -400 186483 240 0 FreeSans 560 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 74728 -400 74784 240 0 FreeSans 560 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 188200 -400 188256 240 0 FreeSans 560 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 189973 -400 190029 240 0 FreeSans 560 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 191746 -400 191802 240 0 FreeSans 560 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 193519 -400 193575 240 0 FreeSans 560 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 195292 -400 195348 240 0 FreeSans 560 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 197065 -400 197121 240 0 FreeSans 560 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 198838 -400 198894 240 0 FreeSans 560 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 200611 -400 200667 240 0 FreeSans 560 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 202384 -400 202440 240 0 FreeSans 560 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 204157 -400 204213 240 0 FreeSans 560 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 76501 -400 76557 240 0 FreeSans 560 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 205930 -400 205986 240 0 FreeSans 560 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 207703 -400 207759 240 0 FreeSans 560 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 209476 -400 209532 240 0 FreeSans 560 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 211249 -400 211305 240 0 FreeSans 560 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 213022 -400 213078 240 0 FreeSans 560 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 214795 -400 214851 240 0 FreeSans 560 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 216568 -400 216624 240 0 FreeSans 560 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 218341 -400 218397 240 0 FreeSans 560 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 220114 -400 220170 240 0 FreeSans 560 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 221887 -400 221943 240 0 FreeSans 560 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 78274 -400 78330 240 0 FreeSans 560 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 223660 -400 223716 240 0 FreeSans 560 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 225433 -400 225489 240 0 FreeSans 560 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 227206 -400 227262 240 0 FreeSans 560 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 228979 -400 229035 240 0 FreeSans 560 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 230752 -400 230808 240 0 FreeSans 560 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 232525 -400 232581 240 0 FreeSans 560 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 234298 -400 234354 240 0 FreeSans 560 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 236071 -400 236127 240 0 FreeSans 560 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 237844 -400 237900 240 0 FreeSans 560 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 239617 -400 239673 240 0 FreeSans 560 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 80047 -400 80103 240 0 FreeSans 560 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 289852 -400 289908 240 0 FreeSans 560 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 290443 -400 290499 240 0 FreeSans 560 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 291034 -400 291090 240 0 FreeSans 560 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 291625 -400 291681 240 0 FreeSans 560 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 291170 319892 292400 322292 0 FreeSans 560 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 291170 314892 292400 317292 0 FreeSans 560 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 321921 830 324321 0 FreeSans 560 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 316921 830 319321 0 FreeSans 560 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 291170 270281 292400 272681 0 FreeSans 560 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 291170 275281 292400 277681 0 FreeSans 560 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 291170 117615 292400 120015 0 FreeSans 560 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 291170 112615 292400 115015 0 FreeSans 560 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 102444 830 104844 0 FreeSans 560 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 107444 830 109844 0 FreeSans 560 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 260297 351170 262697 352400 0 FreeSans 960 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 255297 351170 257697 352400 0 FreeSans 960 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 291170 73415 292400 75815 0 FreeSans 560 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 291170 68415 292400 70815 0 FreeSans 560 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 279721 830 282121 0 FreeSans 560 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 274721 830 277121 0 FreeSans 560 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 291170 95715 292400 98115 0 FreeSans 560 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 291170 90715 292400 93115 0 FreeSans 560 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 86444 830 88844 0 FreeSans 560 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 81444 830 83844 0 FreeSans 560 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 262 -400 318 240 0 FreeSans 560 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 853 -400 909 240 0 FreeSans 560 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 1444 -400 1500 240 0 FreeSans 560 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 3808 -400 3864 240 0 FreeSans 560 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 23902 -400 23958 240 0 FreeSans 560 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 25675 -400 25731 240 0 FreeSans 560 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 27448 -400 27504 240 0 FreeSans 560 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 29221 -400 29277 240 0 FreeSans 560 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 30994 -400 31050 240 0 FreeSans 560 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 32767 -400 32823 240 0 FreeSans 560 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 34540 -400 34596 240 0 FreeSans 560 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 36313 -400 36369 240 0 FreeSans 560 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 38086 -400 38142 240 0 FreeSans 560 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 39859 -400 39915 240 0 FreeSans 560 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 6172 -400 6228 240 0 FreeSans 560 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 41632 -400 41688 240 0 FreeSans 560 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 43405 -400 43461 240 0 FreeSans 560 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 45178 -400 45234 240 0 FreeSans 560 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 46951 -400 47007 240 0 FreeSans 560 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 48724 -400 48780 240 0 FreeSans 560 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 50497 -400 50553 240 0 FreeSans 560 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 52270 -400 52326 240 0 FreeSans 560 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 54043 -400 54099 240 0 FreeSans 560 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 55816 -400 55872 240 0 FreeSans 560 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 57589 -400 57645 240 0 FreeSans 560 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 8536 -400 8592 240 0 FreeSans 560 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 59362 -400 59418 240 0 FreeSans 560 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 61135 -400 61191 240 0 FreeSans 560 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 10900 -400 10956 240 0 FreeSans 560 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 13264 -400 13320 240 0 FreeSans 560 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 15037 -400 15093 240 0 FreeSans 560 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 16810 -400 16866 240 0 FreeSans 560 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 18583 -400 18639 240 0 FreeSans 560 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 20356 -400 20412 240 0 FreeSans 560 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 22129 -400 22185 240 0 FreeSans 560 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 2035 -400 2091 240 0 FreeSans 560 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 4399 -400 4455 240 0 FreeSans 560 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 24493 -400 24549 240 0 FreeSans 560 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 26266 -400 26322 240 0 FreeSans 560 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 28039 -400 28095 240 0 FreeSans 560 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 29812 -400 29868 240 0 FreeSans 560 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 31585 -400 31641 240 0 FreeSans 560 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 33358 -400 33414 240 0 FreeSans 560 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 35131 -400 35187 240 0 FreeSans 560 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 36904 -400 36960 240 0 FreeSans 560 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 38677 -400 38733 240 0 FreeSans 560 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 40450 -400 40506 240 0 FreeSans 560 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 6763 -400 6819 240 0 FreeSans 560 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 42223 -400 42279 240 0 FreeSans 560 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 43996 -400 44052 240 0 FreeSans 560 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 45769 -400 45825 240 0 FreeSans 560 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 47542 -400 47598 240 0 FreeSans 560 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 49315 -400 49371 240 0 FreeSans 560 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 51088 -400 51144 240 0 FreeSans 560 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 52861 -400 52917 240 0 FreeSans 560 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 54634 -400 54690 240 0 FreeSans 560 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 56407 -400 56463 240 0 FreeSans 560 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 58180 -400 58236 240 0 FreeSans 560 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 9127 -400 9183 240 0 FreeSans 560 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 59953 -400 60009 240 0 FreeSans 560 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 61726 -400 61782 240 0 FreeSans 560 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 11491 -400 11547 240 0 FreeSans 560 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 13855 -400 13911 240 0 FreeSans 560 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 15628 -400 15684 240 0 FreeSans 560 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 17401 -400 17457 240 0 FreeSans 560 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 19174 -400 19230 240 0 FreeSans 560 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 20947 -400 21003 240 0 FreeSans 560 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 22720 -400 22776 240 0 FreeSans 560 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 4990 -400 5046 240 0 FreeSans 560 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 25084 -400 25140 240 0 FreeSans 560 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 26857 -400 26913 240 0 FreeSans 560 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 28630 -400 28686 240 0 FreeSans 560 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 30403 -400 30459 240 0 FreeSans 560 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 32176 -400 32232 240 0 FreeSans 560 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 33949 -400 34005 240 0 FreeSans 560 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 35722 -400 35778 240 0 FreeSans 560 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 37495 -400 37551 240 0 FreeSans 560 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 39268 -400 39324 240 0 FreeSans 560 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 41041 -400 41097 240 0 FreeSans 560 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 7354 -400 7410 240 0 FreeSans 560 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 42814 -400 42870 240 0 FreeSans 560 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 44587 -400 44643 240 0 FreeSans 560 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 46360 -400 46416 240 0 FreeSans 560 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 48133 -400 48189 240 0 FreeSans 560 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 49906 -400 49962 240 0 FreeSans 560 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 51679 -400 51735 240 0 FreeSans 560 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 53452 -400 53508 240 0 FreeSans 560 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 55225 -400 55281 240 0 FreeSans 560 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 56998 -400 57054 240 0 FreeSans 560 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 58771 -400 58827 240 0 FreeSans 560 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 9718 -400 9774 240 0 FreeSans 560 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 60544 -400 60600 240 0 FreeSans 560 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 62317 -400 62373 240 0 FreeSans 560 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 12082 -400 12138 240 0 FreeSans 560 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 14446 -400 14502 240 0 FreeSans 560 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 16219 -400 16275 240 0 FreeSans 560 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 17992 -400 18048 240 0 FreeSans 560 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 19765 -400 19821 240 0 FreeSans 560 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 21538 -400 21594 240 0 FreeSans 560 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 23311 -400 23367 240 0 FreeSans 560 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 5581 -400 5637 240 0 FreeSans 560 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 7945 -400 8001 240 0 FreeSans 560 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 10309 -400 10365 240 0 FreeSans 560 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 12673 -400 12729 240 0 FreeSans 560 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 2626 -400 2682 240 0 FreeSans 560 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 3217 -400 3273 240 0 FreeSans 560 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 s 85447 351150 86547 352400 0 FreeSans 960 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 111297 351150 112397 352400 0 FreeSans 960 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 86697 351150 87797 352400 0 FreeSans 960 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 112547 351150 113647 352400 0 FreeSans 960 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal5 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 82797 351150 85297 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 108647 351150 111147 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 34097 351150 36597 352400 0 FreeSans 960 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 60097 351150 62597 352400 0 FreeSans 960 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal5 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 87947 351150 90447 352400 0 FreeSans 960 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 113797 351150 116297 352400 0 FreeSans 960 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 292000 352000
<< end >>
