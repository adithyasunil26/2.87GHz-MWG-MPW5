magic
tech sky130A
magscale 1 2
timestamp 1640959680
<< nwell >>
rect -250 320 6220 1010
rect -120 -750 190 -360
rect 2850 -750 3160 -360
rect 2858 -752 3160 -750
rect 5820 -760 6130 -370
<< nmos >>
rect -110 -20 -50 180
rect 2964 -20 3024 180
rect 6020 -20 6080 180
<< pmos >>
rect -110 360 -50 760
rect 2964 360 3024 760
rect 6020 360 6080 760
<< varactor >>
rect 17 -688 53 -488
rect 2991 -690 3027 -490
rect 5955 -694 5991 -494
<< ndiff >>
rect -210 150 -110 180
rect -210 110 -180 150
rect -140 110 -110 150
rect -210 50 -110 110
rect -210 10 -180 50
rect -140 10 -110 50
rect -210 -20 -110 10
rect -50 150 50 180
rect -50 110 -20 150
rect 20 110 50 150
rect -50 50 50 110
rect -50 10 -20 50
rect 20 10 50 50
rect -50 -20 50 10
rect 2864 150 2964 180
rect 2864 110 2892 150
rect 2932 110 2964 150
rect 2864 50 2964 110
rect 2864 10 2892 50
rect 2932 10 2964 50
rect 2864 -20 2964 10
rect 3024 150 3124 180
rect 3024 110 3052 150
rect 3092 110 3124 150
rect 3024 50 3124 110
rect 3024 10 3052 50
rect 3092 10 3124 50
rect 3024 -20 3124 10
rect 5920 150 6020 180
rect 5920 110 5952 150
rect 5992 110 6020 150
rect 5920 50 6020 110
rect 5920 10 5952 50
rect 5992 10 6020 50
rect 5920 -20 6020 10
rect 6080 150 6180 180
rect 6080 110 6112 150
rect 6152 110 6180 150
rect 6080 50 6180 110
rect 6080 10 6112 50
rect 6152 10 6180 50
rect 6080 -20 6180 10
<< pdiff >>
rect -210 730 -110 760
rect -210 690 -180 730
rect -140 690 -110 730
rect -210 640 -110 690
rect -210 600 -180 640
rect -140 600 -110 640
rect -210 540 -110 600
rect -210 500 -180 540
rect -140 500 -110 540
rect -210 440 -110 500
rect -210 400 -180 440
rect -140 400 -110 440
rect -210 360 -110 400
rect -50 730 50 760
rect -50 690 -20 730
rect 20 690 50 730
rect -50 640 50 690
rect -50 600 -20 640
rect 20 600 50 640
rect -50 540 50 600
rect -50 500 -20 540
rect 20 500 50 540
rect -50 440 50 500
rect -50 400 -20 440
rect 20 400 50 440
rect -50 360 50 400
rect 2864 730 2964 760
rect 2864 690 2892 730
rect 2932 690 2964 730
rect 2864 640 2964 690
rect 2864 600 2892 640
rect 2932 600 2964 640
rect 2864 540 2964 600
rect 2864 500 2892 540
rect 2932 500 2964 540
rect 2864 440 2964 500
rect 2864 400 2892 440
rect 2932 400 2964 440
rect 2864 360 2964 400
rect 3024 730 3124 760
rect 3024 690 3052 730
rect 3092 690 3124 730
rect 3024 640 3124 690
rect 3024 600 3052 640
rect 3092 600 3124 640
rect 3024 540 3124 600
rect 3024 500 3052 540
rect 3092 500 3124 540
rect 3024 440 3124 500
rect 3024 400 3052 440
rect 3092 400 3124 440
rect 3024 360 3124 400
rect 5920 730 6020 760
rect 5920 690 5952 730
rect 5992 690 6020 730
rect 5920 640 6020 690
rect 5920 600 5952 640
rect 5992 600 6020 640
rect 5920 540 6020 600
rect 5920 500 5952 540
rect 5992 500 6020 540
rect 5920 440 6020 500
rect 5920 400 5952 440
rect 5992 400 6020 440
rect 5920 360 6020 400
rect 6080 730 6180 760
rect 6080 690 6112 730
rect 6152 690 6180 730
rect 6080 640 6180 690
rect 6080 600 6112 640
rect 6152 600 6180 640
rect 6080 540 6180 600
rect 6080 500 6112 540
rect 6152 500 6180 540
rect 6080 440 6180 500
rect 6080 400 6112 440
rect 6152 400 6180 440
rect 6080 360 6180 400
<< ndiffc >>
rect -180 110 -140 150
rect -180 10 -140 50
rect -20 110 20 150
rect -20 10 20 50
rect 2892 110 2932 150
rect 2892 10 2932 50
rect 3052 110 3092 150
rect 3052 10 3092 50
rect 5952 110 5992 150
rect 5952 10 5992 50
rect 6112 110 6152 150
rect 6112 10 6152 50
<< pdiffc >>
rect -180 690 -140 730
rect -180 600 -140 640
rect -180 500 -140 540
rect -180 400 -140 440
rect -20 690 20 730
rect -20 600 20 640
rect -20 500 20 540
rect -20 400 20 440
rect 2892 690 2932 730
rect 2892 600 2932 640
rect 2892 500 2932 540
rect 2892 400 2932 440
rect 3052 690 3092 730
rect 3052 600 3092 640
rect 3052 500 3092 540
rect 3052 400 3092 440
rect 5952 690 5992 730
rect 5952 600 5992 640
rect 5952 500 5992 540
rect 5952 400 5992 440
rect 6112 690 6152 730
rect 6112 600 6152 640
rect 6112 500 6152 540
rect 6112 400 6152 440
<< psubdiff >>
rect -350 1470 -90 1500
rect -710 1300 -450 1330
rect -710 1100 -680 1300
rect -480 1100 -450 1300
rect -350 1270 -320 1470
rect -120 1270 -90 1470
rect -350 1240 -90 1270
rect 630 1470 890 1500
rect 630 1270 660 1470
rect 860 1270 890 1470
rect 630 1240 890 1270
rect 1610 1470 1870 1500
rect 1610 1270 1640 1470
rect 1840 1270 1870 1470
rect 1610 1240 1870 1270
rect 2590 1470 2850 1500
rect 2590 1270 2620 1470
rect 2820 1270 2850 1470
rect 2590 1240 2850 1270
rect 3570 1470 3830 1500
rect 3570 1270 3600 1470
rect 3800 1270 3830 1470
rect 3570 1240 3830 1270
rect 4550 1470 4810 1500
rect 4550 1270 4580 1470
rect 4780 1270 4810 1470
rect 4550 1240 4810 1270
rect 5530 1470 5790 1500
rect 5530 1270 5560 1470
rect 5760 1270 5790 1470
rect 5530 1240 5790 1270
rect 6510 1470 6770 1500
rect 6510 1270 6540 1470
rect 6740 1270 6770 1470
rect 6510 1240 6770 1270
rect 7270 1300 7530 1330
rect -710 1070 -450 1100
rect 7270 1100 7300 1300
rect 7500 1100 7530 1300
rect 7270 1070 7530 1100
rect -710 320 -450 350
rect -710 120 -680 320
rect -480 120 -450 320
rect 7270 320 7530 350
rect -710 90 -450 120
rect 7270 120 7300 320
rect 7500 120 7530 320
rect 7270 90 7530 120
rect 0 -120 230 -90
rect 0 -170 30 -120
rect 200 -170 230 -120
rect 0 -200 230 -170
rect 2824 -120 3124 -90
rect 2824 -180 2854 -120
rect 3094 -180 3124 -120
rect 2824 -200 3124 -180
rect 5670 -120 5900 -90
rect 5670 -170 5700 -120
rect 5870 -170 5900 -120
rect 5670 -200 5900 -170
rect 2624 -270 2754 -240
rect 2624 -340 2654 -270
rect 2724 -340 2754 -270
rect 2624 -370 2754 -340
rect -710 -660 -450 -630
rect -710 -860 -680 -660
rect -480 -860 -450 -660
rect 2624 -650 2754 -620
rect 2624 -720 2654 -650
rect 2724 -720 2754 -650
rect 7270 -660 7530 -630
rect 2624 -750 2754 -720
rect -710 -890 -450 -860
rect 7270 -860 7300 -660
rect 7500 -860 7530 -660
rect 7270 -890 7530 -860
rect -320 -920 -60 -890
rect -320 -1120 -290 -920
rect -90 -1120 -60 -920
rect -320 -1150 -60 -1120
rect 660 -920 920 -890
rect 660 -1120 690 -920
rect 890 -1120 920 -920
rect 660 -1150 920 -1120
rect 1640 -920 1900 -890
rect 1640 -1120 1670 -920
rect 1870 -1120 1900 -920
rect 1640 -1150 1900 -1120
rect 2620 -920 2880 -890
rect 2620 -1120 2650 -920
rect 2850 -1120 2880 -920
rect 2620 -1150 2880 -1120
rect 3600 -920 3860 -890
rect 3600 -1120 3630 -920
rect 3830 -1120 3860 -920
rect 3600 -1150 3860 -1120
rect 4580 -920 4840 -890
rect 4580 -1120 4610 -920
rect 4810 -1120 4840 -920
rect 4580 -1150 4840 -1120
rect 5560 -920 5820 -890
rect 5560 -1120 5590 -920
rect 5790 -1120 5820 -920
rect 5560 -1150 5820 -1120
rect 6540 -920 6800 -890
rect 6540 -1120 6570 -920
rect 6770 -1120 6800 -920
rect 6540 -1150 6800 -1120
<< nsubdiff >>
rect 174 950 494 970
rect 174 880 204 950
rect 464 880 494 950
rect 174 860 494 880
rect 2834 950 3154 970
rect 2834 880 2864 950
rect 3124 880 3154 950
rect 2834 860 3154 880
rect 5244 950 5564 970
rect 5244 880 5274 950
rect 5534 880 5564 950
rect 5244 860 5564 880
rect -80 -512 17 -488
rect -80 -664 -68 -512
rect -34 -664 17 -512
rect -80 -688 17 -664
rect 53 -512 150 -488
rect 53 -664 104 -512
rect 138 -664 150 -512
rect 2894 -514 2991 -490
rect 53 -688 150 -664
rect 2894 -666 2906 -514
rect 2940 -666 2991 -514
rect 2894 -690 2991 -666
rect 3027 -514 3124 -490
rect 3027 -666 3078 -514
rect 3112 -666 3124 -514
rect 3027 -690 3124 -666
rect 5858 -518 5955 -494
rect 5858 -670 5870 -518
rect 5904 -670 5955 -518
rect 5858 -694 5955 -670
rect 5991 -518 6088 -494
rect 5991 -670 6042 -518
rect 6076 -670 6088 -518
rect 5991 -694 6088 -670
<< psubdiffcont >>
rect -680 1100 -480 1300
rect -320 1270 -120 1470
rect 660 1270 860 1470
rect 1640 1270 1840 1470
rect 2620 1270 2820 1470
rect 3600 1270 3800 1470
rect 4580 1270 4780 1470
rect 5560 1270 5760 1470
rect 6540 1270 6740 1470
rect 7300 1100 7500 1300
rect -680 120 -480 320
rect 7300 120 7500 320
rect 30 -170 200 -120
rect 2854 -180 3094 -120
rect 5700 -170 5870 -120
rect 2654 -340 2724 -270
rect -680 -860 -480 -660
rect 2654 -720 2724 -650
rect 7300 -860 7500 -660
rect -290 -1120 -90 -920
rect 690 -1120 890 -920
rect 1670 -1120 1870 -920
rect 2650 -1120 2850 -920
rect 3630 -1120 3830 -920
rect 4610 -1120 4810 -920
rect 5590 -1120 5790 -920
rect 6570 -1120 6770 -920
<< nsubdiffcont >>
rect 204 880 464 950
rect 2864 880 3124 950
rect 5274 880 5534 950
rect -68 -664 -34 -512
rect 104 -664 138 -512
rect 2906 -666 2940 -514
rect 3078 -666 3112 -514
rect 5870 -670 5904 -518
rect 6042 -670 6076 -518
<< poly >>
rect -110 760 -50 790
rect 2964 760 3024 790
rect 6020 760 6080 790
rect -110 300 -50 360
rect 2964 300 3024 360
rect 6020 300 6080 360
rect -190 280 -50 300
rect -190 240 -170 280
rect -130 240 -50 280
rect -190 220 -50 240
rect 2884 280 3024 300
rect 2884 240 2904 280
rect 2944 240 3024 280
rect 2884 220 3024 240
rect 5940 280 6080 300
rect 5940 240 5960 280
rect 6000 240 6080 280
rect 5940 220 6080 240
rect -110 180 -50 220
rect 2964 180 3024 220
rect 6020 180 6080 220
rect -110 -50 -50 -20
rect 2964 -50 3024 -20
rect 6020 -50 6080 -20
rect 2 -416 68 -400
rect 2 -450 18 -416
rect 52 -450 68 -416
rect 2 -466 68 -450
rect 2976 -418 3042 -402
rect 2976 -452 2992 -418
rect 3026 -452 3042 -418
rect 17 -488 53 -466
rect 2976 -468 3042 -452
rect 5940 -422 6006 -406
rect 5940 -456 5956 -422
rect 5990 -456 6006 -422
rect 2991 -490 3027 -468
rect 5940 -472 6006 -456
rect 17 -714 53 -688
rect 5955 -494 5991 -472
rect 2991 -716 3027 -690
rect 5955 -720 5991 -694
<< polycont >>
rect -170 240 -130 280
rect 2904 240 2944 280
rect 5960 240 6000 280
rect 18 -450 52 -416
rect 2992 -452 3026 -418
rect 5956 -456 5990 -422
<< locali >>
rect -750 1470 7560 1530
rect -750 1300 -320 1470
rect -750 1100 -680 1300
rect -480 1270 -320 1300
rect -120 1270 660 1470
rect 860 1270 1640 1470
rect 1840 1270 2620 1470
rect 2820 1270 3600 1470
rect 3800 1270 4580 1470
rect 4780 1270 5560 1470
rect 5760 1270 6540 1470
rect 6740 1300 7560 1470
rect 6740 1270 7300 1300
rect -480 1200 7300 1270
rect -480 1100 -420 1200
rect -750 320 -420 1100
rect 7230 1100 7300 1200
rect 7500 1100 7560 1300
rect -250 950 6220 1010
rect -250 880 204 950
rect 464 880 2864 950
rect 3124 880 5274 950
rect 5534 880 6220 950
rect -250 830 6220 880
rect -200 730 -120 830
rect 2874 750 2954 830
rect 5930 750 6010 830
rect -200 690 -180 730
rect -140 690 -120 730
rect -200 640 -120 690
rect -200 600 -180 640
rect -140 600 -120 640
rect -200 540 -120 600
rect -200 500 -180 540
rect -140 500 -120 540
rect -200 440 -120 500
rect -200 400 -180 440
rect -140 400 -120 440
rect -200 370 -120 400
rect -40 730 40 750
rect -40 690 -20 730
rect 20 690 40 730
rect -40 640 40 690
rect -40 600 -20 640
rect 20 600 40 640
rect -40 540 40 600
rect -40 500 -20 540
rect 20 500 40 540
rect -40 440 40 500
rect -40 400 -20 440
rect 20 400 40 440
rect -750 120 -680 320
rect -480 120 -420 320
rect -190 290 -110 300
rect -190 230 -180 290
rect -120 230 -110 290
rect -190 220 -110 230
rect -40 290 40 400
rect 2872 730 2954 750
rect 2872 690 2892 730
rect 2932 690 2954 730
rect 2872 640 2954 690
rect 2872 600 2892 640
rect 2932 600 2954 640
rect 2872 540 2954 600
rect 2872 500 2892 540
rect 2932 500 2954 540
rect 2872 440 2954 500
rect 2872 400 2892 440
rect 2932 400 2954 440
rect 2872 370 2954 400
rect 3032 730 3114 750
rect 3032 690 3052 730
rect 3092 690 3114 730
rect 3032 640 3114 690
rect 3032 600 3052 640
rect 3092 600 3114 640
rect 3032 540 3114 600
rect 3032 500 3052 540
rect 3092 500 3114 540
rect 3032 440 3114 500
rect 3032 400 3052 440
rect 3092 400 3114 440
rect 3032 370 3114 400
rect 5930 730 6012 750
rect 5930 690 5952 730
rect 5992 690 6012 730
rect 5930 640 6012 690
rect 5930 600 5952 640
rect 5992 600 6012 640
rect 5930 540 6012 600
rect 5930 500 5952 540
rect 5992 500 6012 540
rect 5930 440 6012 500
rect 5930 400 5952 440
rect 5992 400 6012 440
rect 5930 370 6012 400
rect 6090 730 6172 750
rect 6090 690 6112 730
rect 6152 690 6172 730
rect 6090 640 6172 690
rect 6090 600 6112 640
rect 6152 600 6172 640
rect 6090 540 6172 600
rect 6090 500 6112 540
rect 6152 500 6172 540
rect 6090 440 6172 500
rect 6090 400 6112 440
rect 6152 400 6172 440
rect 6090 370 6172 400
rect -40 230 2884 290
rect -750 -660 -420 120
rect -200 150 -120 170
rect -200 110 -180 150
rect -140 110 -120 150
rect -200 50 -120 110
rect -200 10 -180 50
rect -140 10 -120 50
rect -200 -80 -120 10
rect -40 150 40 230
rect 3034 290 3114 370
rect 6090 310 6170 370
rect 7230 320 7560 1100
rect 3034 230 5940 290
rect 3034 170 3114 230
rect 6090 210 6190 310
rect 6090 170 6170 210
rect -40 110 -20 150
rect 20 110 40 150
rect -40 50 40 110
rect -40 10 -20 50
rect 20 10 40 50
rect -40 -10 40 10
rect 2872 150 2954 170
rect 2872 110 2892 150
rect 2932 110 2954 150
rect 2872 50 2954 110
rect 2872 10 2892 50
rect 2932 10 2954 50
rect 2872 -10 2954 10
rect 3032 150 3114 170
rect 3032 110 3052 150
rect 3092 110 3114 150
rect 3032 50 3114 110
rect 3032 10 3052 50
rect 3092 10 3114 50
rect 3032 -10 3114 10
rect 5930 150 6012 170
rect 5930 110 5952 150
rect 5992 110 6012 150
rect 5930 50 6012 110
rect 5930 10 5952 50
rect 5992 10 6012 50
rect 5930 -10 6012 10
rect 6090 150 6172 170
rect 6090 110 6112 150
rect 6152 110 6172 150
rect 6090 50 6172 110
rect 6090 10 6112 50
rect 6152 10 6172 50
rect 6090 -10 6172 10
rect 7230 120 7300 320
rect 7500 120 7560 320
rect 2874 -80 2954 -10
rect 5930 -80 6010 -10
rect -230 -120 6220 -80
rect -230 -170 30 -120
rect 200 -170 2854 -120
rect -230 -180 2854 -170
rect 3094 -170 5700 -120
rect 5870 -170 6220 -120
rect 3094 -180 6220 -170
rect -230 -220 6220 -180
rect 2614 -270 2764 -220
rect 2614 -340 2654 -270
rect 2724 -340 2764 -270
rect 2 -450 18 -416
rect 52 -450 68 -416
rect -750 -860 -680 -660
rect -480 -860 -420 -660
rect -68 -512 -34 -496
rect -68 -680 -34 -664
rect 104 -512 138 -496
rect 104 -680 138 -664
rect 2614 -650 2764 -340
rect 2976 -452 2992 -418
rect 3026 -452 3042 -418
rect 5940 -456 5956 -422
rect 5990 -456 6006 -422
rect 2614 -720 2654 -650
rect 2724 -720 2764 -650
rect 2906 -514 2940 -498
rect 2906 -682 2940 -666
rect 3078 -514 3112 -498
rect 3078 -682 3112 -666
rect 5870 -518 5904 -502
rect 5870 -686 5904 -670
rect 6042 -518 6076 -502
rect 6042 -686 6076 -670
rect 6256 -680 6290 -510
rect 7230 -660 7560 120
rect 2614 -800 2764 -720
rect 2620 -860 2750 -800
rect 7230 -860 7300 -660
rect 7500 -860 7560 -660
rect -750 -920 7560 -860
rect -750 -1120 -290 -920
rect -90 -1120 690 -920
rect 890 -1120 1670 -920
rect 1870 -1120 2650 -920
rect 2850 -1120 3630 -920
rect 3830 -1120 4610 -920
rect 4810 -1120 5590 -920
rect 5790 -1120 6570 -920
rect 6770 -1120 7560 -920
rect -750 -1190 7560 -1120
<< viali >>
rect -180 280 -120 290
rect -180 240 -170 280
rect -170 240 -130 280
rect -130 240 -120 280
rect -180 230 -120 240
rect 2884 280 2964 300
rect 2884 240 2904 280
rect 2904 240 2944 280
rect 2944 240 2964 280
rect 2884 220 2964 240
rect 5940 280 6020 300
rect 5940 240 5960 280
rect 5960 240 6000 280
rect 6000 240 6020 280
rect 5940 220 6020 240
rect 6190 230 6250 290
rect 18 -450 52 -416
rect -68 -664 -34 -512
rect 104 -664 138 -512
rect 2992 -452 3026 -418
rect 5956 -456 5990 -422
rect 2906 -666 2940 -514
rect 3078 -666 3112 -514
rect 5870 -670 5904 -518
rect 6042 -670 6076 -518
<< metal1 >>
rect -200 290 -110 310
rect -200 230 -180 290
rect -120 230 -110 290
rect -200 210 -110 230
rect 2594 300 2984 310
rect 2594 220 2884 300
rect 2964 220 2984 300
rect 2594 210 2984 220
rect 5570 300 6040 310
rect 5570 220 5940 300
rect 6020 220 6040 300
rect 5570 210 6040 220
rect 6170 290 6270 310
rect 6170 230 6190 290
rect 6250 230 6270 290
rect 2594 -100 2694 210
rect -10 -200 2694 -100
rect -10 -416 90 -200
rect 5570 -260 5670 210
rect 6170 170 6270 230
rect 6172 -10 6270 170
rect 6170 -100 6270 -10
rect -10 -450 18 -416
rect 52 -450 90 -416
rect -10 -470 90 -450
rect 2964 -308 5670 -260
rect 5920 -200 6270 -100
rect 2964 -418 3064 -308
rect 2964 -452 2992 -418
rect 3026 -452 3064 -418
rect 2964 -470 3064 -452
rect 5920 -422 6020 -200
rect 5920 -456 5956 -422
rect 5990 -456 6020 -422
rect 5920 -470 6020 -456
rect -130 -512 6276 -500
rect -130 -664 -68 -512
rect -34 -664 104 -512
rect 138 -514 6276 -512
rect 138 -664 2906 -514
rect -130 -666 2906 -664
rect 2940 -666 3078 -514
rect 3112 -518 6276 -514
rect 3112 -666 5870 -518
rect -130 -670 5870 -666
rect 5904 -670 6042 -518
rect 6076 -670 6276 -518
rect -130 -680 6276 -670
rect 5864 -682 5910 -680
rect 6036 -682 6082 -680
<< via1 >>
rect -180 230 -120 290
rect 6190 230 6250 290
<< metal2 >>
rect -200 290 6270 310
rect -200 230 -180 290
rect -120 230 6190 290
rect 6250 230 6270 290
rect -200 210 6270 230
<< labels >>
rlabel locali 10 200 10 200 1 out1
rlabel locali 3074 190 3074 190 1 out2
rlabel locali 5980 -160 5980 -160 1 gnd
rlabel viali 6220 260 6220 260 1 out3
rlabel locali 6130 190 6130 190 1 out3
rlabel locali 6286 -610 6286 -610 1 vcont
rlabel locali 6020 900 6020 900 1 vdd
<< end >>
