magic
tech sky130A
timestamp 1643048290
<< nwell >>
rect -3185 7805 -3090 9815
rect -3290 7585 -2985 7805
<< nsubdiff >>
rect -3210 7755 -3065 7770
rect -3210 7645 -3195 7755
rect -3080 7645 -3065 7755
rect -3210 7635 -3065 7645
<< nsubdiffcont >>
rect -3195 7645 -3080 7755
<< locali >>
rect 1861 10772 2085 11271
rect 3136 10783 3360 11282
rect 4565 10810 4789 11309
rect 6163 10788 6387 11287
rect 7803 9114 8347 9515
rect -3205 7755 -3070 7765
rect -3205 7645 -3195 7755
rect -3080 7645 -3070 7755
rect -3205 7640 -3070 7645
rect 7885 6690 8734 6954
rect -5053 5917 -4915 6349
rect -4015 5926 -3823 6332
rect 7861 4862 8710 5126
rect -4902 4072 -4702 4384
rect -4254 4037 -3882 4394
rect -331 3685 129 3956
rect -378 2878 294 3207
rect 7909 3059 8758 3323
rect -331 2025 129 2296
rect 535 -1232 958 -444
rect 1849 -1174 2272 -386
rect 3309 -1203 3732 -415
rect 5047 -1217 5470 -429
rect 6493 -1217 6916 -429
rect -5150 -1610 -5145 -1590
rect -5215 -2120 -5140 -2100
<< viali >>
rect -4970 12335 -4950 12355
rect -4805 7745 -4785 7765
rect -3195 7645 -3080 7755
rect -4805 7395 -4785 7415
rect -515 2395 -490 2420
rect -5170 -1610 -5150 -1590
rect -5235 -2120 -5215 -2100
<< metal1 >>
rect -4980 12360 -4940 12365
rect -4980 12330 -4975 12360
rect -4945 12330 -4940 12360
rect -4980 12325 -4940 12330
rect 380 9245 4010 9380
rect 4015 9245 8130 9370
rect -4815 7770 -4775 7775
rect -4815 7740 -4810 7770
rect -4780 7740 -4775 7770
rect -4815 7735 -4775 7740
rect -3205 7755 -3070 7765
rect -3205 7645 -3195 7755
rect -3080 7645 -3070 7755
rect -3205 7640 -3070 7645
rect 380 7630 460 9245
rect 8055 8900 8130 9245
rect 8055 8810 8565 8900
rect 8055 8805 8130 8810
rect -595 7510 465 7630
rect 380 7505 460 7510
rect -4815 7420 -4775 7425
rect -4815 7390 -4810 7420
rect -4780 7390 -4775 7420
rect -4815 7385 -4775 7390
rect -3320 5535 -3275 5540
rect -3320 5530 -3315 5535
rect -3375 5515 -3315 5530
rect -3320 5500 -3315 5515
rect -3280 5500 -3275 5535
rect -3320 5495 -3275 5500
rect -3320 5405 -3275 5410
rect -3320 5395 -3315 5405
rect -3375 5380 -3315 5395
rect -3320 5370 -3315 5380
rect -3280 5370 -3275 5405
rect -3320 5365 -3275 5370
rect -525 2425 -480 2430
rect -525 2390 -520 2425
rect -485 2390 -480 2425
rect -525 2385 -480 2390
rect -5180 -1585 -5140 -1580
rect -5180 -1615 -5175 -1585
rect -5145 -1615 -5140 -1585
rect -5180 -1620 -5140 -1615
rect -5245 -2095 -5205 -2090
rect -5245 -2125 -5240 -2095
rect -5210 -2125 -5205 -2095
rect -5245 -2130 -5205 -2125
<< via1 >>
rect -4975 12355 -4945 12360
rect -4975 12335 -4970 12355
rect -4970 12335 -4950 12355
rect -4950 12335 -4945 12355
rect -4975 12330 -4945 12335
rect -4810 7765 -4780 7770
rect -4810 7745 -4805 7765
rect -4805 7745 -4785 7765
rect -4785 7745 -4780 7765
rect -4810 7740 -4780 7745
rect -3195 7645 -3080 7755
rect -4810 7415 -4780 7420
rect -4810 7395 -4805 7415
rect -4805 7395 -4785 7415
rect -4785 7395 -4780 7415
rect -4810 7390 -4780 7395
rect -3315 5500 -3280 5535
rect -3315 5370 -3280 5405
rect -520 2420 -485 2425
rect -520 2395 -515 2420
rect -515 2395 -490 2420
rect -490 2395 -485 2420
rect -520 2390 -485 2395
rect -5175 -1590 -5145 -1585
rect -5175 -1610 -5170 -1590
rect -5170 -1610 -5150 -1590
rect -5150 -1610 -5145 -1590
rect -5175 -1615 -5145 -1610
rect -5240 -2100 -5210 -2095
rect -5240 -2120 -5235 -2100
rect -5235 -2120 -5215 -2100
rect -5215 -2120 -5210 -2100
rect -5240 -2125 -5210 -2120
<< metal2 >>
rect -4985 12360 -4935 12370
rect -4985 12355 -4975 12360
rect -5055 12335 -4975 12355
rect -5055 11420 -5025 12335
rect -4985 12330 -4975 12335
rect -4945 12330 -4935 12360
rect -4985 12320 -4935 12330
rect -5055 11395 -4780 11420
rect -4810 8120 -4780 11395
rect -5120 8090 -4780 8120
rect -5120 5590 -5100 8090
rect -4820 7775 -4770 7780
rect -4820 7735 -4815 7775
rect -4775 7735 -4770 7775
rect -4820 7730 -4770 7735
rect -3205 7755 -3070 7765
rect -3205 7645 -3195 7755
rect -3080 7645 -3070 7755
rect -3205 7640 -3070 7645
rect -4820 7420 -4770 7430
rect -4820 7390 -4810 7420
rect -4780 7390 -4770 7420
rect -4820 7380 -4770 7390
rect -4815 6070 -4770 7380
rect -4815 6035 -3270 6070
rect -5120 5575 -4960 5590
rect -3305 5545 -3270 6035
rect -3325 5535 -3270 5545
rect -3325 5500 -3315 5535
rect -3280 5500 -3270 5535
rect -3325 5490 -3270 5500
rect -3325 5405 -3270 5415
rect -3325 5370 -3315 5405
rect -3280 5370 -3270 5405
rect -3325 5360 -3270 5370
rect -5250 4720 -4960 4740
rect -5250 -2095 -5200 4720
rect 12130 4220 12260 4935
rect -5160 4185 12260 4220
rect -5160 2435 -5140 4185
rect -4675 3800 -4625 3810
rect -4675 3770 -4665 3800
rect -4635 3770 -4625 3800
rect -4675 3760 -4625 3770
rect -5160 2415 -5095 2435
rect -530 2425 -475 2435
rect -530 2390 -520 2425
rect -485 2390 -475 2425
rect -530 2380 -475 2390
rect -525 1990 -490 2380
rect -5165 1950 -490 1990
rect -5165 -1575 -5135 1950
rect -5185 -1585 -5135 -1575
rect -5185 -1615 -5175 -1585
rect -5145 -1615 -5135 -1585
rect -5185 -1625 -5135 -1615
rect -5250 -2125 -5240 -2095
rect -5210 -2125 -5200 -2095
rect -5250 -2135 -5200 -2125
<< via2 >>
rect -4815 7770 -4775 7775
rect -4815 7740 -4810 7770
rect -4810 7740 -4780 7770
rect -4780 7740 -4775 7770
rect -4815 7735 -4775 7740
rect -3195 7645 -3080 7755
rect -3315 5370 -3280 5405
rect -4665 3770 -4635 3800
<< metal3 >>
rect -4825 7775 -4765 7785
rect -4825 7735 -4815 7775
rect -4775 7735 -4765 7775
rect -4825 7725 -4765 7735
rect -3290 7755 -2985 7805
rect -4820 7630 -4785 7725
rect -4850 7600 -4785 7630
rect -3290 7645 -3195 7755
rect -3080 7645 -2985 7755
rect -4850 6110 -4815 7600
rect -3290 7585 -2985 7645
rect -4850 6080 -3270 6110
rect -3305 5415 -3270 6080
rect -3325 5405 -3270 5415
rect -3325 5370 -3315 5405
rect -3280 5370 -3270 5405
rect -3325 5360 -3270 5370
rect -4675 3805 -4625 3810
rect -4675 3765 -4670 3805
rect -4630 3765 -4625 3805
rect -4675 3760 -4625 3765
<< via3 >>
rect -3195 7645 -3080 7755
rect -4670 3800 -4630 3805
rect -4670 3770 -4665 3800
rect -4665 3770 -4635 3800
rect -4635 3770 -4630 3800
rect -4670 3765 -4630 3770
<< metal4 >>
rect -4300 11109 -4121 11506
rect -4300 11104 -4118 11109
rect -5794 10779 -5174 10780
rect -4297 10779 -4118 11104
rect -5794 10672 -4118 10779
rect -3896 10672 -3715 10673
rect -5794 10513 -3715 10672
rect -876 10547 -693 11511
rect -876 10528 -692 10547
rect -5794 10509 -4166 10513
rect -5794 10504 -5174 10509
rect -5790 5810 -5439 10504
rect -3896 10488 -3715 10513
rect -3895 10110 -3716 10488
rect -3898 10099 -3716 10110
rect -3898 9708 -3719 10099
rect -3185 7780 -3090 9815
rect -875 9707 -692 10528
rect -3210 7755 -3055 7780
rect -3210 7645 -3195 7755
rect -3080 7645 -3055 7755
rect -3210 7625 -3055 7645
rect -5790 5720 -4891 5810
rect -5790 3260 -5439 5720
rect -4660 3860 -4595 3900
rect -4660 3810 -4625 3860
rect -4675 3805 -4625 3810
rect -4675 3765 -4670 3805
rect -4630 3765 -4625 3805
rect -4675 3760 -4625 3765
rect -5791 3090 -4643 3260
use divider  divider_0
timestamp 1643048290
transform 1 0 -4910 0 1 1985
box -490 -235 4690 2150
use cp  cp_0
timestamp 1640911461
transform 1 0 -4895 0 1 7840
box -415 -1715 4690 2035
use pd  pd_0
timestamp 1643048290
transform 1 0 -4845 0 1 5180
box -215 -855 1685 810
use ro_complete  ro_complete_0
timestamp 1643048290
transform 1 0 8137 0 1 8475
box -57 -5330 4455 1440
use filter  filter_0
timestamp 1640983258
transform 1 0 1800 0 1 10450
box -1800 -11005 6240 390
use divbuf  divbuf_1
timestamp 1641017053
transform 1 0 -4770 0 1 12340
box -460 -1085 31200 495
use divbuf  divbuf_0
timestamp 1641017053
transform 1 0 -4955 0 1 -1605
box -460 -1085 31200 495
<< labels >>
rlabel locali -3140 7755 -3140 7755 1 vdd!
<< end >>
